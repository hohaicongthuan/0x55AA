module layer_10_featuremap_409(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76a662),
	.w1(32'hbbc48830),
	.w2(32'hbbc6542d),
	.w3(32'h3b028d87),
	.w4(32'hbbbee646),
	.w5(32'hbbb1ba8c),
	.w6(32'hbb16ca0a),
	.w7(32'hbb9c760c),
	.w8(32'hbbd968b8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba818f3),
	.w1(32'h3c60da13),
	.w2(32'h3ba9e465),
	.w3(32'h3aad0310),
	.w4(32'h3bc8828d),
	.w5(32'h3c1b2526),
	.w6(32'hbbf6d53c),
	.w7(32'hbae6fb39),
	.w8(32'h3c020bdb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68005a),
	.w1(32'hbb15a191),
	.w2(32'hbbf74ae5),
	.w3(32'hbc4789b3),
	.w4(32'hba27e639),
	.w5(32'hbb2d3c3b),
	.w6(32'hbbcedb64),
	.w7(32'hbb36d88b),
	.w8(32'hbb93667e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba99b7),
	.w1(32'hbc579202),
	.w2(32'h3b5ea3b9),
	.w3(32'hbc265078),
	.w4(32'hbc7f9245),
	.w5(32'h3b159b5e),
	.w6(32'hbc07f3d0),
	.w7(32'hbc284ba1),
	.w8(32'h3b73857b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97584),
	.w1(32'hbbb117dc),
	.w2(32'hbc032ff4),
	.w3(32'hbac2ecf9),
	.w4(32'hbbfe9f8b),
	.w5(32'hbac0a644),
	.w6(32'hbb98bb20),
	.w7(32'hbb2715a8),
	.w8(32'hbad89762),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65af59),
	.w1(32'h3b83f9b1),
	.w2(32'hbb9ddc9f),
	.w3(32'hbb92fc27),
	.w4(32'hba5a8edf),
	.w5(32'h3b6f4a1a),
	.w6(32'h37ff326a),
	.w7(32'h3a19f20e),
	.w8(32'hba580c39),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba723179),
	.w1(32'h3c1552e5),
	.w2(32'hba344ae7),
	.w3(32'h3b15c8dd),
	.w4(32'h3c41c384),
	.w5(32'h3ba08665),
	.w6(32'h3b90ba4a),
	.w7(32'h3ad0a577),
	.w8(32'h3bc14a76),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb399bc8),
	.w1(32'h3b9980d7),
	.w2(32'h3bb72865),
	.w3(32'h3c030c1a),
	.w4(32'h3bbc7960),
	.w5(32'hbc2b329c),
	.w6(32'h3bc442ec),
	.w7(32'h3c03d659),
	.w8(32'h3b1fcdec),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42e56a),
	.w1(32'hbbfb075f),
	.w2(32'h3b28ff5c),
	.w3(32'h3ae4ef15),
	.w4(32'hbc233ab0),
	.w5(32'h3c51d469),
	.w6(32'h3bb4657f),
	.w7(32'h39973e0d),
	.w8(32'h3a6b9c8d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae167af),
	.w1(32'hbc0fd0ec),
	.w2(32'h3ab2a3b8),
	.w3(32'h3affc212),
	.w4(32'hbc039ef4),
	.w5(32'h3ad2f136),
	.w6(32'hbbdecd6d),
	.w7(32'h3b799573),
	.w8(32'h3b50eb66),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046b3b),
	.w1(32'hb9becfa5),
	.w2(32'h3aa86d64),
	.w3(32'h3c336253),
	.w4(32'h3b985350),
	.w5(32'h3c4e9049),
	.w6(32'h3941ac85),
	.w7(32'hbb6a289a),
	.w8(32'hbba0458e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3543b5),
	.w1(32'hbba5fc0d),
	.w2(32'hbbb9255d),
	.w3(32'h3c10f817),
	.w4(32'hbb180b9a),
	.w5(32'hbbf6c539),
	.w6(32'h3bfc724e),
	.w7(32'h3ad3979e),
	.w8(32'h3a5d3458),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37dc26),
	.w1(32'h3c14456c),
	.w2(32'h3cd66da7),
	.w3(32'hbc431678),
	.w4(32'h3c05a1cb),
	.w5(32'h3c18baf8),
	.w6(32'hbb24e9d1),
	.w7(32'h3cae0327),
	.w8(32'h3c949455),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eb916),
	.w1(32'h3b5bd2ca),
	.w2(32'hbb61f87d),
	.w3(32'h3c472324),
	.w4(32'hbb1ad545),
	.w5(32'h3b658dc4),
	.w6(32'h3c5a016c),
	.w7(32'hbb3709cf),
	.w8(32'h3b3669ec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ac54b),
	.w1(32'hb9258272),
	.w2(32'h3ba1a147),
	.w3(32'h3b327a08),
	.w4(32'hbbc20687),
	.w5(32'h3ce1d4ef),
	.w6(32'h3bcfd3a4),
	.w7(32'h3a501cde),
	.w8(32'h3b3ab380),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014721),
	.w1(32'h3aacd2cb),
	.w2(32'h3b923392),
	.w3(32'hbb95f411),
	.w4(32'h3b535eb7),
	.w5(32'h3bfd3f30),
	.w6(32'h3b6f135e),
	.w7(32'h3b1f3a45),
	.w8(32'h3b852bde),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f13bd),
	.w1(32'h3a57e85c),
	.w2(32'h3bf15876),
	.w3(32'h3a355223),
	.w4(32'hbba2bb05),
	.w5(32'hb71ea742),
	.w6(32'h3b0f134b),
	.w7(32'hbb83db26),
	.w8(32'hbb8fa0d6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb39ab),
	.w1(32'hbbd17d2f),
	.w2(32'hbc299553),
	.w3(32'hbac26286),
	.w4(32'hbb691674),
	.w5(32'hbbb3c172),
	.w6(32'hbb5db097),
	.w7(32'hbbec01f3),
	.w8(32'hbc19e055),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50e1d),
	.w1(32'hbbef12c8),
	.w2(32'hbbca1cca),
	.w3(32'hba2484a3),
	.w4(32'hbbffe430),
	.w5(32'h3c6f8db7),
	.w6(32'hbb8217cf),
	.w7(32'hbbbab592),
	.w8(32'hbb2a32be),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6c866),
	.w1(32'h3b9760c8),
	.w2(32'h3c710f7d),
	.w3(32'hbb582edf),
	.w4(32'hbbe945c6),
	.w5(32'h3c61cd42),
	.w6(32'hba349ccf),
	.w7(32'h3aaff42f),
	.w8(32'h3b479cc7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9467fd),
	.w1(32'hba3ee3a5),
	.w2(32'hbaff63ca),
	.w3(32'h3b7b03c2),
	.w4(32'hbb7a62e9),
	.w5(32'hbbb822d6),
	.w6(32'h3ba4f8ba),
	.w7(32'hbb52deb1),
	.w8(32'h3a11f28b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03b48a),
	.w1(32'h3b41a1bc),
	.w2(32'h3c1d0404),
	.w3(32'hba9fdcdd),
	.w4(32'hbc14728d),
	.w5(32'h3ab0b177),
	.w6(32'hb9ceba92),
	.w7(32'h3ad7ccb9),
	.w8(32'h3baf46a7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87e70),
	.w1(32'hbbc229fa),
	.w2(32'hbab51e40),
	.w3(32'h3b7f4ac7),
	.w4(32'hba7cdef6),
	.w5(32'hbc107a20),
	.w6(32'h3bdb69f8),
	.w7(32'h3b38a751),
	.w8(32'hbb811fef),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c92e1),
	.w1(32'hbb5ca10c),
	.w2(32'hbc0a19b3),
	.w3(32'hbb8c9479),
	.w4(32'h3a091d0a),
	.w5(32'hbb34d117),
	.w6(32'hbb80fef3),
	.w7(32'h38b5010c),
	.w8(32'hbbfbb127),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed6495),
	.w1(32'hbae334d3),
	.w2(32'hbba8b167),
	.w3(32'hba9b2b25),
	.w4(32'hbacbb41e),
	.w5(32'hbc15dec6),
	.w6(32'hbbd8a11c),
	.w7(32'h3a5e6d33),
	.w8(32'hb9923970),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17caed),
	.w1(32'h3bb41d81),
	.w2(32'hbb167bb5),
	.w3(32'h3bf39374),
	.w4(32'hba588e10),
	.w5(32'hbc529ae8),
	.w6(32'hba37fad9),
	.w7(32'h3ba0034c),
	.w8(32'hbbdbf04b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a4eb9),
	.w1(32'h3a944750),
	.w2(32'hbb06c4bd),
	.w3(32'h3b3eccf4),
	.w4(32'hbaf4561d),
	.w5(32'h3b1b6661),
	.w6(32'h3b94e906),
	.w7(32'hba9cd64f),
	.w8(32'h3a00577e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb77f4b),
	.w1(32'hba72a788),
	.w2(32'hbb6d9328),
	.w3(32'h3bc593b4),
	.w4(32'h3a0af317),
	.w5(32'hbb9ece5a),
	.w6(32'h3b2ad188),
	.w7(32'hbb6e32e9),
	.w8(32'hbb73eff0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a94b),
	.w1(32'hbc02f1db),
	.w2(32'hbbb2b3a0),
	.w3(32'hbb2b0011),
	.w4(32'hbbbde148),
	.w5(32'hbb90b4b1),
	.w6(32'h38a36cb4),
	.w7(32'h39b5fce8),
	.w8(32'hbb3445cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6af9),
	.w1(32'hbb0a089b),
	.w2(32'h3b6eb6ea),
	.w3(32'hbba9adec),
	.w4(32'hbad02dc1),
	.w5(32'hbb5b0d26),
	.w6(32'hbc00e7da),
	.w7(32'hbae6e8f5),
	.w8(32'h3b4a9de8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18ac78),
	.w1(32'h39f3c592),
	.w2(32'hbb618f9d),
	.w3(32'hba6ddd05),
	.w4(32'hbb01bb6e),
	.w5(32'hbc2a37e3),
	.w6(32'h3b80ee84),
	.w7(32'hb9575f38),
	.w8(32'hbb82eacb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af9f1),
	.w1(32'h3c1575b1),
	.w2(32'h3c999156),
	.w3(32'hba9a277c),
	.w4(32'h3befeead),
	.w5(32'h3cc60598),
	.w6(32'hbc01621d),
	.w7(32'h39b243cf),
	.w8(32'h3c3ac599),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7c75),
	.w1(32'h3aa84e67),
	.w2(32'hba34e58d),
	.w3(32'h3b95c7b9),
	.w4(32'h3c4627e4),
	.w5(32'hbbd26deb),
	.w6(32'h3b984c1e),
	.w7(32'h3c2e9d09),
	.w8(32'h3b00a768),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0ed27),
	.w1(32'h3c09e25b),
	.w2(32'hbabd4f25),
	.w3(32'h394e6ebd),
	.w4(32'h3c9139b3),
	.w5(32'h398af1f7),
	.w6(32'hbb062ff1),
	.w7(32'h3c1ba292),
	.w8(32'h3b777689),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9f15e),
	.w1(32'h3c5d4925),
	.w2(32'h3ae8f9a7),
	.w3(32'hbbcd1f4e),
	.w4(32'h3baf4e2a),
	.w5(32'hbbc447dc),
	.w6(32'h3bbea00a),
	.w7(32'h3ba7e452),
	.w8(32'h3b140869),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7abe80),
	.w1(32'hbb942085),
	.w2(32'hbc1658bc),
	.w3(32'hbb503878),
	.w4(32'hbbe81804),
	.w5(32'hbc280a7e),
	.w6(32'h3c0b8b39),
	.w7(32'hbb6ac50d),
	.w8(32'hbbd36752),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00e11d),
	.w1(32'hbad91a9e),
	.w2(32'hbc055b62),
	.w3(32'hbb88365f),
	.w4(32'hbbbb0af2),
	.w5(32'hb8e322a4),
	.w6(32'hbbb5596c),
	.w7(32'hbc0ac0cc),
	.w8(32'hbc4b8bc5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3bb3),
	.w1(32'h3c175f92),
	.w2(32'h3c7e68e6),
	.w3(32'h3b45f53a),
	.w4(32'h3c0f0e80),
	.w5(32'h3c6e70f2),
	.w6(32'hba9a544c),
	.w7(32'h3b7f7c75),
	.w8(32'h3c855e86),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c751ca0),
	.w1(32'h3bdf99b6),
	.w2(32'hbc1c6579),
	.w3(32'h3c89d343),
	.w4(32'h3b9c58a0),
	.w5(32'hbc1cf26b),
	.w6(32'h3c10bb67),
	.w7(32'h3b206a22),
	.w8(32'hbc2d625b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa0185),
	.w1(32'hbc15e254),
	.w2(32'h3b68c34f),
	.w3(32'h3b9bf56a),
	.w4(32'hbbd58d7f),
	.w5(32'h3aa2ae85),
	.w6(32'hb937a3e1),
	.w7(32'hbb52dee3),
	.w8(32'h3ab721fe),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1f1d),
	.w1(32'hbc435a7f),
	.w2(32'h3b10b1ac),
	.w3(32'h3c432e4b),
	.w4(32'hbb848747),
	.w5(32'hb951df06),
	.w6(32'h3b50c355),
	.w7(32'hbbb13b0b),
	.w8(32'h3bfe4a7e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb7d59),
	.w1(32'hbb812144),
	.w2(32'hba95140a),
	.w3(32'h3b741405),
	.w4(32'hbbb08310),
	.w5(32'h3c154d16),
	.w6(32'hb9bc258b),
	.w7(32'hbb9ddde1),
	.w8(32'hbb6abd64),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e918),
	.w1(32'h3ac24272),
	.w2(32'h3c324eed),
	.w3(32'h3b9d0bee),
	.w4(32'h3bec05cf),
	.w5(32'h3cce1cb3),
	.w6(32'h3af8225a),
	.w7(32'h3b94d145),
	.w8(32'h3c036b6b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21458),
	.w1(32'hbb425a4b),
	.w2(32'hbb905ba6),
	.w3(32'hbbba75c9),
	.w4(32'hb99b9701),
	.w5(32'hbc213c6e),
	.w6(32'hbbb20e47),
	.w7(32'hbb5474f4),
	.w8(32'hbbcb30af),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39615586),
	.w1(32'hbae1697a),
	.w2(32'h3b8fa858),
	.w3(32'h3b8aee6c),
	.w4(32'hbb84c657),
	.w5(32'h3cb1483f),
	.w6(32'h3a7a741e),
	.w7(32'hb977a9c4),
	.w8(32'h39be81b3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796086),
	.w1(32'hbac3759f),
	.w2(32'h3ab2f2f4),
	.w3(32'hbc1af78f),
	.w4(32'h3b981179),
	.w5(32'h3b23de53),
	.w6(32'hbbd20987),
	.w7(32'h3b4d02df),
	.w8(32'h3b92f6ab),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba174a41),
	.w1(32'h3c5228cf),
	.w2(32'h3c825d69),
	.w3(32'hbb94f798),
	.w4(32'h3d049a4d),
	.w5(32'h3cbba731),
	.w6(32'h39987d39),
	.w7(32'h3c44da15),
	.w8(32'hbb0014c5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3428a),
	.w1(32'hbbb20073),
	.w2(32'hbb39e304),
	.w3(32'h3ad12158),
	.w4(32'hbbb32a47),
	.w5(32'hbb857f0a),
	.w6(32'hbc1951a3),
	.w7(32'hbb876561),
	.w8(32'hbb2a95a8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80032b),
	.w1(32'h3b18b97d),
	.w2(32'hbb0ee86f),
	.w3(32'hb94caf39),
	.w4(32'hbbeb05e4),
	.w5(32'hbc436f2e),
	.w6(32'hb86e1041),
	.w7(32'hbad8665b),
	.w8(32'hbb78b451),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d27a),
	.w1(32'h3aa8282e),
	.w2(32'h3b231fe3),
	.w3(32'hbb1fca36),
	.w4(32'hba8a8c41),
	.w5(32'hbc182828),
	.w6(32'hbba153df),
	.w7(32'h3a9ee8f7),
	.w8(32'hbbcb20f4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1133a5),
	.w1(32'hbb897ffd),
	.w2(32'h3ab4a74f),
	.w3(32'h3b1452cb),
	.w4(32'hbb63665c),
	.w5(32'h3bacf6a2),
	.w6(32'hbb9c54cc),
	.w7(32'hbb0b0408),
	.w8(32'hb9740787),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dadd3),
	.w1(32'hbbbd20c5),
	.w2(32'hbb1bd398),
	.w3(32'hbc046263),
	.w4(32'hbb3ce686),
	.w5(32'hbb1262b1),
	.w6(32'hbbbd7e72),
	.w7(32'hb8c01d3c),
	.w8(32'hbbe03aa2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f863),
	.w1(32'h3bbaeef4),
	.w2(32'hbc0b3122),
	.w3(32'h3a258c89),
	.w4(32'h3bead298),
	.w5(32'hbb4bfdb4),
	.w6(32'hbb31976b),
	.w7(32'hbafa1c36),
	.w8(32'hba508ee8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef17dd),
	.w1(32'h3c13e1a1),
	.w2(32'h3bbeeb9c),
	.w3(32'hba67fec9),
	.w4(32'h3b52ca42),
	.w5(32'hbc5948df),
	.w6(32'h38c32c70),
	.w7(32'hbb19e8c7),
	.w8(32'hbb1e9338),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace11ed),
	.w1(32'h3b26da6e),
	.w2(32'h3c3f5467),
	.w3(32'hbb56d2af),
	.w4(32'hbb3d6eba),
	.w5(32'h3c8d4961),
	.w6(32'hbbf291bd),
	.w7(32'hbbf8a783),
	.w8(32'h3c3f124f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfda32f),
	.w1(32'h3bd03c0b),
	.w2(32'h3bbc79b2),
	.w3(32'h3c928c5c),
	.w4(32'h3c46f882),
	.w5(32'h3c90abb6),
	.w6(32'h3c3dbb1c),
	.w7(32'h3b3ad43e),
	.w8(32'h3c6c1a67),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc071ba),
	.w1(32'hba3529e8),
	.w2(32'hbb9cf5bc),
	.w3(32'hbbecaaad),
	.w4(32'h3b08e724),
	.w5(32'hbbac434f),
	.w6(32'hbb722d1b),
	.w7(32'h3bb5c15b),
	.w8(32'hbb8c9536),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0db350),
	.w1(32'h3c7b6e2a),
	.w2(32'h3c166cbc),
	.w3(32'hb8508a1d),
	.w4(32'h3c929096),
	.w5(32'h3c14d6e2),
	.w6(32'hbb146446),
	.w7(32'h3c62574d),
	.w8(32'h3c0d11ed),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d87fd),
	.w1(32'h3aaf5e6f),
	.w2(32'hbb8f578b),
	.w3(32'hbbfaa700),
	.w4(32'h3a5016ae),
	.w5(32'h3b5952d1),
	.w6(32'h3ae1ec99),
	.w7(32'hbb879122),
	.w8(32'hbb282901),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf75517),
	.w1(32'hbb32cbc2),
	.w2(32'hbbcb1c68),
	.w3(32'hbbf5f425),
	.w4(32'hbbee99e3),
	.w5(32'hbcadbcc1),
	.w6(32'hbad6bd0c),
	.w7(32'hbb22ccf2),
	.w8(32'hbbbd7425),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad18c34),
	.w1(32'hbaa98acf),
	.w2(32'hbb6a9f82),
	.w3(32'hbb5f7126),
	.w4(32'h3c43aa20),
	.w5(32'hbc2b41ef),
	.w6(32'hbb9b20fd),
	.w7(32'hbbab6974),
	.w8(32'hbb72314e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91cefb),
	.w1(32'hbad2a03f),
	.w2(32'hbbf3f239),
	.w3(32'hbaa449d2),
	.w4(32'h3afdf0c9),
	.w5(32'h3c284c45),
	.w6(32'hbbcbf3ca),
	.w7(32'h3b811794),
	.w8(32'hbb367a2c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5aba68),
	.w1(32'hbc67e182),
	.w2(32'h3c2b256f),
	.w3(32'hbbe5fd9c),
	.w4(32'hbc124e1b),
	.w5(32'h3cdd264c),
	.w6(32'hb6a66a75),
	.w7(32'hbc323250),
	.w8(32'h3ae6e56b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe92258),
	.w1(32'hbb8911b2),
	.w2(32'hba61683b),
	.w3(32'hbc24c81b),
	.w4(32'hbb303907),
	.w5(32'h3b3ce3a7),
	.w6(32'hbc4bec27),
	.w7(32'hb8ccf1c3),
	.w8(32'hba4ca938),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222359),
	.w1(32'h3ace83eb),
	.w2(32'h3b8aa86c),
	.w3(32'hbc0c2289),
	.w4(32'h3acca9a6),
	.w5(32'hbb5e0971),
	.w6(32'hbbcaed65),
	.w7(32'h3ae5cd3b),
	.w8(32'hbaeb7a5b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd7fe),
	.w1(32'h3b61eade),
	.w2(32'hbc34c5ab),
	.w3(32'h3c26be37),
	.w4(32'h3bd4475c),
	.w5(32'hbb841494),
	.w6(32'h3b41b19f),
	.w7(32'h3bd97d58),
	.w8(32'hbab61430),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce5b5c),
	.w1(32'hbaf5afbc),
	.w2(32'hbbd66c8d),
	.w3(32'h3c118294),
	.w4(32'h3b29068c),
	.w5(32'hbbbefb55),
	.w6(32'h3ab1deda),
	.w7(32'hbb0ba1fe),
	.w8(32'h3b394816),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817555),
	.w1(32'hbba77f3e),
	.w2(32'h3a6f39a9),
	.w3(32'hb9879980),
	.w4(32'hbac4ff77),
	.w5(32'hbba2b622),
	.w6(32'h3b8c95b9),
	.w7(32'hbba27c15),
	.w8(32'hbb83c844),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb172d1),
	.w1(32'hbb0de62c),
	.w2(32'hbb26a63a),
	.w3(32'hbc222146),
	.w4(32'hba80cfdb),
	.w5(32'h3b6c8f22),
	.w6(32'hbafb8218),
	.w7(32'h3a70fc8a),
	.w8(32'h3b20b436),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ecb8),
	.w1(32'h3ac98f1b),
	.w2(32'hba9e1aff),
	.w3(32'h3a221d57),
	.w4(32'hbba41d34),
	.w5(32'hb8a5bfa1),
	.w6(32'hbabfb322),
	.w7(32'h3b0691ac),
	.w8(32'h3b3fea01),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058874),
	.w1(32'hbb58a698),
	.w2(32'hbb394901),
	.w3(32'hbbb0155d),
	.w4(32'hbaa5a969),
	.w5(32'h3a68d2e6),
	.w6(32'hbacabf64),
	.w7(32'hbb854ebc),
	.w8(32'hbad44514),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96998e),
	.w1(32'hbc09b18f),
	.w2(32'hbb81a94f),
	.w3(32'hbb048f1a),
	.w4(32'hba141be5),
	.w5(32'h3c7a98ea),
	.w6(32'h3b5323a4),
	.w7(32'h3b0d520c),
	.w8(32'h3b64ed20),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd5d6),
	.w1(32'h3b1e9569),
	.w2(32'hba70acfd),
	.w3(32'h3c28928c),
	.w4(32'h3981b13f),
	.w5(32'hbb9434e0),
	.w6(32'hbb6aaae6),
	.w7(32'hbb338c7a),
	.w8(32'hbc066f25),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1143f),
	.w1(32'h3aba02d5),
	.w2(32'h3ba5aaec),
	.w3(32'hba9e1c67),
	.w4(32'hba527441),
	.w5(32'hbb264d83),
	.w6(32'hbadd0796),
	.w7(32'hbb968e3b),
	.w8(32'h3862cc2e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab102f4),
	.w1(32'hbc0c6b40),
	.w2(32'hbc16c44c),
	.w3(32'hbba407ea),
	.w4(32'h3af659b2),
	.w5(32'h3b2604af),
	.w6(32'h3a8714c2),
	.w7(32'hbb5e6e87),
	.w8(32'hbb0b19a1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb059d20),
	.w1(32'h3a455edc),
	.w2(32'h3bd44749),
	.w3(32'h3b8e2624),
	.w4(32'h3bc7e460),
	.w5(32'h3c2fabc8),
	.w6(32'hbac78922),
	.w7(32'h3b69b3ed),
	.w8(32'h3b315235),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8aa81),
	.w1(32'hbb791f18),
	.w2(32'hbbaebac6),
	.w3(32'h3bb3aa93),
	.w4(32'hbb8000ec),
	.w5(32'hbb7ada05),
	.w6(32'hbb4011e2),
	.w7(32'hbc09635c),
	.w8(32'hb968f924),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee9b32),
	.w1(32'h3b26915a),
	.w2(32'hbad20c08),
	.w3(32'hbbcd1e66),
	.w4(32'hbb9b7277),
	.w5(32'hbbd46502),
	.w6(32'hbb51c62d),
	.w7(32'hbb804695),
	.w8(32'hbb9e6c54),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbddbe4),
	.w1(32'h3b42264d),
	.w2(32'hbb5ec8fa),
	.w3(32'hbbe419a7),
	.w4(32'h3b9e295a),
	.w5(32'h3bc61a9a),
	.w6(32'h3b1bd7f6),
	.w7(32'h3b8028f5),
	.w8(32'h3b01f05b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60b13a),
	.w1(32'h3b430a87),
	.w2(32'hba988261),
	.w3(32'h3c241c6b),
	.w4(32'hbbc688db),
	.w5(32'h39a23ab3),
	.w6(32'hbaa83643),
	.w7(32'hbb5991b3),
	.w8(32'h3be07721),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172387),
	.w1(32'h3c2c93a7),
	.w2(32'h3b9ecebf),
	.w3(32'hb9a79990),
	.w4(32'h3b9b2b81),
	.w5(32'hbb80e14c),
	.w6(32'hbac8a1ab),
	.w7(32'h3bd79447),
	.w8(32'h3b2355b4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff562),
	.w1(32'hba1d6de3),
	.w2(32'hbb0fded8),
	.w3(32'h3bfc30e9),
	.w4(32'hbaed7bfd),
	.w5(32'hbb10172e),
	.w6(32'h3b436121),
	.w7(32'hbb64ca2f),
	.w8(32'hbb5eb6aa),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadea10),
	.w1(32'hbaa69a41),
	.w2(32'hbb76a75f),
	.w3(32'hb8b4b7ed),
	.w4(32'hbba9f7dd),
	.w5(32'hbabee061),
	.w6(32'hbacf84d3),
	.w7(32'h3c394421),
	.w8(32'h3c1199e6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafd317),
	.w1(32'h3a047a91),
	.w2(32'hb9f0750b),
	.w3(32'h3c4e8094),
	.w4(32'hbb60ac3b),
	.w5(32'h3b06270a),
	.w6(32'h3aa2118a),
	.w7(32'h3a059438),
	.w8(32'h38c079eb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905ea1f),
	.w1(32'hbba615d9),
	.w2(32'hbbd23b9a),
	.w3(32'hbb3be7bf),
	.w4(32'hbb84db62),
	.w5(32'hbba47fad),
	.w6(32'h3b1f3f37),
	.w7(32'hbb4a3e75),
	.w8(32'h394aef65),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ba6bb),
	.w1(32'hbbcbcb06),
	.w2(32'h3b28dcb3),
	.w3(32'hba128b8b),
	.w4(32'h3ab5752f),
	.w5(32'h3bf4266e),
	.w6(32'hb7cbff6f),
	.w7(32'h3bfa9e5b),
	.w8(32'h3bc0348a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced4a5),
	.w1(32'h3b0e1011),
	.w2(32'hbb3d08fe),
	.w3(32'h3b8a928b),
	.w4(32'hbad365ed),
	.w5(32'hbc0c75eb),
	.w6(32'hbb0cde69),
	.w7(32'hba4bdcd3),
	.w8(32'h39c2b43d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4639f),
	.w1(32'hbb8088d0),
	.w2(32'hba7df04a),
	.w3(32'hbbd4fbda),
	.w4(32'hbba7dd49),
	.w5(32'hbb8a590c),
	.w6(32'hbbb88eae),
	.w7(32'hbb8ad177),
	.w8(32'h3a7a22e8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1df7),
	.w1(32'h3a2e875d),
	.w2(32'hb8c58c4b),
	.w3(32'hbbabb490),
	.w4(32'hbbb2519e),
	.w5(32'hbb993f73),
	.w6(32'h3a6b66a9),
	.w7(32'hbb577121),
	.w8(32'h3ac09bd2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee99c),
	.w1(32'hba1644b3),
	.w2(32'hbaf9f387),
	.w3(32'hbb90ec36),
	.w4(32'hbaaceff0),
	.w5(32'hbbaae5d3),
	.w6(32'hb95029f7),
	.w7(32'hbb4da7ce),
	.w8(32'hbac1c55b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da14e),
	.w1(32'hbba8c49d),
	.w2(32'hbb8462c2),
	.w3(32'hbacfb393),
	.w4(32'hbbe33ea2),
	.w5(32'hbb53a0dc),
	.w6(32'hbb87b740),
	.w7(32'hbc1a2ff6),
	.w8(32'hbb2f522d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020675),
	.w1(32'hbb5c12a0),
	.w2(32'hbab8adee),
	.w3(32'hbb6049d8),
	.w4(32'h3b4a2103),
	.w5(32'h3a3ebc7c),
	.w6(32'hbb7fc51a),
	.w7(32'h3b8f3352),
	.w8(32'hbac7c402),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37279),
	.w1(32'hbaf12c0b),
	.w2(32'hbb84f220),
	.w3(32'h3b1941cd),
	.w4(32'hbb7d0d84),
	.w5(32'hb900587d),
	.w6(32'h397c1d02),
	.w7(32'h3bdcde71),
	.w8(32'h3b8bd3cb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0289c7),
	.w1(32'h3b7b4804),
	.w2(32'h3baf2c45),
	.w3(32'h3a849e54),
	.w4(32'h3b3e7070),
	.w5(32'hbb1b3d90),
	.w6(32'hbb98bc02),
	.w7(32'h3a2b99ad),
	.w8(32'hbb165a8d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c93b3),
	.w1(32'hb9e6b02e),
	.w2(32'h3abc32a2),
	.w3(32'hbb0fcbad),
	.w4(32'hbbbd7ea1),
	.w5(32'hbabab852),
	.w6(32'hb97189aa),
	.w7(32'hbb3093a0),
	.w8(32'h39e03860),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274ca9),
	.w1(32'h3a9222b0),
	.w2(32'h3c0485bc),
	.w3(32'hbb1d7737),
	.w4(32'h3b1e275d),
	.w5(32'hbbac866c),
	.w6(32'hbb87edc2),
	.w7(32'hbb8fd73d),
	.w8(32'hba0de938),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7fdb6),
	.w1(32'hbbc22e84),
	.w2(32'hbafcc9d2),
	.w3(32'hbbc32682),
	.w4(32'h3a12f280),
	.w5(32'h37d13d4e),
	.w6(32'h3c43d0cf),
	.w7(32'hbae67afa),
	.w8(32'hba1f02f8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a053c04),
	.w1(32'hbb56af1e),
	.w2(32'h3b3df853),
	.w3(32'hbbd827f7),
	.w4(32'hbad2abd8),
	.w5(32'hba738ffd),
	.w6(32'h389f0240),
	.w7(32'h3a181074),
	.w8(32'h3ac6f9d6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376b3c),
	.w1(32'h3be994cb),
	.w2(32'h39cc50c7),
	.w3(32'hbb7d26ed),
	.w4(32'h3a3b8720),
	.w5(32'hba10926c),
	.w6(32'hbb53cda8),
	.w7(32'hba8abf59),
	.w8(32'h3b574f40),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c41079),
	.w1(32'hbaad6fc2),
	.w2(32'hbb413f52),
	.w3(32'h39a4253b),
	.w4(32'h3a20b04e),
	.w5(32'hbac93465),
	.w6(32'hbb5997a9),
	.w7(32'hbb5e3ded),
	.w8(32'hbc075d7e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f0b1),
	.w1(32'hbb6f6c9b),
	.w2(32'h3a1d8b5e),
	.w3(32'hbb0d6a9b),
	.w4(32'hba947a77),
	.w5(32'h3b6c505c),
	.w6(32'hbbf5fa02),
	.w7(32'hbbdf2a9b),
	.w8(32'h3b26fc22),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5db6),
	.w1(32'hbb715548),
	.w2(32'hbb3a6127),
	.w3(32'hbba596e3),
	.w4(32'hbbae0af7),
	.w5(32'hbc154e6b),
	.w6(32'h3971fee9),
	.w7(32'hb9cfe889),
	.w8(32'hba9966fb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08493e),
	.w1(32'hbb2eef93),
	.w2(32'hbb1449c4),
	.w3(32'hba8c52f8),
	.w4(32'hbbb89c9d),
	.w5(32'hbb333bc8),
	.w6(32'hbae40d1f),
	.w7(32'h3b82eb8d),
	.w8(32'h3c1cff74),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62f361),
	.w1(32'hbb88a76b),
	.w2(32'hbb9af809),
	.w3(32'hba6f4ee4),
	.w4(32'hbadbc2b5),
	.w5(32'hbc0ab26a),
	.w6(32'h3bc58aea),
	.w7(32'h3a9709d2),
	.w8(32'h3a4b35b4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8cb2c),
	.w1(32'hbb66fdee),
	.w2(32'hbbfdb60e),
	.w3(32'hbb4dac15),
	.w4(32'hbb483b89),
	.w5(32'h3c156315),
	.w6(32'h3b6b36e6),
	.w7(32'h3bfd2cdb),
	.w8(32'h3b30b6d7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929796),
	.w1(32'hbb15cd39),
	.w2(32'hbb6b715a),
	.w3(32'h3c5d11d0),
	.w4(32'hbacb84bf),
	.w5(32'hb7e06701),
	.w6(32'hbbd7434a),
	.w7(32'h3aa19944),
	.w8(32'h3aabd791),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff0bb5),
	.w1(32'hbb53221f),
	.w2(32'hbb9d3244),
	.w3(32'h3b532e58),
	.w4(32'h3abf548b),
	.w5(32'h3b95b32e),
	.w6(32'hbb3b9889),
	.w7(32'hba87e00e),
	.w8(32'hb70b5d08),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67eae),
	.w1(32'hb96378e9),
	.w2(32'h39badf58),
	.w3(32'h3b9a9fc5),
	.w4(32'hbb6fc83c),
	.w5(32'hbb390aa0),
	.w6(32'h3acaad7d),
	.w7(32'hbbbadcc2),
	.w8(32'h3a4f6fc0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb719c9d),
	.w1(32'hbb088df9),
	.w2(32'hba2fc6df),
	.w3(32'hbc03167a),
	.w4(32'h3a6eed6b),
	.w5(32'h3c1e6589),
	.w6(32'hbb980a0b),
	.w7(32'h3c000229),
	.w8(32'h3b80c42e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3d914),
	.w1(32'hbbc2859e),
	.w2(32'hbc0db5cd),
	.w3(32'h3c67296c),
	.w4(32'hbba1f403),
	.w5(32'hbc1036f2),
	.w6(32'hbb4682d6),
	.w7(32'h3b4ff7de),
	.w8(32'h3b4c6e28),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94821a),
	.w1(32'h3ba473da),
	.w2(32'h3c192a43),
	.w3(32'h3aa29665),
	.w4(32'h3c18d232),
	.w5(32'h3b71893c),
	.w6(32'h3b20e224),
	.w7(32'h3b358e1c),
	.w8(32'hbac8582a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91352),
	.w1(32'hba4698d4),
	.w2(32'hbbb1473e),
	.w3(32'hb9cda2c7),
	.w4(32'hbb04e3df),
	.w5(32'hbbd18a5e),
	.w6(32'h3b472bfe),
	.w7(32'hbb32ae4c),
	.w8(32'hbb9b4ef3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab68d01),
	.w1(32'h3b91fa68),
	.w2(32'h3bb3a406),
	.w3(32'hba0d568f),
	.w4(32'hbade6547),
	.w5(32'hbbde88e3),
	.w6(32'hbad997ab),
	.w7(32'hba8e5bab),
	.w8(32'hb998985a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193a9c),
	.w1(32'h3a8c2553),
	.w2(32'hbb522a14),
	.w3(32'hbb43a712),
	.w4(32'hbb03f40a),
	.w5(32'h3b5f62e0),
	.w6(32'hba938034),
	.w7(32'h3b449fb8),
	.w8(32'h3c2af6f8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbfcb),
	.w1(32'h3b212a2e),
	.w2(32'hbb5352d4),
	.w3(32'h3bb707d6),
	.w4(32'hbb7fa493),
	.w5(32'hbb02c5d1),
	.w6(32'hbb0f0a7d),
	.w7(32'hb9c03e4b),
	.w8(32'hbb972116),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d99b),
	.w1(32'hbaa23558),
	.w2(32'hbad3d8d2),
	.w3(32'hbb4b4dad),
	.w4(32'h3aa8d48d),
	.w5(32'h3a1c2a34),
	.w6(32'hbb5d9bbb),
	.w7(32'h3b4cc804),
	.w8(32'h3b95ee9d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39217158),
	.w1(32'hbad607b3),
	.w2(32'hbb05cfa1),
	.w3(32'h39bf9e03),
	.w4(32'hbb4730b1),
	.w5(32'hba58210b),
	.w6(32'h3a177c73),
	.w7(32'h3ad1d175),
	.w8(32'h3a65bc52),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2d12),
	.w1(32'hbbf19bd8),
	.w2(32'hbbfa1314),
	.w3(32'hbb8059ca),
	.w4(32'hbb1b0655),
	.w5(32'hbb553f0f),
	.w6(32'hb8919669),
	.w7(32'h3ad526e6),
	.w8(32'hba274a85),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eac19),
	.w1(32'h3989cc80),
	.w2(32'h3b20a43e),
	.w3(32'h3a536c63),
	.w4(32'hbbdabd64),
	.w5(32'hbb9d2fdf),
	.w6(32'hbb214b3a),
	.w7(32'hbb93cb35),
	.w8(32'hb9a62777),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb29c),
	.w1(32'hbc0f1119),
	.w2(32'hbb7dcda5),
	.w3(32'hbc1629f0),
	.w4(32'hbbb316cc),
	.w5(32'hbb2a17f1),
	.w6(32'h3abd0904),
	.w7(32'h3c0ef6a0),
	.w8(32'h3bd6ed8e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb475edf),
	.w1(32'hb9913290),
	.w2(32'hbb2c9c3f),
	.w3(32'hbb386701),
	.w4(32'hbae8c318),
	.w5(32'h3a9dc7c5),
	.w6(32'h3b381624),
	.w7(32'hbb7f5a1b),
	.w8(32'h3b6c27cb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1ef2),
	.w1(32'h3beb3fb9),
	.w2(32'h3b7c84f0),
	.w3(32'h3b3d6f59),
	.w4(32'hb9beff29),
	.w5(32'h3c4c34d4),
	.w6(32'h3b755eae),
	.w7(32'h3b736744),
	.w8(32'h3b87211e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587675),
	.w1(32'hbad0312b),
	.w2(32'h3bc73e6c),
	.w3(32'h3c2ecb77),
	.w4(32'hbb8ca7e9),
	.w5(32'hbb0116c3),
	.w6(32'hbc13b2ee),
	.w7(32'hbadb73b5),
	.w8(32'h3ba5409c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d9e0),
	.w1(32'h3aef89e3),
	.w2(32'h3b1db80e),
	.w3(32'hbb8fe180),
	.w4(32'h3789967f),
	.w5(32'hbc3b6950),
	.w6(32'h3bae3894),
	.w7(32'hba9ce6b0),
	.w8(32'hbb82a82f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaa0a3),
	.w1(32'hbc5959ca),
	.w2(32'hbc06a64d),
	.w3(32'hbb07c056),
	.w4(32'hbab30bb5),
	.w5(32'h3bec31d7),
	.w6(32'hb9c609b6),
	.w7(32'h3b822913),
	.w8(32'h3b3492ee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6078aa),
	.w1(32'hbaed801d),
	.w2(32'hbb821fb5),
	.w3(32'h3bb59de2),
	.w4(32'hba99ec09),
	.w5(32'h3c287d89),
	.w6(32'hbb718975),
	.w7(32'hbaa03074),
	.w8(32'h3b69ebe6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308fb2),
	.w1(32'h3b0c8a25),
	.w2(32'h3a1d8329),
	.w3(32'h3c11b123),
	.w4(32'h3a2343e7),
	.w5(32'h3b697b22),
	.w6(32'hbbb61caf),
	.w7(32'hbb9708c9),
	.w8(32'hbb120e1b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b478a6f),
	.w1(32'hbbe2c1df),
	.w2(32'hbbc10cce),
	.w3(32'hbaee475f),
	.w4(32'hbb028beb),
	.w5(32'h3b056758),
	.w6(32'hbb5e7f49),
	.w7(32'hb9114382),
	.w8(32'hba9c8be3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ef33b),
	.w1(32'hba192691),
	.w2(32'hbb83e347),
	.w3(32'hbb136acf),
	.w4(32'h3a8016f3),
	.w5(32'hbb962e64),
	.w6(32'h39ec87fa),
	.w7(32'hb9ced945),
	.w8(32'hbb5295b6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab7203),
	.w1(32'hbab528e9),
	.w2(32'hbb01efdc),
	.w3(32'h38f1f685),
	.w4(32'hbbafc354),
	.w5(32'hb9dce260),
	.w6(32'hbac0a59f),
	.w7(32'h3b1cc1b4),
	.w8(32'h3bbe1e8c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97efc9),
	.w1(32'hbbe685a3),
	.w2(32'hbc0e30a1),
	.w3(32'h3b3ca604),
	.w4(32'hbc025369),
	.w5(32'hbb89ac91),
	.w6(32'hbb01323a),
	.w7(32'hbb9c49f0),
	.w8(32'hbaf10696),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40e199),
	.w1(32'h3adfdef9),
	.w2(32'hbbac7859),
	.w3(32'hbbb8007a),
	.w4(32'h37a91a21),
	.w5(32'h3c23a464),
	.w6(32'hbba71d5a),
	.w7(32'h3b8d897c),
	.w8(32'h39e004c7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec12f4),
	.w1(32'hbacdf118),
	.w2(32'hba974ac7),
	.w3(32'h3c545ab9),
	.w4(32'hbb2deccc),
	.w5(32'hbbf2793c),
	.w6(32'hbb92976c),
	.w7(32'hba08b47c),
	.w8(32'hb9e21784),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e87af7),
	.w1(32'h3b66926d),
	.w2(32'h3af9b701),
	.w3(32'h38afeac9),
	.w4(32'hbaf247e3),
	.w5(32'hbc2fcedb),
	.w6(32'hb95f1b32),
	.w7(32'hba846b5f),
	.w8(32'hbb534cb3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fb875),
	.w1(32'h3c00b7a7),
	.w2(32'h3c832f2a),
	.w3(32'hbc05ce58),
	.w4(32'h3c11b97b),
	.w5(32'h3bd0317d),
	.w6(32'hbb8fe1e2),
	.w7(32'hbacae027),
	.w8(32'hbb8bc3c0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb125d2),
	.w1(32'h3c40de6d),
	.w2(32'h3bfc77a5),
	.w3(32'hbb6c047e),
	.w4(32'h3b3a62ec),
	.w5(32'hbc258668),
	.w6(32'h3b7c6891),
	.w7(32'hbb9b7a9a),
	.w8(32'hbb4e8194),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85a3a87),
	.w1(32'hbaa86f76),
	.w2(32'hbaca9230),
	.w3(32'hbc359a10),
	.w4(32'h3b1003de),
	.w5(32'h3b1882af),
	.w6(32'hba344da0),
	.w7(32'hb94ea0a4),
	.w8(32'h39e8052b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b2d04),
	.w1(32'hba7e126f),
	.w2(32'hbb590af9),
	.w3(32'hb8dfd854),
	.w4(32'h3b8878d7),
	.w5(32'h3c3ca36a),
	.w6(32'hba9e00f7),
	.w7(32'h398c6cb6),
	.w8(32'hb880455f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58bf59),
	.w1(32'hbb282472),
	.w2(32'h3b35db87),
	.w3(32'h3c3166eb),
	.w4(32'h3c2e1a12),
	.w5(32'h3c6f86b3),
	.w6(32'hbb8d86c8),
	.w7(32'h3b078ce0),
	.w8(32'hb9ebe97f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b67f),
	.w1(32'hbb118619),
	.w2(32'hbb3fc361),
	.w3(32'h3c23bd87),
	.w4(32'h3a2ccbbb),
	.w5(32'h3a211082),
	.w6(32'hba0d187c),
	.w7(32'hbbc16533),
	.w8(32'hbb091b40),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79f5d8),
	.w1(32'h39bd399b),
	.w2(32'hbbe4f044),
	.w3(32'h3a8adec7),
	.w4(32'hbbb7141f),
	.w5(32'hba07463e),
	.w6(32'h3b392fb3),
	.w7(32'hbb140bc0),
	.w8(32'h3b07cadb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ecf0),
	.w1(32'h3a1d0801),
	.w2(32'h3ad62d18),
	.w3(32'h3c00a29d),
	.w4(32'hbba4db56),
	.w5(32'hbb4bdddb),
	.w6(32'hba654449),
	.w7(32'h3bbcf068),
	.w8(32'h3b5cafcb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a196f),
	.w1(32'hbbaa33ca),
	.w2(32'hbb595b8e),
	.w3(32'h3bd483f1),
	.w4(32'h3aa77857),
	.w5(32'hbbafe0cf),
	.w6(32'h3b3a7b04),
	.w7(32'hb7b5c767),
	.w8(32'hbbbc86ce),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482baf),
	.w1(32'hbb45076e),
	.w2(32'hbae50331),
	.w3(32'hbb4f1493),
	.w4(32'hb9e05687),
	.w5(32'hb9754913),
	.w6(32'hba478859),
	.w7(32'hbb01bf10),
	.w8(32'hbb1ec394),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45acfb),
	.w1(32'hba693fbf),
	.w2(32'hba0f76ef),
	.w3(32'hbaa642cd),
	.w4(32'hbb4b6ad0),
	.w5(32'hba7c9326),
	.w6(32'h39e48349),
	.w7(32'h3a9a06de),
	.w8(32'h3bc8dc76),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266689),
	.w1(32'hbba6220d),
	.w2(32'hbbaffbea),
	.w3(32'hbb4494bf),
	.w4(32'h38aa614d),
	.w5(32'h3acd19af),
	.w6(32'h3a259007),
	.w7(32'hbb8ccb15),
	.w8(32'hbb3a17c8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf46f08),
	.w1(32'hbbb4429b),
	.w2(32'hbb23c72e),
	.w3(32'hbb13f2bb),
	.w4(32'hbb4a5bb8),
	.w5(32'hbacfd497),
	.w6(32'hbbb95ee7),
	.w7(32'hbb87ebb5),
	.w8(32'h3b43bcd1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ed59f),
	.w1(32'h3a8929dc),
	.w2(32'hbb9c8ef1),
	.w3(32'hbb8f6bba),
	.w4(32'h3858338c),
	.w5(32'hbb76f977),
	.w6(32'h3ae9eb52),
	.w7(32'h3ada611c),
	.w8(32'hbba2c2b4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b4821),
	.w1(32'h3b2bb89f),
	.w2(32'hba635f4f),
	.w3(32'hba2cfcd0),
	.w4(32'hbb215177),
	.w5(32'hbbb4d114),
	.w6(32'hbb09758d),
	.w7(32'hbb7c96d0),
	.w8(32'hbb87e522),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866f78),
	.w1(32'h3ad09aa8),
	.w2(32'h3b8146de),
	.w3(32'hbc0df2a4),
	.w4(32'hbb529a8d),
	.w5(32'hbb556744),
	.w6(32'hb8c56470),
	.w7(32'h375048d8),
	.w8(32'hbaed82ae),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b546a6e),
	.w1(32'hbbaf9ae1),
	.w2(32'h3b12d83a),
	.w3(32'hbbf98b1d),
	.w4(32'h3ba91667),
	.w5(32'h3c84c7e7),
	.w6(32'h3aa7f70b),
	.w7(32'h3bc9b10b),
	.w8(32'hbbe80ef6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183819),
	.w1(32'hbb07a370),
	.w2(32'hbbb7e9d9),
	.w3(32'hbbd6e809),
	.w4(32'hbb4af8db),
	.w5(32'hbb9e80d2),
	.w6(32'h3b87d9ff),
	.w7(32'hbae7ae1a),
	.w8(32'hba814d80),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8b8b),
	.w1(32'h3aa9286f),
	.w2(32'hbb3c3507),
	.w3(32'hbbc88cbd),
	.w4(32'hbba1b5ce),
	.w5(32'h3abeb18e),
	.w6(32'hbbaaa39f),
	.w7(32'hb7d4b7c5),
	.w8(32'hbbac0266),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97de61),
	.w1(32'h3c161239),
	.w2(32'h3b98a447),
	.w3(32'hbbdae2d6),
	.w4(32'h3b6808b1),
	.w5(32'hbb904911),
	.w6(32'hb7263bc9),
	.w7(32'h3bc2cbde),
	.w8(32'h396ffff3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5d20f),
	.w1(32'h3b2d9b83),
	.w2(32'h3b049a58),
	.w3(32'hbb0e2208),
	.w4(32'h3ac4a3ab),
	.w5(32'h3b0db157),
	.w6(32'hba9da891),
	.w7(32'hbba989c4),
	.w8(32'h3ad40911),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75cd50),
	.w1(32'hb9f09da5),
	.w2(32'hba01f3a6),
	.w3(32'hba0458eb),
	.w4(32'h38d9791d),
	.w5(32'h3957880d),
	.w6(32'h3bcebb5a),
	.w7(32'h3998ff25),
	.w8(32'hbb1d53fe),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaac39),
	.w1(32'hb9fe91f0),
	.w2(32'h3ac9321e),
	.w3(32'hba8280dd),
	.w4(32'h3b012e14),
	.w5(32'hba8a7ce9),
	.w6(32'h3a776266),
	.w7(32'hbbbfc767),
	.w8(32'hbbb8b93b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29234),
	.w1(32'h3a23aed4),
	.w2(32'hbb245f5f),
	.w3(32'hbbc54583),
	.w4(32'hbb60bc35),
	.w5(32'hb9e2052b),
	.w6(32'hbab26211),
	.w7(32'hbc00b0c5),
	.w8(32'hbb9f665c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad151e1),
	.w1(32'h3b8b0b90),
	.w2(32'h3c02f1f3),
	.w3(32'h3b15db3d),
	.w4(32'hbbc598eb),
	.w5(32'hbbd27390),
	.w6(32'hbb72dc75),
	.w7(32'hb9d93937),
	.w8(32'h3a0a8d85),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74c69f),
	.w1(32'hba42fb40),
	.w2(32'hbb170b8d),
	.w3(32'hbbea0635),
	.w4(32'h394a186c),
	.w5(32'hbad071b2),
	.w6(32'h3b2aa595),
	.w7(32'h3ad94cd9),
	.w8(32'hba369212),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f43f1),
	.w1(32'hbb3cc663),
	.w2(32'hba1379c2),
	.w3(32'hbb6ff97d),
	.w4(32'hbc060c3a),
	.w5(32'hbba03930),
	.w6(32'h3b00c9ab),
	.w7(32'hbbe58644),
	.w8(32'h3a7d9b2b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2739df),
	.w1(32'hb93bddfb),
	.w2(32'h3b1f8a5a),
	.w3(32'hbb25ac77),
	.w4(32'hba184715),
	.w5(32'h3ac01fa7),
	.w6(32'h3b60d33f),
	.w7(32'hba5cdcff),
	.w8(32'hbaacabf7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1af6a1),
	.w1(32'hbaf1c112),
	.w2(32'hbb2e21e1),
	.w3(32'hbacd3637),
	.w4(32'h3b08ede0),
	.w5(32'hba890c5c),
	.w6(32'h3ad15abb),
	.w7(32'h3c071ed0),
	.w8(32'h3c279b58),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5d122),
	.w1(32'hb9ae8f5f),
	.w2(32'hbbd1508a),
	.w3(32'h3c261a7c),
	.w4(32'h3a62d830),
	.w5(32'h3c2b1d18),
	.w6(32'h3b1ee67a),
	.w7(32'h3b1b0e90),
	.w8(32'h3ab5ec47),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7acc14),
	.w1(32'hbb224cf8),
	.w2(32'h3a3d16d6),
	.w3(32'h3c077370),
	.w4(32'h3b61e901),
	.w5(32'h3c0bb5ad),
	.w6(32'hbb3f3f13),
	.w7(32'h3ae7e29a),
	.w8(32'h3b2bcc82),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fc407),
	.w1(32'hb8eacf4a),
	.w2(32'hbb6403c8),
	.w3(32'h3ba1d5c9),
	.w4(32'hbb85f8e9),
	.w5(32'hbbba0b0c),
	.w6(32'h3b7b29e9),
	.w7(32'hbb1562ea),
	.w8(32'hbb707b72),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee8395),
	.w1(32'hba1ece7f),
	.w2(32'hba0eba7b),
	.w3(32'h39ae4f6b),
	.w4(32'hba77d915),
	.w5(32'hbc02d461),
	.w6(32'h3901574a),
	.w7(32'hbb600e9d),
	.w8(32'hbb5f6da5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6247b),
	.w1(32'h3bdb3ed5),
	.w2(32'h3ad86fb2),
	.w3(32'hbbe576e7),
	.w4(32'h3b08f828),
	.w5(32'hbaa19b30),
	.w6(32'h3ac4a1eb),
	.w7(32'h3ae8b792),
	.w8(32'h3b298d88),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac94ac8),
	.w1(32'h3b473e69),
	.w2(32'hbb8bf8fc),
	.w3(32'h39c76907),
	.w4(32'hbc05c4d9),
	.w5(32'hbc814b22),
	.w6(32'h396744b3),
	.w7(32'h3b5d1a66),
	.w8(32'h3bb389ce),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f827),
	.w1(32'hbb3d3080),
	.w2(32'h3983352c),
	.w3(32'h3b387de1),
	.w4(32'hbb24922b),
	.w5(32'hbbcefb0b),
	.w6(32'h3bf04c37),
	.w7(32'hbb53455d),
	.w8(32'hbbaca06c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf956e2),
	.w1(32'h3b651902),
	.w2(32'hbb88c949),
	.w3(32'hbbf69ef0),
	.w4(32'h39acfd21),
	.w5(32'h3b1b50c3),
	.w6(32'hbb470f05),
	.w7(32'h3af60a68),
	.w8(32'h3abea1ff),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05b277),
	.w1(32'h3a9a399b),
	.w2(32'hb9873328),
	.w3(32'h3aa66313),
	.w4(32'h3ac5f0bc),
	.w5(32'hbc01b579),
	.w6(32'hbbab0bfa),
	.w7(32'hbb4d43c2),
	.w8(32'hbb5527ef),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233730),
	.w1(32'hbac6aa67),
	.w2(32'hb9c4f622),
	.w3(32'hbb23498e),
	.w4(32'hb98be795),
	.w5(32'hbb177b57),
	.w6(32'hb9b20a1f),
	.w7(32'hba796310),
	.w8(32'hba736374),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857eb99),
	.w1(32'hbbab438f),
	.w2(32'hbb96da3d),
	.w3(32'hbb5d4a87),
	.w4(32'h3b196a1a),
	.w5(32'h3abcdf95),
	.w6(32'hba776add),
	.w7(32'hba2b5403),
	.w8(32'hbb4350f0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48dcb0),
	.w1(32'hbb842331),
	.w2(32'hbbb0bee0),
	.w3(32'hba274d4e),
	.w4(32'hbbc1333a),
	.w5(32'h3b4850f6),
	.w6(32'h3a92ffb5),
	.w7(32'h3bb575c2),
	.w8(32'h3a550f47),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5b04),
	.w1(32'hbb3d4d99),
	.w2(32'hbaa8e901),
	.w3(32'h3c014a14),
	.w4(32'hbb310e00),
	.w5(32'h3a37bf93),
	.w6(32'hbadbf2a2),
	.w7(32'h3b00150c),
	.w8(32'hba8e0063),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8573f1),
	.w1(32'h3c177b86),
	.w2(32'h3b0c0504),
	.w3(32'hbb308195),
	.w4(32'h39c78ac9),
	.w5(32'hbbc8eade),
	.w6(32'hbb87e67e),
	.w7(32'h3a547917),
	.w8(32'h3b731a9c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a5428),
	.w1(32'h3b072304),
	.w2(32'hbae4b0fc),
	.w3(32'hbab7e9b1),
	.w4(32'h3b1644a1),
	.w5(32'h391fefab),
	.w6(32'h3b950ee7),
	.w7(32'h3c18dcfc),
	.w8(32'h3badf4a3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869c5c7),
	.w1(32'hbb111c93),
	.w2(32'hbb327510),
	.w3(32'h3b652bf7),
	.w4(32'hbbd4b400),
	.w5(32'hbb4c22ff),
	.w6(32'h3b3f3ade),
	.w7(32'hbac4e251),
	.w8(32'h3b564634),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034d40),
	.w1(32'hbbe2fe47),
	.w2(32'hbbea8f0d),
	.w3(32'hbb390f56),
	.w4(32'hbc1f38c6),
	.w5(32'hbbd1970e),
	.w6(32'h3adb6eda),
	.w7(32'hbbb2d939),
	.w8(32'hb96d249c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa65a62),
	.w1(32'h3bba33f1),
	.w2(32'h3acd6451),
	.w3(32'hbb4719e9),
	.w4(32'hb9f9f16d),
	.w5(32'hbbcdf744),
	.w6(32'hba68d3c3),
	.w7(32'hbaa88e93),
	.w8(32'hbaeae5fa),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134534),
	.w1(32'h3b8596ee),
	.w2(32'h3ab16c69),
	.w3(32'hbb99bd72),
	.w4(32'h3b945c12),
	.w5(32'hbbd7ad76),
	.w6(32'hbaf9c940),
	.w7(32'hbb52473b),
	.w8(32'hbbe505b4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ed1b),
	.w1(32'h3acdaa1b),
	.w2(32'hbb6c27a8),
	.w3(32'hbc070593),
	.w4(32'hbb11700f),
	.w5(32'hbbd2cf39),
	.w6(32'hbab04847),
	.w7(32'h3b475db4),
	.w8(32'h3a4ed17e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bcead),
	.w1(32'h3b02f99d),
	.w2(32'hbb6a069b),
	.w3(32'hbb920393),
	.w4(32'hbb58d393),
	.w5(32'hbc027402),
	.w6(32'hbab09b81),
	.w7(32'hbac951c2),
	.w8(32'hbb4a2164),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc086764),
	.w1(32'hbb3bf6a7),
	.w2(32'hbb27d0e8),
	.w3(32'hbb830184),
	.w4(32'hba674d38),
	.w5(32'hba598172),
	.w6(32'hbb46676d),
	.w7(32'hba6b3dcb),
	.w8(32'h3ab9a20b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f6535),
	.w1(32'h392324d8),
	.w2(32'h3b44300e),
	.w3(32'h3c05a683),
	.w4(32'hbaae77fd),
	.w5(32'hbb416c41),
	.w6(32'h3b82e465),
	.w7(32'h3ad4f5d3),
	.w8(32'hbb237992),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011f99),
	.w1(32'hb88ff206),
	.w2(32'h396d0441),
	.w3(32'hbc1b1bc3),
	.w4(32'hbbc13e80),
	.w5(32'hbb1048ea),
	.w6(32'h3a7d137e),
	.w7(32'hbb093908),
	.w8(32'h3b89a93e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20a59),
	.w1(32'h3b441eb9),
	.w2(32'hbb1a3bfc),
	.w3(32'hbbbda983),
	.w4(32'hbbb37c7f),
	.w5(32'hbbfe0517),
	.w6(32'h399ccc74),
	.w7(32'hbab3fa4c),
	.w8(32'hba4f67bd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9588e5),
	.w1(32'h3a30fa8e),
	.w2(32'h3b344801),
	.w3(32'hbb4dba7d),
	.w4(32'h3b6d4690),
	.w5(32'h3a8f1dad),
	.w6(32'hbb30381e),
	.w7(32'hbb762f20),
	.w8(32'hba19ce6c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4752),
	.w1(32'hbb35c395),
	.w2(32'hb9dac431),
	.w3(32'hbb81c636),
	.w4(32'hbba39c47),
	.w5(32'hbc2c3957),
	.w6(32'h3a2f9f01),
	.w7(32'hbb64cb52),
	.w8(32'hbb300ff9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad59d86),
	.w1(32'hbb8d6406),
	.w2(32'hbb5e2d7f),
	.w3(32'hbaba1183),
	.w4(32'h3b5cd6da),
	.w5(32'h3bade86a),
	.w6(32'h3b11d210),
	.w7(32'h3a378773),
	.w8(32'h3aa38d38),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69c7b),
	.w1(32'hbab152ed),
	.w2(32'hba5e1977),
	.w3(32'h3ad27cf1),
	.w4(32'hba695eed),
	.w5(32'hba9aa69f),
	.w6(32'hbbc6450a),
	.w7(32'h3a3041b4),
	.w8(32'h3b0e9c39),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad243d1),
	.w1(32'h3b7b0e78),
	.w2(32'h3aa501c7),
	.w3(32'hba96fd0f),
	.w4(32'h3b9166c6),
	.w5(32'h3a2fdfbc),
	.w6(32'h3b0df939),
	.w7(32'h3b9281df),
	.w8(32'h3afb8868),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bf3f4),
	.w1(32'h3adef240),
	.w2(32'h3bbfc091),
	.w3(32'h3c20fc35),
	.w4(32'h3b0bb7a4),
	.w5(32'hbbf8951c),
	.w6(32'h3b22da15),
	.w7(32'hbae9f81c),
	.w8(32'hba2ae2da),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351d48),
	.w1(32'hbb1d31a4),
	.w2(32'hbb1e7fff),
	.w3(32'hbbb8277d),
	.w4(32'hbb534900),
	.w5(32'hba6cf043),
	.w6(32'h3acdd5aa),
	.w7(32'h3b9f01f1),
	.w8(32'h3ba38ba0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ebdd6),
	.w1(32'h3aa75692),
	.w2(32'hbb8cc261),
	.w3(32'hb9b7a886),
	.w4(32'hbb258173),
	.w5(32'hbb88d768),
	.w6(32'h3baa47f3),
	.w7(32'h3a1f34ab),
	.w8(32'h3c1a3ce3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7413d),
	.w1(32'hbbb575e7),
	.w2(32'hbb77ef88),
	.w3(32'h39ad1970),
	.w4(32'hbaf8293c),
	.w5(32'hb9e139df),
	.w6(32'h3b6f3886),
	.w7(32'h3a0ac890),
	.w8(32'h39f879f8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d791),
	.w1(32'hba16b66d),
	.w2(32'hba4f8f5e),
	.w3(32'hbb03a612),
	.w4(32'hba3ebee7),
	.w5(32'hb953004b),
	.w6(32'hbaaf07b0),
	.w7(32'h36ccd1a2),
	.w8(32'hb9d33962),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fcee8),
	.w1(32'hba46c28f),
	.w2(32'hb9e704c8),
	.w3(32'hb9260efa),
	.w4(32'hba14b542),
	.w5(32'hba5fd2cf),
	.w6(32'hb86f67db),
	.w7(32'hb97080cf),
	.w8(32'h399c9bd8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7fab1),
	.w1(32'h3a4190a2),
	.w2(32'h3a3710fb),
	.w3(32'hb90ffc4b),
	.w4(32'hb9e94a9e),
	.w5(32'hb8e32116),
	.w6(32'h3911000f),
	.w7(32'hb8edbeed),
	.w8(32'hb930dd41),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de987e),
	.w1(32'hb4698850),
	.w2(32'h39838270),
	.w3(32'hb9dd576a),
	.w4(32'h39ae392b),
	.w5(32'h39477890),
	.w6(32'h396ea494),
	.w7(32'h39fb962b),
	.w8(32'h39fe4e51),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a712533),
	.w1(32'h3a17f048),
	.w2(32'h3a0c995f),
	.w3(32'h3a13479d),
	.w4(32'h39ae905b),
	.w5(32'h382ba4c8),
	.w6(32'h3a864787),
	.w7(32'hb889d816),
	.w8(32'h389c10d8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba755d79),
	.w1(32'hb98fb91c),
	.w2(32'h3ab5c647),
	.w3(32'hbae8d564),
	.w4(32'hba82e10c),
	.w5(32'hb9fcfb9d),
	.w6(32'hba623867),
	.w7(32'hb638f57a),
	.w8(32'h3abfc5d4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06823d),
	.w1(32'h39870a2c),
	.w2(32'h3a88cf9c),
	.w3(32'hb9821b9a),
	.w4(32'h3a146fb2),
	.w5(32'h38fdfb89),
	.w6(32'hbabf6720),
	.w7(32'hba300817),
	.w8(32'h39a7017c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed5a7c),
	.w1(32'h3a2cd5c9),
	.w2(32'h3a0e8221),
	.w3(32'hb9b6298a),
	.w4(32'h3a1b612b),
	.w5(32'h39f93548),
	.w6(32'hb996a561),
	.w7(32'h3a45343a),
	.w8(32'h3a49cfdd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9754e6d),
	.w1(32'hb9faaf21),
	.w2(32'hb9692c5a),
	.w3(32'h3961568f),
	.w4(32'hb9b769ea),
	.w5(32'hb9df676f),
	.w6(32'hba368819),
	.w7(32'hba0bc818),
	.w8(32'hba19988e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c1d7c),
	.w1(32'hb89d7200),
	.w2(32'h39ca867f),
	.w3(32'hbaaea0b6),
	.w4(32'hb9c1f741),
	.w5(32'hb9c49f2c),
	.w6(32'hbaa6502e),
	.w7(32'hb96f4e38),
	.w8(32'hb8fd5291),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba285521),
	.w1(32'h3a395c7e),
	.w2(32'hba13c893),
	.w3(32'hba043261),
	.w4(32'hb945586e),
	.w5(32'h393c1ff5),
	.w6(32'hb9f4cc7f),
	.w7(32'hb97bde4e),
	.w8(32'hb8099071),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055210),
	.w1(32'h3b0f8a2e),
	.w2(32'hb9ba787d),
	.w3(32'hbb07dcdc),
	.w4(32'h3ac30472),
	.w5(32'h3874742c),
	.w6(32'hbaa54f56),
	.w7(32'h3b3a308e),
	.w8(32'h3af3be60),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1422),
	.w1(32'h39c8cbd1),
	.w2(32'hb7cb1c51),
	.w3(32'h3a981948),
	.w4(32'h38ff3314),
	.w5(32'h37cab914),
	.w6(32'h3abd4bd3),
	.w7(32'hb8c0aab6),
	.w8(32'hb925f004),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39314dd9),
	.w1(32'h39b8e6d2),
	.w2(32'h3994483c),
	.w3(32'h38a0576f),
	.w4(32'h3a3e0477),
	.w5(32'h37eb0bb7),
	.w6(32'h3877eda6),
	.w7(32'h3a44bc1e),
	.w8(32'h3a34f837),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b4beb),
	.w1(32'h3a17ab22),
	.w2(32'hba26f644),
	.w3(32'hb9294cbe),
	.w4(32'h38995098),
	.w5(32'hb90e771e),
	.w6(32'h3a1cc84f),
	.w7(32'h399a4814),
	.w8(32'h39e83f06),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39854565),
	.w1(32'h3a86f3ad),
	.w2(32'hbaccbe53),
	.w3(32'hba3adf5e),
	.w4(32'hba9470ed),
	.w5(32'hba7141f2),
	.w6(32'h389ced8f),
	.w7(32'h383604fc),
	.w8(32'hba3c91a6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2df891),
	.w1(32'h3a625014),
	.w2(32'hbab26fa9),
	.w3(32'hba9fc6e7),
	.w4(32'h39038b8d),
	.w5(32'hba5067eb),
	.w6(32'hb9e13617),
	.w7(32'h39c54ef2),
	.w8(32'hb9ccd65d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998149b),
	.w1(32'hba0600b5),
	.w2(32'hba5f7db4),
	.w3(32'h37d6acbe),
	.w4(32'hb9a92461),
	.w5(32'hba0055b3),
	.w6(32'h38d75e48),
	.w7(32'h39d37a9e),
	.w8(32'h39ce2110),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0e2e9),
	.w1(32'hb98e60da),
	.w2(32'hb8e5d168),
	.w3(32'hba308c82),
	.w4(32'hba434154),
	.w5(32'hba4bed8e),
	.w6(32'hba6d184d),
	.w7(32'hb9c5854d),
	.w8(32'h38b2b632),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecd97d),
	.w1(32'h386ed91f),
	.w2(32'h38538f89),
	.w3(32'hba60867a),
	.w4(32'hb43f831c),
	.w5(32'h39f6be77),
	.w6(32'hb9d28158),
	.w7(32'h3a1d1ed1),
	.w8(32'h3a50068c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99756de),
	.w1(32'h39525316),
	.w2(32'h39518b83),
	.w3(32'h39fd7d63),
	.w4(32'hb8f3dc5f),
	.w5(32'hb9114ada),
	.w6(32'h3a182ff9),
	.w7(32'hb8da53d3),
	.w8(32'h39c11604),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb249de4),
	.w1(32'hba2f5f48),
	.w2(32'hbb595919),
	.w3(32'hbb26267b),
	.w4(32'hba7bc674),
	.w5(32'hbaa8f365),
	.w6(32'hbad0c5db),
	.w7(32'h3a4dee51),
	.w8(32'hb99d388e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0a543),
	.w1(32'hb99ed64e),
	.w2(32'hb9e1fa11),
	.w3(32'hba2ecda8),
	.w4(32'hba4196eb),
	.w5(32'hb934be01),
	.w6(32'hba2fb33f),
	.w7(32'hba6510cb),
	.w8(32'hba3c0f92),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba867ae4),
	.w1(32'h3a27948f),
	.w2(32'h3a89b5f2),
	.w3(32'hba22d977),
	.w4(32'h3a09ded0),
	.w5(32'h39a0884f),
	.w6(32'hbab64c91),
	.w7(32'h394266f8),
	.w8(32'h39cea802),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b28bdd),
	.w1(32'h3a3f88b8),
	.w2(32'h3a889001),
	.w3(32'hba6582f7),
	.w4(32'h396813b4),
	.w5(32'h39deaabc),
	.w6(32'hb944b2f9),
	.w7(32'hb9fb4a70),
	.w8(32'h39125b5f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991f58e),
	.w1(32'h3839653c),
	.w2(32'hba00b0ad),
	.w3(32'h39b47af2),
	.w4(32'hb9e2e7c1),
	.w5(32'h392b711f),
	.w6(32'h398fa3a4),
	.w7(32'hba1d01b8),
	.w8(32'h3940cc22),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934a6c0),
	.w1(32'hb981d39f),
	.w2(32'hb9583c55),
	.w3(32'h39256016),
	.w4(32'h390fc071),
	.w5(32'h3996f1b5),
	.w6(32'hb8f72f92),
	.w7(32'h3a124055),
	.w8(32'h39b237e3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398887f4),
	.w1(32'hb9832ae9),
	.w2(32'hba33a9a3),
	.w3(32'h3987f7f2),
	.w4(32'hba1808bb),
	.w5(32'hb98cf251),
	.w6(32'h39b1f864),
	.w7(32'hba17f467),
	.w8(32'hba0a91ce),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a36d),
	.w1(32'hb8d87856),
	.w2(32'h39879c7a),
	.w3(32'h390555b9),
	.w4(32'h38e484c9),
	.w5(32'h39c2bfca),
	.w6(32'h37e99696),
	.w7(32'hb8f70111),
	.w8(32'h370face7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382109dc),
	.w1(32'hb939abe8),
	.w2(32'hb977a8f5),
	.w3(32'hb88a8dcb),
	.w4(32'h3801a2d7),
	.w5(32'hb9466a18),
	.w6(32'hba511574),
	.w7(32'hba3d1912),
	.w8(32'hb9f1fe09),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7075e),
	.w1(32'hb9cfa0c9),
	.w2(32'hb9f94c90),
	.w3(32'hbacb2610),
	.w4(32'hbaafa8e4),
	.w5(32'hb9a8b302),
	.w6(32'hba9ec825),
	.w7(32'hba261446),
	.w8(32'hb74d9307),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba374ecf),
	.w1(32'h380342ce),
	.w2(32'h3990ecff),
	.w3(32'hba97928f),
	.w4(32'h38d554a9),
	.w5(32'hb94e6291),
	.w6(32'hba9e19c8),
	.w7(32'hb99ca188),
	.w8(32'h37ed1a1e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c8def),
	.w1(32'hb9a4c7db),
	.w2(32'hba3bb7fa),
	.w3(32'h39de55eb),
	.w4(32'hb9239622),
	.w5(32'hb9bc31b7),
	.w6(32'hb9372125),
	.w7(32'h39498d8d),
	.w8(32'hb9abd09e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f77a4),
	.w1(32'hb8aa90b7),
	.w2(32'hba4b0b94),
	.w3(32'hba9bd750),
	.w4(32'hba1b7a1c),
	.w5(32'hbaa9fb3b),
	.w6(32'hba659978),
	.w7(32'h39a17a0d),
	.w8(32'hba064ccd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26c24b),
	.w1(32'hb6f5c999),
	.w2(32'hba9578c1),
	.w3(32'hba37e11f),
	.w4(32'hb99cbc2b),
	.w5(32'hb9b73d38),
	.w6(32'h39627599),
	.w7(32'h3a14ff3b),
	.w8(32'h39a4de29),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa4492),
	.w1(32'hb98705f3),
	.w2(32'h3828dfd9),
	.w3(32'hb951b99c),
	.w4(32'hb701b01c),
	.w5(32'hb9466de6),
	.w6(32'h37ac1ada),
	.w7(32'h391cacdb),
	.w8(32'h39fa410f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51e541),
	.w1(32'h3a0afae9),
	.w2(32'hb9f3b6e3),
	.w3(32'hba4011e4),
	.w4(32'h3940dbc7),
	.w5(32'h3719a6ea),
	.w6(32'hb781cb74),
	.w7(32'h3a033274),
	.w8(32'h381efac5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c738b9),
	.w1(32'h38ebd844),
	.w2(32'hb8782e80),
	.w3(32'hb9802b32),
	.w4(32'h39f19292),
	.w5(32'hb8cc1919),
	.w6(32'h38b92f48),
	.w7(32'h39746531),
	.w8(32'h39ac1bdf),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927462e),
	.w1(32'hba6d98b9),
	.w2(32'hba2a8db7),
	.w3(32'h399d0e3a),
	.w4(32'hba102279),
	.w5(32'hba17a3fa),
	.w6(32'h3a04cecd),
	.w7(32'h389d4f60),
	.w8(32'hba00d087),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a3b95),
	.w1(32'h39567ed5),
	.w2(32'h39986756),
	.w3(32'hb913e929),
	.w4(32'h3871b031),
	.w5(32'hb90d023b),
	.w6(32'hb9145d41),
	.w7(32'hb9b5d265),
	.w8(32'hb9b5ebfa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84bb0d5),
	.w1(32'hba525f00),
	.w2(32'hba054b95),
	.w3(32'hb9f6ad92),
	.w4(32'hb9d2dbee),
	.w5(32'hb9802242),
	.w6(32'hb9af3310),
	.w7(32'h39449091),
	.w8(32'h3958ae4e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba005cb0),
	.w1(32'h35812cc0),
	.w2(32'h39361666),
	.w3(32'hba771377),
	.w4(32'h395cdcd3),
	.w5(32'hb9b44de3),
	.w6(32'hba145ed9),
	.w7(32'h37f67e7a),
	.w8(32'h3766829e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d160b),
	.w1(32'h3a52379c),
	.w2(32'hbb014263),
	.w3(32'hbaadeeed),
	.w4(32'hb9ba59e3),
	.w5(32'hba7fca32),
	.w6(32'hb905e03b),
	.w7(32'h398642af),
	.w8(32'hbaa94286),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b3484),
	.w1(32'h3a18c563),
	.w2(32'hba1ac147),
	.w3(32'hba7fe526),
	.w4(32'h39342917),
	.w5(32'hb8db2a1e),
	.w6(32'hba479b2d),
	.w7(32'h3a66fdb7),
	.w8(32'h38f03e92),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fe576),
	.w1(32'hb8dfc7dd),
	.w2(32'hbaf9d23e),
	.w3(32'hba9f8c3d),
	.w4(32'hba6f4d47),
	.w5(32'hba5a2629),
	.w6(32'hba5d85bd),
	.w7(32'hb96f32b7),
	.w8(32'hba6ccfbd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44a42c),
	.w1(32'h396c508e),
	.w2(32'h392e1b00),
	.w3(32'h3998365d),
	.w4(32'h37ab60ea),
	.w5(32'hb9ad4b42),
	.w6(32'h3991d666),
	.w7(32'hb8aefd89),
	.w8(32'hba013221),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f8e2bf),
	.w1(32'h39a9935e),
	.w2(32'hb8092edb),
	.w3(32'hb9699d80),
	.w4(32'h39dbd889),
	.w5(32'h38b313b5),
	.w6(32'hb94d15a8),
	.w7(32'h39c9c0a0),
	.w8(32'h395c6b37),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393743e3),
	.w1(32'hb9d04828),
	.w2(32'hb9cd630f),
	.w3(32'h391755d0),
	.w4(32'hb9859336),
	.w5(32'h39440ed0),
	.w6(32'h399c2f8f),
	.w7(32'h392bf99a),
	.w8(32'hb86a2438),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8907458),
	.w1(32'h3a246047),
	.w2(32'h3973b2cf),
	.w3(32'hb9943f5c),
	.w4(32'h39b4b157),
	.w5(32'hb9d76ae4),
	.w6(32'hb9d8053b),
	.w7(32'hb9f122ba),
	.w8(32'hb9ff0cad),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23fde1),
	.w1(32'hb9a7b675),
	.w2(32'hb93ffbc0),
	.w3(32'hba9c9069),
	.w4(32'hba2158f4),
	.w5(32'hba425cc9),
	.w6(32'hb880f5d1),
	.w7(32'hb911f1a9),
	.w8(32'hb8bb1f6f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2d513),
	.w1(32'hb9fd8494),
	.w2(32'hba4e2ea9),
	.w3(32'hb9d65c8b),
	.w4(32'hb9faac70),
	.w5(32'h3907a649),
	.w6(32'h39505147),
	.w7(32'hb9efa017),
	.w8(32'hb9aec174),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8294e7),
	.w1(32'h39ba66ea),
	.w2(32'h3a1ad5cd),
	.w3(32'hb9d23c22),
	.w4(32'h38010fae),
	.w5(32'h3a17984a),
	.w6(32'hb9fd4d3c),
	.w7(32'h38b7ba5f),
	.w8(32'h39e64bad),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977ff96),
	.w1(32'hb92c7406),
	.w2(32'h3961f805),
	.w3(32'h3a0ecd82),
	.w4(32'hb966072b),
	.w5(32'h39b72497),
	.w6(32'h38da50c8),
	.w7(32'hb9564c2f),
	.w8(32'h3a02e314),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b8df16),
	.w1(32'hb95f95c0),
	.w2(32'hb9fff973),
	.w3(32'hb908d4e5),
	.w4(32'hb9a66e27),
	.w5(32'hb892a53b),
	.w6(32'hb75a68c9),
	.w7(32'hb80b8f0f),
	.w8(32'h387ccb33),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba394b70),
	.w1(32'h399f910a),
	.w2(32'hba35d8c2),
	.w3(32'hb96be8dc),
	.w4(32'hb907c1b5),
	.w5(32'hb9ea0b60),
	.w6(32'hb9a831d7),
	.w7(32'h36ad9ccf),
	.w8(32'hb989ccd0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b2b68),
	.w1(32'h39b3611c),
	.w2(32'h39f31d39),
	.w3(32'hba17ff53),
	.w4(32'hb99a1766),
	.w5(32'h39574c4d),
	.w6(32'hba582adc),
	.w7(32'h3920437b),
	.w8(32'hb944b221),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38574f83),
	.w1(32'h3a41fef3),
	.w2(32'hbac2fb63),
	.w3(32'hbab03130),
	.w4(32'hb9d1ad2c),
	.w5(32'hba92a246),
	.w6(32'hbaa41a60),
	.w7(32'hb9b24b2e),
	.w8(32'hbaaeaa70),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e89703),
	.w1(32'hba29332b),
	.w2(32'hba53b123),
	.w3(32'hb9ff9772),
	.w4(32'hb98b630b),
	.w5(32'hb97aa2ad),
	.w6(32'h37be89a9),
	.w7(32'hba2d107e),
	.w8(32'hba3a9a88),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac50997),
	.w1(32'h398c7480),
	.w2(32'h3a4bc4a4),
	.w3(32'hbac9e217),
	.w4(32'h3a3e11aa),
	.w5(32'h3a0871a4),
	.w6(32'hbaba9e58),
	.w7(32'h3899011e),
	.w8(32'h3a77cd10),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule