module layer_10_featuremap_391(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31eb89),
	.w1(32'hb96e22f0),
	.w2(32'hba5befc5),
	.w3(32'hbad04bbb),
	.w4(32'hb80b34cf),
	.w5(32'hba4e5072),
	.w6(32'hb9b28f69),
	.w7(32'h3a464f6e),
	.w8(32'hb92d23ec),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387eef20),
	.w1(32'h39ac68d3),
	.w2(32'hbac4f94f),
	.w3(32'hb918a5c7),
	.w4(32'h3a3e17bb),
	.w5(32'h37b57d00),
	.w6(32'hba8cc7f1),
	.w7(32'hb8fff38b),
	.w8(32'hb94a5c9d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169489),
	.w1(32'hb9fea255),
	.w2(32'hba167079),
	.w3(32'hba866036),
	.w4(32'hbaa9a01c),
	.w5(32'hbacb91c5),
	.w6(32'hbaa21d73),
	.w7(32'hbad9d0ba),
	.w8(32'h3978c7f4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3a4d7),
	.w1(32'hba4d8a1d),
	.w2(32'hb9987931),
	.w3(32'h39d649db),
	.w4(32'hba7ac84f),
	.w5(32'hba86a51a),
	.w6(32'h399ac302),
	.w7(32'h3a257dcc),
	.w8(32'h39497a6a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf8bfb),
	.w1(32'hb8cca555),
	.w2(32'hbb117f8b),
	.w3(32'h3a79e10b),
	.w4(32'h37c0cf46),
	.w5(32'hb9517acc),
	.w6(32'h3ae2e091),
	.w7(32'h390e99ad),
	.w8(32'hb99055ad),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42c47c),
	.w1(32'hba39f101),
	.w2(32'h398c852c),
	.w3(32'hb9efcb6e),
	.w4(32'h39f82cef),
	.w5(32'hb99768b8),
	.w6(32'hba92b392),
	.w7(32'h3a4663c8),
	.w8(32'h39173093),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7dd04),
	.w1(32'h3ac2ea94),
	.w2(32'h391a5c3e),
	.w3(32'hbb101b11),
	.w4(32'hba79b323),
	.w5(32'hb9bb5915),
	.w6(32'hbaa9e017),
	.w7(32'h3ab4127c),
	.w8(32'h3ac1aafa),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4b294),
	.w1(32'h39de54d5),
	.w2(32'hba85cf0a),
	.w3(32'hb99368a3),
	.w4(32'hbb0c3e37),
	.w5(32'hbb3362ad),
	.w6(32'h3a074cd3),
	.w7(32'hbad6d8d9),
	.w8(32'hb9ab15ab),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d81c0),
	.w1(32'h3a604817),
	.w2(32'hb9f8822d),
	.w3(32'h3a34c4bb),
	.w4(32'hba4be88f),
	.w5(32'hb990c69a),
	.w6(32'h3a35dbd8),
	.w7(32'h39d6a09e),
	.w8(32'h3a673000),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eee42),
	.w1(32'hbac4e128),
	.w2(32'hba66d2c0),
	.w3(32'hba4bbff9),
	.w4(32'hbae079b7),
	.w5(32'hb9703636),
	.w6(32'hbae51716),
	.w7(32'hba240c1e),
	.w8(32'hba624e26),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7e00),
	.w1(32'hbaae038f),
	.w2(32'hbaa26fe0),
	.w3(32'hba182016),
	.w4(32'hbaa1aa21),
	.w5(32'hb9f84a24),
	.w6(32'hba97283e),
	.w7(32'h396b234b),
	.w8(32'h3991786a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae50877),
	.w1(32'h3aad7d22),
	.w2(32'h3a4513cf),
	.w3(32'hbaed3da7),
	.w4(32'h3a3dd8c1),
	.w5(32'h38bc4de1),
	.w6(32'hba51444b),
	.w7(32'h3a23ee98),
	.w8(32'h3a065a3b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b498308),
	.w1(32'hba446442),
	.w2(32'hbb3155c7),
	.w3(32'h3b3f10c9),
	.w4(32'h39e50bb3),
	.w5(32'hbadb818a),
	.w6(32'h3b3ab1ba),
	.w7(32'hb8be1285),
	.w8(32'hba5ad3c0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca792),
	.w1(32'hba4d34a2),
	.w2(32'hb9ec1415),
	.w3(32'hba13cffd),
	.w4(32'hba90e6a9),
	.w5(32'h393eaa07),
	.w6(32'hb89e6f34),
	.w7(32'hbab89bdd),
	.w8(32'hbaabf5d3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba976d72),
	.w1(32'hba23b12a),
	.w2(32'hbaa156be),
	.w3(32'hbac973ed),
	.w4(32'hba4ca755),
	.w5(32'hbaa4be0b),
	.w6(32'hbb2619c0),
	.w7(32'hba4bbde4),
	.w8(32'h367337e7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977168a),
	.w1(32'hbb12f29e),
	.w2(32'hbb244def),
	.w3(32'hbacf97a6),
	.w4(32'hbb2daca4),
	.w5(32'hbb2f07da),
	.w6(32'hba03a1b2),
	.w7(32'hbb305170),
	.w8(32'hbb1698bf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8030d),
	.w1(32'h3a3e6d47),
	.w2(32'h3a76b672),
	.w3(32'hbae5efd6),
	.w4(32'hb6ecde62),
	.w5(32'h3a8f1f63),
	.w6(32'hba282466),
	.w7(32'hb9fb49e9),
	.w8(32'h387119b0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b4d1),
	.w1(32'h3a8ba8d0),
	.w2(32'h3b190090),
	.w3(32'h3ad70a6d),
	.w4(32'h3abd1023),
	.w5(32'h3ac4a9f0),
	.w6(32'hba589c60),
	.w7(32'h39f6a7ba),
	.w8(32'hba5b220b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a866ced),
	.w1(32'hba5e4ad8),
	.w2(32'hbaddb430),
	.w3(32'h3aafcc11),
	.w4(32'hba954d95),
	.w5(32'hba6c2ea7),
	.w6(32'h3a0cacf3),
	.w7(32'hba5b937f),
	.w8(32'h39ad1e6c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab9112),
	.w1(32'hba8a3c00),
	.w2(32'hba848416),
	.w3(32'h3ad32f09),
	.w4(32'hbabfc5ee),
	.w5(32'hb8e1a0f8),
	.w6(32'h3a634593),
	.w7(32'hbac9e529),
	.w8(32'hbaa745aa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04dcbd),
	.w1(32'h3b0fd332),
	.w2(32'h3ac25c2e),
	.w3(32'hb976717c),
	.w4(32'h3b15edb9),
	.w5(32'hb83076d7),
	.w6(32'h3b15b795),
	.w7(32'h3a305621),
	.w8(32'hb9a27838),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d347ed),
	.w1(32'hbaaee258),
	.w2(32'h3abc1afb),
	.w3(32'hba8ef63c),
	.w4(32'hbb23c41f),
	.w5(32'h3a2a1a71),
	.w6(32'hb9f402aa),
	.w7(32'hba83c03a),
	.w8(32'hba4b46a4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10820e),
	.w1(32'h3a431b5f),
	.w2(32'hba8ed421),
	.w3(32'h39f430c8),
	.w4(32'hb9d7b655),
	.w5(32'h3adc6fca),
	.w6(32'h3ac295ce),
	.w7(32'hba278579),
	.w8(32'hbb46e73d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22613e),
	.w1(32'hbb300c9d),
	.w2(32'hbb841123),
	.w3(32'hbb10b28a),
	.w4(32'hbb1cb10c),
	.w5(32'hbb4e486f),
	.w6(32'hbb41ccc0),
	.w7(32'hb94f5c03),
	.w8(32'hbac8dbeb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8a78e),
	.w1(32'hbad9025a),
	.w2(32'hb9af37ea),
	.w3(32'hb91ec4a9),
	.w4(32'hb9ade022),
	.w5(32'h38f82f55),
	.w6(32'h3ad4f058),
	.w7(32'hba018b06),
	.w8(32'hbb388f6a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e016e),
	.w1(32'h3b27ae05),
	.w2(32'h39e2cd17),
	.w3(32'hb9674f69),
	.w4(32'h3a8ef589),
	.w5(32'h39f44091),
	.w6(32'hbae80ca6),
	.w7(32'h3a875fdd),
	.w8(32'hb9b7c3e4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a184a47),
	.w1(32'hba8c8393),
	.w2(32'hbadcabdb),
	.w3(32'h3a43b48d),
	.w4(32'hbae9b053),
	.w5(32'hba7d5c2b),
	.w6(32'h39818a10),
	.w7(32'hba8c136b),
	.w8(32'h39888dd0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2376),
	.w1(32'hba5b5b23),
	.w2(32'hba33767f),
	.w3(32'hb9de819f),
	.w4(32'hbae8be48),
	.w5(32'hb94ecd68),
	.w6(32'hba38a984),
	.w7(32'hba92d9e9),
	.w8(32'h3a5ca2d6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998bd7a),
	.w1(32'hbb02a606),
	.w2(32'hba040719),
	.w3(32'hba1838d7),
	.w4(32'hb9f7e140),
	.w5(32'h399d23e6),
	.w6(32'hbaa4c65c),
	.w7(32'hbaf042c5),
	.w8(32'hbb3cada5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac33e),
	.w1(32'h3a3e3271),
	.w2(32'h3a09c462),
	.w3(32'hbb1daebe),
	.w4(32'h3ace8f58),
	.w5(32'hba9b353d),
	.w6(32'hbb309114),
	.w7(32'h3a9af8d5),
	.w8(32'hbada1ac2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1068),
	.w1(32'h39f7158f),
	.w2(32'hb823450f),
	.w3(32'h3a094fb2),
	.w4(32'hb90f22d2),
	.w5(32'h3a4fe396),
	.w6(32'hb8f466e1),
	.w7(32'hb9a5dd16),
	.w8(32'hba81a661),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39feb4af),
	.w1(32'hbb003583),
	.w2(32'hba9e3754),
	.w3(32'hb6d93d21),
	.w4(32'hbac3ec3f),
	.w5(32'hb95c2ba8),
	.w6(32'hba517682),
	.w7(32'hbab5956b),
	.w8(32'hb9fd4743),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39859de4),
	.w1(32'hbb47e88b),
	.w2(32'hbb3d3fe6),
	.w3(32'h3a6f5543),
	.w4(32'hba90d6b5),
	.w5(32'hba0d44d2),
	.w6(32'hba25d75d),
	.w7(32'h38ba365b),
	.w8(32'hb960d9d2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310996),
	.w1(32'hba53317b),
	.w2(32'hbae316b2),
	.w3(32'hb990f7f5),
	.w4(32'hba0598d4),
	.w5(32'h3a229787),
	.w6(32'hba839768),
	.w7(32'h3a6fe390),
	.w8(32'h3a9cff3c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820fff),
	.w1(32'h3ae3b55d),
	.w2(32'h3b0dd2be),
	.w3(32'h39aeebd1),
	.w4(32'h3a825d17),
	.w5(32'hba16a651),
	.w6(32'hba18bf42),
	.w7(32'h3a8bb4fe),
	.w8(32'hbb042cb0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b707d1a),
	.w1(32'h3a769121),
	.w2(32'h3a9d2055),
	.w3(32'h3a4b0b64),
	.w4(32'h3ac4cb71),
	.w5(32'hbae3f006),
	.w6(32'hb5038de6),
	.w7(32'h3ae1639b),
	.w8(32'h39b052ca),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f82a),
	.w1(32'h3b009c89),
	.w2(32'h3970604e),
	.w3(32'hb7098896),
	.w4(32'h3af34a28),
	.w5(32'h3a28709c),
	.w6(32'h3a934599),
	.w7(32'h3af9b01e),
	.w8(32'h3a38d80e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2776a0),
	.w1(32'h3b027e7c),
	.w2(32'h39d6e054),
	.w3(32'hb9d6ee1b),
	.w4(32'h3ad2a89a),
	.w5(32'h3ab0d26e),
	.w6(32'hba3251b8),
	.w7(32'h3afb1bba),
	.w8(32'h3a4d9667),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8acc0),
	.w1(32'h3ae90850),
	.w2(32'h39a04587),
	.w3(32'h3aa8b03e),
	.w4(32'h3a3bb0bc),
	.w5(32'h39c29b5d),
	.w6(32'h3a35a46d),
	.w7(32'h3a9e57a6),
	.w8(32'h3ade76c1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837e022),
	.w1(32'hb9a3e439),
	.w2(32'hbaa5042c),
	.w3(32'hbab2b754),
	.w4(32'hbabcd643),
	.w5(32'hb992ef1a),
	.w6(32'hbb19b98f),
	.w7(32'hba6230a9),
	.w8(32'h3963b06e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1b01f),
	.w1(32'hbb494fa1),
	.w2(32'hbac47b9e),
	.w3(32'h3ae9fedc),
	.w4(32'h390a146b),
	.w5(32'h3b05f3d4),
	.w6(32'hba38ec6e),
	.w7(32'h3a4954a3),
	.w8(32'hb944a895),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60160),
	.w1(32'h3949b2d7),
	.w2(32'h39be51bc),
	.w3(32'h3abcdb3c),
	.w4(32'h3aadf065),
	.w5(32'h3abeba0a),
	.w6(32'h39e337a5),
	.w7(32'hb9b775b8),
	.w8(32'h3a16a486),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a669482),
	.w1(32'hba29263d),
	.w2(32'hbacc1d7b),
	.w3(32'h3ad0f9c7),
	.w4(32'hb93335b0),
	.w5(32'hbaa13175),
	.w6(32'h3a9f681a),
	.w7(32'h3963d9f4),
	.w8(32'hb995e3bc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6751e),
	.w1(32'h376e607c),
	.w2(32'hbb46d61f),
	.w3(32'h3851a235),
	.w4(32'h3a4b9196),
	.w5(32'hbafbd3fe),
	.w6(32'h3a088b35),
	.w7(32'h3a561bc2),
	.w8(32'hba8db4b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59de5e),
	.w1(32'hbaa3e003),
	.w2(32'hba14732f),
	.w3(32'h3aebc120),
	.w4(32'hba5336d6),
	.w5(32'h3b026b16),
	.w6(32'h3aab87d8),
	.w7(32'hba6ec0a0),
	.w8(32'h3ab02464),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951cfac),
	.w1(32'hbb103401),
	.w2(32'hbb464db2),
	.w3(32'h397c1e7f),
	.w4(32'hbb37fccc),
	.w5(32'hbb64b080),
	.w6(32'h397b0215),
	.w7(32'hbb462eb6),
	.w8(32'hbb68e5c9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93e32),
	.w1(32'hb8a7a6df),
	.w2(32'h3a94db4d),
	.w3(32'hbb5b0a31),
	.w4(32'hbabae09c),
	.w5(32'hb9c37a98),
	.w6(32'hbaaa3793),
	.w7(32'hba06123b),
	.w8(32'hb9675038),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba793713),
	.w1(32'hbabd4130),
	.w2(32'hb9e68569),
	.w3(32'hba8445db),
	.w4(32'hbb0e7978),
	.w5(32'hb97fe71d),
	.w6(32'hb9ef3f2a),
	.w7(32'hbac6f9f1),
	.w8(32'hb919f30d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ac6f8),
	.w1(32'h3ada3dda),
	.w2(32'h396494db),
	.w3(32'h394b478e),
	.w4(32'h3919067b),
	.w5(32'hbacae583),
	.w6(32'h396637b2),
	.w7(32'h39940030),
	.w8(32'hb9c3d77e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9516510),
	.w1(32'h38a86df0),
	.w2(32'h3b11f510),
	.w3(32'hbab974f2),
	.w4(32'h3aa43bc9),
	.w5(32'hbae836f0),
	.w6(32'hba9b0d3c),
	.w7(32'h3a75aac8),
	.w8(32'h37711edc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b971),
	.w1(32'h3a578d0b),
	.w2(32'hbacef4c9),
	.w3(32'h3b01398a),
	.w4(32'h3a37a881),
	.w5(32'hba3d1e0a),
	.w6(32'h3ab867d2),
	.w7(32'h39b015a0),
	.w8(32'hba9eafa2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0444a0),
	.w1(32'hbb12f4fa),
	.w2(32'h3977d316),
	.w3(32'hbacdd832),
	.w4(32'hbb3126eb),
	.w5(32'hb97138b2),
	.w6(32'hba22ca7e),
	.w7(32'hbb4cdd47),
	.w8(32'hbaa3d1ce),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e0bb),
	.w1(32'h3a8377bd),
	.w2(32'h3ab56aa1),
	.w3(32'hbac23dfc),
	.w4(32'h39b6fc73),
	.w5(32'h3977f843),
	.w6(32'hbb0f6e50),
	.w7(32'h3ac873b8),
	.w8(32'h3a024f20),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2dc7),
	.w1(32'hb9cda835),
	.w2(32'hba7dbe71),
	.w3(32'h3b188ef2),
	.w4(32'hb8e815fe),
	.w5(32'hba9d1f25),
	.w6(32'h3ae251c5),
	.w7(32'h399121fa),
	.w8(32'hbaf3e353),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdd5e0),
	.w1(32'hb9836195),
	.w2(32'hba0d52f4),
	.w3(32'h3ab6b0f9),
	.w4(32'hbab54eb5),
	.w5(32'hba976b9b),
	.w6(32'h3954491f),
	.w7(32'hba87c139),
	.w8(32'hb9d1b471),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f2a89),
	.w1(32'hb9bfbed6),
	.w2(32'hbadfff9d),
	.w3(32'h3a834bc6),
	.w4(32'h39d39af5),
	.w5(32'hba5d99c7),
	.w6(32'hba7e06fe),
	.w7(32'h3adcc083),
	.w8(32'hb9af578d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb035183),
	.w1(32'hba1252ac),
	.w2(32'hbb1aca2a),
	.w3(32'hbaac9208),
	.w4(32'h3a7f1a66),
	.w5(32'hba037467),
	.w6(32'hbac4b26f),
	.w7(32'h3a76b051),
	.w8(32'h394b456a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93c125),
	.w1(32'hb8b1c0aa),
	.w2(32'h3a989e64),
	.w3(32'hba0a7281),
	.w4(32'hba054a8c),
	.w5(32'h3a8869de),
	.w6(32'h39a3ad4c),
	.w7(32'hbabde509),
	.w8(32'h3b396308),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43b8ec),
	.w1(32'hbb0e38be),
	.w2(32'hbaff83be),
	.w3(32'hba68ab84),
	.w4(32'hbb2c925c),
	.w5(32'hba7a8e4d),
	.w6(32'h390a723d),
	.w7(32'hbb3aa543),
	.w8(32'hbabc0fa7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacba4f8),
	.w1(32'hbaadd21f),
	.w2(32'hba1b5925),
	.w3(32'hba7146ca),
	.w4(32'hb9eadad5),
	.w5(32'hbb1e9842),
	.w6(32'hbaa516e7),
	.w7(32'h3a906318),
	.w8(32'hb989785e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a1731),
	.w1(32'h3aad2286),
	.w2(32'h392880c1),
	.w3(32'h3a6b7ca3),
	.w4(32'hb964b349),
	.w5(32'hba9e4910),
	.w6(32'hb9b79c34),
	.w7(32'hba24420d),
	.w8(32'hba53edcf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a250f02),
	.w1(32'hbab1d60d),
	.w2(32'hba86848e),
	.w3(32'hba899756),
	.w4(32'hbb0de472),
	.w5(32'hb91ca065),
	.w6(32'hb9a81892),
	.w7(32'hbb159f15),
	.w8(32'hb97a9f8d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4e59),
	.w1(32'hba320dc7),
	.w2(32'hba4717c1),
	.w3(32'h39317b78),
	.w4(32'h3a02661e),
	.w5(32'h39aa8f4a),
	.w6(32'hbab4ea9f),
	.w7(32'h39d6dc0f),
	.w8(32'hba82ec36),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63100a),
	.w1(32'hba57cf74),
	.w2(32'hba7f7924),
	.w3(32'h3ae0d1ea),
	.w4(32'hba8a3bc8),
	.w5(32'h39e219f5),
	.w6(32'h3a49d2ce),
	.w7(32'h394ce87e),
	.w8(32'h3a8064ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39331e3e),
	.w1(32'h3af2d651),
	.w2(32'h3aa5920e),
	.w3(32'h3b0698aa),
	.w4(32'h3ab7784f),
	.w5(32'h398200c3),
	.w6(32'h3aedbbbb),
	.w7(32'h3ae2df04),
	.w8(32'h385b6d1a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6ab4),
	.w1(32'h3a9d6f42),
	.w2(32'hb913387f),
	.w3(32'h3ad38832),
	.w4(32'h3a6f09c2),
	.w5(32'h3912b98e),
	.w6(32'h3a2ce2e7),
	.w7(32'hba45ee38),
	.w8(32'h3a84fe70),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6eac9),
	.w1(32'hbaa49e13),
	.w2(32'hbabf0608),
	.w3(32'hba8f524c),
	.w4(32'hbab7f88b),
	.w5(32'hb9b52514),
	.w6(32'hb9bc570e),
	.w7(32'hbab09c57),
	.w8(32'hbb04d2d6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f4a70),
	.w1(32'h3a817b49),
	.w2(32'hba893cd0),
	.w3(32'hbae82023),
	.w4(32'h39ab62cb),
	.w5(32'hbb4b271c),
	.w6(32'hbac0b52f),
	.w7(32'hb9be9c64),
	.w8(32'hba490f1e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa53f6e),
	.w1(32'h3a8080f6),
	.w2(32'hba80cb66),
	.w3(32'hbb0a535f),
	.w4(32'hb9c3cfe7),
	.w5(32'hb9a0030e),
	.w6(32'h37be59b6),
	.w7(32'hba584806),
	.w8(32'h39deed01),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb085ccf),
	.w1(32'hb732338d),
	.w2(32'hba225a86),
	.w3(32'hbaddbcbf),
	.w4(32'hbab29fda),
	.w5(32'h39cf04a0),
	.w6(32'hbb065a19),
	.w7(32'hba9aee4c),
	.w8(32'h3a713e4e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4680ef),
	.w1(32'h3aa75b43),
	.w2(32'hbba2593e),
	.w3(32'hba10ad70),
	.w4(32'h3ae0adb3),
	.w5(32'h3a5ebc94),
	.w6(32'hbb427e22),
	.w7(32'h3bd06ac1),
	.w8(32'h3ba3645c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2fbf),
	.w1(32'h3b3a3d37),
	.w2(32'h3c03be60),
	.w3(32'hbb12a2f1),
	.w4(32'h3b10b3c7),
	.w5(32'h3aec8e9a),
	.w6(32'h3b8c457f),
	.w7(32'hbadef791),
	.w8(32'h3b1264f2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bcb16),
	.w1(32'hbb346466),
	.w2(32'hbb4aa8c2),
	.w3(32'hbb02bd44),
	.w4(32'hbb5bd619),
	.w5(32'hba4f21f2),
	.w6(32'hbb284650),
	.w7(32'hbb55b071),
	.w8(32'hba6953ca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedce82),
	.w1(32'hb95c2ab4),
	.w2(32'h3c0dea11),
	.w3(32'h3aafcdfe),
	.w4(32'hbc0fb7b9),
	.w5(32'h3a82bee7),
	.w6(32'h3c0533a8),
	.w7(32'hbc0540de),
	.w8(32'hba5c98a2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3b7e0),
	.w1(32'hbb22108d),
	.w2(32'hbb40d0f3),
	.w3(32'h3af07391),
	.w4(32'hbb93bddc),
	.w5(32'hbc137fa2),
	.w6(32'h3ace1896),
	.w7(32'h3a156bf9),
	.w8(32'hba1e925a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9e86),
	.w1(32'hbb78229b),
	.w2(32'hbbde4077),
	.w3(32'hbc1c7854),
	.w4(32'hbbecf477),
	.w5(32'hbb69bc1e),
	.w6(32'hbb8ae3a7),
	.w7(32'hbb90555d),
	.w8(32'hbba2f01f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb874631),
	.w1(32'h3a5a9ad2),
	.w2(32'h3aecc5e1),
	.w3(32'hbba5bfc1),
	.w4(32'h3b8c34f2),
	.w5(32'h3b482523),
	.w6(32'hba085c87),
	.w7(32'hbaaabf19),
	.w8(32'hbaf7c80e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9b28f),
	.w1(32'h3b41e874),
	.w2(32'h3c4ef39e),
	.w3(32'h3b6264a2),
	.w4(32'h3c877a7e),
	.w5(32'h3ca7692c),
	.w6(32'hbb2fb5ce),
	.w7(32'h3c36751a),
	.w8(32'h3c24b85b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf90b0d),
	.w1(32'h3b344d4a),
	.w2(32'h3b5bf57d),
	.w3(32'h3c730e5f),
	.w4(32'h3ab24b8d),
	.w5(32'h39c229ae),
	.w6(32'h3c1d75df),
	.w7(32'h3b65e3d9),
	.w8(32'hb8848dc2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b787254),
	.w1(32'hb8c52c1e),
	.w2(32'hbad7bd03),
	.w3(32'h3a091600),
	.w4(32'h3b4813f9),
	.w5(32'hb9cb89e4),
	.w6(32'hbb25ce7e),
	.w7(32'h3b7ea9df),
	.w8(32'h3b8df61c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f19ea),
	.w1(32'h3be15f41),
	.w2(32'h3c418029),
	.w3(32'h3aabb607),
	.w4(32'h3beb25cb),
	.w5(32'h3c3d018b),
	.w6(32'h3a5028d9),
	.w7(32'h3a9d3a3c),
	.w8(32'h3b4417c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf292f2),
	.w1(32'hbb83146c),
	.w2(32'hbb478b9d),
	.w3(32'h3bfabc1b),
	.w4(32'hbbc5bad6),
	.w5(32'hbb5c1ebb),
	.w6(32'h39fc6863),
	.w7(32'hbbb1f896),
	.w8(32'hbb308879),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922aa6),
	.w1(32'hbc80cb67),
	.w2(32'hbc322009),
	.w3(32'hbaba30df),
	.w4(32'hbc0e1e9f),
	.w5(32'hbc092dde),
	.w6(32'hba7366eb),
	.w7(32'hbc51c18c),
	.w8(32'hbc1ccfd8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e999e),
	.w1(32'h3b355d24),
	.w2(32'hbb5867a1),
	.w3(32'hbb982327),
	.w4(32'h3a8d5957),
	.w5(32'hbac34215),
	.w6(32'hbc33400e),
	.w7(32'h3b088a2d),
	.w8(32'hbbd19187),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e4c5),
	.w1(32'h3ad92199),
	.w2(32'h3b4e6801),
	.w3(32'hbc13c629),
	.w4(32'h3abd4e80),
	.w5(32'hbb19ef2f),
	.w6(32'hbbdd57d1),
	.w7(32'hbb6b9870),
	.w8(32'hbbd335dc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf21bee),
	.w1(32'h3b23a4ab),
	.w2(32'hbb1cc21f),
	.w3(32'h395b6ad7),
	.w4(32'h3b625d2a),
	.w5(32'hbb252a11),
	.w6(32'hbb8a53a2),
	.w7(32'hbb8936bf),
	.w8(32'hbbf550d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcffe2),
	.w1(32'hbad6653c),
	.w2(32'h3bfd91da),
	.w3(32'hbb6fe27d),
	.w4(32'h3b126891),
	.w5(32'h3b536f6d),
	.w6(32'hbb15fac0),
	.w7(32'h3a9cd149),
	.w8(32'h3b3202be),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066a88),
	.w1(32'h3aa6482b),
	.w2(32'h3b37592f),
	.w3(32'h3bd6db8d),
	.w4(32'h3bf0a8aa),
	.w5(32'h3b429dd0),
	.w6(32'h3b54789b),
	.w7(32'hbba0c657),
	.w8(32'hbc20eeb5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a935a6c),
	.w1(32'hbb96562f),
	.w2(32'hbbc18fbe),
	.w3(32'h3a5569f9),
	.w4(32'hbb7062e3),
	.w5(32'hb95994f7),
	.w6(32'hbbd714de),
	.w7(32'hbbdd17d0),
	.w8(32'hbb97ee1f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe89c23),
	.w1(32'hbb4ae213),
	.w2(32'hbb6c3e3f),
	.w3(32'hbbb760a2),
	.w4(32'hbba19008),
	.w5(32'hbb90a3ef),
	.w6(32'hbbf40a70),
	.w7(32'hbbce12f7),
	.w8(32'hbc3d81f7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bdf521),
	.w1(32'h3a5103b2),
	.w2(32'h39422e88),
	.w3(32'hbb7cc837),
	.w4(32'h3b8eba77),
	.w5(32'h3aab8afb),
	.w6(32'hbc0d7aef),
	.w7(32'h3c050460),
	.w8(32'h3ba4118b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0391d0),
	.w1(32'h3bcd53e8),
	.w2(32'h3bdc5e61),
	.w3(32'hb9cd05b8),
	.w4(32'h3aa212d2),
	.w5(32'hbac44eb7),
	.w6(32'hbb6afde2),
	.w7(32'h39cf9bf0),
	.w8(32'hba8f510a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74ba11),
	.w1(32'hbbaf7530),
	.w2(32'hbbc98a75),
	.w3(32'hba45c17f),
	.w4(32'hbbc7f856),
	.w5(32'hbbfc5ebd),
	.w6(32'h3a89ee4a),
	.w7(32'hbc03a07f),
	.w8(32'hbc66a275),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f6f6),
	.w1(32'h3bc446a9),
	.w2(32'h3b6b2cee),
	.w3(32'hbbcb6486),
	.w4(32'hbbdb59fc),
	.w5(32'hbb2d6d25),
	.w6(32'hbc1c4aaf),
	.w7(32'h3b2e5d84),
	.w8(32'h3b01fa36),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075ab5),
	.w1(32'hbb79f080),
	.w2(32'hbbde764f),
	.w3(32'h3ab5dba9),
	.w4(32'h3b5a563f),
	.w5(32'h3b8ec08b),
	.w6(32'h3c680f42),
	.w7(32'h3b1da453),
	.w8(32'hbb13808f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c7f5c),
	.w1(32'h3b9b5d2d),
	.w2(32'h3b500164),
	.w3(32'hb99e45a1),
	.w4(32'h3b2527c2),
	.w5(32'h3b923e6a),
	.w6(32'hbb5e2b88),
	.w7(32'h3adc4e40),
	.w8(32'h3b35bdda),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c6dea),
	.w1(32'h3b090fec),
	.w2(32'hb6e356cf),
	.w3(32'h3bb401b4),
	.w4(32'h3b203b0a),
	.w5(32'hba8e4985),
	.w6(32'h3b3b699c),
	.w7(32'h3b75dce2),
	.w8(32'h3b357d2d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90eae45),
	.w1(32'h3b3e8e53),
	.w2(32'h3b5b6d08),
	.w3(32'h3a2e6b1a),
	.w4(32'hbb131749),
	.w5(32'hbaba77a4),
	.w6(32'h3b930ca1),
	.w7(32'hbba366ab),
	.w8(32'hbbbf6ec6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31de95),
	.w1(32'hbbc49794),
	.w2(32'hb995f5df),
	.w3(32'h39e21cd6),
	.w4(32'hbbbdd1cc),
	.w5(32'hbbb24181),
	.w6(32'hbbbeedb6),
	.w7(32'hb9ee455b),
	.w8(32'hbaf52966),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace4dd),
	.w1(32'hb81d0a75),
	.w2(32'h3bb0ba20),
	.w3(32'h3b45ad3d),
	.w4(32'hbbbb1d80),
	.w5(32'h3ac95a04),
	.w6(32'hba03d72f),
	.w7(32'hbaf4b318),
	.w8(32'hbc59f044),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f8e7),
	.w1(32'h3bcb1e01),
	.w2(32'h3bb4ea7e),
	.w3(32'hbbb23537),
	.w4(32'hbb0d6fcd),
	.w5(32'hbab98f75),
	.w6(32'hbbf2bf0a),
	.w7(32'h3a40527f),
	.w8(32'hbb7cfb2d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcade7f),
	.w1(32'hbbe22799),
	.w2(32'hbb8ac14d),
	.w3(32'hbae3a680),
	.w4(32'hbbfbd2d4),
	.w5(32'hbbe50edf),
	.w6(32'hba9b2f77),
	.w7(32'hbc73149c),
	.w8(32'hbc7daf44),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ddef),
	.w1(32'h3c02bd80),
	.w2(32'h3c205800),
	.w3(32'hbbb80eac),
	.w4(32'h3c87be18),
	.w5(32'h3c25ddf1),
	.w6(32'hbc15f9ba),
	.w7(32'h3bf0b89b),
	.w8(32'hbb8eecfe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b941b0e),
	.w1(32'h3af31059),
	.w2(32'h3b69e5c2),
	.w3(32'h3bf792be),
	.w4(32'h3b0d5010),
	.w5(32'hb9600a12),
	.w6(32'hbbc55719),
	.w7(32'hbb824e5a),
	.w8(32'hba5f36b9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b8f11),
	.w1(32'hbc40e9da),
	.w2(32'hbc5c99df),
	.w3(32'h3bb2a0c4),
	.w4(32'hbb9058f6),
	.w5(32'hbbb9f4a1),
	.w6(32'h395d0ef2),
	.w7(32'hbbea84a5),
	.w8(32'hbc0b0645),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e430e),
	.w1(32'hbb24314f),
	.w2(32'h3a16eb71),
	.w3(32'hbba17b3e),
	.w4(32'h3b234a80),
	.w5(32'h3a9136a4),
	.w6(32'hbbfa9d0f),
	.w7(32'hb7afbe49),
	.w8(32'hba876af2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06d98d),
	.w1(32'hbbc81656),
	.w2(32'hbbc3675f),
	.w3(32'hbb1d6ace),
	.w4(32'hbbe9b085),
	.w5(32'h398cf502),
	.w6(32'hbb31abd9),
	.w7(32'hbc05c97a),
	.w8(32'hbb354c0e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079a4e),
	.w1(32'hbacb6e1c),
	.w2(32'hbaa88c43),
	.w3(32'h3ba91eff),
	.w4(32'hbae0b4f1),
	.w5(32'hbb199c96),
	.w6(32'hba9398a1),
	.w7(32'h3a83e9bd),
	.w8(32'hbbd54f9a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12d839),
	.w1(32'hba48442f),
	.w2(32'hba76b996),
	.w3(32'hbbed6c4b),
	.w4(32'hb7c826cd),
	.w5(32'hba902f66),
	.w6(32'hbbe81330),
	.w7(32'hbb6fad43),
	.w8(32'hbb07687c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24bc49),
	.w1(32'h3b16cfd5),
	.w2(32'hbb6a4a9b),
	.w3(32'h3ad3c952),
	.w4(32'h3a75c117),
	.w5(32'hbb2cb446),
	.w6(32'h3b905a5a),
	.w7(32'h3bb3356e),
	.w8(32'hbc053d95),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4172b),
	.w1(32'h3a85d72c),
	.w2(32'hbb1c0713),
	.w3(32'hbb59ab91),
	.w4(32'hbbe560ce),
	.w5(32'hbb512c7d),
	.w6(32'hba631d38),
	.w7(32'h3a48c5a3),
	.w8(32'hba2f4f4d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaa623),
	.w1(32'h3b538c20),
	.w2(32'h3bd63a16),
	.w3(32'hbb79bc51),
	.w4(32'h3c0ad5a3),
	.w5(32'h3c402461),
	.w6(32'h393c8904),
	.w7(32'h3c08f228),
	.w8(32'h3c08778e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d689f),
	.w1(32'h3b82e43c),
	.w2(32'h3c175aa7),
	.w3(32'h3b928946),
	.w4(32'h3b87f666),
	.w5(32'h3bad7512),
	.w6(32'h3bb2b4fb),
	.w7(32'hbbb86571),
	.w8(32'hbb28cde0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b1d4),
	.w1(32'hbae2173a),
	.w2(32'hbb91c773),
	.w3(32'h3b820bb7),
	.w4(32'hbb769a36),
	.w5(32'hbbab62fe),
	.w6(32'hbb50b2ea),
	.w7(32'hbbf5a1d2),
	.w8(32'hbb30e676),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb492cd9),
	.w1(32'hbad36dd4),
	.w2(32'hba0ef1fc),
	.w3(32'hbae5ff67),
	.w4(32'h3ab94b32),
	.w5(32'h383ccd6c),
	.w6(32'h3ae95857),
	.w7(32'h3a06937d),
	.w8(32'h3ae0c1e9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2eaa),
	.w1(32'hbb97cc65),
	.w2(32'hbb08ac76),
	.w3(32'hbafd6ca7),
	.w4(32'h3b15d249),
	.w5(32'h3a912ecf),
	.w6(32'hbb90d268),
	.w7(32'h3a9a069d),
	.w8(32'h3a8b915c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb816c38),
	.w1(32'h3a826fef),
	.w2(32'h3a8bae68),
	.w3(32'hbb9f665d),
	.w4(32'h3b701809),
	.w5(32'h3b618c6a),
	.w6(32'hbad82f1e),
	.w7(32'h3af00ee9),
	.w8(32'h3b75ec10),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e59278),
	.w1(32'hbbde5810),
	.w2(32'hbb87cee3),
	.w3(32'h3a961066),
	.w4(32'hbc4bc53c),
	.w5(32'hbbe1d8c3),
	.w6(32'h3b286e21),
	.w7(32'hbb9d3ceb),
	.w8(32'hbb90c11f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54ddcb),
	.w1(32'h3b17b64b),
	.w2(32'h3c283236),
	.w3(32'hbbaec584),
	.w4(32'h3b4e8279),
	.w5(32'h3bace0a7),
	.w6(32'h3a622528),
	.w7(32'h3b882214),
	.w8(32'h3bd34fd7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ce8f),
	.w1(32'h3acf5e0b),
	.w2(32'hbbb1efb3),
	.w3(32'h3c2d1442),
	.w4(32'h3ad2c3a3),
	.w5(32'hbb853d7f),
	.w6(32'h3bc1e2e3),
	.w7(32'h399fb285),
	.w8(32'hbc119b35),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91a041),
	.w1(32'h3b779b1f),
	.w2(32'h3bd30ffc),
	.w3(32'hbb2ef5b9),
	.w4(32'h3b5c30e1),
	.w5(32'h3b62142d),
	.w6(32'hbbab531c),
	.w7(32'h3b0be8fd),
	.w8(32'h3b8cb04e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958f3e),
	.w1(32'h3c49b6bd),
	.w2(32'h3b9a19dd),
	.w3(32'h3bedef4a),
	.w4(32'h3b10f1c2),
	.w5(32'h3b2b4a63),
	.w6(32'h3b5cf9dc),
	.w7(32'h3b7384f0),
	.w8(32'h3b927084),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc14ff5),
	.w1(32'hbb84c2e3),
	.w2(32'hbb8c192a),
	.w3(32'hbb409bb8),
	.w4(32'h3b5328af),
	.w5(32'h3a43e83c),
	.w6(32'hba05ee02),
	.w7(32'hbb8f87f1),
	.w8(32'hbb6974d0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1a82),
	.w1(32'h39dca524),
	.w2(32'h3af6cba6),
	.w3(32'h3b6887a6),
	.w4(32'h3a23841e),
	.w5(32'h3b486fc1),
	.w6(32'hbb18a801),
	.w7(32'hbb23182b),
	.w8(32'hbb7d42e0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf12df),
	.w1(32'h3ad27ee3),
	.w2(32'hb99c59a3),
	.w3(32'h3b0d8cd5),
	.w4(32'hbb931ae6),
	.w5(32'hbb42d4ad),
	.w6(32'hba8b38b5),
	.w7(32'h3b114162),
	.w8(32'h3a9f242f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af12bc9),
	.w1(32'h3bece86f),
	.w2(32'h3b9c0859),
	.w3(32'hbaae15dc),
	.w4(32'hbb7e5ae3),
	.w5(32'h37a0e2b8),
	.w6(32'h3b02467d),
	.w7(32'h3bb31edb),
	.w8(32'h3b9d3fd4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348eb7),
	.w1(32'hbadfb3f8),
	.w2(32'h3b50d83f),
	.w3(32'h3c0ac421),
	.w4(32'h3b168fd5),
	.w5(32'h3be0e24a),
	.w6(32'h3c314586),
	.w7(32'h3b3f0cc4),
	.w8(32'hbb023422),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2e3db),
	.w1(32'h3a003434),
	.w2(32'hbbb2e457),
	.w3(32'h3c13e0bf),
	.w4(32'hbb8e41ac),
	.w5(32'hbbeb3a77),
	.w6(32'hba47dc72),
	.w7(32'hbc00c9a6),
	.w8(32'hbbe129fb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dcc52),
	.w1(32'hbbba9cac),
	.w2(32'hbb17cd74),
	.w3(32'hbbaaeb0c),
	.w4(32'hbb028d46),
	.w5(32'hbb5532f5),
	.w6(32'hba249eff),
	.w7(32'hbb4e1855),
	.w8(32'hbb168d1e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd3db8),
	.w1(32'h3a609c74),
	.w2(32'h3b2ce29f),
	.w3(32'hbb7aceda),
	.w4(32'h3b0198f7),
	.w5(32'h3b3c5b23),
	.w6(32'hbb185697),
	.w7(32'h3b8c3e2e),
	.w8(32'h3b7c97be),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfdb04),
	.w1(32'h3c10f3c8),
	.w2(32'hbb4430b0),
	.w3(32'h3bb0b2b3),
	.w4(32'hbbba8af8),
	.w5(32'hbb82c4e0),
	.w6(32'h3c1a9912),
	.w7(32'hbb5dac32),
	.w8(32'hbc81350c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32831b),
	.w1(32'h3b95b406),
	.w2(32'h3aae2738),
	.w3(32'hbbc17187),
	.w4(32'h3a060e98),
	.w5(32'hbbc92875),
	.w6(32'hbaebc9d4),
	.w7(32'hba2d9bee),
	.w8(32'hbbe0244f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3871a),
	.w1(32'hbb6873d9),
	.w2(32'hbb11d544),
	.w3(32'hbb2f9e67),
	.w4(32'hbb1a3ac9),
	.w5(32'hb9b49e16),
	.w6(32'hbc134172),
	.w7(32'hbb4bfd42),
	.w8(32'hba8aa649),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21899),
	.w1(32'hba667212),
	.w2(32'h3af4d414),
	.w3(32'hb8b69c81),
	.w4(32'hbb2b5784),
	.w5(32'h3b3b40d4),
	.w6(32'h397fca35),
	.w7(32'h395d4b05),
	.w8(32'hbb072a61),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9a56f),
	.w1(32'hbbea64ec),
	.w2(32'hbb381390),
	.w3(32'hbb887ced),
	.w4(32'hbc16da48),
	.w5(32'hbad6063e),
	.w6(32'hb9d840bf),
	.w7(32'hbbeb2b4b),
	.w8(32'hbadd7b24),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291394),
	.w1(32'h3c13fe58),
	.w2(32'h3c6f91d1),
	.w3(32'hbbc90d57),
	.w4(32'hbaf80bd9),
	.w5(32'h3be17497),
	.w6(32'hbad60200),
	.w7(32'h3ca9502c),
	.w8(32'h3ca3bf77),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e6aaf),
	.w1(32'hbbfaaeff),
	.w2(32'hbbddfb2c),
	.w3(32'h3c41ed66),
	.w4(32'hbc84faef),
	.w5(32'hbcaed69f),
	.w6(32'h3cea817e),
	.w7(32'hbc8cad07),
	.w8(32'hbc9081ad),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9a140),
	.w1(32'hba9e3ef1),
	.w2(32'hbab1f3d7),
	.w3(32'hbc7ec73c),
	.w4(32'hbb970b21),
	.w5(32'hbb5df505),
	.w6(32'hbccd2c87),
	.w7(32'hbb12c04a),
	.w8(32'h3a6bd597),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c9aec),
	.w1(32'hb8e07bb5),
	.w2(32'hbb411a10),
	.w3(32'hb98d8bf5),
	.w4(32'h3b585773),
	.w5(32'hbb1bd163),
	.w6(32'h3b9969aa),
	.w7(32'h3c004bc0),
	.w8(32'h39891ccd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90cd85),
	.w1(32'hbb59b749),
	.w2(32'h3b292f92),
	.w3(32'hbac10ae9),
	.w4(32'hbb241b51),
	.w5(32'hbaf23b71),
	.w6(32'hba639458),
	.w7(32'hbbb1d9dc),
	.w8(32'hbb7aa272),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a2feb),
	.w1(32'hb9f98a71),
	.w2(32'hba78fb22),
	.w3(32'hbb087543),
	.w4(32'hbb0b5411),
	.w5(32'h39c38b9b),
	.w6(32'hbb73e9ef),
	.w7(32'h3a5e864c),
	.w8(32'hbbbc0826),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb502525),
	.w1(32'hbc42ec54),
	.w2(32'hbc130521),
	.w3(32'hbb367651),
	.w4(32'hbc2cb501),
	.w5(32'hbc6e4e41),
	.w6(32'hbbec04ed),
	.w7(32'hbc926fda),
	.w8(32'hbc8a8295),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39f44d),
	.w1(32'hbb15cd05),
	.w2(32'hbbb7a22c),
	.w3(32'hbc51e0b0),
	.w4(32'hbbba3490),
	.w5(32'hbb87b31b),
	.w6(32'hbc860c33),
	.w7(32'hb97721c6),
	.w8(32'hb8d5d79c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2789),
	.w1(32'hbbb89244),
	.w2(32'hbbe68fa3),
	.w3(32'hbbaf971d),
	.w4(32'hb9d6933a),
	.w5(32'hba9b1a84),
	.w6(32'h3aa334e8),
	.w7(32'h3ae1abc3),
	.w8(32'h3af728d1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd5684),
	.w1(32'h3ab6955d),
	.w2(32'h3bade4b5),
	.w3(32'hbb10975e),
	.w4(32'h394b1803),
	.w5(32'hba6342f8),
	.w6(32'h3aa13d45),
	.w7(32'h3b7e0f9a),
	.w8(32'h3bbf23ad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44057c),
	.w1(32'hbb467a85),
	.w2(32'hbb0cb7cf),
	.w3(32'hb99fdace),
	.w4(32'hba16401e),
	.w5(32'hbb472e7f),
	.w6(32'h3a5abf42),
	.w7(32'hbb50c50b),
	.w8(32'hbb22a961),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb549367),
	.w1(32'h3c0d622f),
	.w2(32'h3bc32ede),
	.w3(32'h39c9f108),
	.w4(32'h3c1eaf04),
	.w5(32'h3c10822d),
	.w6(32'hba1de4b9),
	.w7(32'h3c1b9a84),
	.w8(32'h3c12a15e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40fb29),
	.w1(32'hba697b56),
	.w2(32'h3b83773e),
	.w3(32'h3be54d74),
	.w4(32'hbb3a00d8),
	.w5(32'hbb849b8e),
	.w6(32'h3b80ae9b),
	.w7(32'h3a807439),
	.w8(32'hbb70cf44),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58849d),
	.w1(32'hbaf606b6),
	.w2(32'hbaece126),
	.w3(32'h3b3c3078),
	.w4(32'hbac82265),
	.w5(32'hbaae1504),
	.w6(32'hbb8abae7),
	.w7(32'hbb746d61),
	.w8(32'hbae40eae),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa058b),
	.w1(32'h3ae35aab),
	.w2(32'h3b642227),
	.w3(32'hbb1a394b),
	.w4(32'hba2a17ac),
	.w5(32'hb93c8ef4),
	.w6(32'h3a97eb94),
	.w7(32'h3910bd39),
	.w8(32'hbb26dd76),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b200988),
	.w1(32'hbb1283dd),
	.w2(32'h3acd06a6),
	.w3(32'h3b180ee1),
	.w4(32'hbaf48898),
	.w5(32'hbb512e01),
	.w6(32'hbb5ff710),
	.w7(32'hbc26d1cd),
	.w8(32'hb93214e5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af8e81),
	.w1(32'hba2c6706),
	.w2(32'hb9d6f78b),
	.w3(32'hb84ddff6),
	.w4(32'h3b8b7247),
	.w5(32'h3c0bfd89),
	.w6(32'h3b0c8f7a),
	.w7(32'h3c318d11),
	.w8(32'h3c288933),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bf7d9),
	.w1(32'hbb53e9b0),
	.w2(32'hbb8d1889),
	.w3(32'h3c2141f2),
	.w4(32'hbaebab19),
	.w5(32'h3b88a405),
	.w6(32'h3c652096),
	.w7(32'hbb053c70),
	.w8(32'h3bba84c8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d4cc1),
	.w1(32'h3b9b27fd),
	.w2(32'h3c305aef),
	.w3(32'h3b429e8b),
	.w4(32'hba775381),
	.w5(32'h3be891be),
	.w6(32'hbaac921a),
	.w7(32'hbbb48e83),
	.w8(32'hbb200bcc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b717fef),
	.w1(32'h3b35cfea),
	.w2(32'h3bec58c9),
	.w3(32'hba8f9937),
	.w4(32'h3b0e1d49),
	.w5(32'h3b1b151c),
	.w6(32'hbb970d4a),
	.w7(32'h3b3cded7),
	.w8(32'h3b1e2844),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6993),
	.w1(32'h3b8ba3f3),
	.w2(32'h3b38318f),
	.w3(32'hbad5a3e4),
	.w4(32'h3b131c84),
	.w5(32'h3b1d42ef),
	.w6(32'hb9ede40c),
	.w7(32'h3a68a8e3),
	.w8(32'h3ab559b0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd0a4),
	.w1(32'h3b3377f4),
	.w2(32'h3bc76a21),
	.w3(32'h3af2851d),
	.w4(32'h3bd34834),
	.w5(32'hbae8cd7e),
	.w6(32'h3b99d68b),
	.w7(32'hbb070034),
	.w8(32'hba87cb44),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac36fdb),
	.w1(32'hbb23204e),
	.w2(32'h3a12a5b4),
	.w3(32'hba8444b2),
	.w4(32'hbba71ea5),
	.w5(32'hb9ca8d53),
	.w6(32'h38194ee4),
	.w7(32'hbb46547b),
	.w8(32'hba6e664f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a325d2a),
	.w1(32'h3b0129d1),
	.w2(32'h3bd7530f),
	.w3(32'h3afb3955),
	.w4(32'h39e30f1d),
	.w5(32'hba162e26),
	.w6(32'h3a577377),
	.w7(32'hbbcb2ee0),
	.w8(32'hbae601d7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd344a8),
	.w1(32'hbc2fb5cf),
	.w2(32'hbc17e661),
	.w3(32'h3a705381),
	.w4(32'hbc80ba18),
	.w5(32'hbc451783),
	.w6(32'hbb99c628),
	.w7(32'hbc77b861),
	.w8(32'hbc856bcd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb47fd),
	.w1(32'h3bc1c498),
	.w2(32'h3bfac5ba),
	.w3(32'hbc1eb6d5),
	.w4(32'h3b175e6a),
	.w5(32'hbaa28c73),
	.w6(32'hbc38060d),
	.w7(32'hbacb56c5),
	.w8(32'hbab8ada2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f3275),
	.w1(32'h3995dda8),
	.w2(32'h3b793441),
	.w3(32'hba37381a),
	.w4(32'hbab9a2a8),
	.w5(32'h3bb6c1ae),
	.w6(32'hbb2ee5a7),
	.w7(32'hbb366074),
	.w8(32'h3b7c5728),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa24a39),
	.w1(32'hbb9c849f),
	.w2(32'h3c006656),
	.w3(32'h3bc7990a),
	.w4(32'h3c067ef4),
	.w5(32'h3bf62fe9),
	.w6(32'h3b65f35b),
	.w7(32'hbb82a78f),
	.w8(32'h374d01a7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f448),
	.w1(32'hbac1b369),
	.w2(32'h3ae4aa49),
	.w3(32'h3c07988a),
	.w4(32'hbb1c5c75),
	.w5(32'hbac8f77a),
	.w6(32'hbbd1b351),
	.w7(32'hbabcff79),
	.w8(32'h3b75deb2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76bdb2),
	.w1(32'hbb193c79),
	.w2(32'hbc03b23e),
	.w3(32'hb965e282),
	.w4(32'hbadf7ac4),
	.w5(32'hbc29b592),
	.w6(32'hbad8fe0d),
	.w7(32'h3bb467a6),
	.w8(32'hbacc07e4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a5f9),
	.w1(32'hbc0d76c8),
	.w2(32'hbc05b55d),
	.w3(32'hbc72eb24),
	.w4(32'hbb9e9a27),
	.w5(32'hbbe2046d),
	.w6(32'hbc60b8dd),
	.w7(32'hbb39e5aa),
	.w8(32'hbb5f1951),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46107),
	.w1(32'hbbde3655),
	.w2(32'hbb61725f),
	.w3(32'hbb049530),
	.w4(32'hbb74d3e4),
	.w5(32'hbb2562cb),
	.w6(32'hbae366da),
	.w7(32'hbb81a7dd),
	.w8(32'hbbe4025f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61032f),
	.w1(32'h3b0177c7),
	.w2(32'h3bdead56),
	.w3(32'hbb47c5cc),
	.w4(32'h3af16f83),
	.w5(32'h3b49a6d1),
	.w6(32'hbb1de62a),
	.w7(32'h3a45aad0),
	.w8(32'h3ad4a5b5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d73d6f),
	.w1(32'h3b980851),
	.w2(32'h3c15f5b2),
	.w3(32'h3b171317),
	.w4(32'hbc35c6cd),
	.w5(32'hbc3fbbda),
	.w6(32'h3b2f93e2),
	.w7(32'hbc5c9fcd),
	.w8(32'hbcb59746),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8c95),
	.w1(32'hbb2bd4b8),
	.w2(32'hbb623acf),
	.w3(32'hbc8156fa),
	.w4(32'hbaf9e83a),
	.w5(32'hbb7e19fb),
	.w6(32'hbca25ce2),
	.w7(32'hbb8bee14),
	.w8(32'hbbda857b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da1e8b),
	.w1(32'h3a85b429),
	.w2(32'h3a491b7c),
	.w3(32'hbb4cc83a),
	.w4(32'hbac1207c),
	.w5(32'hbb8b2bcd),
	.w6(32'hbb93b5ee),
	.w7(32'hbb1362f4),
	.w8(32'hbc159277),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c78bc2),
	.w1(32'hbb8835c1),
	.w2(32'hbb08c451),
	.w3(32'hbb0ebcc9),
	.w4(32'hbab980aa),
	.w5(32'hbab4f0b1),
	.w6(32'hbc5584fd),
	.w7(32'hbacc39c0),
	.w8(32'hba587c52),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1a068),
	.w1(32'h3b9bd218),
	.w2(32'h3b6407cd),
	.w3(32'hba1367f9),
	.w4(32'h3af68631),
	.w5(32'h3accab76),
	.w6(32'hbaf9883f),
	.w7(32'h3b6e5c02),
	.w8(32'h3abc0d40),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49b88a),
	.w1(32'hbb6396c2),
	.w2(32'hbb8eee9a),
	.w3(32'h3aa28db9),
	.w4(32'h3ad78ef9),
	.w5(32'hba72b95d),
	.w6(32'h3b579367),
	.w7(32'h3bd4bac7),
	.w8(32'h3af6786e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc969),
	.w1(32'hbb8b148c),
	.w2(32'hbbaf0232),
	.w3(32'hbafd4673),
	.w4(32'hbbfd64f6),
	.w5(32'hbbda25c8),
	.w6(32'h3b333837),
	.w7(32'hbc05e242),
	.w8(32'hbc15c202),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf05a),
	.w1(32'hbb955ec6),
	.w2(32'h3aae9f85),
	.w3(32'hbc050f46),
	.w4(32'h39ba2521),
	.w5(32'hbb2fb2d8),
	.w6(32'hbbd4e38f),
	.w7(32'hbade9104),
	.w8(32'hbb27e75b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84235a),
	.w1(32'h3a2b3480),
	.w2(32'h3b4dc26d),
	.w3(32'h3aefa513),
	.w4(32'h3a40a018),
	.w5(32'h3b4c77bd),
	.w6(32'h3a9a9b24),
	.w7(32'h393e1f22),
	.w8(32'h3ba7d0d1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbe686),
	.w1(32'h3a956e54),
	.w2(32'h3c060116),
	.w3(32'h3a6189e0),
	.w4(32'h3b8ae501),
	.w5(32'h3c087d22),
	.w6(32'h38c1724e),
	.w7(32'h3c0a0a95),
	.w8(32'h3b061e05),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14c727),
	.w1(32'h3b3c390e),
	.w2(32'h3b24ed0e),
	.w3(32'h3b84c4e7),
	.w4(32'h3aba6f52),
	.w5(32'hbb886028),
	.w6(32'hbb93512c),
	.w7(32'h38aeca48),
	.w8(32'h399db5f9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99b097),
	.w1(32'hbbda15ec),
	.w2(32'hbba1c4a7),
	.w3(32'hbb78b20e),
	.w4(32'hbbb5b8f1),
	.w5(32'h3b02ac4e),
	.w6(32'hba328174),
	.w7(32'h3b130ad3),
	.w8(32'h3b56a205),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77a2ba),
	.w1(32'h3b9fd785),
	.w2(32'h3c606c94),
	.w3(32'hb9cc1916),
	.w4(32'h3c13627d),
	.w5(32'h3c7956a2),
	.w6(32'h3a0974c3),
	.w7(32'hba18a535),
	.w8(32'h3b2de57f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9661),
	.w1(32'h3bf68927),
	.w2(32'h3c554923),
	.w3(32'h3c4425f2),
	.w4(32'h3c87f9ab),
	.w5(32'h3c8a9995),
	.w6(32'h3ac08319),
	.w7(32'h3bafdb50),
	.w8(32'h3b6c5339),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07f007),
	.w1(32'hbb2cbacc),
	.w2(32'hba647469),
	.w3(32'h3c210ead),
	.w4(32'hb98d6262),
	.w5(32'hbb34a848),
	.w6(32'h3b979119),
	.w7(32'h3ad1ad8d),
	.w8(32'hbab9b329),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d3c58),
	.w1(32'h3c4c9454),
	.w2(32'h3c94401e),
	.w3(32'hbb9a318e),
	.w4(32'h3c909d5e),
	.w5(32'h3c83e7ab),
	.w6(32'hba8e141c),
	.w7(32'h3c41e035),
	.w8(32'h3c6108c0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fd205),
	.w1(32'hbb395817),
	.w2(32'hbb44a673),
	.w3(32'h3c924035),
	.w4(32'hbba4789d),
	.w5(32'hbb362744),
	.w6(32'h3c83b687),
	.w7(32'hbb917f0d),
	.w8(32'hb83e6197),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9be47d),
	.w1(32'hbb39c168),
	.w2(32'h39874201),
	.w3(32'hb981c2d7),
	.w4(32'hbbaf9653),
	.w5(32'h3b84d51a),
	.w6(32'h3a8b319a),
	.w7(32'hbb85f1c8),
	.w8(32'hbb3ab885),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecf14),
	.w1(32'h3ba23c3d),
	.w2(32'h3a88c16b),
	.w3(32'h3ac61ae1),
	.w4(32'hbae25eb8),
	.w5(32'hba25638d),
	.w6(32'h3b7dbdd2),
	.w7(32'hbbd4fd19),
	.w8(32'hbbda86a0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c063169),
	.w1(32'h3ae22997),
	.w2(32'h3b77d3ef),
	.w3(32'h3bef9922),
	.w4(32'h3a7f64e2),
	.w5(32'h3b0eb993),
	.w6(32'h3a145cab),
	.w7(32'h3b71ba1b),
	.w8(32'h3b03a326),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64abf2),
	.w1(32'h3bab1254),
	.w2(32'h3c702203),
	.w3(32'h3ac3887d),
	.w4(32'h38b47244),
	.w5(32'h3b16c921),
	.w6(32'hbb651e35),
	.w7(32'hbb8a726d),
	.w8(32'h38dd1ed8),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3de428),
	.w1(32'h3bc7ba9d),
	.w2(32'h3b99423f),
	.w3(32'h3bd30e1d),
	.w4(32'h3b83d95b),
	.w5(32'h3b65da5f),
	.w6(32'h3b27b446),
	.w7(32'h3b283aa4),
	.w8(32'h3b1189b5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c1882),
	.w1(32'hbbacc8de),
	.w2(32'hbb48f200),
	.w3(32'hba903f2b),
	.w4(32'h3ade66a5),
	.w5(32'hbba6b46a),
	.w6(32'h3aa82b35),
	.w7(32'hba36a69c),
	.w8(32'hbc13e2f0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b919472),
	.w1(32'hbb0d4a94),
	.w2(32'hbaf6c8b9),
	.w3(32'h3b240eca),
	.w4(32'hbb474c28),
	.w5(32'hbb6310c1),
	.w6(32'hbb47d4ff),
	.w7(32'hbb816e5a),
	.w8(32'hbacfe332),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4f67),
	.w1(32'h3b4a53d7),
	.w2(32'h3bffd17c),
	.w3(32'h3ac1ae0b),
	.w4(32'hb92243b0),
	.w5(32'h3be02a8b),
	.w6(32'hbb3293dd),
	.w7(32'hbb23851a),
	.w8(32'h3b205736),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf3347),
	.w1(32'hbb7eb079),
	.w2(32'hbb91c5b8),
	.w3(32'h3bca0ece),
	.w4(32'hbba3e388),
	.w5(32'hbb061be5),
	.w6(32'h399e1960),
	.w7(32'hbc73141b),
	.w8(32'hbc3343e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0643f3),
	.w1(32'hbb842f15),
	.w2(32'hbb06c9d7),
	.w3(32'hbb979335),
	.w4(32'hbb132ba3),
	.w5(32'hbb9440f9),
	.w6(32'hbc0ca038),
	.w7(32'hba8c1a99),
	.w8(32'hbbbf0f0c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab6fc6),
	.w1(32'hbb677883),
	.w2(32'h3bb6e678),
	.w3(32'hbbbf1420),
	.w4(32'h3bda7ef7),
	.w5(32'h3a087f5e),
	.w6(32'hbbb7b5c0),
	.w7(32'h3bd43b62),
	.w8(32'h3b975f11),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b33a),
	.w1(32'hbb673248),
	.w2(32'hbac15ead),
	.w3(32'hbb48d7f3),
	.w4(32'h3b6de654),
	.w5(32'hbb8259a3),
	.w6(32'hbb63081a),
	.w7(32'h3c014cb5),
	.w8(32'h3ba85bf7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ae31),
	.w1(32'h395970e2),
	.w2(32'hb8247672),
	.w3(32'h3b96ac51),
	.w4(32'h3935ea1f),
	.w5(32'hb90d7d49),
	.w6(32'h3bd660b9),
	.w7(32'h39ae835a),
	.w8(32'hb8f89f80),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c07e7),
	.w1(32'h3793a240),
	.w2(32'h388c0521),
	.w3(32'h3790e50c),
	.w4(32'h3909b918),
	.w5(32'h3939df5f),
	.w6(32'hb7f92d9e),
	.w7(32'h38193084),
	.w8(32'h383fd0cc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6430917),
	.w1(32'h36c7a077),
	.w2(32'h37506010),
	.w3(32'h3548d063),
	.w4(32'h37480800),
	.w5(32'h376a36d3),
	.w6(32'hb6dffe15),
	.w7(32'h350a46cf),
	.w8(32'h36d3a135),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370879a0),
	.w1(32'hb899804f),
	.w2(32'hb7f74da5),
	.w3(32'hb5f2465f),
	.w4(32'hb876c02e),
	.w5(32'hb8241634),
	.w6(32'hb792e800),
	.w7(32'hb87516f1),
	.w8(32'hb835b24d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3703acb5),
	.w1(32'hb6893149),
	.w2(32'h3764f97f),
	.w3(32'h3766ab22),
	.w4(32'hb6055ea2),
	.w5(32'h37a36512),
	.w6(32'hb63b1384),
	.w7(32'hb751e275),
	.w8(32'h3688caa2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b6f7d),
	.w1(32'h38707f13),
	.w2(32'hb7fc35b1),
	.w3(32'h389e2a86),
	.w4(32'h38a0088f),
	.w5(32'hb7a0239b),
	.w6(32'h38ff2392),
	.w7(32'h391e5628),
	.w8(32'h38711db3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38772992),
	.w1(32'h387d9d43),
	.w2(32'hb836b6af),
	.w3(32'hb8f3459f),
	.w4(32'hb835ff98),
	.w5(32'hb9122b2d),
	.w6(32'h382c1e83),
	.w7(32'h38a4028b),
	.w8(32'hb8495daa),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9065369),
	.w1(32'hb8064f3d),
	.w2(32'hb902b189),
	.w3(32'hb93ce2e0),
	.w4(32'hb88a9fe1),
	.w5(32'hb9087056),
	.w6(32'h371fde4f),
	.w7(32'h38748f58),
	.w8(32'hb8829952),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8286eb6),
	.w1(32'hb8be1a8a),
	.w2(32'hb93496dc),
	.w3(32'hb7f8e001),
	.w4(32'hb878e8ba),
	.w5(32'hb91d5bce),
	.w6(32'hb7a9da68),
	.w7(32'hb80c7e06),
	.w8(32'hb8d634d4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9548046),
	.w1(32'hb8e4555c),
	.w2(32'hb817023e),
	.w3(32'hb983c10d),
	.w4(32'hb96dbb54),
	.w5(32'hb92227fa),
	.w6(32'hb9228c51),
	.w7(32'hb90150c9),
	.w8(32'hb8c1efcf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8a848),
	.w1(32'h399a5b87),
	.w2(32'hb88a0393),
	.w3(32'h39989168),
	.w4(32'h38fc593b),
	.w5(32'hb9930db4),
	.w6(32'h39c13ea0),
	.w7(32'h398959b4),
	.w8(32'hb85a6cf6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdcf26),
	.w1(32'hb9968508),
	.w2(32'hb976270f),
	.w3(32'hb9991c00),
	.w4(32'hb93f2984),
	.w5(32'hb984c1b0),
	.w6(32'hb96b975b),
	.w7(32'hb8e32b64),
	.w8(32'hb93b43bb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36827141),
	.w1(32'hb6649edd),
	.w2(32'h37048800),
	.w3(32'h3710dd25),
	.w4(32'h35cc224c),
	.w5(32'h3746ff0e),
	.w6(32'h35ef80ea),
	.w7(32'hb6924b4b),
	.w8(32'h3643ced4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34a85423),
	.w1(32'h36392475),
	.w2(32'h368faab9),
	.w3(32'hb5e188ce),
	.w4(32'hb6b13962),
	.w5(32'hb6bb943c),
	.w6(32'h3680a696),
	.w7(32'hb594d233),
	.w8(32'hb66f49c7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7171731),
	.w1(32'h381f4f45),
	.w2(32'hb9534cac),
	.w3(32'hb7e971cc),
	.w4(32'h384d3792),
	.w5(32'hb94c6c35),
	.w6(32'h38765141),
	.w7(32'h3933e6ae),
	.w8(32'hb7d364ff),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fbddc5),
	.w1(32'hb8d38d55),
	.w2(32'hb9885c4b),
	.w3(32'hb966e6ee),
	.w4(32'hb8d69706),
	.w5(32'hb9b47049),
	.w6(32'h3780af5e),
	.w7(32'h36f52b28),
	.w8(32'hb9251aea),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85c6e26),
	.w1(32'hb916f1dd),
	.w2(32'hb9cfa451),
	.w3(32'hb7f82678),
	.w4(32'hb887f1e0),
	.w5(32'hb9d6c525),
	.w6(32'h38d2b7da),
	.w7(32'h389d7362),
	.w8(32'hb98863f1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed027c),
	.w1(32'h37c9e1de),
	.w2(32'hb89fe2fc),
	.w3(32'h388db891),
	.w4(32'hb8901dea),
	.w5(32'hb98481cb),
	.w6(32'h383fa142),
	.w7(32'hb8606fe2),
	.w8(32'hb93cb5ef),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3764faf0),
	.w1(32'hb74ed12e),
	.w2(32'hb79dbfd4),
	.w3(32'h36b661bb),
	.w4(32'hb77566d1),
	.w5(32'hb79e77a9),
	.w6(32'hb44a043f),
	.w7(32'hb797ab3a),
	.w8(32'hb7a1ba9c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cd05a9),
	.w1(32'hb83c1581),
	.w2(32'hb820a7fb),
	.w3(32'hb74bec75),
	.w4(32'hb824127a),
	.w5(32'hb80a144d),
	.w6(32'hb886606b),
	.w7(32'hb79142c5),
	.w8(32'hb76956ac),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cdcea),
	.w1(32'h395790d8),
	.w2(32'h391f84aa),
	.w3(32'h3900aaf3),
	.w4(32'h399ed3e6),
	.w5(32'h38ff2993),
	.w6(32'h35b10e1f),
	.w7(32'h392791d1),
	.w8(32'h39249aca),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0ef23),
	.w1(32'hb89526a6),
	.w2(32'hb96c4df0),
	.w3(32'h397d60fd),
	.w4(32'h389d424b),
	.w5(32'hb8d1f8aa),
	.w6(32'h39215eba),
	.w7(32'h38f0f8b1),
	.w8(32'hb8723db8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904675f),
	.w1(32'hb83d0765),
	.w2(32'hb8f04d93),
	.w3(32'h38852770),
	.w4(32'h3767e6c2),
	.w5(32'hb8e19c72),
	.w6(32'h380036cb),
	.w7(32'h37dc6ac1),
	.w8(32'hb5a0e78b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e67911),
	.w1(32'h379cb2d6),
	.w2(32'hb819115d),
	.w3(32'hb8e7386f),
	.w4(32'h384486a5),
	.w5(32'h37627afe),
	.w6(32'hb7d50182),
	.w7(32'h386157ff),
	.w8(32'h36ada6af),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ea379f),
	.w1(32'hb84de04a),
	.w2(32'hb906937c),
	.w3(32'hb8b2660b),
	.w4(32'hb93bca53),
	.w5(32'hb984862d),
	.w6(32'h383e037d),
	.w7(32'hb862a2e0),
	.w8(32'hb941ac91),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb600b3c3),
	.w1(32'h369e7ea2),
	.w2(32'h373bb4e6),
	.w3(32'h3646d2f5),
	.w4(32'h36fcd03d),
	.w5(32'h3735f5b4),
	.w6(32'hb5f7d24f),
	.w7(32'h36894fdd),
	.w8(32'h36be9343),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b235a0),
	.w1(32'hb511b8fc),
	.w2(32'hb350c8db),
	.w3(32'h35d30bc7),
	.w4(32'hb62efd62),
	.w5(32'h364577df),
	.w6(32'hb60fcd4d),
	.w7(32'hb63026cb),
	.w8(32'h34d27892),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376417f0),
	.w1(32'h34e31520),
	.w2(32'hb6c433f3),
	.w3(32'h37e68a51),
	.w4(32'hb67f3cac),
	.w5(32'hb789f2e8),
	.w6(32'h3704574a),
	.w7(32'hb63b4aa7),
	.w8(32'hb6900325),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351c9dee),
	.w1(32'h34a1062d),
	.w2(32'h373d2c23),
	.w3(32'h33d6febf),
	.w4(32'h36dc72e3),
	.w5(32'h37453b2e),
	.w6(32'h3636faa9),
	.w7(32'h34a2429f),
	.w8(32'h365f6549),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381562b4),
	.w1(32'h37feab07),
	.w2(32'hb81c72f6),
	.w3(32'h38109f13),
	.w4(32'h37ecd39f),
	.w5(32'hb7d39c18),
	.w6(32'h37c81a39),
	.w7(32'h36b1193e),
	.w8(32'hb7bad361),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4f460),
	.w1(32'hb9834bb7),
	.w2(32'hba0605ab),
	.w3(32'hb987f34e),
	.w4(32'hb9a43fae),
	.w5(32'hb9fc9dea),
	.w6(32'h3743264c),
	.w7(32'hb8f89b0c),
	.w8(32'hb98afd34),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c5dcb7),
	.w1(32'hb8a180e0),
	.w2(32'hb921bf08),
	.w3(32'hb8a07817),
	.w4(32'hb8d3184a),
	.w5(32'hb9309eb6),
	.w6(32'hb759f074),
	.w7(32'hb88eaa1a),
	.w8(32'hb8e93e4b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1ffe8),
	.w1(32'hb6a0d008),
	.w2(32'h368c1cbd),
	.w3(32'hb77e67c6),
	.w4(32'hb64aeab4),
	.w5(32'hb35fc511),
	.w6(32'hb75365ce),
	.w7(32'hb75c5475),
	.w8(32'hb6f40a4b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e30fd7),
	.w1(32'hb955e7c9),
	.w2(32'hb9bc7941),
	.w3(32'hb84faacc),
	.w4(32'hb914b914),
	.w5(32'hb9d777f6),
	.w6(32'h38727181),
	.w7(32'hb7a2abc3),
	.w8(32'hb92bd7a9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6a3bf),
	.w1(32'h37bc709e),
	.w2(32'hb880e324),
	.w3(32'h3867bc67),
	.w4(32'hb760d0a2),
	.w5(32'hb90042cd),
	.w6(32'h3819713c),
	.w7(32'h37ddefed),
	.w8(32'hb8b06c89),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb44d9cb6),
	.w1(32'hb63e1d8d),
	.w2(32'h34fb2211),
	.w3(32'h35aee20e),
	.w4(32'hb56e2f7a),
	.w5(32'hb58445c9),
	.w6(32'hb68c71cd),
	.w7(32'hb69532df),
	.w8(32'hb59743f1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3df7b),
	.w1(32'hb700dfe2),
	.w2(32'hb8e9532f),
	.w3(32'hb83052c6),
	.w4(32'h37d7dd07),
	.w5(32'hb8d8558e),
	.w6(32'h3755d5c0),
	.w7(32'h38a9005a),
	.w8(32'hb88a2dad),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3239f),
	.w1(32'h38ea3399),
	.w2(32'h38e05ef2),
	.w3(32'h38036a2f),
	.w4(32'h382c94af),
	.w5(32'h38636dec),
	.w6(32'h38267d27),
	.w7(32'h3868b1e4),
	.w8(32'h389584ce),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916ea0e),
	.w1(32'hb8d36406),
	.w2(32'hb8ad192b),
	.w3(32'hb9278113),
	.w4(32'hb900c0f2),
	.w5(32'hb8fa53e8),
	.w6(32'hb8d94ae2),
	.w7(32'hb8e113d1),
	.w8(32'hb8cc834b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354dbe1a),
	.w1(32'h36324938),
	.w2(32'hb5ef2cd8),
	.w3(32'hb5bf800a),
	.w4(32'hb63ee51a),
	.w5(32'hb6b519aa),
	.w6(32'hb65c8fee),
	.w7(32'hb69461bf),
	.w8(32'hb684b02b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7087ed4),
	.w1(32'hb6e9ceae),
	.w2(32'h370bddd9),
	.w3(32'hb660cfde),
	.w4(32'hb5f022ad),
	.w5(32'h36f8f169),
	.w6(32'h3510a948),
	.w7(32'h33ada8d8),
	.w8(32'h36cdfc74),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793e7f7),
	.w1(32'h387e614f),
	.w2(32'hb8350cc2),
	.w3(32'hb84d87ec),
	.w4(32'h379c5f86),
	.w5(32'hb8560e63),
	.w6(32'h3618d0cb),
	.w7(32'h3821e7d2),
	.w8(32'hb756bf52),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92986f9),
	.w1(32'hb92fa75d),
	.w2(32'hb9a68d83),
	.w3(32'hb869695a),
	.w4(32'hb94c2eb0),
	.w5(32'hb9e38115),
	.w6(32'h37dc4ae5),
	.w7(32'hb8df2215),
	.w8(32'hb9a2a147),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd18ad),
	.w1(32'hb7aa7ded),
	.w2(32'hb940336b),
	.w3(32'h37d1ee68),
	.w4(32'hb7e85ed5),
	.w5(32'hb95667c3),
	.w6(32'h38ee5ea5),
	.w7(32'h388996f2),
	.w8(32'hb92ab02b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a16deb),
	.w1(32'hb971165d),
	.w2(32'hb9a84ede),
	.w3(32'hb93de315),
	.w4(32'hb93803de),
	.w5(32'hb9c7c690),
	.w6(32'hb9258754),
	.w7(32'hb8edc714),
	.w8(32'hb98e68f7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca589d),
	.w1(32'h3770fec6),
	.w2(32'h36167009),
	.w3(32'hb65512cd),
	.w4(32'h380f6390),
	.w5(32'h37effffc),
	.w6(32'hb754172a),
	.w7(32'h37bb8e78),
	.w8(32'h371df4c0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67e94b6),
	.w1(32'hb75db334),
	.w2(32'hb779a362),
	.w3(32'hb60d581b),
	.w4(32'hb700160e),
	.w5(32'hb73ffae6),
	.w6(32'hb61241f6),
	.w7(32'hb603040a),
	.w8(32'hb6e233cb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5874e98),
	.w1(32'hb796443e),
	.w2(32'hb7b91bc9),
	.w3(32'h36634e67),
	.w4(32'hb78f9630),
	.w5(32'hb7b69ac9),
	.w6(32'h35665270),
	.w7(32'hb6610e75),
	.w8(32'hb7be19e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361132fd),
	.w1(32'h327a49a3),
	.w2(32'h363d7f28),
	.w3(32'h3650350c),
	.w4(32'h366df75f),
	.w5(32'h35ac8dba),
	.w6(32'h3596029e),
	.w7(32'hb63ce48b),
	.w8(32'hb6801df4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccf594),
	.w1(32'hb8f10174),
	.w2(32'hb960262e),
	.w3(32'h38c968ca),
	.w4(32'hb9126800),
	.w5(32'hb9659821),
	.w6(32'h38dafaca),
	.w7(32'hb75438de),
	.w8(32'hb8dcaf37),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b03e8),
	.w1(32'hb95312af),
	.w2(32'hb98b11d9),
	.w3(32'hb87038d5),
	.w4(32'hb98a39ed),
	.w5(32'hb9a9c7fb),
	.w6(32'h381349da),
	.w7(32'hb8c33a0b),
	.w8(32'hb90bb6ce),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394443b4),
	.w1(32'h3939f0cc),
	.w2(32'h39358b40),
	.w3(32'h39160220),
	.w4(32'h395c3fa3),
	.w5(32'h39688a2b),
	.w6(32'h391c348e),
	.w7(32'h39689a32),
	.w8(32'h39248b3d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79540d7),
	.w1(32'h37a7925e),
	.w2(32'h386c17a1),
	.w3(32'hb8199664),
	.w4(32'h3789efbe),
	.w5(32'h37dd25d3),
	.w6(32'hb77c8e1e),
	.w7(32'h38139b6c),
	.w8(32'h3879ef47),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38833b21),
	.w1(32'hb78bd344),
	.w2(32'hb7e57bd4),
	.w3(32'h382f2fc5),
	.w4(32'h359207ad),
	.w5(32'hb7aeb859),
	.w6(32'h37f4537b),
	.w7(32'h3723ca01),
	.w8(32'h36289937),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4016c),
	.w1(32'hb6240de3),
	.w2(32'hb71ab3bc),
	.w3(32'h37f315ab),
	.w4(32'hb686b9a6),
	.w5(32'hb76be0c0),
	.w6(32'h37ed87c7),
	.w7(32'h37b36e4b),
	.w8(32'hb5b76d22),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793799d),
	.w1(32'hb7b9d33c),
	.w2(32'hb78b5166),
	.w3(32'hb79b02b0),
	.w4(32'hb7147364),
	.w5(32'hb6f1dbc6),
	.w6(32'hb7bc4848),
	.w7(32'hb7175e37),
	.w8(32'hb6e49b0c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f6849),
	.w1(32'hb9208d4d),
	.w2(32'hb960cd39),
	.w3(32'hb9061a8c),
	.w4(32'hb9848e9d),
	.w5(32'hb9950357),
	.w6(32'hb8bfb1cd),
	.w7(32'hb94f3fde),
	.w8(32'hb96069aa),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5f432),
	.w1(32'hb7f7fe13),
	.w2(32'hb80acc57),
	.w3(32'hb7406027),
	.w4(32'hb7a3bdce),
	.w5(32'hb7c43f6d),
	.w6(32'hb61e7197),
	.w7(32'hb727e1dd),
	.w8(32'hb70ef892),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970b19c),
	.w1(32'hb9693cac),
	.w2(32'hb9570aea),
	.w3(32'hb9591fc7),
	.w4(32'hb8b538ea),
	.w5(32'hb90e5ea7),
	.w6(32'hb8dc77ad),
	.w7(32'hb869ab40),
	.w8(32'hb91cf51d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule