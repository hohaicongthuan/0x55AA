module layer_10_featuremap_308(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a7d4f),
	.w1(32'h3c88507a),
	.w2(32'hbb243231),
	.w3(32'h3ca5fa29),
	.w4(32'h3b6477f8),
	.w5(32'hbbc9bb5b),
	.w6(32'h3d019897),
	.w7(32'h3c051d29),
	.w8(32'hbc175bfa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59d99b),
	.w1(32'hbc2dda68),
	.w2(32'hbbde4fb3),
	.w3(32'hbc088828),
	.w4(32'hbc7fb133),
	.w5(32'hbb919fac),
	.w6(32'hbb517d3f),
	.w7(32'hbc20833b),
	.w8(32'hbb82ae3b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399edfab),
	.w1(32'h3b983b66),
	.w2(32'h3b4e2a2b),
	.w3(32'hbba88456),
	.w4(32'hba087f76),
	.w5(32'h3c3c493c),
	.w6(32'hbba6cd91),
	.w7(32'h3a8ca46f),
	.w8(32'h3c397f1b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35d22c),
	.w1(32'h3c16e55d),
	.w2(32'h3c2a27d7),
	.w3(32'h3c06ce7f),
	.w4(32'h3c1d3f0a),
	.w5(32'h3b850550),
	.w6(32'h3c654a61),
	.w7(32'h3c2a8aba),
	.w8(32'h3c12d29d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18453a),
	.w1(32'hbafb0dae),
	.w2(32'h3b930067),
	.w3(32'h3b8bea31),
	.w4(32'hb9c89e52),
	.w5(32'h3b516fc8),
	.w6(32'h3bdf4558),
	.w7(32'h3c54ba89),
	.w8(32'h3bdc0f7c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb0ad),
	.w1(32'h3c4fd288),
	.w2(32'h3aa02801),
	.w3(32'h3c2df76f),
	.w4(32'h3a88695c),
	.w5(32'hbc40aefb),
	.w6(32'h3cb56798),
	.w7(32'h3c0ab9a7),
	.w8(32'hbb7308c6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9c22),
	.w1(32'h3b9d93a1),
	.w2(32'hbc0cc2a2),
	.w3(32'h3995cb49),
	.w4(32'hbc0549a3),
	.w5(32'hbba268f1),
	.w6(32'h3c57bd28),
	.w7(32'hbb133c25),
	.w8(32'hbb91a932),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299e76),
	.w1(32'h3bc99e44),
	.w2(32'hbc48f395),
	.w3(32'h3bc8fdff),
	.w4(32'h3b05d482),
	.w5(32'hbbb1e8d1),
	.w6(32'h3c9bc20c),
	.w7(32'h3b7afde3),
	.w8(32'hb9f486f5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6521b),
	.w1(32'h3c59cc76),
	.w2(32'h3b233611),
	.w3(32'h3c0a12d8),
	.w4(32'h3b799ba5),
	.w5(32'h3be6d47c),
	.w6(32'h3c88805f),
	.w7(32'h3c235f2c),
	.w8(32'h3c172fb5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf7d7b),
	.w1(32'h3c2b0555),
	.w2(32'hba893243),
	.w3(32'h3c6ed531),
	.w4(32'h3b56cc3b),
	.w5(32'hba9eb8bf),
	.w6(32'h3cc46141),
	.w7(32'h3bfc4a11),
	.w8(32'hb8f84b14),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334bda),
	.w1(32'h3c60bc38),
	.w2(32'h3be2ff03),
	.w3(32'h3c1a9886),
	.w4(32'h3bc8c09f),
	.w5(32'h39c9dd0d),
	.w6(32'h3cbae6ca),
	.w7(32'h3c805b1b),
	.w8(32'hbbaec713),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbbd35),
	.w1(32'h3b5fab8f),
	.w2(32'hbc00c018),
	.w3(32'hba87ec9f),
	.w4(32'h3b1427f3),
	.w5(32'h3b1a1e12),
	.w6(32'hbbc10304),
	.w7(32'hb9587f80),
	.w8(32'h3bcbcc04),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93beec),
	.w1(32'h3c118552),
	.w2(32'hbad76c6e),
	.w3(32'h3bfa7c75),
	.w4(32'h3aa5e36c),
	.w5(32'hbbea9830),
	.w6(32'h3c7eb285),
	.w7(32'h3c30fea5),
	.w8(32'hbc0c8aed),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee1ba),
	.w1(32'h39d2b373),
	.w2(32'hbbda8936),
	.w3(32'hbb73863a),
	.w4(32'hbc12e20c),
	.w5(32'hbc35969b),
	.w6(32'hbba23a34),
	.w7(32'hbc17863a),
	.w8(32'hbba656ba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0855c2),
	.w1(32'h3916812c),
	.w2(32'hbb8c7645),
	.w3(32'hbac8b0ba),
	.w4(32'hbae03a49),
	.w5(32'h3b0b3ea6),
	.w6(32'h3c0607b7),
	.w7(32'h3aefbe5a),
	.w8(32'h3c1e1390),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119532),
	.w1(32'h3c1f3700),
	.w2(32'hbbb43322),
	.w3(32'h3b8b3481),
	.w4(32'h3b4335b1),
	.w5(32'h3b4268a2),
	.w6(32'h3c969a1e),
	.w7(32'hbb111b1d),
	.w8(32'h3bffc701),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174590),
	.w1(32'h3bf0df0b),
	.w2(32'hb9621cea),
	.w3(32'h3c1fa3f6),
	.w4(32'hba835e6b),
	.w5(32'hbb60c19a),
	.w6(32'h3c9b197b),
	.w7(32'h3c126863),
	.w8(32'hba09b7f1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c51d3),
	.w1(32'h3aedaa5f),
	.w2(32'hbb6feb4a),
	.w3(32'hbb8796c6),
	.w4(32'hbc074b4d),
	.w5(32'hbc6f1654),
	.w6(32'hbab1cdd9),
	.w7(32'hbb1f8e4f),
	.w8(32'hbca00cc0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84564),
	.w1(32'hbbeef2bf),
	.w2(32'hbbce8d2e),
	.w3(32'hbbe0e885),
	.w4(32'hbc2bc52a),
	.w5(32'hb8d47154),
	.w6(32'hbc1f2154),
	.w7(32'hbc746d2f),
	.w8(32'hbb263a8b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7deb),
	.w1(32'hbb75b740),
	.w2(32'h3aed76c6),
	.w3(32'hb946811b),
	.w4(32'hba132e50),
	.w5(32'hbb9f0100),
	.w6(32'hbb248a54),
	.w7(32'hbb508738),
	.w8(32'h39d0bcba),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb690638),
	.w1(32'h3ba511b4),
	.w2(32'hbb88263f),
	.w3(32'hbb39ee90),
	.w4(32'hbb88aa1b),
	.w5(32'h3b69c4ce),
	.w6(32'h3c1ae8e8),
	.w7(32'hbc2329a5),
	.w8(32'h3999f108),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7bd59),
	.w1(32'hbb301c3b),
	.w2(32'hbae594d7),
	.w3(32'hba6217b4),
	.w4(32'hba65c629),
	.w5(32'h3a8f1c35),
	.w6(32'hbbad4e0c),
	.w7(32'hbb7b44b9),
	.w8(32'hbaccb572),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf009b9),
	.w1(32'h3c13a0c8),
	.w2(32'h3bc68658),
	.w3(32'h3b3ca682),
	.w4(32'h3aa0238b),
	.w5(32'hbb68eccf),
	.w6(32'hbba35df0),
	.w7(32'hba5ce669),
	.w8(32'h3acdf1a9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2acb),
	.w1(32'hb946c397),
	.w2(32'hbb9647dc),
	.w3(32'hba6790db),
	.w4(32'hbb8166f5),
	.w5(32'hbb024a5c),
	.w6(32'h3a8954f0),
	.w7(32'hbb93aacf),
	.w8(32'h3adb3283),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b7ef),
	.w1(32'hba79cba0),
	.w2(32'h3badf617),
	.w3(32'hbb2741d0),
	.w4(32'hba908620),
	.w5(32'hbba060a0),
	.w6(32'h3b5e5129),
	.w7(32'h3b88a81c),
	.w8(32'h3b80ded1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36709b),
	.w1(32'h3b682511),
	.w2(32'hbbdf28b7),
	.w3(32'h3b9a99bc),
	.w4(32'hbc0d3eda),
	.w5(32'hbba294e4),
	.w6(32'h3cbc4c42),
	.w7(32'h3b148436),
	.w8(32'hbc01f1e3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd92bc4),
	.w1(32'hbbca2da5),
	.w2(32'hbac70a78),
	.w3(32'hbba6e19b),
	.w4(32'hbb56647a),
	.w5(32'h3b5bc55d),
	.w6(32'hbb8ea318),
	.w7(32'hbab0686b),
	.w8(32'h3c09efa7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14daf0),
	.w1(32'h3c98b9cd),
	.w2(32'h388e7ff4),
	.w3(32'h3cb28d5c),
	.w4(32'h3c173df4),
	.w5(32'hb9f9cd50),
	.w6(32'h3ce46a1d),
	.w7(32'h3c485f39),
	.w8(32'hbbf2bb0c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba704a43),
	.w1(32'hbb1ec6a4),
	.w2(32'h3b157777),
	.w3(32'h3b21b458),
	.w4(32'hbb15898b),
	.w5(32'hbc03f9d3),
	.w6(32'hbb7c4c97),
	.w7(32'hbab3cf68),
	.w8(32'hbc154435),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03eef),
	.w1(32'hb97c68a3),
	.w2(32'h3b419a71),
	.w3(32'hbbd524b5),
	.w4(32'hbb761778),
	.w5(32'h3c248b40),
	.w6(32'hbb6f642d),
	.w7(32'hbb567aa0),
	.w8(32'h3c24ff81),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a88ac),
	.w1(32'h3bdd44d2),
	.w2(32'h3c2b2018),
	.w3(32'h3c30b82c),
	.w4(32'h3c0b8e9a),
	.w5(32'h3b821e30),
	.w6(32'h39bfdf43),
	.w7(32'h3ac1fafa),
	.w8(32'hba1e403d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f699),
	.w1(32'h3a2eee92),
	.w2(32'h3ae000ac),
	.w3(32'hbb7c1734),
	.w4(32'h3b364f8b),
	.w5(32'hbbb3ff77),
	.w6(32'hbcb2a0ca),
	.w7(32'hbc2d3353),
	.w8(32'hbba1f59a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd806),
	.w1(32'hbbb86272),
	.w2(32'hbae55b4b),
	.w3(32'hbb85832f),
	.w4(32'hbbaf223d),
	.w5(32'hbb3e5db3),
	.w6(32'hbc025006),
	.w7(32'hbbe382df),
	.w8(32'hba367190),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a489),
	.w1(32'h384bca52),
	.w2(32'h3b6884ef),
	.w3(32'hba072df3),
	.w4(32'hba03d291),
	.w5(32'h3bbd30f8),
	.w6(32'hba430084),
	.w7(32'h3babb78f),
	.w8(32'hba078ad7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8da2a8),
	.w1(32'hbbf3e21c),
	.w2(32'hbc0752ef),
	.w3(32'h3bc96ade),
	.w4(32'hbb3d9ae3),
	.w5(32'hbb464e43),
	.w6(32'hbb300ee7),
	.w7(32'hbb9b7b90),
	.w8(32'h3bcfef84),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbf1c1),
	.w1(32'h3be096c3),
	.w2(32'h3b01d6e1),
	.w3(32'h3b901d6d),
	.w4(32'hb80c9742),
	.w5(32'hbaf4792b),
	.w6(32'h3c8db4bd),
	.w7(32'h3a89784a),
	.w8(32'hbb9be167),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574861),
	.w1(32'h3beb54e9),
	.w2(32'hba465126),
	.w3(32'h3a73c989),
	.w4(32'hb97ffe58),
	.w5(32'hbbc3aa7d),
	.w6(32'h3b34cacb),
	.w7(32'h3b93134b),
	.w8(32'h3a81eca2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d63da),
	.w1(32'h3c218d6c),
	.w2(32'hb9b90630),
	.w3(32'h3bfa6692),
	.w4(32'hbb968ca9),
	.w5(32'h3c20bc0f),
	.w6(32'h3c93dd1f),
	.w7(32'hbad0aa0b),
	.w8(32'h3bc46d3a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1e200),
	.w1(32'hbc0e4666),
	.w2(32'h3baea982),
	.w3(32'hbbafbaa4),
	.w4(32'hbc2e9192),
	.w5(32'h3c7ecc49),
	.w6(32'hbc61b821),
	.w7(32'hbbaa1406),
	.w8(32'h3c910b00),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4504fe),
	.w1(32'h3aeec1f0),
	.w2(32'h3aca34d7),
	.w3(32'h3b732370),
	.w4(32'h3b503e1a),
	.w5(32'h3bece532),
	.w6(32'h3a3d60be),
	.w7(32'hbb63564d),
	.w8(32'h3acaf407),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dfae9),
	.w1(32'h3c39b558),
	.w2(32'h38db9a46),
	.w3(32'h3aa80998),
	.w4(32'h3ad20690),
	.w5(32'hbbf8b0db),
	.w6(32'h3b7400c5),
	.w7(32'h3b7e2df7),
	.w8(32'h39eb0f3d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14c37e),
	.w1(32'h3ada0404),
	.w2(32'hbc03a0f8),
	.w3(32'h3956c28d),
	.w4(32'hbc275c42),
	.w5(32'hbb2ab318),
	.w6(32'h3ca99dfa),
	.w7(32'h3a766de6),
	.w8(32'hbb21052e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5865a),
	.w1(32'hbb6810c2),
	.w2(32'hbbf6b5e3),
	.w3(32'h390991c5),
	.w4(32'hbb8569fe),
	.w5(32'h3c2aa945),
	.w6(32'h3bd19e3c),
	.w7(32'hbb0c487f),
	.w8(32'h3c283479),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c119e26),
	.w1(32'h3c26829c),
	.w2(32'h3bad1ee8),
	.w3(32'h3c5baa95),
	.w4(32'h3bd4904c),
	.w5(32'h3b1f3982),
	.w6(32'h3c7ee817),
	.w7(32'h3c0e16ca),
	.w8(32'h3b93eab9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfacb34),
	.w1(32'h3c406015),
	.w2(32'h3c48051c),
	.w3(32'h3c199260),
	.w4(32'h3c0c52da),
	.w5(32'hbbb737ef),
	.w6(32'h3c9cf8a9),
	.w7(32'h3c8f401e),
	.w8(32'hbaaa79bc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c65f),
	.w1(32'hbb9c9fff),
	.w2(32'hbbf1e1d8),
	.w3(32'hbc27f172),
	.w4(32'hbc21239e),
	.w5(32'hbb4d8291),
	.w6(32'hbb384b0f),
	.w7(32'hba080d13),
	.w8(32'hbb864a49),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25d65),
	.w1(32'hbc4fdaa2),
	.w2(32'hbbe819cd),
	.w3(32'hbc1f62e2),
	.w4(32'hbbb1bd75),
	.w5(32'h3c17c7d3),
	.w6(32'hbbf4ef6c),
	.w7(32'hbb87be16),
	.w8(32'h3c071b79),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca4d38),
	.w1(32'h3bdf6142),
	.w2(32'hba8fca82),
	.w3(32'h3c780364),
	.w4(32'h3bdd90e5),
	.w5(32'hbc9f6131),
	.w6(32'h3bda6884),
	.w7(32'h3b0b9160),
	.w8(32'hbc48ea3d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c023),
	.w1(32'hba81e779),
	.w2(32'hbba39ebc),
	.w3(32'hbb94e922),
	.w4(32'hbc140dc4),
	.w5(32'hbb32bb17),
	.w6(32'h3b27d03b),
	.w7(32'h3adbdc72),
	.w8(32'h394748d2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba145f5),
	.w1(32'hb9ee1fa6),
	.w2(32'hbc04fae6),
	.w3(32'h3ad46a30),
	.w4(32'hbbdd1384),
	.w5(32'h3b2e8282),
	.w6(32'h3bbc4fd4),
	.w7(32'hbbab6d1b),
	.w8(32'hbb3c30a5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb541282),
	.w1(32'hbbcbc398),
	.w2(32'h39ae2185),
	.w3(32'hbb5bc22f),
	.w4(32'hb8d6b26d),
	.w5(32'hbb9e65ce),
	.w6(32'hbc1bde75),
	.w7(32'hba00562e),
	.w8(32'hbc1c9af1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefdbfc),
	.w1(32'hbc56dc86),
	.w2(32'hbc358c86),
	.w3(32'hbc016bf4),
	.w4(32'hbb926d93),
	.w5(32'hbb1c499f),
	.w6(32'hbc053c43),
	.w7(32'hbc425f49),
	.w8(32'hbbaefd6f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831878),
	.w1(32'h3b8e1292),
	.w2(32'hbafd79bf),
	.w3(32'hbb886dc2),
	.w4(32'h3b987a3c),
	.w5(32'hbaef9b70),
	.w6(32'hba9abcc5),
	.w7(32'h3989c4ce),
	.w8(32'h3a300269),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5d6d1),
	.w1(32'hbbc26534),
	.w2(32'hbb40034c),
	.w3(32'hbbeffb42),
	.w4(32'h3b228db1),
	.w5(32'hb9af7830),
	.w6(32'hbc19f9ff),
	.w7(32'hbaa07e8a),
	.w8(32'hbbc78d57),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2742),
	.w1(32'hbad35ee9),
	.w2(32'h3b51b47f),
	.w3(32'h3aed4c59),
	.w4(32'h3b82cf40),
	.w5(32'h3b190ac2),
	.w6(32'h3b2dbbb1),
	.w7(32'h3b1893ec),
	.w8(32'h3b93c0f9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5101),
	.w1(32'h3bbb00d3),
	.w2(32'hbabc2355),
	.w3(32'hbb5cdc7d),
	.w4(32'hbbf39edc),
	.w5(32'h3bffd630),
	.w6(32'h3b2b42dc),
	.w7(32'hbb86b50f),
	.w8(32'h3b10ddc4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a6c6),
	.w1(32'h3b9282db),
	.w2(32'h3bb25776),
	.w3(32'h3aece021),
	.w4(32'h39c67f9d),
	.w5(32'h3b2c02a1),
	.w6(32'h3a07bd4f),
	.w7(32'h3b138a03),
	.w8(32'hbb101250),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6afbd),
	.w1(32'h3b3153a4),
	.w2(32'hbaa561c5),
	.w3(32'h3b8340f8),
	.w4(32'h3c026d14),
	.w5(32'hbc433bdf),
	.w6(32'h3bfef12b),
	.w7(32'h3b612aee),
	.w8(32'hbbe40187),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc381c83),
	.w1(32'hbaa12c02),
	.w2(32'hbbdf2c36),
	.w3(32'hba99187c),
	.w4(32'hbc0020b9),
	.w5(32'hbb877ee9),
	.w6(32'h3bdfb730),
	.w7(32'hbb831320),
	.w8(32'hbc3e4312),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2165ab),
	.w1(32'hbc42fc11),
	.w2(32'hbc13ec1f),
	.w3(32'hbb8dc4a2),
	.w4(32'hbbf3eab6),
	.w5(32'h38b0447c),
	.w6(32'hbc46244a),
	.w7(32'hbc32eb0c),
	.w8(32'h39293f19),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4751fe),
	.w1(32'hba4e349f),
	.w2(32'hbb68f475),
	.w3(32'h3bde51dc),
	.w4(32'hbb464eff),
	.w5(32'h3a05868e),
	.w6(32'h3afc5dad),
	.w7(32'hbb71a64a),
	.w8(32'h3b64d591),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f187d6),
	.w1(32'hba9ef82d),
	.w2(32'hbbd35f99),
	.w3(32'h3b76262f),
	.w4(32'hba7dd131),
	.w5(32'hbb523232),
	.w6(32'h3cc2746a),
	.w7(32'h3b8a42b5),
	.w8(32'h3b5705e4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ca795),
	.w1(32'hbb6e52d6),
	.w2(32'h39b4d784),
	.w3(32'hbb262119),
	.w4(32'hbb90518e),
	.w5(32'hba1b3a10),
	.w6(32'hbb60d347),
	.w7(32'h3acddb31),
	.w8(32'hbbc8ceaa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494fb1),
	.w1(32'h3a052e2d),
	.w2(32'hbb2dd568),
	.w3(32'hbabce4e9),
	.w4(32'hbb97e3ea),
	.w5(32'h3bd0f919),
	.w6(32'hba996296),
	.w7(32'hbb080c9b),
	.w8(32'h3ad94652),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb81e),
	.w1(32'hbbd2b3f4),
	.w2(32'h3a1bc2cf),
	.w3(32'hbb409529),
	.w4(32'hba9e3581),
	.w5(32'h3a4a78ed),
	.w6(32'hbb817643),
	.w7(32'hba012858),
	.w8(32'h3a59e9ca),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38683f0f),
	.w1(32'hba0c3c34),
	.w2(32'hba2efd29),
	.w3(32'hbb0b8343),
	.w4(32'h3afa0d93),
	.w5(32'hbb1520c1),
	.w6(32'h3ad0010f),
	.w7(32'h3a9743d8),
	.w8(32'h3bc98707),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d92f2),
	.w1(32'h3c2a1a0e),
	.w2(32'hbc9a7b27),
	.w3(32'h3bbd9a9d),
	.w4(32'h3bf0f893),
	.w5(32'h3b87978e),
	.w6(32'h3c75401e),
	.w7(32'h3b4d7f9e),
	.w8(32'h3ba8018c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c116f),
	.w1(32'h3c81d24b),
	.w2(32'h3c492874),
	.w3(32'h3c88022f),
	.w4(32'h3c720d31),
	.w5(32'hbbc2a961),
	.w6(32'h3cb21009),
	.w7(32'h3c8cd86e),
	.w8(32'hbaf1e779),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecd0c0),
	.w1(32'hbbcc8b41),
	.w2(32'hbb2ec832),
	.w3(32'hbbaa53f0),
	.w4(32'hba6c6504),
	.w5(32'hbbb55560),
	.w6(32'hbbb04c38),
	.w7(32'hbae1d0eb),
	.w8(32'h3b125599),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba4890),
	.w1(32'h3ad2e062),
	.w2(32'h3bfe5fdc),
	.w3(32'hbbd1d083),
	.w4(32'h3ac4cf3a),
	.w5(32'h3bbddbb2),
	.w6(32'h3ae1152d),
	.w7(32'h3c6298b7),
	.w8(32'h3bbccea2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0a71e),
	.w1(32'h3b21b547),
	.w2(32'hbb03a7a1),
	.w3(32'h3b974234),
	.w4(32'hbb06beb2),
	.w5(32'hbb29e512),
	.w6(32'h3b6d44aa),
	.w7(32'hbb4f0af3),
	.w8(32'hb733200a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af924d3),
	.w1(32'hb9fb9d73),
	.w2(32'hbbb4ca79),
	.w3(32'h3b94c07a),
	.w4(32'h3ba56334),
	.w5(32'hbb1489b4),
	.w6(32'h3c04b730),
	.w7(32'hbbe4211d),
	.w8(32'h3a86ccce),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eeb41),
	.w1(32'hbc2db40b),
	.w2(32'hbb0a9758),
	.w3(32'hbaedb712),
	.w4(32'hbace6bc2),
	.w5(32'hbbbbdaba),
	.w6(32'h3c5cc2d6),
	.w7(32'h3b5d5243),
	.w8(32'hbc54e77d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f9f7),
	.w1(32'hbc672609),
	.w2(32'hbb99aca8),
	.w3(32'hba994c5b),
	.w4(32'hbc316440),
	.w5(32'h3bcf901c),
	.w6(32'hbb1e54a6),
	.w7(32'hb9bce94e),
	.w8(32'h3c0c1d50),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39c9a),
	.w1(32'h3c608c8c),
	.w2(32'hbb8081ab),
	.w3(32'h3c135a2b),
	.w4(32'h39cc211a),
	.w5(32'hb9da8a35),
	.w6(32'h3c7df29b),
	.w7(32'h3c140e70),
	.w8(32'h38b31d83),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac228d7),
	.w1(32'h3a3281f9),
	.w2(32'hbb95c145),
	.w3(32'h3a9e1f55),
	.w4(32'hba90193e),
	.w5(32'hbbd70660),
	.w6(32'h3a50805c),
	.w7(32'hbab55fc7),
	.w8(32'hbc1469d5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5903b0),
	.w1(32'h3c11a59a),
	.w2(32'hbb8e6067),
	.w3(32'hba2426b6),
	.w4(32'h3ad52f3f),
	.w5(32'hbbd3a4f5),
	.w6(32'h3b8d9344),
	.w7(32'hbb6aeb5b),
	.w8(32'hbc1ebb22),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3b3d),
	.w1(32'hbc2ce894),
	.w2(32'hbb7d7e65),
	.w3(32'hbc00f734),
	.w4(32'h3b1125c7),
	.w5(32'h3bd3966d),
	.w6(32'hbc32a9f4),
	.w7(32'hbb89a8c4),
	.w8(32'h3bcd8eab),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc0841),
	.w1(32'h3b8c61d4),
	.w2(32'h3b2c9f49),
	.w3(32'h3b255325),
	.w4(32'h3c172e5e),
	.w5(32'hbb35d552),
	.w6(32'h3bc113d1),
	.w7(32'h3bca8d32),
	.w8(32'h3ba1edb4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1c200),
	.w1(32'h3c3e895c),
	.w2(32'hbbb3235a),
	.w3(32'h3c31bc9a),
	.w4(32'h3bbf1091),
	.w5(32'hbc3cdbd7),
	.w6(32'h3caf16a7),
	.w7(32'h3c554bfa),
	.w8(32'hbc8736e0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b50ad),
	.w1(32'hbc77afb9),
	.w2(32'hbc827c16),
	.w3(32'hbc34910e),
	.w4(32'hbc1fd195),
	.w5(32'hbbbf0983),
	.w6(32'hbc6f82b9),
	.w7(32'hbc64120f),
	.w8(32'h3ada1eb0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba371a8),
	.w1(32'hbb5460a9),
	.w2(32'hbbeccfca),
	.w3(32'h3a4858c0),
	.w4(32'hbba4638e),
	.w5(32'hbbbf4a4e),
	.w6(32'h3c0e3272),
	.w7(32'h39bc53a4),
	.w8(32'hbbcaa7de),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b714096),
	.w1(32'hba33195a),
	.w2(32'hbba3337a),
	.w3(32'hbb2e0115),
	.w4(32'h3bb52521),
	.w5(32'h3c5f085f),
	.w6(32'hbb9ea5f7),
	.w7(32'h3aa5315d),
	.w8(32'h3be06e1f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29060d),
	.w1(32'h3baf969e),
	.w2(32'h3c97973d),
	.w3(32'h3bfa07be),
	.w4(32'h3cad2b0c),
	.w5(32'h3b374698),
	.w6(32'h3acfdc47),
	.w7(32'h3c6e4193),
	.w8(32'h3ab941e4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b2ea),
	.w1(32'h3b84009d),
	.w2(32'h3b4b4c85),
	.w3(32'h3ae184f1),
	.w4(32'h3be4ae98),
	.w5(32'h3ae8fda5),
	.w6(32'hbad93121),
	.w7(32'h3baf8f0b),
	.w8(32'h3b68acff),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ea3d),
	.w1(32'h3b355d59),
	.w2(32'h3b2e0cf1),
	.w3(32'h3a5ec7c2),
	.w4(32'h3b600a2c),
	.w5(32'hbbd6688b),
	.w6(32'h3c0dad18),
	.w7(32'h3c3defa9),
	.w8(32'hbb845c31),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f816),
	.w1(32'hbb1d20e5),
	.w2(32'hbb8b30e0),
	.w3(32'hbbb9ac57),
	.w4(32'hbb8618a9),
	.w5(32'h3be60299),
	.w6(32'h3b807893),
	.w7(32'hbaff4a9e),
	.w8(32'h3b35c3c2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3084ed),
	.w1(32'hbb68764e),
	.w2(32'hbb2e5cee),
	.w3(32'hb9a77bf6),
	.w4(32'hba712bac),
	.w5(32'hbba00a7a),
	.w6(32'hbbcad88d),
	.w7(32'hbb70c717),
	.w8(32'h3b24c63e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5d8c),
	.w1(32'h3c01df26),
	.w2(32'hbb29032e),
	.w3(32'h3bcecc69),
	.w4(32'hbb92cded),
	.w5(32'hbb9c63a2),
	.w6(32'h3c97447f),
	.w7(32'h3b9c6b8f),
	.w8(32'hbbd6a334),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affb863),
	.w1(32'h3bb83f50),
	.w2(32'hbc015f17),
	.w3(32'h3baecec8),
	.w4(32'hbc0af958),
	.w5(32'hbc6ae7d0),
	.w6(32'h3cadbe86),
	.w7(32'hbb8aa1a8),
	.w8(32'hbb0419ea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a21d),
	.w1(32'hbb2cefde),
	.w2(32'hb9d9c6e2),
	.w3(32'hbbf81be3),
	.w4(32'hbace5a05),
	.w5(32'h3ac9d814),
	.w6(32'hbc83fa82),
	.w7(32'h3ae92e87),
	.w8(32'h3b32a7f2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1ebf),
	.w1(32'h3b79b2c5),
	.w2(32'hbc15ed38),
	.w3(32'h3c2da6ab),
	.w4(32'h3bab49c4),
	.w5(32'h39e5378f),
	.w6(32'h3c6dcf63),
	.w7(32'h3a63352f),
	.w8(32'hbb334c83),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a54e3),
	.w1(32'h3be83626),
	.w2(32'h3be8e87c),
	.w3(32'h3bae4bd4),
	.w4(32'h3ba744f6),
	.w5(32'h399f7a46),
	.w6(32'hbb06003a),
	.w7(32'hba520f33),
	.w8(32'hb999f130),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb8b5d),
	.w1(32'hb8204d02),
	.w2(32'hbc5f4dbc),
	.w3(32'h3a3b61a3),
	.w4(32'hbc1d2db9),
	.w5(32'hbb874708),
	.w6(32'h3b6f5eed),
	.w7(32'hbc57372f),
	.w8(32'hbaba63a5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52cb07),
	.w1(32'h3c30dfe9),
	.w2(32'hbc23f7b2),
	.w3(32'h3c707516),
	.w4(32'h3b1d3115),
	.w5(32'hbb1320ae),
	.w6(32'h3cd01c86),
	.w7(32'hbb11aa48),
	.w8(32'hbbd24e54),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c520),
	.w1(32'h3b216eb0),
	.w2(32'hbbb05a9d),
	.w3(32'hbade9cea),
	.w4(32'hbbedcafe),
	.w5(32'h3c62bed6),
	.w6(32'hbaf72d78),
	.w7(32'hbc4dc740),
	.w8(32'h3bce9525),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103f0e),
	.w1(32'h3b520251),
	.w2(32'h3c03fff3),
	.w3(32'h3bab3a97),
	.w4(32'h3c1a886a),
	.w5(32'h3a91900f),
	.w6(32'hba276354),
	.w7(32'h3aa0534c),
	.w8(32'hbb8350bd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824b75),
	.w1(32'h3b27dcc4),
	.w2(32'hbb285d27),
	.w3(32'h3b0748bb),
	.w4(32'hbab5adc9),
	.w5(32'h3b428dcf),
	.w6(32'hbc35b91b),
	.w7(32'hbb73941c),
	.w8(32'h3af2374f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61ae8d),
	.w1(32'h3c1a39a1),
	.w2(32'hbb0b2751),
	.w3(32'h3bcbe3b5),
	.w4(32'h3b5b693e),
	.w5(32'hbb343a74),
	.w6(32'h3ba86089),
	.w7(32'h3aa1713d),
	.w8(32'hbb575b34),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9d70d),
	.w1(32'h3bc6248e),
	.w2(32'h3ad19b54),
	.w3(32'h3afbff1b),
	.w4(32'hbb3442e0),
	.w5(32'h3ba14984),
	.w6(32'h3c18f805),
	.w7(32'h3b5e0933),
	.w8(32'h3bb7d473),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c221ba7),
	.w1(32'h3b87b34d),
	.w2(32'h3c564c34),
	.w3(32'hbc11b67a),
	.w4(32'h3ba01761),
	.w5(32'h3c8afa54),
	.w6(32'hbc00a8e0),
	.w7(32'h3ab6c162),
	.w8(32'h3c78c3ed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf12de),
	.w1(32'hbba7c531),
	.w2(32'hbbd4c034),
	.w3(32'h3af89f13),
	.w4(32'h39003cc4),
	.w5(32'h3a235007),
	.w6(32'hbaf7cca4),
	.w7(32'hbb36c676),
	.w8(32'h3b88faa0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d640),
	.w1(32'h3b63ea1a),
	.w2(32'hbbb8a906),
	.w3(32'h3a5c1be0),
	.w4(32'hba9b1efd),
	.w5(32'hbb8551fe),
	.w6(32'hb9cb7041),
	.w7(32'hbb7a8884),
	.w8(32'hbbd9c812),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5256),
	.w1(32'hbb5c8c2b),
	.w2(32'hbba1f78d),
	.w3(32'hbbe987a4),
	.w4(32'hbc3091fe),
	.w5(32'hbb242428),
	.w6(32'hbb41d011),
	.w7(32'hbbe65126),
	.w8(32'h3b0b5d28),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d96f),
	.w1(32'h3a0360ed),
	.w2(32'hbae09195),
	.w3(32'hbb5fe52a),
	.w4(32'hbb8863fa),
	.w5(32'h3b623577),
	.w6(32'h3c051476),
	.w7(32'hbb9da873),
	.w8(32'h3b89b826),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17c282),
	.w1(32'h3b937a97),
	.w2(32'h3ab06db3),
	.w3(32'h3bbce2d9),
	.w4(32'h3bfa35fe),
	.w5(32'h3b0324a5),
	.w6(32'h3adf194c),
	.w7(32'h3b32310a),
	.w8(32'hb9cce68e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f30cb),
	.w1(32'h3b136f19),
	.w2(32'h3a82865b),
	.w3(32'h3b66daf5),
	.w4(32'h3a8855f3),
	.w5(32'hbb0b9c10),
	.w6(32'hb9e265ef),
	.w7(32'hbbc49194),
	.w8(32'hbb57dfeb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76a37c),
	.w1(32'hbaef5937),
	.w2(32'hbb924330),
	.w3(32'h3bdc9b42),
	.w4(32'h3b8bde4f),
	.w5(32'h3b0ba216),
	.w6(32'h3bf8c9bf),
	.w7(32'h3b7e18dc),
	.w8(32'h3b6372bf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091955),
	.w1(32'h3b9fa8fc),
	.w2(32'h3b1fa132),
	.w3(32'h39f9eeae),
	.w4(32'hbaacc4a7),
	.w5(32'h3c3aff7a),
	.w6(32'h3929b7b4),
	.w7(32'hbb0d4ab5),
	.w8(32'h3bb0eec8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9452e2),
	.w1(32'hbb403237),
	.w2(32'hba02b352),
	.w3(32'h3bf309bc),
	.w4(32'h3c30113b),
	.w5(32'h3aaaabf9),
	.w6(32'h3b142f1b),
	.w7(32'h3beaec0f),
	.w8(32'h3ae2dd98),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bb92),
	.w1(32'hbb848b80),
	.w2(32'h3b9e3182),
	.w3(32'hbb9497c1),
	.w4(32'hbb908d60),
	.w5(32'hbba29a8e),
	.w6(32'hbbc746da),
	.w7(32'hbb0cac0c),
	.w8(32'hbb338ead),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4e16d),
	.w1(32'hbb187e08),
	.w2(32'hbb28f9cb),
	.w3(32'hbb17d08a),
	.w4(32'hba9d5de0),
	.w5(32'h3c77db34),
	.w6(32'hbb8a0b00),
	.w7(32'hbb87d909),
	.w8(32'h3c148065),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f63a8),
	.w1(32'h392df474),
	.w2(32'h3b913082),
	.w3(32'h3ba63171),
	.w4(32'h3bce413e),
	.w5(32'hbb7b0778),
	.w6(32'h3ae5d3a4),
	.w7(32'h3bfbbfda),
	.w8(32'h3aeeaf8d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac79276),
	.w1(32'h3ab39317),
	.w2(32'hba9b53e8),
	.w3(32'hbb204ad9),
	.w4(32'hbb86911c),
	.w5(32'hba18dfe6),
	.w6(32'h3bb388c7),
	.w7(32'hbafa55b3),
	.w8(32'hbb279cc4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a1c1f),
	.w1(32'hbb013014),
	.w2(32'h3a90db92),
	.w3(32'hbb5cbb10),
	.w4(32'hbb2b1f23),
	.w5(32'hbb6988b8),
	.w6(32'h3a9bb051),
	.w7(32'hb9b5b9ab),
	.w8(32'hbab14edc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c3dd1),
	.w1(32'hbb6e151d),
	.w2(32'hbb71f899),
	.w3(32'hbb138be5),
	.w4(32'hb9c80358),
	.w5(32'h393c05c2),
	.w6(32'hbb8c4214),
	.w7(32'hbb81f852),
	.w8(32'h3c283e20),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd80dc3),
	.w1(32'h3bef9a6a),
	.w2(32'h3be6b8cb),
	.w3(32'hb9fe2c1c),
	.w4(32'h3b190eb4),
	.w5(32'hbac8da6c),
	.w6(32'h3c0c4b42),
	.w7(32'h3bb9c8ca),
	.w8(32'h3b13682c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eda378),
	.w1(32'h3b7e1d88),
	.w2(32'hbad41823),
	.w3(32'hbb0b2310),
	.w4(32'hbba775e5),
	.w5(32'hbb835c64),
	.w6(32'h3b03695e),
	.w7(32'h3b17bd0b),
	.w8(32'h3b33d9f1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e49634),
	.w1(32'h3b9826f9),
	.w2(32'hbad59681),
	.w3(32'hbacb23e7),
	.w4(32'hbbec0e3e),
	.w5(32'h3b2f5138),
	.w6(32'h3be64753),
	.w7(32'h3a7cfa71),
	.w8(32'h3b927b2b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdba32b),
	.w1(32'h3b715489),
	.w2(32'hba410f37),
	.w3(32'hb937a088),
	.w4(32'hbb6e019b),
	.w5(32'h3ab04ebb),
	.w6(32'h394a1cc8),
	.w7(32'hbb197d9f),
	.w8(32'h3bcd1092),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45e4b0),
	.w1(32'hbb82b511),
	.w2(32'hbb9147ff),
	.w3(32'h3b03dc9a),
	.w4(32'h3a2f30a4),
	.w5(32'hbb71959e),
	.w6(32'h3b5bde8e),
	.w7(32'hba9a3da6),
	.w8(32'hbb9b8133),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e8c06),
	.w1(32'hbc116796),
	.w2(32'hbc1f11af),
	.w3(32'hbb5c3110),
	.w4(32'h3a1e4da7),
	.w5(32'h3a4c77f5),
	.w6(32'hbc65388b),
	.w7(32'hbbd492b6),
	.w8(32'hbb86a80d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04fd09),
	.w1(32'h39bc94f7),
	.w2(32'h3b74ef8e),
	.w3(32'h3bb6bc6b),
	.w4(32'h3bcd4e77),
	.w5(32'h3bcc9308),
	.w6(32'hba27da60),
	.w7(32'h3c119651),
	.w8(32'h3b902545),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47e1c),
	.w1(32'hbbbfe9f1),
	.w2(32'h3ad0278b),
	.w3(32'h3b185ace),
	.w4(32'h3ba61c1f),
	.w5(32'h3b798412),
	.w6(32'hbaca93c2),
	.w7(32'h39d1d8bc),
	.w8(32'hba1cc9fe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f18fb),
	.w1(32'hbc10a69e),
	.w2(32'hbaadbe84),
	.w3(32'hba96c8fb),
	.w4(32'hbabc408c),
	.w5(32'h3b9c53a6),
	.w6(32'h3bcb8548),
	.w7(32'h3bbd2173),
	.w8(32'h3b0d666d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a164e),
	.w1(32'hbac49ea7),
	.w2(32'hbb59ce43),
	.w3(32'h3b7b7eef),
	.w4(32'hba41785d),
	.w5(32'h3ba1e759),
	.w6(32'h3ba6233f),
	.w7(32'h3b507199),
	.w8(32'h3b312257),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f79e9),
	.w1(32'hbbeb5b3f),
	.w2(32'hbb8ec14d),
	.w3(32'h3b761740),
	.w4(32'h3b750486),
	.w5(32'hba2d379e),
	.w6(32'h3b06f792),
	.w7(32'hba506547),
	.w8(32'hba8675c4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978d144),
	.w1(32'h38f2b165),
	.w2(32'hbbab0e7d),
	.w3(32'h3a83fdb2),
	.w4(32'hbbc165a2),
	.w5(32'h3c318d5e),
	.w6(32'h3bcefa4a),
	.w7(32'hbb71574e),
	.w8(32'h3b6cc270),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095d7a),
	.w1(32'hbc11daf3),
	.w2(32'hb9b45605),
	.w3(32'h3c0d9d3f),
	.w4(32'h3c48c328),
	.w5(32'hb9dcddc2),
	.w6(32'hbbff2ba8),
	.w7(32'h3b92b779),
	.w8(32'hbc1f694f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255e78),
	.w1(32'hbb1edca6),
	.w2(32'h3ab36187),
	.w3(32'h3a6ba2b6),
	.w4(32'hbb530630),
	.w5(32'hbbdf4013),
	.w6(32'hbb329f84),
	.w7(32'h3ac99b2b),
	.w8(32'h3b1bf9d3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba105d3),
	.w1(32'hbb22d694),
	.w2(32'hb817bc57),
	.w3(32'hbbf41df9),
	.w4(32'hbb37a92f),
	.w5(32'hbb8f7af2),
	.w6(32'h3b000592),
	.w7(32'hbb4bf1a2),
	.w8(32'hba171c88),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2fef8),
	.w1(32'hba1fccf0),
	.w2(32'hba64839f),
	.w3(32'hbc010d6a),
	.w4(32'hbba2001e),
	.w5(32'h3ba94326),
	.w6(32'hbb8a6290),
	.w7(32'hbb952478),
	.w8(32'h3abc7676),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d1d07),
	.w1(32'hbac9105d),
	.w2(32'h3b88da7c),
	.w3(32'hbb297cc6),
	.w4(32'hbbaf9128),
	.w5(32'h3b9efb7a),
	.w6(32'hbb1c7988),
	.w7(32'h3b44a6c9),
	.w8(32'h387d625d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88519d),
	.w1(32'hbbba3677),
	.w2(32'hbbb5cdcd),
	.w3(32'hbb588182),
	.w4(32'hbadcbd8d),
	.w5(32'h3b0e8611),
	.w6(32'hbb40ad44),
	.w7(32'hbb1f1ed7),
	.w8(32'h3b156e8a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e9241),
	.w1(32'h3aa01495),
	.w2(32'hba4debc6),
	.w3(32'hbaa538f6),
	.w4(32'hbb19687e),
	.w5(32'hbb8879ba),
	.w6(32'hbbb33de6),
	.w7(32'hbbb70d33),
	.w8(32'hbb865fb9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94131bd),
	.w1(32'h3c0225e3),
	.w2(32'h3c28689a),
	.w3(32'hbadb2404),
	.w4(32'h3ba37dd4),
	.w5(32'h3c3a2d4b),
	.w6(32'h3a9c13da),
	.w7(32'h3bc7c50c),
	.w8(32'h3c3b8855),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab5fa),
	.w1(32'h3abe0704),
	.w2(32'h3bc3543e),
	.w3(32'h3b918573),
	.w4(32'h3bcf10c5),
	.w5(32'h3c058098),
	.w6(32'h3b9dd57d),
	.w7(32'h3bfe8c7f),
	.w8(32'h3a43380b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a051d),
	.w1(32'hbb36e4c7),
	.w2(32'hbb9e8410),
	.w3(32'h3af3105f),
	.w4(32'hba481a33),
	.w5(32'hbb32ad2b),
	.w6(32'hbb8c0c50),
	.w7(32'hbba82ec5),
	.w8(32'hbb277161),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ab68),
	.w1(32'hbb60ae17),
	.w2(32'h39a85ad0),
	.w3(32'hbc16afea),
	.w4(32'hbba3b89c),
	.w5(32'hbac02603),
	.w6(32'hbb990c4d),
	.w7(32'hbaaf366f),
	.w8(32'h39723498),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe5380),
	.w1(32'h3a42c8cc),
	.w2(32'hbb49e20d),
	.w3(32'hbaa0f551),
	.w4(32'hb91edd9c),
	.w5(32'h3bd8eb31),
	.w6(32'hbb396948),
	.w7(32'hbbf0d666),
	.w8(32'hbc125d29),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50e979),
	.w1(32'hbc1cb6b3),
	.w2(32'hbb8ce6b6),
	.w3(32'h3b9cc17c),
	.w4(32'h3c7310eb),
	.w5(32'h3ad6c178),
	.w6(32'hbb5359df),
	.w7(32'h3bbe5b2b),
	.w8(32'hba83ef4b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbad84),
	.w1(32'hbb15e3cc),
	.w2(32'h3b9d7156),
	.w3(32'h3a14c5d7),
	.w4(32'h3bbff079),
	.w5(32'h38ba3c22),
	.w6(32'hbc029b38),
	.w7(32'h3bd6a7bb),
	.w8(32'hb9b007c6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e47ec),
	.w1(32'hbb97e34f),
	.w2(32'hbbb901e8),
	.w3(32'hbc166d23),
	.w4(32'hbbef00c2),
	.w5(32'h3b9feeac),
	.w6(32'hbc07e71a),
	.w7(32'hbc199f7e),
	.w8(32'hbbf02deb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93fc3e),
	.w1(32'hbbc31759),
	.w2(32'hbb994ba0),
	.w3(32'h3b5198cb),
	.w4(32'hbbd44023),
	.w5(32'h3b431293),
	.w6(32'hbc31d624),
	.w7(32'hbba424c4),
	.w8(32'hbba2f749),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf66e37),
	.w1(32'hbbc287b9),
	.w2(32'hbc19b494),
	.w3(32'h3b1abc4b),
	.w4(32'h3b6cf674),
	.w5(32'hb9c7f9a0),
	.w6(32'hbb228e3f),
	.w7(32'hbbacfc6a),
	.w8(32'h39dcfeb9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e34c5),
	.w1(32'h3aa46229),
	.w2(32'hb9bed81d),
	.w3(32'hb9fb2cd8),
	.w4(32'h3b2d6d46),
	.w5(32'hbbbca5dc),
	.w6(32'h3a87e4ff),
	.w7(32'h3b1180ed),
	.w8(32'h3b28ad87),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a39d5),
	.w1(32'h3a592cbe),
	.w2(32'hb796a2ce),
	.w3(32'hbbd262ab),
	.w4(32'hbb7f7844),
	.w5(32'h3b8497cb),
	.w6(32'h3b0d803f),
	.w7(32'h3b34263c),
	.w8(32'h3b9a4e32),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59db09),
	.w1(32'h3aa36526),
	.w2(32'hbadd995f),
	.w3(32'h399f3292),
	.w4(32'hbbe18b68),
	.w5(32'hba824e1d),
	.w6(32'h3adf3a66),
	.w7(32'hba4dfbe9),
	.w8(32'hbc48e9a3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9461),
	.w1(32'hbc16fca4),
	.w2(32'hbbe11fe3),
	.w3(32'h3b1e6926),
	.w4(32'hbb9ab423),
	.w5(32'h39ef351d),
	.w6(32'hbc795ce0),
	.w7(32'hbbd79af8),
	.w8(32'h3b51b62a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45bdad),
	.w1(32'hbac318d9),
	.w2(32'hbb8dc57c),
	.w3(32'hba77b3a5),
	.w4(32'hbabf43ff),
	.w5(32'hbba0f819),
	.w6(32'h3b29decd),
	.w7(32'hbb62320e),
	.w8(32'hbb4f0a9c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af49acb),
	.w1(32'hba6879a2),
	.w2(32'hbb9fbe22),
	.w3(32'hbb89bd7d),
	.w4(32'hbb890729),
	.w5(32'hbba8ea6a),
	.w6(32'hba66775a),
	.w7(32'hbb954250),
	.w8(32'hbc70028f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fd320),
	.w1(32'hbb85f235),
	.w2(32'hbb447ac8),
	.w3(32'h3aed4478),
	.w4(32'h3931eb12),
	.w5(32'hbb2acd27),
	.w6(32'hbc901d34),
	.w7(32'hbb4e0c71),
	.w8(32'hbc008363),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9fec),
	.w1(32'hbb73cc82),
	.w2(32'hbc01e3ec),
	.w3(32'hba2bd06d),
	.w4(32'hbaed7048),
	.w5(32'hbad44e09),
	.w6(32'hb793a09e),
	.w7(32'hbbaaab99),
	.w8(32'hbb4e96b1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22025c),
	.w1(32'hbba1fa4f),
	.w2(32'hbb92559a),
	.w3(32'hbb5c4292),
	.w4(32'h3b4cc145),
	.w5(32'hbaa2eb5c),
	.w6(32'hbb51051f),
	.w7(32'hbaff1789),
	.w8(32'h3a4701cc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e391e9),
	.w1(32'hbb6e4f60),
	.w2(32'hb95a2ae4),
	.w3(32'hbbb036a8),
	.w4(32'hba5e90d3),
	.w5(32'h3c890e52),
	.w6(32'hbb7fa6c3),
	.w7(32'hbae5bba9),
	.w8(32'h3c3fd6fc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1f5b1),
	.w1(32'h39ece91e),
	.w2(32'h3ba21c9d),
	.w3(32'h3c3f25d8),
	.w4(32'h3c36a268),
	.w5(32'h3c08caa3),
	.w6(32'h3b86849d),
	.w7(32'h3c398e3a),
	.w8(32'h3b89bc06),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc697b),
	.w1(32'hba578723),
	.w2(32'h3a903276),
	.w3(32'h3bdc87f4),
	.w4(32'h39e92b17),
	.w5(32'h3aa2b8f2),
	.w6(32'h3aa3f295),
	.w7(32'h3bf2fe27),
	.w8(32'h397dde1a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7b573),
	.w1(32'hbb8ec5af),
	.w2(32'hb8945cec),
	.w3(32'h3a192594),
	.w4(32'h3a8f91b0),
	.w5(32'hbb9ba930),
	.w6(32'hbc3cea8e),
	.w7(32'hbbd5677d),
	.w8(32'h3b52f52a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c387c3c),
	.w1(32'h3c0895ed),
	.w2(32'h3c3d6eb8),
	.w3(32'h3a38d21e),
	.w4(32'h3bc5c800),
	.w5(32'h3bf88376),
	.w6(32'h3b39df61),
	.w7(32'h3c27dd06),
	.w8(32'h3bc4c8a8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d9a19),
	.w1(32'h3ba36a60),
	.w2(32'h3bf33e9e),
	.w3(32'h3b623a7e),
	.w4(32'hbae4ef4c),
	.w5(32'h3a9b451e),
	.w6(32'h3c16c168),
	.w7(32'h3b1ed1ee),
	.w8(32'h3ae6a93b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffa10b),
	.w1(32'h3b63a932),
	.w2(32'hbbfe707a),
	.w3(32'h3b315d1b),
	.w4(32'hbab16619),
	.w5(32'h3a79e583),
	.w6(32'h37fbc16c),
	.w7(32'hbbac64a1),
	.w8(32'hbb97a186),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d3bd2),
	.w1(32'h3b56775e),
	.w2(32'h39cbb96a),
	.w3(32'h39569d38),
	.w4(32'h3a710aed),
	.w5(32'h3ba08ac2),
	.w6(32'h3ae0a6a9),
	.w7(32'h3b781b92),
	.w8(32'h3b420077),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4c6a7),
	.w1(32'h3b4e634c),
	.w2(32'hbaf4c916),
	.w3(32'h3ac45234),
	.w4(32'hbb50f902),
	.w5(32'hba74f462),
	.w6(32'hb9e082e1),
	.w7(32'hba77f52e),
	.w8(32'h3b91ebf8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b203085),
	.w1(32'h3b18f156),
	.w2(32'h3b3d5152),
	.w3(32'hba97520a),
	.w4(32'hbac2b776),
	.w5(32'hb9a5acd1),
	.w6(32'hba2bd7c6),
	.w7(32'h3a8bbb41),
	.w8(32'h3b3e8b12),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acacee9),
	.w1(32'h3b7e9fcb),
	.w2(32'hbab5d287),
	.w3(32'h3ad545f3),
	.w4(32'h3b2da6dd),
	.w5(32'h3bb67999),
	.w6(32'h37d02374),
	.w7(32'hb7ee8317),
	.w8(32'h3bde369a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c086e41),
	.w1(32'hbbbb76fd),
	.w2(32'h3c18c2b5),
	.w3(32'hbc4c5394),
	.w4(32'hbb3d611c),
	.w5(32'h3af69ca8),
	.w6(32'hbc020f42),
	.w7(32'h3bd32c28),
	.w8(32'hbba378c6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795406),
	.w1(32'hba5fc720),
	.w2(32'h3bd7f83d),
	.w3(32'h3b32e83a),
	.w4(32'hbae22272),
	.w5(32'h3abb9076),
	.w6(32'hbb2c69ca),
	.w7(32'h38911569),
	.w8(32'hb9e3b68c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18bd86),
	.w1(32'hbb2bc24d),
	.w2(32'h3b2cc856),
	.w3(32'hbbbb7e3c),
	.w4(32'h3abc03d3),
	.w5(32'h3b431be1),
	.w6(32'hbc16ec5e),
	.w7(32'hba942b55),
	.w8(32'h3b83a8b3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab62fcb),
	.w1(32'h3aadb226),
	.w2(32'hbb397f5f),
	.w3(32'h3baa4bf6),
	.w4(32'hbad6d603),
	.w5(32'h3b14546c),
	.w6(32'h3b8cfc48),
	.w7(32'hbbb7671a),
	.w8(32'hbaa47fb7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ccb7b),
	.w1(32'hbb38e260),
	.w2(32'hbafec168),
	.w3(32'hba7dd393),
	.w4(32'h3baf7081),
	.w5(32'h3bf3a26d),
	.w6(32'hbafa6da8),
	.w7(32'hbb5d5084),
	.w8(32'h3c0511b8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92b9a7),
	.w1(32'h3b981977),
	.w2(32'h3c2c13cc),
	.w3(32'hbac86525),
	.w4(32'hba3012ad),
	.w5(32'h3a9903f7),
	.w6(32'h3af507e3),
	.w7(32'h3c13f86a),
	.w8(32'hbbb77a42),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226988),
	.w1(32'hbb50b816),
	.w2(32'hbbbc2f99),
	.w3(32'hbbb52999),
	.w4(32'hbb6602f2),
	.w5(32'h39ddaf7b),
	.w6(32'hbbf60ab8),
	.w7(32'hbb756717),
	.w8(32'hba47c79f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babc7c9),
	.w1(32'hbadc19cb),
	.w2(32'hbbc39c82),
	.w3(32'h3876a294),
	.w4(32'hba3d5f74),
	.w5(32'hbbb66b9d),
	.w6(32'hbb7f0af8),
	.w7(32'hbc093557),
	.w8(32'hbbb022dd),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2961b2),
	.w1(32'hbc2c3c5b),
	.w2(32'hbc3a8c32),
	.w3(32'h3be8e87e),
	.w4(32'h3ba72ebd),
	.w5(32'hba4a3455),
	.w6(32'h3c4c8f79),
	.w7(32'h3a8b5bd2),
	.w8(32'hbae446de),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e517a),
	.w1(32'hbaa6d1f9),
	.w2(32'hbb95a5c3),
	.w3(32'h3ab03350),
	.w4(32'hbae8ca4a),
	.w5(32'h3ab33b2c),
	.w6(32'h39eb14bd),
	.w7(32'hbb7652bc),
	.w8(32'hbb1b198e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b3f67),
	.w1(32'hbb850738),
	.w2(32'hb9d17fc9),
	.w3(32'h3b8657a5),
	.w4(32'h3bd37ee8),
	.w5(32'h391ac29f),
	.w6(32'h3a9cb81e),
	.w7(32'h3b1530c6),
	.w8(32'hbc3ef377),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18a5f1),
	.w1(32'hbc162660),
	.w2(32'hb9d7dd37),
	.w3(32'hbb1e56f5),
	.w4(32'h3bee4997),
	.w5(32'h3b5441f5),
	.w6(32'hbc734d02),
	.w7(32'h396d7508),
	.w8(32'h3b813ff6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a985d),
	.w1(32'hbb654471),
	.w2(32'h3ae54dd1),
	.w3(32'hbb75d286),
	.w4(32'hba9bff21),
	.w5(32'h39a24f46),
	.w6(32'hbb149a8f),
	.w7(32'hbaf92cef),
	.w8(32'hb945c952),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8969a1),
	.w1(32'h3bcc499a),
	.w2(32'hbb13ae5d),
	.w3(32'h3b9ca8cc),
	.w4(32'hba134b9f),
	.w5(32'hbb99c482),
	.w6(32'h3a9ef268),
	.w7(32'hbbb1bea6),
	.w8(32'hba81b2af),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0485eb),
	.w1(32'h39a4f3f8),
	.w2(32'hbb021939),
	.w3(32'hbbd2abe6),
	.w4(32'hbbe570f2),
	.w5(32'h3981a342),
	.w6(32'h39f46e1f),
	.w7(32'hb99a701e),
	.w8(32'h3bc5fa67),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a38bd),
	.w1(32'hbb991ebe),
	.w2(32'hba09a82b),
	.w3(32'h3ac13ce3),
	.w4(32'h3b8ed737),
	.w5(32'hbb26ef2b),
	.w6(32'h3aa16f39),
	.w7(32'hbae7f648),
	.w8(32'hbb2efd2a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91f54),
	.w1(32'hbb2c4177),
	.w2(32'hbbacd163),
	.w3(32'h3a31d7b6),
	.w4(32'h3b9c9a9f),
	.w5(32'hbaf05b71),
	.w6(32'hbbbde5d1),
	.w7(32'hbb37f86d),
	.w8(32'hb9f29afc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0232eb),
	.w1(32'hba074a4d),
	.w2(32'hba6478cb),
	.w3(32'hb9d31fec),
	.w4(32'hbb87c1fe),
	.w5(32'h3be7c454),
	.w6(32'h39749150),
	.w7(32'h39683245),
	.w8(32'hbb330a0d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba785aec),
	.w1(32'hbb08ca28),
	.w2(32'hbb15c2cb),
	.w3(32'h3b150983),
	.w4(32'hbbfabb4d),
	.w5(32'h3b726b69),
	.w6(32'hb94310ba),
	.w7(32'h3ad4a8ec),
	.w8(32'h3b5a8b6c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb753b1a),
	.w1(32'h3a297af4),
	.w2(32'hba3ae41d),
	.w3(32'h3af5e065),
	.w4(32'hbaa75c79),
	.w5(32'h3ab0c507),
	.w6(32'h3bebee9e),
	.w7(32'h3a189dbf),
	.w8(32'h3b33f71a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f91d8b),
	.w1(32'h3bacf422),
	.w2(32'h39b9d888),
	.w3(32'h3b8e88da),
	.w4(32'h3a06eb65),
	.w5(32'h3bd5df24),
	.w6(32'hbb473453),
	.w7(32'hbb2ceccc),
	.w8(32'h3c4e9738),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfedf3d),
	.w1(32'hba262519),
	.w2(32'h3bad0640),
	.w3(32'hbb4a3c6b),
	.w4(32'h3ae5a88e),
	.w5(32'hbbe8561e),
	.w6(32'hbb5cad7d),
	.w7(32'h3b4ddf69),
	.w8(32'h3c5ca624),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf03e2f),
	.w1(32'h3c27f7c1),
	.w2(32'hbb92e88c),
	.w3(32'h39bce752),
	.w4(32'hbba78f86),
	.w5(32'hbba2a3ea),
	.w6(32'h3cd9033e),
	.w7(32'h3c53e040),
	.w8(32'hbc1f485c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab427a3),
	.w1(32'hbb005aa9),
	.w2(32'h3aa11dc6),
	.w3(32'h3bf5f74d),
	.w4(32'h3b978466),
	.w5(32'h3b941846),
	.w6(32'hb95b06f0),
	.w7(32'h3aac735d),
	.w8(32'h3b3cae87),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978028),
	.w1(32'hbad13f25),
	.w2(32'hbb901043),
	.w3(32'h3b4e69c4),
	.w4(32'h3afa002c),
	.w5(32'h3c1f5018),
	.w6(32'h3b96512e),
	.w7(32'hbac845ef),
	.w8(32'h3a5b1f3a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23138a),
	.w1(32'h3a710819),
	.w2(32'h3b208cb3),
	.w3(32'h3c15b9a1),
	.w4(32'h3beb35bb),
	.w5(32'hbab71265),
	.w6(32'h3acba77c),
	.w7(32'h3b34852b),
	.w8(32'hbb14bf20),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa30c21),
	.w1(32'hbb77352d),
	.w2(32'hbbbe5ed9),
	.w3(32'hbae7c73b),
	.w4(32'hbb9ca18a),
	.w5(32'hb95a77cb),
	.w6(32'hbbb307ed),
	.w7(32'hbb891736),
	.w8(32'hb9d86e68),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b362ada),
	.w1(32'h3b048fdc),
	.w2(32'h39dc1f0f),
	.w3(32'h3ada3c6d),
	.w4(32'hbb6a8196),
	.w5(32'h38fa64c0),
	.w6(32'hb9eced74),
	.w7(32'h3b9857d2),
	.w8(32'h3bc68cef),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb049732),
	.w1(32'hba5e4afc),
	.w2(32'hbb25a60c),
	.w3(32'h3ac0ca81),
	.w4(32'hba94bb36),
	.w5(32'h3acdfee5),
	.w6(32'h3bce6f67),
	.w7(32'hb9b94024),
	.w8(32'h3ae5fb0b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec03a0),
	.w1(32'hbbe83cc5),
	.w2(32'hba959781),
	.w3(32'h39805aee),
	.w4(32'h3bb31f25),
	.w5(32'hbb2588e4),
	.w6(32'h3b537a39),
	.w7(32'h3a89d18e),
	.w8(32'hbbeb0172),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e44a),
	.w1(32'hbb85fa8a),
	.w2(32'hba40c9e3),
	.w3(32'hbb9046b6),
	.w4(32'h39ba4353),
	.w5(32'hbb1cf2e5),
	.w6(32'hbbf24a54),
	.w7(32'hbb15f64a),
	.w8(32'hbb80d176),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96e4ac),
	.w1(32'hba603c78),
	.w2(32'hba922602),
	.w3(32'hba50fcb9),
	.w4(32'hbc282ba3),
	.w5(32'h3ab6f8da),
	.w6(32'hbbcab9be),
	.w7(32'hbb7ef6ce),
	.w8(32'hbb51c87a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1c40),
	.w1(32'hbb1ec922),
	.w2(32'hbbb69b2e),
	.w3(32'hbb028e30),
	.w4(32'hbb16ab0f),
	.w5(32'hbb58d627),
	.w6(32'hbad37d75),
	.w7(32'hbbcc3ba1),
	.w8(32'h3a6e0770),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41a620),
	.w1(32'h3b493273),
	.w2(32'h3b6798a4),
	.w3(32'hbb9b7d77),
	.w4(32'h3a1b61c2),
	.w5(32'hbbda3e7d),
	.w6(32'hb8f24edc),
	.w7(32'h3ba0c448),
	.w8(32'hbc509f83),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b702),
	.w1(32'hbc3a32a3),
	.w2(32'hba91d0ea),
	.w3(32'hbb800f27),
	.w4(32'hba44bdb3),
	.w5(32'hba8fb14a),
	.w6(32'hbc5439e8),
	.w7(32'hbc0e9524),
	.w8(32'h3b8ce0ce),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c759),
	.w1(32'hbbe842f0),
	.w2(32'h3b88a22f),
	.w3(32'hbb329035),
	.w4(32'h3b3e8d7e),
	.w5(32'hba209cd3),
	.w6(32'hb94f3ed5),
	.w7(32'h399c3cb8),
	.w8(32'h39a4030e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11dcc1),
	.w1(32'h3b88c7f9),
	.w2(32'hb9ec1bab),
	.w3(32'h3a290c3d),
	.w4(32'h39a35bb2),
	.w5(32'h3c15d74d),
	.w6(32'hb997962b),
	.w7(32'hbaf23507),
	.w8(32'h3ba4cbaa),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3feda9),
	.w1(32'hbbbc4970),
	.w2(32'h3aaa2894),
	.w3(32'h3a8f0030),
	.w4(32'h3b7e2d2e),
	.w5(32'h3ba002dd),
	.w6(32'h399d1bb2),
	.w7(32'h3b871aba),
	.w8(32'hbb48bcfe),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a3bb),
	.w1(32'hbb14e992),
	.w2(32'h3b106ed2),
	.w3(32'h3bdc0119),
	.w4(32'h3c2cf06d),
	.w5(32'hb82c8790),
	.w6(32'h3b576a8d),
	.w7(32'h3becc641),
	.w8(32'h3bce4e3a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da1c18),
	.w1(32'h38843580),
	.w2(32'h3a4694a3),
	.w3(32'hba826a7c),
	.w4(32'h3b1bfba5),
	.w5(32'hbaa13397),
	.w6(32'h3b1cc38a),
	.w7(32'h3ab251ea),
	.w8(32'h395328b1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cca211),
	.w1(32'h3a27ebf0),
	.w2(32'hba8d4d94),
	.w3(32'hbb992bee),
	.w4(32'hbbc5b211),
	.w5(32'h3ad40371),
	.w6(32'hbb570002),
	.w7(32'hbbc6a398),
	.w8(32'hbb1dcc80),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcbf3f),
	.w1(32'hba7e9b3d),
	.w2(32'h3bd7d01b),
	.w3(32'hbb40bdac),
	.w4(32'hba5793cd),
	.w5(32'h3c14cc37),
	.w6(32'hbb6e8597),
	.w7(32'h39c0e42c),
	.w8(32'h3a1da487),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30160c),
	.w1(32'hbbddf644),
	.w2(32'hbbe32fea),
	.w3(32'h3b2ee210),
	.w4(32'h3b7df997),
	.w5(32'hbbedadf7),
	.w6(32'hbafd106b),
	.w7(32'hbb87b7c7),
	.w8(32'hbc21af48),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc265671),
	.w1(32'h3902ad32),
	.w2(32'h3b45dfcd),
	.w3(32'hb99c264b),
	.w4(32'hb9ec0936),
	.w5(32'hb7dbe384),
	.w6(32'h3adbc318),
	.w7(32'h3b65a0a3),
	.w8(32'hbbb28338),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a9fb0),
	.w1(32'h3ab2a4c8),
	.w2(32'h3b7a9443),
	.w3(32'h3a427fe7),
	.w4(32'h3b22b124),
	.w5(32'hbaff8514),
	.w6(32'hbb4045f4),
	.w7(32'h3b1615f4),
	.w8(32'h39429344),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a1407),
	.w1(32'h3aa90ed0),
	.w2(32'h3b3c1577),
	.w3(32'h3aabd9b8),
	.w4(32'hbb11199d),
	.w5(32'hbc063509),
	.w6(32'hbb85e8d2),
	.w7(32'hbb6a0a60),
	.w8(32'hbbd7338a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb982999),
	.w1(32'hbb713b0f),
	.w2(32'hbbd07f7d),
	.w3(32'hbb1d38a9),
	.w4(32'hbba967f8),
	.w5(32'hbb8ac217),
	.w6(32'h39bb9572),
	.w7(32'hbbcf176f),
	.w8(32'hba8eb0d2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5115e),
	.w1(32'hbb35f814),
	.w2(32'hbbbc6c27),
	.w3(32'hba21d325),
	.w4(32'hbb029a87),
	.w5(32'hba92ed60),
	.w6(32'h3b1170fb),
	.w7(32'hbb4ffff3),
	.w8(32'h3a795d2e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53595f),
	.w1(32'hbb4190c3),
	.w2(32'hbb700e63),
	.w3(32'h3ab3afd6),
	.w4(32'h3aeaf16f),
	.w5(32'hb9ef4b12),
	.w6(32'h3b9f7db9),
	.w7(32'h3bb5478d),
	.w8(32'hbb3519ca),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077e13),
	.w1(32'h3b918481),
	.w2(32'hbb94f420),
	.w3(32'h3b2c0651),
	.w4(32'h3bed3458),
	.w5(32'h3ba1a797),
	.w6(32'hbb630be1),
	.w7(32'hbb048f08),
	.w8(32'h3acdb601),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9642871),
	.w1(32'h3a0db8d4),
	.w2(32'h3ab5b826),
	.w3(32'h3b8cb872),
	.w4(32'h3b273e11),
	.w5(32'h3bc02bb8),
	.w6(32'h3bd8dadc),
	.w7(32'h3be4b1af),
	.w8(32'h3b9923e4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacdab5),
	.w1(32'hba5f22c2),
	.w2(32'hbab8f103),
	.w3(32'hba04cd5d),
	.w4(32'hba265df2),
	.w5(32'hbc0dd0f7),
	.w6(32'h3b0deb27),
	.w7(32'hba0af898),
	.w8(32'hbc285d56),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd058ad),
	.w1(32'hbb804b07),
	.w2(32'hba5167ae),
	.w3(32'h3a13d569),
	.w4(32'h3c1edf1b),
	.w5(32'h399884ac),
	.w6(32'hbc351479),
	.w7(32'hbafc2104),
	.w8(32'hbc206ccb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1a1d1),
	.w1(32'hbc52152d),
	.w2(32'hbbef6965),
	.w3(32'hba449c5e),
	.w4(32'h3ad6a831),
	.w5(32'hbc0e5d9d),
	.w6(32'hbb6c159f),
	.w7(32'h3ae5ec57),
	.w8(32'hbbc38f64),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be62948),
	.w1(32'h3ba23099),
	.w2(32'hba2fec9c),
	.w3(32'h3b5de36b),
	.w4(32'hbbbb900b),
	.w5(32'h3bbec9f6),
	.w6(32'h3adc6fa8),
	.w7(32'hbbddf3b9),
	.w8(32'hbb5329dc),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b774696),
	.w1(32'hb99261fd),
	.w2(32'h3c144dda),
	.w3(32'hbba7d356),
	.w4(32'hbbb18767),
	.w5(32'hbb876b13),
	.w6(32'hbc381c60),
	.w7(32'hbbb5e462),
	.w8(32'h3c0593b3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f5e1),
	.w1(32'h3ba181c1),
	.w2(32'h3b4929c0),
	.w3(32'hbaef045c),
	.w4(32'hbbbdd570),
	.w5(32'h3c31762c),
	.w6(32'h3bceb83f),
	.w7(32'h3ba4ad6a),
	.w8(32'h3c2a3d06),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc86876),
	.w1(32'hbbeaa259),
	.w2(32'h3b930424),
	.w3(32'hbacf702d),
	.w4(32'h3b587f67),
	.w5(32'h3aeced0d),
	.w6(32'hbc3b50bb),
	.w7(32'h3b22cfde),
	.w8(32'h3befb1bb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c010f),
	.w1(32'hbb5b7fba),
	.w2(32'h3b445942),
	.w3(32'hbc15a24c),
	.w4(32'hbb274a8a),
	.w5(32'h3b13e550),
	.w6(32'hba4b227d),
	.w7(32'h3b75f6b1),
	.w8(32'h3b27adbb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e7c85),
	.w1(32'h3b4d352d),
	.w2(32'hb9246947),
	.w3(32'h3aa3aa80),
	.w4(32'hbbb203f4),
	.w5(32'hbae3783b),
	.w6(32'h3c1bde0b),
	.w7(32'hbaf962dd),
	.w8(32'h3ac3150d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bc168),
	.w1(32'h3c355938),
	.w2(32'h38ab7d8c),
	.w3(32'h3bd3f6ef),
	.w4(32'h3b3eb08e),
	.w5(32'h3aed3285),
	.w6(32'h3b2ee7df),
	.w7(32'hbb057e50),
	.w8(32'h3ae5b4fa),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad14d28),
	.w1(32'h39eb832a),
	.w2(32'hb94a42b7),
	.w3(32'h3b0e2d7a),
	.w4(32'h3a400e24),
	.w5(32'hba809fa8),
	.w6(32'h3a8d218e),
	.w7(32'hb995b02e),
	.w8(32'hba3e8e31),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac43fae),
	.w1(32'hbab6bab4),
	.w2(32'hbab41ba4),
	.w3(32'hba5a334c),
	.w4(32'hba9d509f),
	.w5(32'hbaa4cd71),
	.w6(32'hba8d2bed),
	.w7(32'hba20221b),
	.w8(32'h3a2575a3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af5b9b),
	.w1(32'hb9b42e31),
	.w2(32'h3a2b9dfd),
	.w3(32'hbad1437b),
	.w4(32'hb90c3a36),
	.w5(32'h3b1d7630),
	.w6(32'h3abd86e6),
	.w7(32'h3a494277),
	.w8(32'h3b044fbe),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac52fbb),
	.w1(32'h3b1a297e),
	.w2(32'h3b14d64d),
	.w3(32'h3ae9a153),
	.w4(32'h3aacb69d),
	.w5(32'h37f4ff97),
	.w6(32'h3aa1aa42),
	.w7(32'h3b0b37a4),
	.w8(32'hb9e22a11),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7791f2),
	.w1(32'h3b738d01),
	.w2(32'h3adfe3b9),
	.w3(32'h3b2b6b5d),
	.w4(32'h3aa5eaa7),
	.w5(32'hbabb3210),
	.w6(32'h3bc74236),
	.w7(32'hb7bf778c),
	.w8(32'hbb9f78d7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39138054),
	.w1(32'hbaf457b1),
	.w2(32'hbbd6ba19),
	.w3(32'hba523e72),
	.w4(32'hbb93ec3d),
	.w5(32'hbaadaac2),
	.w6(32'hbb37ca4c),
	.w7(32'hbba2ae8f),
	.w8(32'h39254908),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368e96),
	.w1(32'h3b193b98),
	.w2(32'h3b75a9a2),
	.w3(32'h3af6725f),
	.w4(32'h3b1451cb),
	.w5(32'hba808347),
	.w6(32'h3b7a80a3),
	.w7(32'h3b96a797),
	.w8(32'hbb33a2d0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b59f8),
	.w1(32'hbae05ad5),
	.w2(32'hbb858034),
	.w3(32'h3aa9a8f2),
	.w4(32'hbac498d4),
	.w5(32'hbae9192f),
	.w6(32'h3a8b6ab7),
	.w7(32'hbb287296),
	.w8(32'hbb2b3586),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade7303),
	.w1(32'hba6452b6),
	.w2(32'h3a38ef0d),
	.w3(32'h3a963164),
	.w4(32'hba71befb),
	.w5(32'h3aa20e4e),
	.w6(32'h3b804d26),
	.w7(32'hba21e83c),
	.w8(32'h3afa856b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0344df),
	.w1(32'h3a8fdc45),
	.w2(32'h3a467a6d),
	.w3(32'h3ae179a3),
	.w4(32'h3ac31ad3),
	.w5(32'h3acae8cb),
	.w6(32'h3b3116e1),
	.w7(32'h3ac1142a),
	.w8(32'h3abb245b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c64f65),
	.w1(32'hba597744),
	.w2(32'h36d307e0),
	.w3(32'h3aea6c33),
	.w4(32'h3a6f0340),
	.w5(32'h3a470130),
	.w6(32'hba2eaa46),
	.w7(32'h39ec636c),
	.w8(32'h3b164172),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a860dcc),
	.w1(32'hb789e92e),
	.w2(32'hba3a2989),
	.w3(32'h3b1444cf),
	.w4(32'h3a8633c5),
	.w5(32'hbae4846b),
	.w6(32'h3b119840),
	.w7(32'h3974b688),
	.w8(32'hb9d0b3d0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38520528),
	.w1(32'hb96fdd73),
	.w2(32'h3a01bfd8),
	.w3(32'hba639c44),
	.w4(32'h3a0119b4),
	.w5(32'h3a264e74),
	.w6(32'hba4761a5),
	.w7(32'h380826f8),
	.w8(32'h3abfff6d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a02b0),
	.w1(32'hbb1b63d7),
	.w2(32'hbbfc2d27),
	.w3(32'h3a9f0e0d),
	.w4(32'hbad76c79),
	.w5(32'hbb42aeae),
	.w6(32'h3b0384a5),
	.w7(32'hbb6f6b2d),
	.w8(32'hbb7f02dd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b1a53),
	.w1(32'hba1fc19b),
	.w2(32'hbb1d12cd),
	.w3(32'hb9c93416),
	.w4(32'hba8c82e9),
	.w5(32'hbb353d7d),
	.w6(32'h37e4093a),
	.w7(32'hbac0e295),
	.w8(32'hbbcd5131),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1870c4),
	.w1(32'hba87ac0e),
	.w2(32'hbb6bf3d6),
	.w3(32'h3b0bfe93),
	.w4(32'h3a5d5fad),
	.w5(32'hbae06cbd),
	.w6(32'hba442d36),
	.w7(32'hbb393a73),
	.w8(32'hbbb3cec4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20bbac),
	.w1(32'h39fa77cb),
	.w2(32'hb9a3b436),
	.w3(32'h3aa38a39),
	.w4(32'h3b127df8),
	.w5(32'hb9f8e2a6),
	.w6(32'h3b23e5be),
	.w7(32'h3a8250ad),
	.w8(32'h3a3c5645),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b49f80),
	.w1(32'h3a2c2b58),
	.w2(32'hba8f31e3),
	.w3(32'h3a348c78),
	.w4(32'hbaa6d37a),
	.w5(32'h3abc70ee),
	.w6(32'h3b5657b6),
	.w7(32'h383c5407),
	.w8(32'h3aaab653),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063d59),
	.w1(32'h3aac0385),
	.w2(32'h3ac71610),
	.w3(32'h39d180a2),
	.w4(32'h3a9c2fbe),
	.w5(32'hbaabd5f9),
	.w6(32'hba0e291d),
	.w7(32'h3a642b98),
	.w8(32'hba3538b9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa424f8),
	.w1(32'hba68ac5d),
	.w2(32'h391354ce),
	.w3(32'hba6553ae),
	.w4(32'hba6af294),
	.w5(32'h3a11260c),
	.w6(32'h39e77cc0),
	.w7(32'h3a3dd16f),
	.w8(32'hb9b92e38),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac50634),
	.w1(32'hbb1093d3),
	.w2(32'hbaf6ef1e),
	.w3(32'h3a3230ce),
	.w4(32'h3a269dd0),
	.w5(32'h37a64a34),
	.w6(32'hba719787),
	.w7(32'hba8a11a9),
	.w8(32'hba8e879c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9abb66),
	.w1(32'h3af3c05e),
	.w2(32'h3aa94ac6),
	.w3(32'h3ad246e3),
	.w4(32'h3ac408d9),
	.w5(32'h3b0ba760),
	.w6(32'h3b042148),
	.w7(32'h3b56fa06),
	.w8(32'hba35d842),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02059b),
	.w1(32'h3a3a2acd),
	.w2(32'hb92d6345),
	.w3(32'h393e49d7),
	.w4(32'hb808cb60),
	.w5(32'hb974ae7f),
	.w6(32'h3a74b734),
	.w7(32'h390fe9d0),
	.w8(32'hb917dc67),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba2e6c),
	.w1(32'hb9410236),
	.w2(32'h3a97ac55),
	.w3(32'hbaac6aeb),
	.w4(32'h3902cf7c),
	.w5(32'hba89dce7),
	.w6(32'hba4c76e1),
	.w7(32'h3ac1d1ab),
	.w8(32'hba54ce27),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5e3d2),
	.w1(32'hba91d63a),
	.w2(32'hbae2ec6f),
	.w3(32'hbab9a6f6),
	.w4(32'hba801bad),
	.w5(32'hba8c07a6),
	.w6(32'hb9bf8d2e),
	.w7(32'hbaab4e90),
	.w8(32'hbadc2db3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba4c7c),
	.w1(32'hbb0ec890),
	.w2(32'hbae599b1),
	.w3(32'hba9b7df0),
	.w4(32'hba704e25),
	.w5(32'hbab01a8f),
	.w6(32'hbb35d8e3),
	.w7(32'hbb084ad0),
	.w8(32'hbaad0552),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad52526),
	.w1(32'hb9f67b96),
	.w2(32'hbb2fac6a),
	.w3(32'hbb1b7e5f),
	.w4(32'hba7a431a),
	.w5(32'hb9fe0482),
	.w6(32'h394c9d53),
	.w7(32'hba9c88d9),
	.w8(32'hbafcf5dd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad11225),
	.w1(32'hbb17ccad),
	.w2(32'hbbd86282),
	.w3(32'h3b242d50),
	.w4(32'hba36e22c),
	.w5(32'hba3c4be9),
	.w6(32'hba46a2d4),
	.w7(32'hbb6ec926),
	.w8(32'hbb0eac3d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2942bb),
	.w1(32'hb911c4e4),
	.w2(32'hb9160bca),
	.w3(32'h3b1fc593),
	.w4(32'h3a9d732c),
	.w5(32'h39906355),
	.w6(32'h3ad87546),
	.w7(32'h3a682264),
	.w8(32'hba0d9f19),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73b23c),
	.w1(32'h3ac7cad0),
	.w2(32'hb93437d9),
	.w3(32'h3aa9fd44),
	.w4(32'h39079539),
	.w5(32'hb9a03950),
	.w6(32'h3b2814ff),
	.w7(32'h3b01e937),
	.w8(32'h3b7fa182),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule