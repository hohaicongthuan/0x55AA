module layer_10_featuremap_445(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2928a),
	.w1(32'h3a201f9c),
	.w2(32'h3b70da44),
	.w3(32'h3b0c38fe),
	.w4(32'h3b100e59),
	.w5(32'h3c181d62),
	.w6(32'h3b15ce70),
	.w7(32'h3b0c6afb),
	.w8(32'h3c0e6e07),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57cae8),
	.w1(32'hbc383337),
	.w2(32'hbbceb71a),
	.w3(32'h3c08216d),
	.w4(32'hbbd9e44c),
	.w5(32'hbc012aab),
	.w6(32'h3bb04b00),
	.w7(32'hbc729b87),
	.w8(32'hbc31db27),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e1d4),
	.w1(32'hbc0a1c17),
	.w2(32'hbcb9c5aa),
	.w3(32'h3b4fae7d),
	.w4(32'hb9128d94),
	.w5(32'h3d1f757a),
	.w6(32'hbbb1376e),
	.w7(32'hbbd95708),
	.w8(32'hbc880163),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62dcbd),
	.w1(32'hbb482ebe),
	.w2(32'hb960db4f),
	.w3(32'h3b5c0cbd),
	.w4(32'h3bf73c3f),
	.w5(32'h3c8f8d31),
	.w6(32'hbc00b7b4),
	.w7(32'hbc16650a),
	.w8(32'hbc011977),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf32013),
	.w1(32'h3bae440c),
	.w2(32'h3b6dc279),
	.w3(32'h3c43aa0c),
	.w4(32'h3acd76a7),
	.w5(32'h3c2858d7),
	.w6(32'h3bb4495f),
	.w7(32'hbb8ebccb),
	.w8(32'hbbcea1c7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b751c61),
	.w1(32'h3b7da4e3),
	.w2(32'h3bb86d89),
	.w3(32'h3b5b338c),
	.w4(32'hbb69571e),
	.w5(32'h3913147f),
	.w6(32'h3a48e0e7),
	.w7(32'h3b36598b),
	.w8(32'h3abdd990),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d6eb),
	.w1(32'hbb501729),
	.w2(32'h3b8068c5),
	.w3(32'hbb2e6715),
	.w4(32'h3a3b17ae),
	.w5(32'hbc10d8d3),
	.w6(32'hba665e98),
	.w7(32'h39c35d7a),
	.w8(32'h3c4979e1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09a874),
	.w1(32'h3bc37fb1),
	.w2(32'h3c688406),
	.w3(32'hbae1c4ee),
	.w4(32'h3bdefe2f),
	.w5(32'h3ba0ccd9),
	.w6(32'h3c0dde4b),
	.w7(32'hbc383446),
	.w8(32'hbc17e632),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba529bc8),
	.w1(32'hbc0d014b),
	.w2(32'hbbdbfe3a),
	.w3(32'hbb865f32),
	.w4(32'h3a6e7ab0),
	.w5(32'hbc10684c),
	.w6(32'hbbd9bb44),
	.w7(32'hbc7a765e),
	.w8(32'hbc38bd6f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015dbe),
	.w1(32'h3b460d73),
	.w2(32'hbbab76a2),
	.w3(32'hb9e3084e),
	.w4(32'h3b9ac2e5),
	.w5(32'h3cb54a83),
	.w6(32'hbae5d328),
	.w7(32'h3bad46d4),
	.w8(32'hbb9edf00),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa320e5),
	.w1(32'h3b956e9c),
	.w2(32'h3b418484),
	.w3(32'hbb15e851),
	.w4(32'hbc0f9da3),
	.w5(32'h3c2528ad),
	.w6(32'h3b2fefd2),
	.w7(32'hba333953),
	.w8(32'hbba89c5f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6abd6c),
	.w1(32'h3a893a09),
	.w2(32'h392bc0ef),
	.w3(32'hbaa63b39),
	.w4(32'h3b7dbf96),
	.w5(32'h3b79821f),
	.w6(32'hbb92d074),
	.w7(32'h3b8e38b3),
	.w8(32'h3bbb163e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64495),
	.w1(32'hba9a5f97),
	.w2(32'hbb9d7fee),
	.w3(32'h3aebaf4b),
	.w4(32'h3adbdf43),
	.w5(32'h3b8b3c87),
	.w6(32'h3bd41474),
	.w7(32'hbb60ef08),
	.w8(32'hbb828759),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3349),
	.w1(32'h3b9e4e84),
	.w2(32'h39d1f80d),
	.w3(32'hbb8c46ce),
	.w4(32'h3a9a9f6b),
	.w5(32'h3c309253),
	.w6(32'h3a75d29a),
	.w7(32'h3a1e947e),
	.w8(32'h3aa39ffa),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88d348),
	.w1(32'hba5f5f4c),
	.w2(32'hbbac94be),
	.w3(32'hbb13574d),
	.w4(32'hbb17c65e),
	.w5(32'h3c7812e2),
	.w6(32'h3a0826fc),
	.w7(32'h3b26dfd8),
	.w8(32'hbc5002e5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763bb3),
	.w1(32'hbbefc07b),
	.w2(32'hbbe3e116),
	.w3(32'h3beafc93),
	.w4(32'hbabf3276),
	.w5(32'h3a138be4),
	.w6(32'hba8aa595),
	.w7(32'h3b429425),
	.w8(32'hbad554eb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe39634),
	.w1(32'h3ab0273e),
	.w2(32'hbb3e2eb6),
	.w3(32'h3a58390b),
	.w4(32'h3a504ee6),
	.w5(32'hbab67d97),
	.w6(32'h3a62c6a5),
	.w7(32'hba11a535),
	.w8(32'hbb7d3a39),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cee5),
	.w1(32'h3b94c4c7),
	.w2(32'h3af50c1a),
	.w3(32'hbad707d3),
	.w4(32'hbb1c31dc),
	.w5(32'h3a4ccb8a),
	.w6(32'hbb5732d0),
	.w7(32'hb95f730e),
	.w8(32'hb98f33c4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b689a98),
	.w1(32'hbb8ba408),
	.w2(32'hbbb52bd5),
	.w3(32'hbb97d9e4),
	.w4(32'hbb99f9a8),
	.w5(32'hbb0e94e1),
	.w6(32'h3b136544),
	.w7(32'hbb0372c2),
	.w8(32'hbbb04b7b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72f6f0),
	.w1(32'h3c157009),
	.w2(32'h3a2a02f6),
	.w3(32'h3a95aecd),
	.w4(32'hb51f04f9),
	.w5(32'hbb5663c5),
	.w6(32'hbbd13954),
	.w7(32'h3b075362),
	.w8(32'h3b66120b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd015),
	.w1(32'h3b618794),
	.w2(32'h3adb1e1a),
	.w3(32'hbb6067da),
	.w4(32'h3b393e80),
	.w5(32'h3b95d868),
	.w6(32'hbbb63904),
	.w7(32'h3af3b3e0),
	.w8(32'h3a1a42f5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0efd5a),
	.w1(32'h3bda1d6c),
	.w2(32'h3bcf0d8c),
	.w3(32'h39b21adf),
	.w4(32'h3b60907f),
	.w5(32'h3bdeca63),
	.w6(32'h3a9f137c),
	.w7(32'h3c0e36b4),
	.w8(32'hbb25c0b0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c01f7),
	.w1(32'hbb960b9f),
	.w2(32'hbbd24b76),
	.w3(32'h3af4af40),
	.w4(32'hbb9e9f6c),
	.w5(32'hbc236311),
	.w6(32'hb9232df6),
	.w7(32'h3aaac1b3),
	.w8(32'hbb243698),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa9015),
	.w1(32'h3ae0f483),
	.w2(32'hbba46acd),
	.w3(32'hbc0d3607),
	.w4(32'h3b3f5e4f),
	.w5(32'hba473a80),
	.w6(32'hbc102c37),
	.w7(32'h3b3b0e98),
	.w8(32'hbb1e600f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4acb08),
	.w1(32'h3ba58192),
	.w2(32'h3981aa5f),
	.w3(32'hbb478343),
	.w4(32'h3b86419f),
	.w5(32'h3b5b355a),
	.w6(32'hbb084f79),
	.w7(32'h3a98658c),
	.w8(32'h3ae7c6a2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f860),
	.w1(32'hb982e993),
	.w2(32'h3b9cea70),
	.w3(32'h3b339afc),
	.w4(32'h3bfc9a5d),
	.w5(32'h3b20c83f),
	.w6(32'h3b4ab30e),
	.w7(32'h3b1d9583),
	.w8(32'hba94cce2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b702a8e),
	.w1(32'h3ae1a850),
	.w2(32'h3bd378fb),
	.w3(32'h3b5a0dab),
	.w4(32'h3c2ff50c),
	.w5(32'h3baa90b8),
	.w6(32'h3a9ef974),
	.w7(32'h3bbe5538),
	.w8(32'h3c09a319),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf85715),
	.w1(32'h3ad1b511),
	.w2(32'hba1290a6),
	.w3(32'hbbf09714),
	.w4(32'hba39ff9a),
	.w5(32'hbb52db64),
	.w6(32'h3c0cbcba),
	.w7(32'hbade2382),
	.w8(32'hbb5bf1b6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63afab),
	.w1(32'hbc03d993),
	.w2(32'hbc6325ba),
	.w3(32'hbba0edac),
	.w4(32'hbba442f3),
	.w5(32'hbbbccd92),
	.w6(32'hbbb5497a),
	.w7(32'hbbde72ed),
	.w8(32'hbb42bd75),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4b08),
	.w1(32'h3afe1f15),
	.w2(32'h3b952305),
	.w3(32'hb98bdc82),
	.w4(32'hbb9403c3),
	.w5(32'h3b201604),
	.w6(32'h3b1d000f),
	.w7(32'hbae83322),
	.w8(32'h3ade8da1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a76d3),
	.w1(32'h3bc5b32c),
	.w2(32'hbb53bcbb),
	.w3(32'h3ad90f1a),
	.w4(32'h39e281b7),
	.w5(32'hbba6a739),
	.w6(32'h3b6028ce),
	.w7(32'hbb914ad3),
	.w8(32'hbafee374),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af11dff),
	.w1(32'h3b5fd3c6),
	.w2(32'h3b572b0d),
	.w3(32'h39251f73),
	.w4(32'hbbabd99a),
	.w5(32'h3b15856d),
	.w6(32'h3bbcfd8a),
	.w7(32'hbaf13e5d),
	.w8(32'hbb448223),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a58f),
	.w1(32'h3c0f59f9),
	.w2(32'h3c99291d),
	.w3(32'hba2dabd5),
	.w4(32'h3bd65839),
	.w5(32'hbbdaad63),
	.w6(32'hbbaa17bb),
	.w7(32'h3c197987),
	.w8(32'h3c82dbb2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25fd93),
	.w1(32'hbb244c20),
	.w2(32'h3c543f4d),
	.w3(32'hba2bc070),
	.w4(32'hbbe3bf79),
	.w5(32'hbc6f21a1),
	.w6(32'h3bede4f9),
	.w7(32'h3c42f823),
	.w8(32'h3cd20da7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb790903f),
	.w1(32'h3b28ea96),
	.w2(32'h3bf90950),
	.w3(32'h3a272f61),
	.w4(32'hbbf75920),
	.w5(32'hbc9c5f6f),
	.w6(32'h3bfb1a79),
	.w7(32'h39d2c58b),
	.w8(32'h3c64841f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf60b5),
	.w1(32'hb99cfc73),
	.w2(32'hbb8eb248),
	.w3(32'hbb8f0895),
	.w4(32'h3b5b338e),
	.w5(32'h3ba0f8ff),
	.w6(32'h3b4228b0),
	.w7(32'hbabfb295),
	.w8(32'hbbd6ff22),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc327a),
	.w1(32'h3c448890),
	.w2(32'hbb14bf19),
	.w3(32'hba2b6892),
	.w4(32'h3b89b913),
	.w5(32'hbab833d4),
	.w6(32'hbb5c5684),
	.w7(32'h3be82150),
	.w8(32'h3ad980fa),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399186aa),
	.w1(32'h3bc722cb),
	.w2(32'h3c5765a8),
	.w3(32'h39b84a9d),
	.w4(32'h3af6e7d8),
	.w5(32'hbc5c6d09),
	.w6(32'h3b0475aa),
	.w7(32'hbaa46371),
	.w8(32'h3bb34675),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f29a),
	.w1(32'h3b6dc051),
	.w2(32'hbb9c46f9),
	.w3(32'hbbb2c290),
	.w4(32'hbbbac00f),
	.w5(32'h3a3eb969),
	.w6(32'h3ba47ba0),
	.w7(32'hba144d6c),
	.w8(32'hbb05dd31),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6499cf),
	.w1(32'h3bd1ba93),
	.w2(32'h3be34ed3),
	.w3(32'h3bf76174),
	.w4(32'h3ace3879),
	.w5(32'hbc111254),
	.w6(32'h394b3353),
	.w7(32'hbb2f90ee),
	.w8(32'h3b3ef5fd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f65c5),
	.w1(32'h3c6670b7),
	.w2(32'h3c7dafd4),
	.w3(32'hbb8cc396),
	.w4(32'hbba785e2),
	.w5(32'hbc6b4a65),
	.w6(32'hbb40b229),
	.w7(32'hbbb74f22),
	.w8(32'hbbc087e0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e4efb),
	.w1(32'hba95162b),
	.w2(32'h3ab91c49),
	.w3(32'hba273e92),
	.w4(32'hbbe2ee45),
	.w5(32'hbc89f0c3),
	.w6(32'hbbcd84f3),
	.w7(32'hbb4c3ae2),
	.w8(32'hbc1beafd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050ed2),
	.w1(32'h3ae92f38),
	.w2(32'hbb5e27eb),
	.w3(32'hbad8faee),
	.w4(32'hbba7b9e9),
	.w5(32'h3b6202e3),
	.w6(32'hbb907f12),
	.w7(32'h3a0ad93b),
	.w8(32'h3af84450),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac289),
	.w1(32'h3bb49a72),
	.w2(32'h3c46f161),
	.w3(32'h3b6e1719),
	.w4(32'h3bae59eb),
	.w5(32'h3ba0a956),
	.w6(32'h3b1cf94f),
	.w7(32'h3b778ff8),
	.w8(32'h3bf8ab9b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdcabd),
	.w1(32'h3bad45fa),
	.w2(32'h3ac4a741),
	.w3(32'h3c217015),
	.w4(32'h3a153e5f),
	.w5(32'hbb4863d2),
	.w6(32'h3c19d81d),
	.w7(32'hb6396f73),
	.w8(32'hba795382),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53272),
	.w1(32'hbc41616a),
	.w2(32'hbc7b2d4d),
	.w3(32'hba964bb4),
	.w4(32'h3a8eafe6),
	.w5(32'hbafe8faf),
	.w6(32'hbbbdec61),
	.w7(32'h3b216a1d),
	.w8(32'hbb10de23),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1db13),
	.w1(32'hbbd0b2a0),
	.w2(32'hbc5d30e2),
	.w3(32'hbb56394e),
	.w4(32'hba663ecc),
	.w5(32'h3d1d1f39),
	.w6(32'h3ba6435e),
	.w7(32'hbc1571b7),
	.w8(32'hbc8939e9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67c6bb),
	.w1(32'hbb96cf1d),
	.w2(32'h3a48893e),
	.w3(32'h3c216658),
	.w4(32'hbc014b36),
	.w5(32'hbc2c7729),
	.w6(32'hbbd5a2e5),
	.w7(32'hbb13da5a),
	.w8(32'hbba991be),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a149418),
	.w1(32'hbbd87c7d),
	.w2(32'hbbd80e65),
	.w3(32'hbae1d6e4),
	.w4(32'hb98e1edd),
	.w5(32'hba012b18),
	.w6(32'hbad5e031),
	.w7(32'hbb78e5db),
	.w8(32'hbbd3c79a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be285),
	.w1(32'h3b9a5188),
	.w2(32'hbb9c342f),
	.w3(32'hbb8a4a8d),
	.w4(32'hbbd24533),
	.w5(32'h3be6935a),
	.w6(32'hbc1f5b3e),
	.w7(32'hbb81c7c9),
	.w8(32'hbba02fe3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd463ee),
	.w1(32'hbb770c86),
	.w2(32'h3a99c350),
	.w3(32'h3bb176c7),
	.w4(32'h3afe9a7a),
	.w5(32'hbacb295d),
	.w6(32'hbb8c710f),
	.w7(32'h3aac7b96),
	.w8(32'h3ba95fbe),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fbde7),
	.w1(32'h3b30f7f0),
	.w2(32'hbb50bd58),
	.w3(32'h3b9ecad8),
	.w4(32'h3ba6fc23),
	.w5(32'h3a63f56b),
	.w6(32'h3afb0b26),
	.w7(32'hbaaeaab0),
	.w8(32'hbaa68b50),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d3f68),
	.w1(32'hbba308aa),
	.w2(32'hb910d905),
	.w3(32'hbbd577c5),
	.w4(32'hbbced5ab),
	.w5(32'hbc990c7c),
	.w6(32'h3a99811e),
	.w7(32'h3b41062f),
	.w8(32'h3c822592),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911342),
	.w1(32'hbbc987ad),
	.w2(32'h3aeff430),
	.w3(32'hbc1ed3de),
	.w4(32'hbc236d71),
	.w5(32'hbd055656),
	.w6(32'h3bd44c3b),
	.w7(32'h3c0fab69),
	.w8(32'h3ccfef38),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf052),
	.w1(32'h3b1f3793),
	.w2(32'h3adc2cf3),
	.w3(32'hbcbfa439),
	.w4(32'h39b5b796),
	.w5(32'hbc1eb88b),
	.w6(32'h3b240b83),
	.w7(32'h3b89ad1d),
	.w8(32'h3b87c637),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0192a3),
	.w1(32'h396c2308),
	.w2(32'hb98a0dab),
	.w3(32'hbbac422f),
	.w4(32'h3b805827),
	.w5(32'hbc98c6b8),
	.w6(32'h3b8b845c),
	.w7(32'hbaf54587),
	.w8(32'h3ba2aab8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3850ca),
	.w1(32'h3b57f80b),
	.w2(32'h3be31d84),
	.w3(32'h3ac3c716),
	.w4(32'h39f2e6d3),
	.w5(32'h3baf2717),
	.w6(32'h3b174c41),
	.w7(32'h3a844f81),
	.w8(32'h3bd25810),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10bc6c),
	.w1(32'h3b1ccb5e),
	.w2(32'hbbb0b1cc),
	.w3(32'h3b1d2d64),
	.w4(32'h3ba2f485),
	.w5(32'hbb90e82a),
	.w6(32'h3b62677c),
	.w7(32'h39d3f8d8),
	.w8(32'hbb74b6ee),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ed6d),
	.w1(32'h3b1eeab6),
	.w2(32'h3b96f9ee),
	.w3(32'hbb39f54b),
	.w4(32'h3b066b72),
	.w5(32'hba6b3b0c),
	.w6(32'h3ac639fb),
	.w7(32'hbbf4c78e),
	.w8(32'h38da7504),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb33c8),
	.w1(32'hbb6c4571),
	.w2(32'hbba9a69a),
	.w3(32'h3aa3bdaf),
	.w4(32'h3ba1c4de),
	.w5(32'h3b3d5c4d),
	.w6(32'hb9fdbe15),
	.w7(32'h39e425de),
	.w8(32'hbb96a3d2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee2729),
	.w1(32'hb99397fb),
	.w2(32'hbbe0705f),
	.w3(32'hbb03c08d),
	.w4(32'h3bc0a669),
	.w5(32'h3bfcaa1f),
	.w6(32'hbb57197f),
	.w7(32'h3b4d9773),
	.w8(32'h3a7f44d1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ec32),
	.w1(32'hbb81e440),
	.w2(32'hbb2e5dd1),
	.w3(32'h3b796ee1),
	.w4(32'hba1418de),
	.w5(32'h3b8a2a53),
	.w6(32'h3b257a39),
	.w7(32'h3a85d35f),
	.w8(32'hbbed4ce4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1583f),
	.w1(32'h3a31e985),
	.w2(32'h3aeaa947),
	.w3(32'h3be6e18b),
	.w4(32'h3b67a5cd),
	.w5(32'hbbbbe40a),
	.w6(32'hbb8307ca),
	.w7(32'h3ac63987),
	.w8(32'h3ab1e7e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0791a),
	.w1(32'h3b014ff4),
	.w2(32'h3b536271),
	.w3(32'hbc092ba8),
	.w4(32'hba8f8ca2),
	.w5(32'h3a4b90e1),
	.w6(32'hba890475),
	.w7(32'h3bcd22a5),
	.w8(32'h3bfebeb6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d347a),
	.w1(32'h3c493075),
	.w2(32'h3c72b79a),
	.w3(32'hbbbee147),
	.w4(32'h3bc8746a),
	.w5(32'h3ba1448c),
	.w6(32'h3b3b3aba),
	.w7(32'h3ac304fa),
	.w8(32'hb927bd33),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fcfcb),
	.w1(32'h3b9baf64),
	.w2(32'hbb4fb0b0),
	.w3(32'h3be69e8d),
	.w4(32'h3bb26a07),
	.w5(32'hbbd140b4),
	.w6(32'hb83bf3e5),
	.w7(32'h3ad4b9de),
	.w8(32'hbb6aafa9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a47e),
	.w1(32'hbc117ba3),
	.w2(32'hbbb31e99),
	.w3(32'hbaa67f19),
	.w4(32'h3b64f6d5),
	.w5(32'h3ba23789),
	.w6(32'hbbeb6dc2),
	.w7(32'h3b6f98ed),
	.w8(32'h3b850fa1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb379185),
	.w1(32'hbbe8589a),
	.w2(32'hbc2f7a83),
	.w3(32'h3bc3e830),
	.w4(32'hbc1656cf),
	.w5(32'hba678b2a),
	.w6(32'h3b918673),
	.w7(32'hbadc250b),
	.w8(32'hbb611742),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6fd6),
	.w1(32'hbbbec765),
	.w2(32'hbaba2847),
	.w3(32'hbb9dac03),
	.w4(32'h3881d441),
	.w5(32'hbb666783),
	.w6(32'hba6b8f49),
	.w7(32'hbb63e1ce),
	.w8(32'hbbac7e34),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11fa52),
	.w1(32'hbb5080d4),
	.w2(32'hbc07da64),
	.w3(32'h3ab91410),
	.w4(32'hba974648),
	.w5(32'hbab7c67f),
	.w6(32'hbb92e1fb),
	.w7(32'hba045750),
	.w8(32'h3b5752fe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16bedc),
	.w1(32'h39f051d1),
	.w2(32'h3b051c43),
	.w3(32'hbb0374c2),
	.w4(32'hb9a5abf3),
	.w5(32'h3b006335),
	.w6(32'hbad079dc),
	.w7(32'hbade2211),
	.w8(32'hbb97ad25),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985b1ca),
	.w1(32'hba6880c5),
	.w2(32'hbb1283ee),
	.w3(32'h39fd5e50),
	.w4(32'hbbdc4c6e),
	.w5(32'h39f30c60),
	.w6(32'hbbb5d333),
	.w7(32'h3c13d41f),
	.w8(32'h3c0abdc3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0513b6),
	.w1(32'h39e1e914),
	.w2(32'hba0a6db2),
	.w3(32'h3aa11043),
	.w4(32'hbb331115),
	.w5(32'hbafd55d1),
	.w6(32'h3c344423),
	.w7(32'h3b0738d0),
	.w8(32'h3b7e567e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50b5bb),
	.w1(32'hba41e9c0),
	.w2(32'h3b73d683),
	.w3(32'hbb21e073),
	.w4(32'h3c60c326),
	.w5(32'h3d068430),
	.w6(32'h3a823b0a),
	.w7(32'h37147981),
	.w8(32'h3aa5b0be),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c208cb4),
	.w1(32'h3b9fc057),
	.w2(32'h3c1c7f96),
	.w3(32'h3c674046),
	.w4(32'hbadbff88),
	.w5(32'hbb4eca56),
	.w6(32'hbb0158db),
	.w7(32'h3b8dcbe9),
	.w8(32'h3b8f91e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbd28e),
	.w1(32'h38f52922),
	.w2(32'hbb6079d9),
	.w3(32'hbafdce4a),
	.w4(32'hbb816d28),
	.w5(32'h3be069da),
	.w6(32'h3bb770f9),
	.w7(32'hba8032f4),
	.w8(32'h3a831459),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fff0f),
	.w1(32'hb9b5cd20),
	.w2(32'h3a5460a7),
	.w3(32'hb9d08705),
	.w4(32'hbb6837dc),
	.w5(32'hbb86099c),
	.w6(32'h3ab3998f),
	.w7(32'hbbfcd0ab),
	.w8(32'hbb9c19eb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2895ab),
	.w1(32'h3b8b0d3a),
	.w2(32'hbaf82d97),
	.w3(32'hbb67b4af),
	.w4(32'hbb4be197),
	.w5(32'h39c936e6),
	.w6(32'hbb30b446),
	.w7(32'hbb0a8408),
	.w8(32'hbba827e4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b164b19),
	.w1(32'hbb57b585),
	.w2(32'hbb0112f5),
	.w3(32'h3b914c9c),
	.w4(32'hbb6668ce),
	.w5(32'hbb4b9880),
	.w6(32'hba989a76),
	.w7(32'h3beeaf4d),
	.w8(32'h3b753b49),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b163299),
	.w1(32'hbb8a4ca4),
	.w2(32'hbb8d6666),
	.w3(32'h38ccb275),
	.w4(32'h39cd5094),
	.w5(32'hb9a39671),
	.w6(32'h3b3df8aa),
	.w7(32'h3931d431),
	.w8(32'hbba3c76b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7907b3),
	.w1(32'h3b11cc83),
	.w2(32'hbb1f616e),
	.w3(32'hbb0d5f54),
	.w4(32'h3a3b386c),
	.w5(32'hbb6b9955),
	.w6(32'hbb13945f),
	.w7(32'h3b159181),
	.w8(32'h3be907c0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e813e),
	.w1(32'hbba379b6),
	.w2(32'hbb33dcf5),
	.w3(32'h39fa4166),
	.w4(32'hbba0ab6a),
	.w5(32'hbb8b404c),
	.w6(32'h3bbddc15),
	.w7(32'hbb4aa357),
	.w8(32'hbb2c94f0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82f6c0),
	.w1(32'hb9b68267),
	.w2(32'hbbc70d24),
	.w3(32'hbbe1d1a3),
	.w4(32'hbc5d5854),
	.w5(32'hbc71706b),
	.w6(32'hbb4912c4),
	.w7(32'h3b3dbd5d),
	.w8(32'h3ba06e31),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa5433),
	.w1(32'hba595380),
	.w2(32'hbb3a1c45),
	.w3(32'hbc00f691),
	.w4(32'h380da578),
	.w5(32'h3a0bb829),
	.w6(32'h3c268915),
	.w7(32'hb9876b8b),
	.w8(32'h3aa73c7f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9849),
	.w1(32'hbb541d9b),
	.w2(32'h3bde727b),
	.w3(32'hba44b9a5),
	.w4(32'hba908ac6),
	.w5(32'h3b158106),
	.w6(32'hb993541b),
	.w7(32'h3bc68d8b),
	.w8(32'h3c464d47),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842a91),
	.w1(32'hbbe7cea4),
	.w2(32'hbb46e6b9),
	.w3(32'hbb19d9a4),
	.w4(32'h3ac1d82e),
	.w5(32'hba8cadf8),
	.w6(32'h3bd00c06),
	.w7(32'h3ae3c268),
	.w8(32'hba0b38a0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc8bdb),
	.w1(32'hba5e9087),
	.w2(32'h3ab6361f),
	.w3(32'hbb3c35b9),
	.w4(32'hba1d241a),
	.w5(32'hbb3249d1),
	.w6(32'hba3bd357),
	.w7(32'hbb741350),
	.w8(32'hbb8cbcf4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f756),
	.w1(32'hba58d27c),
	.w2(32'h3b34f1c2),
	.w3(32'hbbbec5b6),
	.w4(32'hbbdacff5),
	.w5(32'hbacb3d5a),
	.w6(32'hbb6eb1af),
	.w7(32'hbc1788a0),
	.w8(32'hbb537ba3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75d517),
	.w1(32'h3a87031c),
	.w2(32'h3b26d529),
	.w3(32'hbb710d8b),
	.w4(32'hbbc4dd89),
	.w5(32'hbbde2fe5),
	.w6(32'hbb2f5ae8),
	.w7(32'hbaeff97c),
	.w8(32'hbae65917),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc892c),
	.w1(32'hbb08c679),
	.w2(32'hbb003b08),
	.w3(32'hbadd7fc1),
	.w4(32'hbb51c517),
	.w5(32'hbc0b8fb6),
	.w6(32'h3a01a843),
	.w7(32'hbb0e279f),
	.w8(32'hbb76538d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb415fc8),
	.w1(32'h3b2a99b2),
	.w2(32'h3bb9f4f3),
	.w3(32'hbbc8f8a5),
	.w4(32'hbad9cec3),
	.w5(32'h3b6b4f51),
	.w6(32'hbb9c5d6c),
	.w7(32'hbbda3cf2),
	.w8(32'hbafe85fc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7df440),
	.w1(32'hbb508b67),
	.w2(32'hbab4fd32),
	.w3(32'hba9d4bbc),
	.w4(32'h3b6a7e99),
	.w5(32'hbbdcf036),
	.w6(32'hbb96231a),
	.w7(32'hbb85c749),
	.w8(32'hbb24d623),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990348),
	.w1(32'hbbb3187b),
	.w2(32'hbb6c8449),
	.w3(32'hb981831f),
	.w4(32'hbbb89a66),
	.w5(32'hbc04e7cb),
	.w6(32'hb9ea7d70),
	.w7(32'h3b497b9e),
	.w8(32'h3a6d8491),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0dfb),
	.w1(32'h3b3ead94),
	.w2(32'h3b93a351),
	.w3(32'hbb1e3c21),
	.w4(32'h3c354cf4),
	.w5(32'h3c613a94),
	.w6(32'h3bee6ab4),
	.w7(32'h3b4b93be),
	.w8(32'h3be1d38e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72eeb),
	.w1(32'hbbb8f4c7),
	.w2(32'hbbfc488b),
	.w3(32'h3c260869),
	.w4(32'h3ba4c08d),
	.w5(32'hbab013dc),
	.w6(32'h3aae87fa),
	.w7(32'h3af10f22),
	.w8(32'hbb9e4837),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb634f93),
	.w1(32'h3b0accc5),
	.w2(32'h3b8c15ed),
	.w3(32'hb9b80c5f),
	.w4(32'h3bc37a76),
	.w5(32'h3c0244a4),
	.w6(32'h3a9cdbd3),
	.w7(32'hb961303e),
	.w8(32'hbbfb6f35),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c105899),
	.w1(32'hbab69e45),
	.w2(32'hba0979b4),
	.w3(32'h39abc869),
	.w4(32'h3ad64a10),
	.w5(32'h3c85f708),
	.w6(32'hbc02067c),
	.w7(32'h3ab2d936),
	.w8(32'hb78b4b69),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3a7f6),
	.w1(32'hb9f89d5f),
	.w2(32'hbb3e3268),
	.w3(32'h3b8610c1),
	.w4(32'h3b84d5ab),
	.w5(32'hba63208b),
	.w6(32'hba5aad38),
	.w7(32'h3bc9c687),
	.w8(32'h3bd0a46c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad497b4),
	.w1(32'hbb9eb169),
	.w2(32'hbbd40513),
	.w3(32'h3ab8cf4a),
	.w4(32'hba846cd9),
	.w5(32'hbbc7fdc8),
	.w6(32'h3b2cba1b),
	.w7(32'h3b843eb2),
	.w8(32'h3b8d3fb0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b81d3),
	.w1(32'h396fb3f8),
	.w2(32'hbb3ac5ea),
	.w3(32'hbbeb0b42),
	.w4(32'h3bb7edf5),
	.w5(32'h3bc5ce02),
	.w6(32'h3b308cdd),
	.w7(32'h3bbc443f),
	.w8(32'h3a3e06c1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb060844),
	.w1(32'h3a9bafa2),
	.w2(32'hbb430483),
	.w3(32'h3b06e2a8),
	.w4(32'h3c7826cd),
	.w5(32'h3cec9199),
	.w6(32'h3916a90e),
	.w7(32'h3bdeb8d2),
	.w8(32'h3bba8fbf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f039a),
	.w1(32'hbbb21a12),
	.w2(32'h3b9db4a5),
	.w3(32'h3c8e020a),
	.w4(32'hba5910d2),
	.w5(32'h39d472f6),
	.w6(32'h3afa9168),
	.w7(32'hba78db8e),
	.w8(32'hbafc9853),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08c986),
	.w1(32'h3c7db7dd),
	.w2(32'h3c14922f),
	.w3(32'h3aa67237),
	.w4(32'hbbc9bd18),
	.w5(32'hb8305431),
	.w6(32'h3a7a90ef),
	.w7(32'h3be1604d),
	.w8(32'h3b6f7147),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be83952),
	.w1(32'h3ab3f0cf),
	.w2(32'h3c7bde02),
	.w3(32'h3a7c3236),
	.w4(32'h3b4cd1df),
	.w5(32'h3af40299),
	.w6(32'h3bef1841),
	.w7(32'h3c32a971),
	.w8(32'h3aa7f143),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cdf8e),
	.w1(32'h3b97210f),
	.w2(32'h3bcf06e3),
	.w3(32'h371d9da2),
	.w4(32'h3b56ea2e),
	.w5(32'h38aff581),
	.w6(32'hbb91f9ff),
	.w7(32'hb99cd6be),
	.w8(32'hbbd234bd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9006fb),
	.w1(32'hba11159e),
	.w2(32'h3ade4e19),
	.w3(32'hbba26914),
	.w4(32'h3b96adf1),
	.w5(32'h3bf82d86),
	.w6(32'hbb451c1a),
	.w7(32'h3bb32343),
	.w8(32'h3bd45482),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48eada),
	.w1(32'hbb7a447c),
	.w2(32'hbc1a4bdb),
	.w3(32'h3a60a65e),
	.w4(32'hbb463742),
	.w5(32'hbb85f22c),
	.w6(32'h3a8b5df5),
	.w7(32'hbb7a50b1),
	.w8(32'h3abadc1f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7f6ea),
	.w1(32'h3b3c7dbd),
	.w2(32'hbb8cf28a),
	.w3(32'h3b42c357),
	.w4(32'h3b170404),
	.w5(32'hba60b580),
	.w6(32'h3bea9886),
	.w7(32'h3c02fa54),
	.w8(32'h3bf5a116),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92215f),
	.w1(32'h3ac91a87),
	.w2(32'h3b4ebb6c),
	.w3(32'hba2738e6),
	.w4(32'hbbad4128),
	.w5(32'hbb82f4fa),
	.w6(32'h3ac0e234),
	.w7(32'hb9613649),
	.w8(32'h39005641),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52d3bf),
	.w1(32'h3a869d25),
	.w2(32'h3bbc3cae),
	.w3(32'hbbb91573),
	.w4(32'hbabbe4cd),
	.w5(32'hbb153d3a),
	.w6(32'h3b3a44e1),
	.w7(32'hbc32f1d4),
	.w8(32'hbc7d0321),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38698c44),
	.w1(32'hbb525a2a),
	.w2(32'h3b0408b8),
	.w3(32'hba9f32a6),
	.w4(32'hbaeab049),
	.w5(32'hba7ec651),
	.w6(32'hbb8a1200),
	.w7(32'h3a352d33),
	.w8(32'h3b8d877a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38513f),
	.w1(32'hbb562733),
	.w2(32'hbb602218),
	.w3(32'hbab10429),
	.w4(32'h3a03244a),
	.w5(32'h3b44ac74),
	.w6(32'hba50632a),
	.w7(32'h3aeb6ebe),
	.w8(32'h38aa3ea4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b026dd8),
	.w1(32'hba4047a1),
	.w2(32'hba462901),
	.w3(32'hbad41d4d),
	.w4(32'hb8b34528),
	.w5(32'h3b414eef),
	.w6(32'hbbb10d00),
	.w7(32'hbb86fb52),
	.w8(32'hbb8f0306),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c3881),
	.w1(32'hba9004be),
	.w2(32'hbbc2792d),
	.w3(32'hba389771),
	.w4(32'h3aca960a),
	.w5(32'h3c7d5626),
	.w6(32'hbbc45440),
	.w7(32'hbc458268),
	.w8(32'hbc60e47d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0387a),
	.w1(32'hbb430f92),
	.w2(32'hbb875c48),
	.w3(32'h3af06bf8),
	.w4(32'hbbf57dc6),
	.w5(32'hbad1fc2d),
	.w6(32'hbc97b272),
	.w7(32'hbb340ea4),
	.w8(32'hbaf39a7c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d00e1),
	.w1(32'h3b1c359b),
	.w2(32'h3a549bca),
	.w3(32'h3b2a9532),
	.w4(32'h3ae189c8),
	.w5(32'hbad54c37),
	.w6(32'h3aaf2d83),
	.w7(32'h3adc71b9),
	.w8(32'hba7d3d29),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897d805),
	.w1(32'hbb3ba4f2),
	.w2(32'hbbea15b5),
	.w3(32'hbbbe2524),
	.w4(32'hbaaa5aec),
	.w5(32'hbb271050),
	.w6(32'hbbb5c0ab),
	.w7(32'hbb805acf),
	.w8(32'hbb933e74),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b31cb),
	.w1(32'hbaad9408),
	.w2(32'h3ab8975f),
	.w3(32'hbab43bcf),
	.w4(32'h3c28ff93),
	.w5(32'h3c5323bd),
	.w6(32'hbae9e32b),
	.w7(32'h3a87f2af),
	.w8(32'h3b9b4780),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8b54),
	.w1(32'h3bf52da3),
	.w2(32'h3bcc403e),
	.w3(32'h3b999851),
	.w4(32'h3ba2e217),
	.w5(32'h3c15b58f),
	.w6(32'h3b9c424f),
	.w7(32'hbbab5fcf),
	.w8(32'hbbbde54c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb237a),
	.w1(32'h3c4be1f2),
	.w2(32'h3b2e6a85),
	.w3(32'h3b813f44),
	.w4(32'h3b42ab5f),
	.w5(32'h39de8ac6),
	.w6(32'hbbb6fc6d),
	.w7(32'hbb0c1032),
	.w8(32'h3b4e288a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe0e00),
	.w1(32'h3bcd5b50),
	.w2(32'h3ba62f43),
	.w3(32'h3bd18dfd),
	.w4(32'h3afb7954),
	.w5(32'h395ca6f6),
	.w6(32'h3c179363),
	.w7(32'hbaa9ac8f),
	.w8(32'h3ab5139f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5af8),
	.w1(32'h3a1cc927),
	.w2(32'hba945ace),
	.w3(32'hb9cab35d),
	.w4(32'hbb935028),
	.w5(32'hb9509c73),
	.w6(32'hba314d5c),
	.w7(32'h3b563623),
	.w8(32'hba9533d2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce74a0),
	.w1(32'h3b26d51c),
	.w2(32'hbaa3cdb9),
	.w3(32'hbb8541ca),
	.w4(32'hbba7e5e4),
	.w5(32'hbbbc99af),
	.w6(32'hbac55ca5),
	.w7(32'hbb57b191),
	.w8(32'hbb96bb0c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba52b1),
	.w1(32'hba9eaa42),
	.w2(32'hbb180a1d),
	.w3(32'hbb4d4772),
	.w4(32'h3beecfd2),
	.w5(32'hba6bf3ae),
	.w6(32'hbb2b30c0),
	.w7(32'h3b038718),
	.w8(32'hbba733d9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39950ce8),
	.w1(32'hbb53ef51),
	.w2(32'hbb34f961),
	.w3(32'hbaf85bfd),
	.w4(32'hbb9b080d),
	.w5(32'hbb723549),
	.w6(32'hbbae2416),
	.w7(32'hbbe04e53),
	.w8(32'hbc13af6f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7cce0),
	.w1(32'h3b7cf1e8),
	.w2(32'h3c345cee),
	.w3(32'hbbd06bf4),
	.w4(32'h3ba46e6a),
	.w5(32'h3c82a86e),
	.w6(32'hbbb2f696),
	.w7(32'hbb3b4184),
	.w8(32'hbc0fc9ef),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f9b2),
	.w1(32'h3b855f26),
	.w2(32'h391729f0),
	.w3(32'h3abe756c),
	.w4(32'h3bb40c6e),
	.w5(32'h3bd23755),
	.w6(32'hbc1edb6a),
	.w7(32'h3be11ee4),
	.w8(32'h3b9e2197),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021ce0),
	.w1(32'hbb2ae749),
	.w2(32'hbb6e8ec5),
	.w3(32'h3bdb85b2),
	.w4(32'hbc2809b3),
	.w5(32'hbc1b60a5),
	.w6(32'h3bcad1cd),
	.w7(32'hbb711cab),
	.w8(32'hba642136),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb47bef),
	.w1(32'h3b91864e),
	.w2(32'h3b6a4d2e),
	.w3(32'hbbc4f4e8),
	.w4(32'h3ad852d0),
	.w5(32'hbb65561c),
	.w6(32'h3ad4e317),
	.w7(32'hba38b230),
	.w8(32'hbb173a2e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b150dff),
	.w1(32'h3c15c4b1),
	.w2(32'h3c36b7f1),
	.w3(32'hb9d54816),
	.w4(32'h3ad7ffb9),
	.w5(32'h3b2c0d6f),
	.w6(32'h3b13a80f),
	.w7(32'hbaad9942),
	.w8(32'hbbd9c0b9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c232c6d),
	.w1(32'h3c2bd854),
	.w2(32'h3b0f14f7),
	.w3(32'h3b2e08c6),
	.w4(32'h3cb0fc2e),
	.w5(32'h3cf5d92c),
	.w6(32'hbba9fd34),
	.w7(32'h3963aea6),
	.w8(32'h3b0bcd40),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f833),
	.w1(32'hbbc46b0d),
	.w2(32'hbbccbb9a),
	.w3(32'h3c807640),
	.w4(32'hbbd8a168),
	.w5(32'hba4c422e),
	.w6(32'h3b4299b7),
	.w7(32'h3b6547cc),
	.w8(32'hb9cd44c0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bcd84),
	.w1(32'h3ae79883),
	.w2(32'h3bbb7c11),
	.w3(32'hbb292d5d),
	.w4(32'h3a4264fd),
	.w5(32'hbaf38a6a),
	.w6(32'hbbbccc4f),
	.w7(32'h3b298f25),
	.w8(32'hbad9bd07),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9621d2),
	.w1(32'hbc1be69f),
	.w2(32'hbbd3d1f9),
	.w3(32'hba3180eb),
	.w4(32'hbb16b6d7),
	.w5(32'hbbca46ab),
	.w6(32'h3a4dd949),
	.w7(32'hbb319791),
	.w8(32'hba711f3b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad86ea6),
	.w1(32'hbb00d4fc),
	.w2(32'hbc2fc764),
	.w3(32'hbb79f407),
	.w4(32'hbba01d5e),
	.w5(32'h3a3965ed),
	.w6(32'h39e9681c),
	.w7(32'hbc3cf84b),
	.w8(32'hbc55b187),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadff93b),
	.w1(32'h3be26cf3),
	.w2(32'h3c286d06),
	.w3(32'hbb970c43),
	.w4(32'h3c53f7a8),
	.w5(32'h3caa851e),
	.w6(32'hbc521daf),
	.w7(32'hbc2e8bec),
	.w8(32'hbb946ecc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29ce84),
	.w1(32'h3a78724f),
	.w2(32'h3ba75cc0),
	.w3(32'h3c789c41),
	.w4(32'h3c4cbe93),
	.w5(32'h3d06e433),
	.w6(32'hbc11b01e),
	.w7(32'h3c5f130f),
	.w8(32'h3c822bd7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f8122),
	.w1(32'h3c4e84e8),
	.w2(32'h3bf99152),
	.w3(32'h3c7a29d1),
	.w4(32'h3a900de8),
	.w5(32'h3b90e940),
	.w6(32'h3adcc5c1),
	.w7(32'h3b0eeaca),
	.w8(32'h3a422578),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1266a6),
	.w1(32'hb93afcee),
	.w2(32'h3b6a8379),
	.w3(32'h3b801f19),
	.w4(32'hbb037a48),
	.w5(32'hbb87717f),
	.w6(32'hbac95f4a),
	.w7(32'hbabbab0a),
	.w8(32'hbbafeceb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7e61),
	.w1(32'h3b9ea0c9),
	.w2(32'h3bfd6094),
	.w3(32'hbb1acb8b),
	.w4(32'h3aaa1e08),
	.w5(32'h3b158450),
	.w6(32'hbbd9c7a9),
	.w7(32'hbb1c7170),
	.w8(32'hbacd397e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf54fe8),
	.w1(32'h3b88a87f),
	.w2(32'h3ba850a9),
	.w3(32'h3ad18d00),
	.w4(32'h3ba2291b),
	.w5(32'h3a325687),
	.w6(32'hbb91a28b),
	.w7(32'h3c00741c),
	.w8(32'hbb047454),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8125a3),
	.w1(32'hbb636619),
	.w2(32'h39ae31c9),
	.w3(32'hba9237e2),
	.w4(32'hbbcb252a),
	.w5(32'hbc39c5b5),
	.w6(32'hbb5815de),
	.w7(32'h3c11a418),
	.w8(32'h3b8c79ea),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb72e0),
	.w1(32'h39913068),
	.w2(32'hbbb36a07),
	.w3(32'hbc2a1dc8),
	.w4(32'hbbf811d2),
	.w5(32'hbc322e8a),
	.w6(32'h3ba39c99),
	.w7(32'hbc34dc48),
	.w8(32'hbc6689e3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb40751),
	.w1(32'hba067ed9),
	.w2(32'hbb8b03f6),
	.w3(32'hbc2f8ed8),
	.w4(32'hbbc3234f),
	.w5(32'hbab6e4e6),
	.w6(32'hbc05d580),
	.w7(32'hbbf20ce8),
	.w8(32'hbb7df51f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48eec7),
	.w1(32'hbba42e25),
	.w2(32'hbb95e095),
	.w3(32'hbb53ee38),
	.w4(32'hbae13976),
	.w5(32'hbbb51543),
	.w6(32'hbbb4f3dd),
	.w7(32'hba4ca061),
	.w8(32'h3a3baad4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876dd5),
	.w1(32'hba5cad57),
	.w2(32'h39d78efa),
	.w3(32'hbbd02827),
	.w4(32'hbbbfa234),
	.w5(32'hbb19fa90),
	.w6(32'hbad8c077),
	.w7(32'hbb8a56f9),
	.w8(32'hb933df1b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4f4a),
	.w1(32'h3a1bc23a),
	.w2(32'hba96f41f),
	.w3(32'hbb6f3447),
	.w4(32'h3baebcb1),
	.w5(32'h3bedf8b0),
	.w6(32'h3ba46467),
	.w7(32'h3b7aecb6),
	.w8(32'h3ba77508),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7576c),
	.w1(32'h3ad6acb5),
	.w2(32'h3b8c924c),
	.w3(32'h3b8d1441),
	.w4(32'hba7bf1b3),
	.w5(32'hbb33b530),
	.w6(32'hb9f52c15),
	.w7(32'h3ac46568),
	.w8(32'hbbc0d89d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce79b),
	.w1(32'h3a910073),
	.w2(32'h3b350682),
	.w3(32'hba9afae6),
	.w4(32'h3b9af6c9),
	.w5(32'h3b66467e),
	.w6(32'hbb80558d),
	.w7(32'hba9c8f04),
	.w8(32'hbb96363d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76241d),
	.w1(32'h3b69050a),
	.w2(32'h3b357c58),
	.w3(32'h3b685773),
	.w4(32'h3b0c56ca),
	.w5(32'hba141f0f),
	.w6(32'hbb91c55e),
	.w7(32'h3a0f500b),
	.w8(32'hbaf0bca4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812a1f),
	.w1(32'h3b533cb2),
	.w2(32'hbbf417b3),
	.w3(32'hbacaf13b),
	.w4(32'hbb627bb6),
	.w5(32'hba8a0280),
	.w6(32'hba735217),
	.w7(32'hbac1f3ce),
	.w8(32'hbafa4cbf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbc53a),
	.w1(32'h3afb5cbc),
	.w2(32'hbaeceeb9),
	.w3(32'hbb02d422),
	.w4(32'hbba3f08b),
	.w5(32'hbbb3694d),
	.w6(32'hbb1ee890),
	.w7(32'hbb6451b2),
	.w8(32'hbbba38ca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78aa93),
	.w1(32'hb9cc301c),
	.w2(32'hbc3ac54f),
	.w3(32'hbbebb81b),
	.w4(32'hbb3eefbd),
	.w5(32'h3b27b771),
	.w6(32'hbc015e30),
	.w7(32'h3b022d2a),
	.w8(32'hb891e2f8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0dc8),
	.w1(32'h3bccc97e),
	.w2(32'hbbf2ee1a),
	.w3(32'h3ae3d046),
	.w4(32'hbb128bd3),
	.w5(32'hbbe0d52a),
	.w6(32'h3b0f534e),
	.w7(32'h3b80133f),
	.w8(32'h3a4efe3d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0ba21),
	.w1(32'h3a5a581d),
	.w2(32'h3acce590),
	.w3(32'hbad675e2),
	.w4(32'h3a8700a8),
	.w5(32'hb92a6c45),
	.w6(32'h3b301c15),
	.w7(32'h397cb494),
	.w8(32'hba856552),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5f35),
	.w1(32'h3bcffcfb),
	.w2(32'h3b0cbfa5),
	.w3(32'hbb207323),
	.w4(32'hbab7485e),
	.w5(32'hb985803f),
	.w6(32'h39f4a417),
	.w7(32'hbb2c9350),
	.w8(32'hb88317da),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802dd2),
	.w1(32'h3bbfdafc),
	.w2(32'h3aee208f),
	.w3(32'hbacd222c),
	.w4(32'h3bb65830),
	.w5(32'h3ab2269b),
	.w6(32'hbb22f8a6),
	.w7(32'h3ba0c7ec),
	.w8(32'h3b1ae494),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d6416),
	.w1(32'hbb1f8780),
	.w2(32'h3a7db351),
	.w3(32'hbbaa5ca1),
	.w4(32'hbb154bb5),
	.w5(32'hba352d4e),
	.w6(32'h3bdf7fd7),
	.w7(32'h3b05832f),
	.w8(32'h3ae0ee75),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92fbdd),
	.w1(32'h3b8f340c),
	.w2(32'h3b7810eb),
	.w3(32'h3acc763b),
	.w4(32'hbb2bb664),
	.w5(32'hbbb8ba7b),
	.w6(32'h3b5577c1),
	.w7(32'h3b28cb93),
	.w8(32'hbb9d02d3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4cb35),
	.w1(32'h3c25b6e7),
	.w2(32'hb787f081),
	.w3(32'hbb716b21),
	.w4(32'h3c118934),
	.w5(32'h3b40753c),
	.w6(32'hbb27c302),
	.w7(32'hbb222573),
	.w8(32'h3a7863dc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1b139),
	.w1(32'hb8582bd5),
	.w2(32'h3b540687),
	.w3(32'h3c07e411),
	.w4(32'hbb573498),
	.w5(32'h380694f0),
	.w6(32'h3b051328),
	.w7(32'hbb7813bd),
	.w8(32'hbb3b50a3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969892e),
	.w1(32'h3b1289aa),
	.w2(32'hba2d6e6f),
	.w3(32'hbbf17a90),
	.w4(32'h3bbc5666),
	.w5(32'h3bbf3978),
	.w6(32'h39fdbcc0),
	.w7(32'h3ba61327),
	.w8(32'h3b5140c4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d6c1),
	.w1(32'hbbca94ae),
	.w2(32'hbc1b721a),
	.w3(32'hba20b200),
	.w4(32'hbc976998),
	.w5(32'hbcb830e3),
	.w6(32'h394d4b7c),
	.w7(32'h3bc5a4b2),
	.w8(32'h3c0d3a79),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4710e),
	.w1(32'hba13518d),
	.w2(32'hbae2eee1),
	.w3(32'hbc22fa81),
	.w4(32'hbb6d5559),
	.w5(32'h39a517b8),
	.w6(32'h3c7d39df),
	.w7(32'hbac7173e),
	.w8(32'hbae9e820),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd77df),
	.w1(32'hbc1cae1e),
	.w2(32'hbc483398),
	.w3(32'h3a99fddf),
	.w4(32'hbc56d0f5),
	.w5(32'hbc722850),
	.w6(32'hbb5d65b1),
	.w7(32'hbc03d5af),
	.w8(32'hbc3ee1f7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d53a),
	.w1(32'h3bbd27b2),
	.w2(32'hbb315565),
	.w3(32'hbc09f378),
	.w4(32'hbbaba5f9),
	.w5(32'hbc11128c),
	.w6(32'hbc3445a2),
	.w7(32'hbb624f93),
	.w8(32'hbba5a1f9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe468),
	.w1(32'h3ab67e1c),
	.w2(32'hbb991905),
	.w3(32'hbbb470ee),
	.w4(32'hba652329),
	.w5(32'hbad79113),
	.w6(32'hbbb9293c),
	.w7(32'h3b0157f9),
	.w8(32'hbb6964b5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0071),
	.w1(32'hbb41a477),
	.w2(32'hbae5e874),
	.w3(32'hba7c49b7),
	.w4(32'hbb9fddcf),
	.w5(32'hbbc83229),
	.w6(32'hba896b11),
	.w7(32'hbb46de2a),
	.w8(32'h3b73e5b0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb48d6),
	.w1(32'h389f9aa6),
	.w2(32'h3c5e62f8),
	.w3(32'hbb8a46a2),
	.w4(32'hbc220e53),
	.w5(32'hbc3f0b12),
	.w6(32'hba67527a),
	.w7(32'h3b80dafb),
	.w8(32'h3ab30e08),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2430d),
	.w1(32'h3b36c276),
	.w2(32'h3a524e2c),
	.w3(32'h3ac43a34),
	.w4(32'hbaf2e7b8),
	.w5(32'hbbe7749f),
	.w6(32'h3c5ff4de),
	.w7(32'hbb7bd1a6),
	.w8(32'hbba8acc2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f48a),
	.w1(32'hbad9e03f),
	.w2(32'h3a7b11aa),
	.w3(32'hbb0b789e),
	.w4(32'hbbe8a1af),
	.w5(32'hbb211857),
	.w6(32'hbb671dd3),
	.w7(32'hbac16dad),
	.w8(32'hba9a902f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3caa66),
	.w1(32'h3ae376bc),
	.w2(32'hbabce317),
	.w3(32'hbb21bbde),
	.w4(32'h3b3196ee),
	.w5(32'hbbc1df91),
	.w6(32'hb9985dad),
	.w7(32'h3b4627b9),
	.w8(32'h3a7d80f8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205372),
	.w1(32'h3b2ae794),
	.w2(32'h3b7a4cb6),
	.w3(32'h397c4575),
	.w4(32'h3b8669c5),
	.w5(32'h3c2b9c0a),
	.w6(32'h3a077473),
	.w7(32'h3b6092e1),
	.w8(32'h3ab655c9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfa806),
	.w1(32'hbba8da56),
	.w2(32'hbbbbe88b),
	.w3(32'h3b2c62df),
	.w4(32'hbbc88caa),
	.w5(32'hbb4b18c7),
	.w6(32'hbb5e7af3),
	.w7(32'hba9fc3da),
	.w8(32'hbb9e95b8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75b21d),
	.w1(32'hbad4cb2b),
	.w2(32'hbbbcd40f),
	.w3(32'h39555828),
	.w4(32'hb90930b8),
	.w5(32'hbaa5475f),
	.w6(32'hbb9ff59c),
	.w7(32'h39da1b5f),
	.w8(32'h39f8d1e0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeaa62),
	.w1(32'hbb1784a9),
	.w2(32'hbb1ce783),
	.w3(32'hbafdd4ca),
	.w4(32'hbaba3205),
	.w5(32'hba911f5e),
	.w6(32'h3b421ab3),
	.w7(32'hbb2742e2),
	.w8(32'h3af5291f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0bc05),
	.w1(32'h3b913a5e),
	.w2(32'h3b8f75e0),
	.w3(32'hbb383aa9),
	.w4(32'h3b515ff2),
	.w5(32'h3bcf7242),
	.w6(32'h3bc6b1e7),
	.w7(32'h3bf1114e),
	.w8(32'h3b15f4ee),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c285da5),
	.w1(32'h3c15e254),
	.w2(32'hba92baf3),
	.w3(32'h3bfd89fb),
	.w4(32'hbbfa6146),
	.w5(32'hbc6890c4),
	.w6(32'hba90c8cf),
	.w7(32'hbc5213b8),
	.w8(32'hbbad44f3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0c4b),
	.w1(32'h3b18e314),
	.w2(32'hbaadf37d),
	.w3(32'hbbe10b21),
	.w4(32'h3be4b277),
	.w5(32'h3bdee04d),
	.w6(32'h37f288e9),
	.w7(32'h3bc13742),
	.w8(32'h3b20433e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88df10),
	.w1(32'hbbaffd42),
	.w2(32'hbbc92ad3),
	.w3(32'h3aef3619),
	.w4(32'hb8925729),
	.w5(32'hb93e8674),
	.w6(32'h3b0dd26e),
	.w7(32'hbb0e2299),
	.w8(32'h398d0479),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170cc2),
	.w1(32'hbc02beec),
	.w2(32'hbbe03b7a),
	.w3(32'hbad87952),
	.w4(32'hbb083d73),
	.w5(32'hbab32c19),
	.w6(32'hb9d4d03e),
	.w7(32'h39490d9a),
	.w8(32'hbada94fb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4c5f9),
	.w1(32'hbb8e2bd8),
	.w2(32'hbb4ea985),
	.w3(32'h3b5ff824),
	.w4(32'hbbdeef79),
	.w5(32'hbc17470d),
	.w6(32'h3a69ad01),
	.w7(32'hbb9cbb7a),
	.w8(32'hbb717dd1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3ef2c),
	.w1(32'h3baed560),
	.w2(32'h3b89ddbb),
	.w3(32'hba489962),
	.w4(32'h3999f352),
	.w5(32'hba26b541),
	.w6(32'hba053175),
	.w7(32'h3aa79aa1),
	.w8(32'h3be69269),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397db1),
	.w1(32'h3bc19a4a),
	.w2(32'h3c2bf311),
	.w3(32'h3b1809cf),
	.w4(32'hbb9f8b68),
	.w5(32'hbb41c2a4),
	.w6(32'h3b7c2494),
	.w7(32'h39bc3802),
	.w8(32'hbbeec086),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67a1e0),
	.w1(32'hbb270105),
	.w2(32'hbb979d0b),
	.w3(32'hbb5ecfc5),
	.w4(32'h3a6d57d0),
	.w5(32'hbb6ab7a7),
	.w6(32'hbbd085bd),
	.w7(32'h3b26295f),
	.w8(32'h3a5088be),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc531a4),
	.w1(32'hba9cdd38),
	.w2(32'h3b765c27),
	.w3(32'hbba8e420),
	.w4(32'h3b12995a),
	.w5(32'h3b359b4a),
	.w6(32'hbaa0955d),
	.w7(32'hb98b4917),
	.w8(32'hbb987e69),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c6c13),
	.w1(32'h3aed4227),
	.w2(32'h3b3a90b6),
	.w3(32'hbaab673e),
	.w4(32'h3b6326ad),
	.w5(32'hbba71e65),
	.w6(32'hbad20ce2),
	.w7(32'hbb8c7bff),
	.w8(32'hbc04889f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b64ad),
	.w1(32'hbb9794d5),
	.w2(32'hbba2406f),
	.w3(32'h3be219a0),
	.w4(32'h3a46939f),
	.w5(32'hb9d99dc6),
	.w6(32'hba12775f),
	.w7(32'h3adcd6c7),
	.w8(32'h3b346e25),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbadff6),
	.w1(32'h3b9774ee),
	.w2(32'h3b0ce7ad),
	.w3(32'h3b9ecf7b),
	.w4(32'h3c229681),
	.w5(32'h3a2e84ea),
	.w6(32'h3b689b31),
	.w7(32'h3bc82e93),
	.w8(32'h3c19d59f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f21e4),
	.w1(32'h3c0111a9),
	.w2(32'h3ba061d7),
	.w3(32'h3afe5131),
	.w4(32'h3a8b0109),
	.w5(32'hbb441904),
	.w6(32'h3c001ead),
	.w7(32'hbc020951),
	.w8(32'hbc30f71c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae44b32),
	.w1(32'h3b849b28),
	.w2(32'h3a093c7c),
	.w3(32'hba9a5266),
	.w4(32'hbc1ad676),
	.w5(32'hbbcc3554),
	.w6(32'hbc000132),
	.w7(32'hbbc9e2df),
	.w8(32'hbb4ef0b5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4bea9),
	.w1(32'h3b6f803a),
	.w2(32'h3a9714ed),
	.w3(32'hbb1171d4),
	.w4(32'h3b10b630),
	.w5(32'hbb8862cd),
	.w6(32'h3a5c6894),
	.w7(32'h3b218ce0),
	.w8(32'h3a095c35),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3c04a),
	.w1(32'hbb0177da),
	.w2(32'hbb7f0a39),
	.w3(32'hbb69dd70),
	.w4(32'h3ac0c414),
	.w5(32'hbac2a392),
	.w6(32'hb9304d86),
	.w7(32'h3be36768),
	.w8(32'h3c113b87),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c1d0),
	.w1(32'h3a92a171),
	.w2(32'hb91b63c1),
	.w3(32'h3ab357b0),
	.w4(32'hb9d55357),
	.w5(32'hba4bc7ae),
	.w6(32'h3c254b8a),
	.w7(32'h3b6d283d),
	.w8(32'hbbc33c60),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905ddbd),
	.w1(32'h3ad3747b),
	.w2(32'h3bce1227),
	.w3(32'hb9a9c0e9),
	.w4(32'hbbd38b7e),
	.w5(32'h3bd98f74),
	.w6(32'hbb997393),
	.w7(32'hbc9f1b34),
	.w8(32'hbc7dc7da),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c6bae),
	.w1(32'h3b71efef),
	.w2(32'h3b7dad6a),
	.w3(32'hbb09df25),
	.w4(32'hbb6fa1a0),
	.w5(32'h3a6818d1),
	.w6(32'hbc7499c5),
	.w7(32'hbbd721e8),
	.w8(32'hb7ae1aec),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8dd9),
	.w1(32'h3b619158),
	.w2(32'hbb250c7c),
	.w3(32'hbbbd4d73),
	.w4(32'h397f25cf),
	.w5(32'hba7eb22e),
	.w6(32'hbb86765f),
	.w7(32'h3aacb9c9),
	.w8(32'hbb8b61bc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e927d),
	.w1(32'h39bf41d8),
	.w2(32'hbb47a690),
	.w3(32'hbb5d76e0),
	.w4(32'h39993976),
	.w5(32'hbba70ff5),
	.w6(32'hbb097c00),
	.w7(32'h392defc4),
	.w8(32'hbb6ec886),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7942c7),
	.w1(32'h3b0f2e04),
	.w2(32'h3b0adbf3),
	.w3(32'hbb49bb28),
	.w4(32'hb9bc15e5),
	.w5(32'hbb509e88),
	.w6(32'hbb38be60),
	.w7(32'hbba73e27),
	.w8(32'hbb903868),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29216e),
	.w1(32'hbb8a4156),
	.w2(32'hba02bb14),
	.w3(32'hbbffb781),
	.w4(32'h3b92fb47),
	.w5(32'h3c4ed073),
	.w6(32'hbb990f67),
	.w7(32'h3c43b977),
	.w8(32'h3bb4cca2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a8c4),
	.w1(32'h3b941131),
	.w2(32'h3b2f6cbe),
	.w3(32'h3b95ad6a),
	.w4(32'h3b83a501),
	.w5(32'hb9f685b6),
	.w6(32'hbab5cc71),
	.w7(32'h3b97c93a),
	.w8(32'h3a470951),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463f50),
	.w1(32'h3b1d9327),
	.w2(32'h3b05cf92),
	.w3(32'h3b9123c0),
	.w4(32'hbacfa53e),
	.w5(32'hbb82576a),
	.w6(32'h3adcaded),
	.w7(32'hba996310),
	.w8(32'hba83a306),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08403),
	.w1(32'h3bb0e1ae),
	.w2(32'hbb75b0da),
	.w3(32'hbb86718a),
	.w4(32'hbb961c88),
	.w5(32'hbaa59c50),
	.w6(32'hbb08c19e),
	.w7(32'hbb2e600e),
	.w8(32'hbbdf66fd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab452c1),
	.w1(32'h3b3892cc),
	.w2(32'h3bd08935),
	.w3(32'hba9205c7),
	.w4(32'h3c0e9647),
	.w5(32'h3c5d36ff),
	.w6(32'hbbb0c1a4),
	.w7(32'h3bad6161),
	.w8(32'h3b811294),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e505d),
	.w1(32'h3b0ef9d5),
	.w2(32'h3b396785),
	.w3(32'h3c0b15d3),
	.w4(32'hba2eaed0),
	.w5(32'hbb64ceb9),
	.w6(32'h3bcab983),
	.w7(32'hba0a4a83),
	.w8(32'h3a791203),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f5357),
	.w1(32'h397bb66c),
	.w2(32'hbb8223c6),
	.w3(32'h3bb250c0),
	.w4(32'hbb47243c),
	.w5(32'hbb23d197),
	.w6(32'h3b658ca9),
	.w7(32'hbbe86c32),
	.w8(32'hbb595eaf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d17f),
	.w1(32'h3be8f925),
	.w2(32'h3b0258aa),
	.w3(32'hbb866ac4),
	.w4(32'h3a937045),
	.w5(32'h3c00cbe0),
	.w6(32'hb9f89e51),
	.w7(32'hba914c26),
	.w8(32'hbb287537),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cbe1a),
	.w1(32'hbb57bc52),
	.w2(32'h3b7539b7),
	.w3(32'h3ab616f1),
	.w4(32'hbb295bd3),
	.w5(32'hbaebd13b),
	.w6(32'h39da7752),
	.w7(32'h3aff2ff3),
	.w8(32'hba821491),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae30125),
	.w1(32'h3ab7d72d),
	.w2(32'h3b533dbf),
	.w3(32'h3adf08e6),
	.w4(32'h3a99ce75),
	.w5(32'h3b898261),
	.w6(32'h39da6831),
	.w7(32'h3b661722),
	.w8(32'h3add0852),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92521f),
	.w1(32'h3a8fa5bb),
	.w2(32'h3ae33f74),
	.w3(32'h3b872ad8),
	.w4(32'h3b040dad),
	.w5(32'h3a7f89f2),
	.w6(32'h3b9e6b7b),
	.w7(32'h3a8174a4),
	.w8(32'h3b099da9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fc6fd),
	.w1(32'hbbf506d4),
	.w2(32'hbb4cb008),
	.w3(32'h3b67e10c),
	.w4(32'h39942e22),
	.w5(32'h3be1b924),
	.w6(32'h3b33d92d),
	.w7(32'h3b2bd439),
	.w8(32'h3ab37daf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d7983),
	.w1(32'h3a1dbe81),
	.w2(32'h3b876c7a),
	.w3(32'h3b797f7c),
	.w4(32'h3b7d75a1),
	.w5(32'hbbd73a83),
	.w6(32'hbb33bed3),
	.w7(32'hbad1fe42),
	.w8(32'h3b88a4f9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba923942),
	.w1(32'h3b5c161a),
	.w2(32'h3b3f01ed),
	.w3(32'h3aca9b25),
	.w4(32'h3a0adfcd),
	.w5(32'hbb2414fe),
	.w6(32'h3a2bff2b),
	.w7(32'h3b432374),
	.w8(32'h3a9459e5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b572b1f),
	.w1(32'h3b38f01d),
	.w2(32'hbb58a8b0),
	.w3(32'h3ba8ab13),
	.w4(32'hb9a1cb24),
	.w5(32'h3b6c4b97),
	.w6(32'h3b67f7ed),
	.w7(32'h39792a5b),
	.w8(32'h3a23738e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9629f2),
	.w1(32'h3b1df1e0),
	.w2(32'hba52cbb3),
	.w3(32'hb98d8e8b),
	.w4(32'hbba91d39),
	.w5(32'hbbc8be97),
	.w6(32'hbb4eb3ac),
	.w7(32'hbaf27bc3),
	.w8(32'hbb45bb1b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec02f1),
	.w1(32'h3bc21024),
	.w2(32'hbaa45bac),
	.w3(32'hbb4cd874),
	.w4(32'hbad22db6),
	.w5(32'h3a8884d1),
	.w6(32'h3a549260),
	.w7(32'hbb70b4a7),
	.w8(32'hba7aa563),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857270),
	.w1(32'hba35aace),
	.w2(32'h3adf0d9b),
	.w3(32'hbaa5a21a),
	.w4(32'hba8eb75d),
	.w5(32'hbb6ff5b0),
	.w6(32'hba0a58eb),
	.w7(32'hbb9931e6),
	.w8(32'hbbfac7a2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30719f),
	.w1(32'h3afead84),
	.w2(32'hb9a24dac),
	.w3(32'hbb223d83),
	.w4(32'hbb182b35),
	.w5(32'hbba1d524),
	.w6(32'h39ff60d4),
	.w7(32'hba975e31),
	.w8(32'hbb5b15a4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e1f15),
	.w1(32'hba6e0764),
	.w2(32'h3b527f15),
	.w3(32'hbb1caa94),
	.w4(32'hb9c9a701),
	.w5(32'hbad89689),
	.w6(32'hbba5b2f8),
	.w7(32'hbb6a2064),
	.w8(32'hb9da0f40),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0970e),
	.w1(32'h3a4ff1d8),
	.w2(32'hbb9c2cb3),
	.w3(32'h39fc035c),
	.w4(32'hbc22fc68),
	.w5(32'hbc3d8494),
	.w6(32'hbaca12ef),
	.w7(32'h3bbe013b),
	.w8(32'h3a2d5a35),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8841a9),
	.w1(32'hbb35487a),
	.w2(32'hbb0a4bc4),
	.w3(32'hbc059c96),
	.w4(32'h3ba3e759),
	.w5(32'h3c6f9939),
	.w6(32'h3b2db803),
	.w7(32'h3b96d578),
	.w8(32'h3aaedc7c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbea69c),
	.w1(32'h3a1d8970),
	.w2(32'hba4989f1),
	.w3(32'h3c43da4c),
	.w4(32'h3a14c04d),
	.w5(32'h3a920c93),
	.w6(32'h3b00013f),
	.w7(32'hba84b8dd),
	.w8(32'h3a38b760),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba587e25),
	.w1(32'h3b077766),
	.w2(32'h38d359b3),
	.w3(32'h3af78967),
	.w4(32'hbbb9b68f),
	.w5(32'hbbb99015),
	.w6(32'h3b41a41b),
	.w7(32'hbb0ad445),
	.w8(32'hba90b31d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d938),
	.w1(32'h3ba080ed),
	.w2(32'h3b9f156a),
	.w3(32'hbb6f807f),
	.w4(32'h3aeaf46c),
	.w5(32'hbc0bfb45),
	.w6(32'hba4ee7b0),
	.w7(32'hbb098810),
	.w8(32'hbbb057ce),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b716),
	.w1(32'hb9c173d5),
	.w2(32'hbacd9ad8),
	.w3(32'hbbbcb2ea),
	.w4(32'hba095b6f),
	.w5(32'hbb5cad61),
	.w6(32'hbbc28d8f),
	.w7(32'h3b6f49ea),
	.w8(32'h3b182ebf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a9ac0),
	.w1(32'hbaf56446),
	.w2(32'hba08bc77),
	.w3(32'hbaca63db),
	.w4(32'h3a806eeb),
	.w5(32'hbab03342),
	.w6(32'h3ad420ca),
	.w7(32'hbb08b19e),
	.w8(32'hbadaaa78),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aab56),
	.w1(32'hbb05232a),
	.w2(32'h3a871be3),
	.w3(32'h3ae3ebfd),
	.w4(32'hbb1afc3e),
	.w5(32'hbb53999a),
	.w6(32'h3953f55e),
	.w7(32'hbb2ad51b),
	.w8(32'hbb5744c4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90368a),
	.w1(32'h3a4755f4),
	.w2(32'hba80ccbe),
	.w3(32'hbb29c342),
	.w4(32'hbb02ef05),
	.w5(32'hbb844562),
	.w6(32'hbb8cef79),
	.w7(32'hbb7144ef),
	.w8(32'hbb26aa5f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5d668),
	.w1(32'h3aba4b43),
	.w2(32'h39e296dd),
	.w3(32'hba96e22f),
	.w4(32'hba9f4598),
	.w5(32'h3a87d39b),
	.w6(32'hbb7c9730),
	.w7(32'hbac29994),
	.w8(32'h3b501daf),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c309),
	.w1(32'hbae9c01f),
	.w2(32'hbb82f2c9),
	.w3(32'hbb7c143a),
	.w4(32'hbb9c735a),
	.w5(32'hbbdf0fd7),
	.w6(32'hb71bb795),
	.w7(32'hbb6e79a0),
	.w8(32'hbbf9519f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123e7b),
	.w1(32'h3a1f93d7),
	.w2(32'hbb2d56ed),
	.w3(32'hbb48b77d),
	.w4(32'hbada343d),
	.w5(32'hbba11794),
	.w6(32'hbb8861a3),
	.w7(32'hbab4800d),
	.w8(32'hba223779),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ccc27),
	.w1(32'h3b07ee4a),
	.w2(32'h3a5ca5ac),
	.w3(32'hbbc34ce9),
	.w4(32'hbb4aaca6),
	.w5(32'hbbd584d5),
	.w6(32'hbb701f57),
	.w7(32'h3aea355a),
	.w8(32'h38441c63),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98161e4),
	.w1(32'h38c5da6c),
	.w2(32'h3a0ab0e8),
	.w3(32'hb9f566b8),
	.w4(32'h3baeb2b7),
	.w5(32'h3c749d66),
	.w6(32'h3b6c73ac),
	.w7(32'h3af5804f),
	.w8(32'h3a7d8b6f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4e20d),
	.w1(32'h3b24f185),
	.w2(32'h3a9563b6),
	.w3(32'h3c56634d),
	.w4(32'h3a9328b2),
	.w5(32'h3afa4062),
	.w6(32'h3a422551),
	.w7(32'h3b093c62),
	.w8(32'h3b864e6b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b024799),
	.w1(32'hbaef8ae0),
	.w2(32'hbb674f7b),
	.w3(32'h3b09913a),
	.w4(32'hba87d441),
	.w5(32'h3afdf23c),
	.w6(32'h3aa3e2b3),
	.w7(32'hbb434769),
	.w8(32'hbb474412),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb527c27),
	.w1(32'hbb1e31eb),
	.w2(32'hba74a56e),
	.w3(32'hbaadf532),
	.w4(32'hbb96c9e8),
	.w5(32'hbb3768f4),
	.w6(32'hba135755),
	.w7(32'hb9a73410),
	.w8(32'hb9963516),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e968d),
	.w1(32'h3a8b4cc9),
	.w2(32'h3a5b11e3),
	.w3(32'hbaeb8f1e),
	.w4(32'h3be902a0),
	.w5(32'h3c746fff),
	.w6(32'hbb673b07),
	.w7(32'h3b82e4c6),
	.w8(32'h3aefe91f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac9c7b),
	.w1(32'hbb2d1ed5),
	.w2(32'hbb8bc60c),
	.w3(32'h3c3020b0),
	.w4(32'h3b8297e6),
	.w5(32'h3ab09de4),
	.w6(32'h3a49b78b),
	.w7(32'h3a310171),
	.w8(32'hbba3afca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525ff0),
	.w1(32'h3afb2c8d),
	.w2(32'h3b86964f),
	.w3(32'h3bddb2ba),
	.w4(32'h3b998845),
	.w5(32'h3c063f2b),
	.w6(32'hbad60f59),
	.w7(32'h3ba1e01f),
	.w8(32'h3bafc089),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09ee97),
	.w1(32'h3ab8f058),
	.w2(32'hbab69ff1),
	.w3(32'h3b8322ea),
	.w4(32'h3b0d1f4a),
	.w5(32'hbb20fbeb),
	.w6(32'h3aa86d7c),
	.w7(32'h3aeac79a),
	.w8(32'h3afbc246),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c6b3),
	.w1(32'h3a07bdef),
	.w2(32'h3ac3059f),
	.w3(32'h3ad96f1e),
	.w4(32'hbbe64f9f),
	.w5(32'hbbd3c6ff),
	.w6(32'hba2886f1),
	.w7(32'hbb803da7),
	.w8(32'hbb2ffc88),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46c04),
	.w1(32'hba11efcf),
	.w2(32'hbbf86335),
	.w3(32'hbbd16d42),
	.w4(32'hbb632a2c),
	.w5(32'h3a91af65),
	.w6(32'hba711b30),
	.w7(32'hbbbbcdbb),
	.w8(32'hbc16536a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4f0fd),
	.w1(32'h3a463502),
	.w2(32'h3b6378f0),
	.w3(32'hbbb63dc3),
	.w4(32'h3a4c7578),
	.w5(32'h3b35a87c),
	.w6(32'hbb2dad7a),
	.w7(32'h3b2ddb7c),
	.w8(32'h3aaf96a5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92dab0),
	.w1(32'h3b565f2a),
	.w2(32'h3ae1753c),
	.w3(32'h397e138e),
	.w4(32'h3a662829),
	.w5(32'h3a3c5a0e),
	.w6(32'h39e25989),
	.w7(32'h3ae3595e),
	.w8(32'hb9a296c4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137b53),
	.w1(32'hb93fa37b),
	.w2(32'h3b7f1d5b),
	.w3(32'h3a4ed44c),
	.w4(32'h3b67b343),
	.w5(32'h3ad5b977),
	.w6(32'hba44a2a7),
	.w7(32'h3afc0b6f),
	.w8(32'h3ba5612a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f15ac),
	.w1(32'h3a9effc7),
	.w2(32'h3b1b634c),
	.w3(32'h3b192410),
	.w4(32'h3c37552f),
	.w5(32'h3bfb8a98),
	.w6(32'h3b0d797c),
	.w7(32'h3ba08cfa),
	.w8(32'h3b2ac40a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0b576),
	.w1(32'hbb092e0a),
	.w2(32'hbb597e64),
	.w3(32'h3c263c51),
	.w4(32'hbb624d4c),
	.w5(32'hbb151d9f),
	.w6(32'h3b0499e5),
	.w7(32'hbc036c14),
	.w8(32'hbbe97cd7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71df59),
	.w1(32'hbb3f428a),
	.w2(32'hba6d208c),
	.w3(32'hbbe11b68),
	.w4(32'hbae17dfe),
	.w5(32'hbbea03dd),
	.w6(32'hbbaee3c8),
	.w7(32'h3b8a80a8),
	.w8(32'h3b49f368),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b92690),
	.w1(32'hb8c5eb69),
	.w2(32'h3748bcd4),
	.w3(32'hbb65e983),
	.w4(32'h3b093bbf),
	.w5(32'hb9d093c2),
	.w6(32'hbaf45645),
	.w7(32'h3afc38df),
	.w8(32'hb9bc293c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b904),
	.w1(32'h3b6edcb6),
	.w2(32'h3a858b66),
	.w3(32'h3b81d8d0),
	.w4(32'h3b62cdc4),
	.w5(32'h3b0a8798),
	.w6(32'h3b851f29),
	.w7(32'hbb0ad800),
	.w8(32'hbba2ee4b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21ff7),
	.w1(32'h3a348973),
	.w2(32'hba69c8bd),
	.w3(32'hbb466ea1),
	.w4(32'hba9752cc),
	.w5(32'hbad8ffde),
	.w6(32'h3b156852),
	.w7(32'h3b631a7c),
	.w8(32'h3bac22de),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a5d6),
	.w1(32'hbab87139),
	.w2(32'h3a2d850f),
	.w3(32'hbb7565d5),
	.w4(32'hba812e40),
	.w5(32'hbb74108d),
	.w6(32'hba9c25c8),
	.w7(32'h39fbfc8c),
	.w8(32'h3949cd50),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bf3bb),
	.w1(32'hbb9dc9c8),
	.w2(32'hbb56ab5b),
	.w3(32'hbb450fec),
	.w4(32'h3c1725a9),
	.w5(32'h3c498c86),
	.w6(32'hbadf143a),
	.w7(32'h3c3bb7a6),
	.w8(32'h3b68720b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd107ac),
	.w1(32'hbb24782f),
	.w2(32'hbbc7121f),
	.w3(32'h3c220816),
	.w4(32'h3af7cb9e),
	.w5(32'h3c16d6a4),
	.w6(32'h3b4de2d6),
	.w7(32'hb91fda1d),
	.w8(32'hbb0e6c90),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f1384),
	.w1(32'hbbe2abe2),
	.w2(32'hbb8603d8),
	.w3(32'h3bb1f126),
	.w4(32'hbbef65d3),
	.w5(32'hbbf3c782),
	.w6(32'h39f2fb3b),
	.w7(32'hbb615a78),
	.w8(32'hba999342),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11404b),
	.w1(32'h3b1e2717),
	.w2(32'hba0e301b),
	.w3(32'hbbb38ea7),
	.w4(32'h3ad03934),
	.w5(32'h39ba0300),
	.w6(32'hbb076892),
	.w7(32'h3ad7e640),
	.w8(32'h3aa6e162),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule