module layer_6_featuremap_7(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3fded8),
	.w1(32'hbc747355),
	.w2(32'hbd0ba3c3),
	.w3(32'hbc24db77),
	.w4(32'h3d0048e3),
	.w5(32'h3c994e82),
	.w6(32'h3b4eecac),
	.w7(32'h3cce89a1),
	.w8(32'hbd21f019),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27976),
	.w1(32'h3bfd861f),
	.w2(32'h3c533123),
	.w3(32'hbd50b3cd),
	.w4(32'h3be8468a),
	.w5(32'h3c97a41d),
	.w6(32'hbc4bb0d2),
	.w7(32'hb9e05088),
	.w8(32'hbbc1124a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ce592),
	.w1(32'h3a837dca),
	.w2(32'hbc2d08b7),
	.w3(32'h3c8b3910),
	.w4(32'h3c4dc131),
	.w5(32'hbccbe4ff),
	.w6(32'hbc1a78bf),
	.w7(32'h3cb1c40a),
	.w8(32'h3a35b7c7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7d353),
	.w1(32'h3c0458b8),
	.w2(32'hbde263e0),
	.w3(32'h3c5984da),
	.w4(32'hbc1d8df4),
	.w5(32'h3d50fe5b),
	.w6(32'h3ccfc4d9),
	.w7(32'h3cf6c2a9),
	.w8(32'h3c57eb57),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5aacc3),
	.w1(32'hbab30787),
	.w2(32'hbc137b37),
	.w3(32'h3cb9b460),
	.w4(32'h3ab95aa2),
	.w5(32'h3b323b2c),
	.w6(32'hbba87619),
	.w7(32'h3943d872),
	.w8(32'hbb5ef84e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a476),
	.w1(32'hbcbda026),
	.w2(32'h3d06dc8b),
	.w3(32'h3b1c3b1f),
	.w4(32'hbd2ff8b9),
	.w5(32'h3d936353),
	.w6(32'hbccf617c),
	.w7(32'h3cbdae20),
	.w8(32'h3cfd317c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83bf78),
	.w1(32'hbc388e01),
	.w2(32'hbc85185f),
	.w3(32'hbbf633f7),
	.w4(32'hbc515854),
	.w5(32'hbc862026),
	.w6(32'hbc942afe),
	.w7(32'hbcaeb1f0),
	.w8(32'hbd024959),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b654e),
	.w1(32'hbc5aeb6c),
	.w2(32'hbd2f3f5c),
	.w3(32'hb9849fda),
	.w4(32'h3b8a9ba1),
	.w5(32'h3d340f28),
	.w6(32'h3c927b26),
	.w7(32'h3c679c19),
	.w8(32'h3b34f167),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcee15),
	.w1(32'h3ac61929),
	.w2(32'hbcb4329d),
	.w3(32'h3c6d8fe7),
	.w4(32'h3bf1f90e),
	.w5(32'h3b5d1de7),
	.w6(32'h3b78f973),
	.w7(32'hbb9ce179),
	.w8(32'h3b9a716c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef136f),
	.w1(32'h393918d4),
	.w2(32'hbad6e95a),
	.w3(32'h3c10a729),
	.w4(32'h3b0f7777),
	.w5(32'h3b46edca),
	.w6(32'h394035dd),
	.w7(32'h3b09c226),
	.w8(32'hbb8c2cfa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a38ef),
	.w1(32'hbd396013),
	.w2(32'hbdd7b651),
	.w3(32'hbc73b90c),
	.w4(32'hbd16fa54),
	.w5(32'hbcc79592),
	.w6(32'hbcbe03f4),
	.w7(32'h3be6803f),
	.w8(32'hbc8d8cfb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd89a750),
	.w1(32'h3c5e7e9c),
	.w2(32'hbc970ba5),
	.w3(32'hbc6b96f5),
	.w4(32'h3ba2b423),
	.w5(32'hbc02c11c),
	.w6(32'h3aab479c),
	.w7(32'hbb961246),
	.w8(32'hbc09dcdf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc52418),
	.w1(32'h3be48cf9),
	.w2(32'h3d43ce78),
	.w3(32'h3a2013f9),
	.w4(32'h3b89ea9e),
	.w5(32'hbca38664),
	.w6(32'h3c2a0567),
	.w7(32'h3bf23244),
	.w8(32'h3a8fe085),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b21a9),
	.w1(32'hbba91fb5),
	.w2(32'hbd5f3604),
	.w3(32'hbcac130c),
	.w4(32'hbc1d111f),
	.w5(32'hbd31fc41),
	.w6(32'hb9b80215),
	.w7(32'hbc8be081),
	.w8(32'hbd338946),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d7172),
	.w1(32'h3d5731e6),
	.w2(32'hbd7a5056),
	.w3(32'hbb813af3),
	.w4(32'hbbb2e0fb),
	.w5(32'hbdab2aec),
	.w6(32'h3c3ec3d9),
	.w7(32'hbd28b30a),
	.w8(32'hbcdacbfe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670f03),
	.w1(32'h3ba2abae),
	.w2(32'hbd3e40ff),
	.w3(32'h3c2c1f4d),
	.w4(32'hbab32499),
	.w5(32'hbd980c6b),
	.w6(32'hbcb1f82c),
	.w7(32'hbd3b42ac),
	.w8(32'hbcc13346),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0910),
	.w1(32'hbc423546),
	.w2(32'h3bf71b6b),
	.w3(32'h3c07a485),
	.w4(32'h3cd0c854),
	.w5(32'hbcb47a3f),
	.w6(32'h3c625064),
	.w7(32'h3b991d8f),
	.w8(32'h3bc1f255),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb7b82),
	.w1(32'h3c98fe0a),
	.w2(32'hb9fb46e5),
	.w3(32'h3c04ca49),
	.w4(32'h3c5cd1fb),
	.w5(32'hba1778a5),
	.w6(32'h3b4f7155),
	.w7(32'h3c8496b7),
	.w8(32'hbc7c9358),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd297040),
	.w1(32'h39f46ef8),
	.w2(32'hbb9ffe78),
	.w3(32'h3ba023b7),
	.w4(32'hbb2935d9),
	.w5(32'h3bdd12bd),
	.w6(32'hbb30ca37),
	.w7(32'hbb1b3b4c),
	.w8(32'hbb7ca9c8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b85c31),
	.w1(32'h3ccedd23),
	.w2(32'h3d044ed8),
	.w3(32'h3bbc30af),
	.w4(32'h3c988a08),
	.w5(32'hbdbacd92),
	.w6(32'hbbdd8773),
	.w7(32'h3c7f334b),
	.w8(32'h3c16b8d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd29b3),
	.w1(32'hbcb28b72),
	.w2(32'hbd30a22a),
	.w3(32'hbd07122d),
	.w4(32'h3b9bb157),
	.w5(32'hbca5b819),
	.w6(32'h3aeb4086),
	.w7(32'hbba8dec7),
	.w8(32'hbc223458),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3813b9),
	.w1(32'h3c429f6a),
	.w2(32'hbcd68c38),
	.w3(32'h3ae16bf0),
	.w4(32'h3c912310),
	.w5(32'h3c50c510),
	.w6(32'h3ca6c254),
	.w7(32'h3cc6e97f),
	.w8(32'h3c28b04c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa775bc),
	.w1(32'h3c222d48),
	.w2(32'h3bec390b),
	.w3(32'h3c38239f),
	.w4(32'h3c28dbfa),
	.w5(32'hbd704aab),
	.w6(32'hba9813be),
	.w7(32'hbc7e280d),
	.w8(32'h3c945e09),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3cede),
	.w1(32'hbcb46537),
	.w2(32'hbd432203),
	.w3(32'hbcf2c596),
	.w4(32'hbc559a29),
	.w5(32'hba7e3466),
	.w6(32'hbcd5e3ad),
	.w7(32'hbced7ffe),
	.w8(32'hbcf873f6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc554eb9),
	.w1(32'h3d90b222),
	.w2(32'hbe1e9b49),
	.w3(32'hbc155676),
	.w4(32'hbcb4163f),
	.w5(32'hbe2a43ff),
	.w6(32'h3d8f07e2),
	.w7(32'h3dc382d2),
	.w8(32'h3d22aeb6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcbef5e),
	.w1(32'hbc925e7e),
	.w2(32'hbc8ec3aa),
	.w3(32'hb9505b3c),
	.w4(32'hbb34b79f),
	.w5(32'hbc2ffda2),
	.w6(32'h3b2a8dbc),
	.w7(32'hbb8ecfde),
	.w8(32'h3b7840ab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c996c62),
	.w1(32'hbd365042),
	.w2(32'hbcf8c756),
	.w3(32'hbc180f15),
	.w4(32'hbc5fb398),
	.w5(32'hbd063ccb),
	.w6(32'h3b1c008e),
	.w7(32'h3ca7d9dd),
	.w8(32'h3bde68cf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd365222),
	.w1(32'hbcca16ad),
	.w2(32'h3d54ed5e),
	.w3(32'h3c410d6e),
	.w4(32'hbd3d0fb4),
	.w5(32'h3d36d098),
	.w6(32'hbd076fc2),
	.w7(32'hbccff1d9),
	.w8(32'hbc4d9351),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d017da4),
	.w1(32'h3a4970b0),
	.w2(32'h3cc683d9),
	.w3(32'h3b5d85da),
	.w4(32'hba7de57c),
	.w5(32'hbd3d4a8a),
	.w6(32'h3a88dffc),
	.w7(32'h3c81b2a3),
	.w8(32'h3b99cd98),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581918),
	.w1(32'hbca50f4d),
	.w2(32'hbc7e3106),
	.w3(32'h3c4c5577),
	.w4(32'hba29c6f5),
	.w5(32'h3c0a2e2b),
	.w6(32'hbc1bce1e),
	.w7(32'hbc33f7cc),
	.w8(32'h3ca64b3a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d178735),
	.w1(32'h3c024ac4),
	.w2(32'h3be70509),
	.w3(32'h3c39f076),
	.w4(32'hbbd9d246),
	.w5(32'h3a33efbe),
	.w6(32'h3c064012),
	.w7(32'h3c204515),
	.w8(32'h3b542902),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909651),
	.w1(32'h3ac1f953),
	.w2(32'hbc2bb2ea),
	.w3(32'h3cafadea),
	.w4(32'hbbb9ee78),
	.w5(32'hbc1e4c34),
	.w6(32'h3cdae7e6),
	.w7(32'h3c86c28e),
	.w8(32'h3c503286),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1645c),
	.w1(32'hbba431c5),
	.w2(32'h3b6bd108),
	.w3(32'h3b75f97e),
	.w4(32'hba6cc680),
	.w5(32'hbc036949),
	.w6(32'hbb9f09cf),
	.w7(32'h3be88b79),
	.w8(32'h3b10dba2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6c94),
	.w1(32'h3c19c762),
	.w2(32'h3c3554c0),
	.w3(32'hbbeae855),
	.w4(32'hbad9c28c),
	.w5(32'h3b85f065),
	.w6(32'h3b5144a1),
	.w7(32'h3bad6bff),
	.w8(32'h3b90169a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39f868),
	.w1(32'hbbe2dd8f),
	.w2(32'hbc33fd4c),
	.w3(32'h3bc348df),
	.w4(32'hbbc88f19),
	.w5(32'hbca07345),
	.w6(32'hbc384a30),
	.w7(32'hbc73f747),
	.w8(32'h3abce0b1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca39c1),
	.w1(32'hbc13da13),
	.w2(32'hbc815d17),
	.w3(32'hbb68cdb0),
	.w4(32'hbc8c35f6),
	.w5(32'hbc4b7852),
	.w6(32'hbc000d71),
	.w7(32'hbc13d58f),
	.w8(32'hbc549bb5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd44a95),
	.w1(32'hbb41b91e),
	.w2(32'h3b111531),
	.w3(32'hbc3b5c92),
	.w4(32'hbb27d0e5),
	.w5(32'h3b022b03),
	.w6(32'hbba53456),
	.w7(32'hbabeb36c),
	.w8(32'hbb79584a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab32005),
	.w1(32'hbcb527a2),
	.w2(32'h3ac21bc9),
	.w3(32'hbb0c3173),
	.w4(32'hbc908a4e),
	.w5(32'hbc073961),
	.w6(32'hbb280ffc),
	.w7(32'h3c15aeba),
	.w8(32'h3c96c5d5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47ea80),
	.w1(32'h3c89cb5a),
	.w2(32'h3cc7055f),
	.w3(32'hbc2105be),
	.w4(32'h3c4fc16d),
	.w5(32'h3ca0b5e3),
	.w6(32'h3c4d5433),
	.w7(32'h3c977dc1),
	.w8(32'h3c5809a2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6df97),
	.w1(32'hbd1b0b5a),
	.w2(32'hbd32a04b),
	.w3(32'h3c8976e6),
	.w4(32'hbc48cffb),
	.w5(32'hbcd0ab9b),
	.w6(32'hbbb317be),
	.w7(32'hbc9b146c),
	.w8(32'hbcae661b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1c51),
	.w1(32'hbb0011f7),
	.w2(32'h3bc93c48),
	.w3(32'hbc4a6efc),
	.w4(32'hbbbe2d86),
	.w5(32'hba6ad8de),
	.w6(32'hb8ba7623),
	.w7(32'h3ade83b0),
	.w8(32'hbbe8f0ea),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e4b0),
	.w1(32'h3b8df2a2),
	.w2(32'h3c249821),
	.w3(32'hbbd6dcf4),
	.w4(32'h3a6d47f3),
	.w5(32'h3bbec2e0),
	.w6(32'h3ac2b920),
	.w7(32'h3b823751),
	.w8(32'h3af50685),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f9554),
	.w1(32'hbc5d12dd),
	.w2(32'hbc52dd09),
	.w3(32'h3c23fef0),
	.w4(32'hbc1ed36e),
	.w5(32'hbbec342d),
	.w6(32'hbb881d3a),
	.w7(32'hbc2ecee7),
	.w8(32'hbc323be4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a04d3),
	.w1(32'hbb52bfc1),
	.w2(32'hbc78dc91),
	.w3(32'hbaca5384),
	.w4(32'hbc3a3531),
	.w5(32'hb9a378d2),
	.w6(32'h3be24e0f),
	.w7(32'h3b3cf092),
	.w8(32'hbc18f0d8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0745),
	.w1(32'h3c9480ab),
	.w2(32'h3d41b79e),
	.w3(32'h3bc431d9),
	.w4(32'h3c7c4f6e),
	.w5(32'h3c8a75a0),
	.w6(32'h3bca2e39),
	.w7(32'h3c82f539),
	.w8(32'h3c1a0ced),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca38001),
	.w1(32'h3ad4e003),
	.w2(32'h3b9421ae),
	.w3(32'h3a629ded),
	.w4(32'hbbc70614),
	.w5(32'hbb9b040d),
	.w6(32'h3c0f113f),
	.w7(32'h3c83a64f),
	.w8(32'h3a867cd1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae27f4),
	.w1(32'hbcb3f269),
	.w2(32'hbcb0faaf),
	.w3(32'hbbef7e16),
	.w4(32'h3c4ac397),
	.w5(32'hbc3368cf),
	.w6(32'hbc167597),
	.w7(32'h3bb141e2),
	.w8(32'h3cb17d24),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0960a1),
	.w1(32'hbbf027d7),
	.w2(32'h3bee8f20),
	.w3(32'hbccd06ad),
	.w4(32'hbc789e60),
	.w5(32'h3baf62d0),
	.w6(32'h3caeb2a5),
	.w7(32'h3cbc5f31),
	.w8(32'h3cc0ab8e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffc3f2),
	.w1(32'h3b10ffbd),
	.w2(32'hbc5de600),
	.w3(32'hbb1b5142),
	.w4(32'h3ac119c7),
	.w5(32'hbc1eb26d),
	.w6(32'h3bca17f9),
	.w7(32'hbb83b6be),
	.w8(32'hbc495d53),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb4d9e1),
	.w1(32'h3b8ecec4),
	.w2(32'hbb1dd99e),
	.w3(32'hbc01053e),
	.w4(32'h3c55f17e),
	.w5(32'h3bbd17b3),
	.w6(32'h3c9bbedc),
	.w7(32'h3c884f46),
	.w8(32'h3b64bdca),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69a756),
	.w1(32'hbbdcd3aa),
	.w2(32'hbb82ff52),
	.w3(32'hbc8812bc),
	.w4(32'hbc0925dd),
	.w5(32'hbb4addca),
	.w6(32'hbaef2858),
	.w7(32'hb9ce7c5b),
	.w8(32'hbb1c7975),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc976295),
	.w1(32'hbcc02112),
	.w2(32'h3c9780fb),
	.w3(32'hbc92fdc8),
	.w4(32'hbc8c1412),
	.w5(32'h3ab75e20),
	.w6(32'hbc83b88d),
	.w7(32'hba051677),
	.w8(32'hbc956619),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd90d8b),
	.w1(32'hbceb2183),
	.w2(32'hbd08c8a2),
	.w3(32'hbb5b1ec4),
	.w4(32'hbb1ccb20),
	.w5(32'hbcac26d2),
	.w6(32'hba4128ee),
	.w7(32'hbc2beeee),
	.w8(32'hbbc0cf23),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ae0a8),
	.w1(32'hbc1e72d7),
	.w2(32'h3bb56f28),
	.w3(32'hbc5e7758),
	.w4(32'hbc4f1356),
	.w5(32'hba9081b8),
	.w6(32'hb90d6f86),
	.w7(32'h3bd830ec),
	.w8(32'h3ad68167),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f24d),
	.w1(32'h3c0d3b12),
	.w2(32'hb99ff8d5),
	.w3(32'hb8805faf),
	.w4(32'h3b0cc7a6),
	.w5(32'hba92c001),
	.w6(32'h3bdbd534),
	.w7(32'h3bf66f36),
	.w8(32'h3b3476bd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cd482),
	.w1(32'h3ca23d62),
	.w2(32'h3c6037f9),
	.w3(32'h3c47295f),
	.w4(32'h3c5fedff),
	.w5(32'h3bc44952),
	.w6(32'h3d019cc7),
	.w7(32'h3c926584),
	.w8(32'h3c80621d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53644c),
	.w1(32'hbca9a7d8),
	.w2(32'hbc7fbc06),
	.w3(32'hbc13a8ab),
	.w4(32'hbbb52c48),
	.w5(32'hbb911e38),
	.w6(32'hbcaa8ffc),
	.w7(32'hbc5ebbb0),
	.w8(32'hbca1cc5a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4da069),
	.w1(32'h3b7a546b),
	.w2(32'hbbc914b9),
	.w3(32'hb94d8c1f),
	.w4(32'hbbc121bd),
	.w5(32'hbc4ba049),
	.w6(32'hbbd1c0fa),
	.w7(32'hbc98a6e7),
	.w8(32'hba7adc18),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5837f6),
	.w1(32'h3c745c59),
	.w2(32'h3bd41878),
	.w3(32'h3c7d3005),
	.w4(32'h3a4945dd),
	.w5(32'hbbc4736b),
	.w6(32'h3c0a57dc),
	.w7(32'hba504b36),
	.w8(32'h3c174da4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1ea63),
	.w1(32'hba5c950e),
	.w2(32'h3ba99e5a),
	.w3(32'h3cfb3176),
	.w4(32'hba0c665c),
	.w5(32'h3c2ea785),
	.w6(32'h3d00ed09),
	.w7(32'h3d17ef9e),
	.w8(32'h3ce0b025),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d104b),
	.w1(32'hbc89ba79),
	.w2(32'h3b2ec65d),
	.w3(32'hbc08c98c),
	.w4(32'h3a434d46),
	.w5(32'h3c672925),
	.w6(32'hbc83a9f3),
	.w7(32'hbc261cd6),
	.w8(32'h3bdf938a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca93cd0),
	.w1(32'h3c3e2c34),
	.w2(32'hbbba45ed),
	.w3(32'h3c4ffac0),
	.w4(32'h3c0d59e5),
	.w5(32'hbb6dfe4d),
	.w6(32'h3cc0d714),
	.w7(32'h3c605ceb),
	.w8(32'h3cd850be),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30d913),
	.w1(32'h3d19264a),
	.w2(32'h3cad117b),
	.w3(32'h3cce1cd7),
	.w4(32'h3cc2b0ae),
	.w5(32'hb9bd8517),
	.w6(32'h3c9ac406),
	.w7(32'h3c7f9d18),
	.w8(32'h3bb123e9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5b36),
	.w1(32'hbba4d231),
	.w2(32'hbbc5e88e),
	.w3(32'hbb7a89e2),
	.w4(32'hbb910fd0),
	.w5(32'hbbcdae57),
	.w6(32'hbb9f080b),
	.w7(32'hbbba4a32),
	.w8(32'hbbd00e68),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule