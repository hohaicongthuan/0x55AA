module layer_10_featuremap_141(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb694f2a),
	.w1(32'h3b2df4a2),
	.w2(32'hbbbfd05b),
	.w3(32'hbb54068d),
	.w4(32'h3be76563),
	.w5(32'hbb432a01),
	.w6(32'h3aff6921),
	.w7(32'hba860e7e),
	.w8(32'hba0351f7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc255a01),
	.w1(32'h3b5539b3),
	.w2(32'hba3b1811),
	.w3(32'hbb86095f),
	.w4(32'h3b9e1065),
	.w5(32'h3ac694dd),
	.w6(32'hbb42fc87),
	.w7(32'h3bafce63),
	.w8(32'hbb334d44),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215a5d),
	.w1(32'hb8a81221),
	.w2(32'h3a18bd4c),
	.w3(32'h3a320417),
	.w4(32'hbac0bf95),
	.w5(32'hba5ce414),
	.w6(32'hba878e02),
	.w7(32'hba400acc),
	.w8(32'hba612108),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398aaaaa),
	.w1(32'h3b44ccab),
	.w2(32'h3a178f55),
	.w3(32'hbaff8d05),
	.w4(32'hb89d5fd7),
	.w5(32'h3b0deb62),
	.w6(32'h3b845a9e),
	.w7(32'h3b70e6f4),
	.w8(32'h3bbf2f95),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2cd5),
	.w1(32'h3a28ae88),
	.w2(32'h3a1b4776),
	.w3(32'h3ad6d95d),
	.w4(32'h3924a590),
	.w5(32'h3ac5484b),
	.w6(32'h3b14bbaf),
	.w7(32'h3ad702bc),
	.w8(32'hb96b469d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500ac9),
	.w1(32'hbad06bcd),
	.w2(32'hbb1a81ec),
	.w3(32'h3a541de5),
	.w4(32'hbb2ed8ea),
	.w5(32'hbaf9711c),
	.w6(32'hbadeb61b),
	.w7(32'hbaff084d),
	.w8(32'hbb11418c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0d338),
	.w1(32'hbb9f8700),
	.w2(32'hbb8b6d13),
	.w3(32'hba8bf444),
	.w4(32'hbc10ee9d),
	.w5(32'hbbd111a0),
	.w6(32'hb886bba9),
	.w7(32'hbb83f0ba),
	.w8(32'hbc1787fd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69b634),
	.w1(32'hbc512459),
	.w2(32'hbc0478f6),
	.w3(32'hbcbeeb54),
	.w4(32'hbca76b9d),
	.w5(32'hbc384f7c),
	.w6(32'hbc96e463),
	.w7(32'hbc872385),
	.w8(32'hbc706836),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698e6b),
	.w1(32'hbad4f041),
	.w2(32'hbadc7c1f),
	.w3(32'hb81f160c),
	.w4(32'hb983a279),
	.w5(32'hbadc187e),
	.w6(32'hbadad6de),
	.w7(32'hbb219956),
	.w8(32'hbb801a94),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b18f),
	.w1(32'hbbca7bd7),
	.w2(32'hbc800df4),
	.w3(32'hbc1c1d26),
	.w4(32'hbb49b3ac),
	.w5(32'hbc45e34f),
	.w6(32'hbb2f5ade),
	.w7(32'hb9c9be13),
	.w8(32'hbc8bea3b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8584a7),
	.w1(32'h3abf89dc),
	.w2(32'hb9ea248f),
	.w3(32'hba151ee9),
	.w4(32'h3a249481),
	.w5(32'hba687652),
	.w6(32'h3b034b43),
	.w7(32'h3b77b00d),
	.w8(32'h3b91ccaf),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2b37d),
	.w1(32'h3c1bb4f6),
	.w2(32'hbc0be2e6),
	.w3(32'h3b81a548),
	.w4(32'h3bd156ab),
	.w5(32'hbbccb973),
	.w6(32'h3bd53aa2),
	.w7(32'h3c0aeb02),
	.w8(32'hbb83e6e9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36424e),
	.w1(32'hbbe01876),
	.w2(32'hbc372aa2),
	.w3(32'hbc6f8fa4),
	.w4(32'hbc4a4031),
	.w5(32'hbc60cb55),
	.w6(32'hbbede6d6),
	.w7(32'hbc1b79a7),
	.w8(32'hbca7f551),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c17e6),
	.w1(32'hbb9d0f72),
	.w2(32'hbc12563f),
	.w3(32'hbb4cbfcd),
	.w4(32'hba6eb03d),
	.w5(32'hbba57621),
	.w6(32'hbb1bf2cd),
	.w7(32'hbb947bff),
	.w8(32'hb9f4082c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf59817),
	.w1(32'hb8e52a78),
	.w2(32'hbc244177),
	.w3(32'hbb067a1c),
	.w4(32'h3b43fbb7),
	.w5(32'hbb142292),
	.w6(32'h3b514bd6),
	.w7(32'h3b04ffb9),
	.w8(32'hbbd48fad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5406c4),
	.w1(32'hbc4d3d5d),
	.w2(32'hbc9adf37),
	.w3(32'hbbbfb25e),
	.w4(32'hbb93d69b),
	.w5(32'hbc54b357),
	.w6(32'hbc218875),
	.w7(32'hbc0d8c8b),
	.w8(32'hbc99b72c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb503886),
	.w1(32'hbad5b252),
	.w2(32'hbaa29db2),
	.w3(32'hbb2139fc),
	.w4(32'hba750a58),
	.w5(32'hb9bcaa50),
	.w6(32'hbb3b6cab),
	.w7(32'hba1cb0ac),
	.w8(32'h3b0754a6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e64f2),
	.w1(32'hbbfd9d71),
	.w2(32'hbba2e981),
	.w3(32'hbc202d2d),
	.w4(32'hbb95973b),
	.w5(32'hbbcdc1e3),
	.w6(32'hbc703d06),
	.w7(32'hbc3f18f3),
	.w8(32'hbc6e362c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55863f),
	.w1(32'hbc04a98a),
	.w2(32'hbbf7294d),
	.w3(32'hbc252f69),
	.w4(32'hbc375948),
	.w5(32'hbc23e3a3),
	.w6(32'hbc291516),
	.w7(32'hbc471d40),
	.w8(32'hbc7b9e0e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987ae7e),
	.w1(32'hba9dcfb1),
	.w2(32'hbac3afc7),
	.w3(32'hba71b611),
	.w4(32'hba1c5ee2),
	.w5(32'hbaa9d4d0),
	.w6(32'hbaa9ced6),
	.w7(32'hbaa88b8a),
	.w8(32'hbad48afe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8606ae),
	.w1(32'hb906237d),
	.w2(32'hb9b6cc76),
	.w3(32'hba7a117f),
	.w4(32'hb96e8af6),
	.w5(32'hb9b5af5d),
	.w6(32'h39befa02),
	.w7(32'hba030bd6),
	.w8(32'hb8c3d553),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a202),
	.w1(32'h3b755589),
	.w2(32'hbbc86f91),
	.w3(32'h39e49cfa),
	.w4(32'h3bfcd0fa),
	.w5(32'hbb2f1ab1),
	.w6(32'hba4c7ecb),
	.w7(32'h3affca83),
	.w8(32'hba66cc01),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63187d),
	.w1(32'hbb9da33b),
	.w2(32'hbd07c595),
	.w3(32'hbb1a0dcd),
	.w4(32'h3bccefe9),
	.w5(32'hbcc4d12b),
	.w6(32'hbc2e8e1c),
	.w7(32'hbb6c1f32),
	.w8(32'hbd0aaea3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03310),
	.w1(32'hba4ed806),
	.w2(32'hbc922910),
	.w3(32'h3ba1b655),
	.w4(32'h3c16e512),
	.w5(32'hbc29308c),
	.w6(32'h3b1045d0),
	.w7(32'h3bec088e),
	.w8(32'hbc74f55e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40fe48),
	.w1(32'h3bc928c3),
	.w2(32'hbc6e53f8),
	.w3(32'hbc157d4b),
	.w4(32'h3c1dc0f4),
	.w5(32'hbc1a890a),
	.w6(32'hbc522013),
	.w7(32'hba69116b),
	.w8(32'hbc9baa45),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215cd7),
	.w1(32'hba04af3d),
	.w2(32'hb9cf4ed8),
	.w3(32'h3aa7871f),
	.w4(32'h3a44b1ea),
	.w5(32'h3a1058ce),
	.w6(32'h3ae41622),
	.w7(32'hba50a8cd),
	.w8(32'hb9b5c0b9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac768e7),
	.w1(32'h384a36c6),
	.w2(32'h3a45a341),
	.w3(32'h3aea8794),
	.w4(32'h38bc9e5c),
	.w5(32'h39cdde01),
	.w6(32'hb9add180),
	.w7(32'hb8ae6f01),
	.w8(32'h3977a19b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a1a5b),
	.w1(32'h3c00dfb1),
	.w2(32'hbb505544),
	.w3(32'hba43c94f),
	.w4(32'h3c0d7c09),
	.w5(32'h3b48eb2d),
	.w6(32'hbb7daaea),
	.w7(32'h3a3d939b),
	.w8(32'hba415068),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdcacb),
	.w1(32'h3c1f9d9a),
	.w2(32'hbb865eb2),
	.w3(32'h3b63852d),
	.w4(32'h3c3544ab),
	.w5(32'hbb6c2529),
	.w6(32'h3bbcf52d),
	.w7(32'h3c049081),
	.w8(32'h3ad80b11),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d85a1),
	.w1(32'h3b872cea),
	.w2(32'hbc22256a),
	.w3(32'hb9f2610c),
	.w4(32'h3bda4cd5),
	.w5(32'hbbe1841a),
	.w6(32'hbb61efe8),
	.w7(32'h3b4b6679),
	.w8(32'hbc0a1dbc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98746b0),
	.w1(32'hb67a0903),
	.w2(32'hb83dc765),
	.w3(32'hba251140),
	.w4(32'h38dd2050),
	.w5(32'hb959cced),
	.w6(32'h38f53a4c),
	.w7(32'hb86feee6),
	.w8(32'h3916d6d5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06af5e),
	.w1(32'hb98cec81),
	.w2(32'h38118941),
	.w3(32'hb9e5b611),
	.w4(32'hb8425460),
	.w5(32'h391b1cbe),
	.w6(32'hb9843f23),
	.w7(32'hb97ed9e2),
	.w8(32'h383a20da),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c010),
	.w1(32'h3a16aa9d),
	.w2(32'hbbeebe91),
	.w3(32'h3ab97236),
	.w4(32'h3bd913e0),
	.w5(32'hbb7058cf),
	.w6(32'h3bb0864d),
	.w7(32'h3bed91b1),
	.w8(32'hbb3d17eb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78080a),
	.w1(32'h3afef927),
	.w2(32'hbb2b0793),
	.w3(32'hba0c4bd9),
	.w4(32'h3ba55208),
	.w5(32'hbab6019e),
	.w6(32'hbb1201d6),
	.w7(32'h3ade41d2),
	.w8(32'hbbdfac5b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9c94),
	.w1(32'h3affc8f1),
	.w2(32'h3b0fd207),
	.w3(32'hbb9a0754),
	.w4(32'h3890f53a),
	.w5(32'h3aff3f3b),
	.w6(32'h39ede532),
	.w7(32'h3a9148a5),
	.w8(32'hbb4e7828),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa89756),
	.w1(32'hbb5e2cd3),
	.w2(32'hbba13ac3),
	.w3(32'h396e6545),
	.w4(32'hbb834b36),
	.w5(32'hbb93abcc),
	.w6(32'h3aac140e),
	.w7(32'hbb25eadf),
	.w8(32'hbb71b867),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5836e9),
	.w1(32'h3b9ff7ef),
	.w2(32'hbc3b48d9),
	.w3(32'h3bab0d99),
	.w4(32'h3c216722),
	.w5(32'hbaa7b702),
	.w6(32'h3c328d9e),
	.w7(32'h3ca22697),
	.w8(32'hbbec05af),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ffca),
	.w1(32'h3cb5cb83),
	.w2(32'hbc04b0a8),
	.w3(32'h3a261e38),
	.w4(32'h3d0b5bbf),
	.w5(32'h3a922cd8),
	.w6(32'hbc6a193a),
	.w7(32'h3ce2c7cf),
	.w8(32'hba302f28),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39921621),
	.w1(32'h3ca40203),
	.w2(32'hbc82c66e),
	.w3(32'h3ba54e10),
	.w4(32'h3cd5a4a9),
	.w5(32'hbbe5061a),
	.w6(32'hbc64c859),
	.w7(32'h3c30e598),
	.w8(32'hbc437c8f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1e9f),
	.w1(32'h3a03abfb),
	.w2(32'h3a090e37),
	.w3(32'hbb8e8795),
	.w4(32'h3a736ee7),
	.w5(32'h3aec40db),
	.w6(32'hbbc39d41),
	.w7(32'hb832a92c),
	.w8(32'hbb364c5a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf18aa8),
	.w1(32'hbb8613e2),
	.w2(32'hbb55098d),
	.w3(32'hbb1e3ac8),
	.w4(32'hbb83eede),
	.w5(32'hbb5be815),
	.w6(32'hbb1f11d8),
	.w7(32'hbb2899a3),
	.w8(32'hbb094086),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb201fad),
	.w1(32'hbb4cbd10),
	.w2(32'hbbd93cfc),
	.w3(32'hbb475625),
	.w4(32'hbb610891),
	.w5(32'hbba265ed),
	.w6(32'hbab9a01e),
	.w7(32'hbb20c667),
	.w8(32'hbaec78ca),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042c97),
	.w1(32'h3ba048a6),
	.w2(32'hbb297160),
	.w3(32'hbc0f3556),
	.w4(32'h3bd73b40),
	.w5(32'hbb32e9b4),
	.w6(32'h3a575cd7),
	.w7(32'h3c33c9ae),
	.w8(32'h39b89e80),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b0ad1),
	.w1(32'hbaa609d0),
	.w2(32'hbc1bf78a),
	.w3(32'hbc0d4e11),
	.w4(32'hbad08e57),
	.w5(32'hbbec5a60),
	.w6(32'hbbf53497),
	.w7(32'hbb44b3ed),
	.w8(32'hbca44b93),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcfc3b),
	.w1(32'hba111eba),
	.w2(32'hbc9a81dc),
	.w3(32'h378247fd),
	.w4(32'h3c2c0455),
	.w5(32'hbc37b743),
	.w6(32'hba8b3b66),
	.w7(32'h3c0f4128),
	.w8(32'hbc536678),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5359f2),
	.w1(32'hbb0e7463),
	.w2(32'hbc962262),
	.w3(32'hbba67889),
	.w4(32'h3bc689c6),
	.w5(32'hbc530539),
	.w6(32'hbb2cbaff),
	.w7(32'h3b96b4b1),
	.w8(32'hbca453bf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9da082),
	.w1(32'hbb6f8995),
	.w2(32'hbc875165),
	.w3(32'hbc3aa6ea),
	.w4(32'h3b26fe98),
	.w5(32'hbc291e2d),
	.w6(32'h3aeea6b8),
	.w7(32'h3a948fae),
	.w8(32'hbc41896b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894619),
	.w1(32'hbc800b2f),
	.w2(32'hbc800352),
	.w3(32'hbcb018ca),
	.w4(32'hbcd5644e),
	.w5(32'hbcb49825),
	.w6(32'hbcd1f0d3),
	.w7(32'hbd208923),
	.w8(32'hbcf67e55),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad555c9),
	.w1(32'h3a65f951),
	.w2(32'h39cd29e5),
	.w3(32'h3b09ed0d),
	.w4(32'h3a27a95f),
	.w5(32'hb94407be),
	.w6(32'h3a73b4e9),
	.w7(32'hb93144cc),
	.w8(32'hba6951f3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b6407),
	.w1(32'hbb7006c8),
	.w2(32'hbb95c55e),
	.w3(32'hb99f8de7),
	.w4(32'hbb5bc4e3),
	.w5(32'hbba29b95),
	.w6(32'hbacdcc40),
	.w7(32'hbb9044e8),
	.w8(32'hbbd416a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a910e9f),
	.w1(32'hbb5a3089),
	.w2(32'hbb351193),
	.w3(32'h3aacf67a),
	.w4(32'hbb875f95),
	.w5(32'hbb9afba0),
	.w6(32'hb81e7d8c),
	.w7(32'hba3653da),
	.w8(32'hbb25379c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0dea),
	.w1(32'hbae7dcca),
	.w2(32'hbc822a54),
	.w3(32'hbc02fa80),
	.w4(32'h3c02135f),
	.w5(32'hbbbcc713),
	.w6(32'h3baa695b),
	.w7(32'h3b781483),
	.w8(32'hbbb2f48b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39808d90),
	.w1(32'hba1bfb6c),
	.w2(32'hbb32d2ab),
	.w3(32'hbac0b22e),
	.w4(32'h3850c5dd),
	.w5(32'hbac72ae3),
	.w6(32'hb863eba1),
	.w7(32'h3ad24dda),
	.w8(32'hbb044ea4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2339),
	.w1(32'hbb84343c),
	.w2(32'hbc164237),
	.w3(32'hbb1ebcc5),
	.w4(32'hbb1acbb4),
	.w5(32'hbbca2c79),
	.w6(32'hbb2780a9),
	.w7(32'hbbb2af98),
	.w8(32'hbc854750),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ab8a),
	.w1(32'h3bdadd5c),
	.w2(32'h3bacd59a),
	.w3(32'h3af984b0),
	.w4(32'h3ba67f11),
	.w5(32'h3ba68eb1),
	.w6(32'h3b4cbc3a),
	.w7(32'h3bb11ae8),
	.w8(32'h3b718355),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed8076),
	.w1(32'hbb60809d),
	.w2(32'hbb2381e5),
	.w3(32'h3bf27444),
	.w4(32'hbb104088),
	.w5(32'hbaea52b5),
	.w6(32'hbb2f0edb),
	.w7(32'hbace8d0f),
	.w8(32'h39084d09),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb108725),
	.w1(32'h3aa49674),
	.w2(32'h3a7ab0f4),
	.w3(32'hbb04cc65),
	.w4(32'h3a827ec0),
	.w5(32'h3a1170e4),
	.w6(32'h3aa43389),
	.w7(32'h3af3817a),
	.w8(32'h3b0263bf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9918db),
	.w1(32'h39eaf389),
	.w2(32'h3a2c825f),
	.w3(32'h38775871),
	.w4(32'hba22d50d),
	.w5(32'h3ac871fd),
	.w6(32'h3b5530e0),
	.w7(32'h3b8c8d71),
	.w8(32'h3b2e638b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebf839),
	.w1(32'h3bc0d690),
	.w2(32'h3aa2c38e),
	.w3(32'h3b3f21da),
	.w4(32'h3baeddab),
	.w5(32'h3b19a570),
	.w6(32'hb847286b),
	.w7(32'h3ba864f7),
	.w8(32'hba151fe9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d2127),
	.w1(32'hbac4ab7e),
	.w2(32'hbacc510f),
	.w3(32'hbae8b231),
	.w4(32'hba45b348),
	.w5(32'hba47ce1f),
	.w6(32'hbab5280a),
	.w7(32'hb885324f),
	.w8(32'hba36fd0d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd2d95),
	.w1(32'hbb6fa61a),
	.w2(32'hbc0de9ed),
	.w3(32'hbbde8e47),
	.w4(32'hbb9a660c),
	.w5(32'hbbe3a225),
	.w6(32'hbb845cc6),
	.w7(32'hbb4ff0ce),
	.w8(32'hbc26a25b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1876d2),
	.w1(32'hbb79d74c),
	.w2(32'hbb947ee8),
	.w3(32'hbc209726),
	.w4(32'hbaa204a3),
	.w5(32'hbb19a48a),
	.w6(32'hbbb23b49),
	.w7(32'hbafa257c),
	.w8(32'hba5e22a0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f0f7b),
	.w1(32'h3ba9bf73),
	.w2(32'h3b15d6fd),
	.w3(32'hba290ed2),
	.w4(32'h3be40884),
	.w5(32'h3b0e1c7a),
	.w6(32'h3c05b918),
	.w7(32'h3b9307c7),
	.w8(32'h3b237bb2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22f765),
	.w1(32'h3b185ec1),
	.w2(32'h3b407df4),
	.w3(32'h3b20284a),
	.w4(32'h3a8027ad),
	.w5(32'h3b12bd11),
	.w6(32'h3ad849cc),
	.w7(32'h3b24b232),
	.w8(32'hb829c895),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3b20c),
	.w1(32'hba222c64),
	.w2(32'hb968ab48),
	.w3(32'hba31c85d),
	.w4(32'hbb0f85f6),
	.w5(32'hba08f4b6),
	.w6(32'hba7a8c36),
	.w7(32'h38310cb9),
	.w8(32'hba20a6e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97badb7),
	.w1(32'hba40c4d0),
	.w2(32'hbaa336fe),
	.w3(32'hbacfca72),
	.w4(32'hba99e013),
	.w5(32'hb8c512c3),
	.w6(32'h3a424695),
	.w7(32'h3a4d026b),
	.w8(32'h3ac1ab8b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fb018),
	.w1(32'hbc439a68),
	.w2(32'hbc2d842c),
	.w3(32'hbc1c8c33),
	.w4(32'hbc3bf8d9),
	.w5(32'hbba36e89),
	.w6(32'hbc2360aa),
	.w7(32'hbc380cfe),
	.w8(32'hbbf818c7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc16b8),
	.w1(32'hbb1f69a5),
	.w2(32'hbcad5865),
	.w3(32'h3b7a06a1),
	.w4(32'h3bdcec48),
	.w5(32'hbc7ed093),
	.w6(32'h3ade9684),
	.w7(32'h3bb841f5),
	.w8(32'hbc8dad6b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f176a),
	.w1(32'hbb015faf),
	.w2(32'hbc8fdce7),
	.w3(32'h3a04cb5b),
	.w4(32'h3c014f10),
	.w5(32'hbc31dbfb),
	.w6(32'hbbf56660),
	.w7(32'h3aef4653),
	.w8(32'hbc94899c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc724920),
	.w1(32'h3b7d00cc),
	.w2(32'hbcf30020),
	.w3(32'hbc00fbf7),
	.w4(32'h3c3bc225),
	.w5(32'hbcbc81cd),
	.w6(32'hbc51d229),
	.w7(32'h3c35ead8),
	.w8(32'hbcc7f770),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15e626),
	.w1(32'h3b81d151),
	.w2(32'h3b891ef5),
	.w3(32'hbb36d785),
	.w4(32'h3afaf11a),
	.w5(32'h3b5cbc6e),
	.w6(32'h3b3c964a),
	.w7(32'h3b6ad1f3),
	.w8(32'h3a8e8578),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1821aa),
	.w1(32'hba94de4f),
	.w2(32'hba398070),
	.w3(32'h3724e287),
	.w4(32'hbae5cb3f),
	.w5(32'hba83446a),
	.w6(32'hba882ae7),
	.w7(32'hbaa904cb),
	.w8(32'hba942105),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad96355),
	.w1(32'hbad7b080),
	.w2(32'hbab527b8),
	.w3(32'hbaeb2d25),
	.w4(32'hbae7a90e),
	.w5(32'hbab0c4a4),
	.w6(32'hba93c810),
	.w7(32'hbacff4d9),
	.w8(32'hbaafb369),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892360),
	.w1(32'hb978f251),
	.w2(32'hbaf38131),
	.w3(32'hbbb27992),
	.w4(32'h3a64ff63),
	.w5(32'hba4734b1),
	.w6(32'hbba1636a),
	.w7(32'hbab65cba),
	.w8(32'hbabc96f6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92145ac),
	.w1(32'hbae2a2b3),
	.w2(32'hbb197994),
	.w3(32'hb9e27293),
	.w4(32'hbb034b72),
	.w5(32'hbad9c04a),
	.w6(32'hbb138315),
	.w7(32'hbb2dffa7),
	.w8(32'hbb485e8a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813deb),
	.w1(32'hbbce5755),
	.w2(32'hbc12adb2),
	.w3(32'hbc135cbe),
	.w4(32'hbbcc4584),
	.w5(32'hbb94a2fb),
	.w6(32'hbb6555a7),
	.w7(32'hbbefe6b3),
	.w8(32'hbb76a665),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca11556),
	.w1(32'hbc2b1c18),
	.w2(32'hbc855341),
	.w3(32'hbc0f768b),
	.w4(32'hbc245158),
	.w5(32'hbc5db95d),
	.w6(32'hbbfe3792),
	.w7(32'hbbd1e4db),
	.w8(32'hbc84f288),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d8a47),
	.w1(32'hbb70760f),
	.w2(32'hbc4b5d77),
	.w3(32'hbc910cc7),
	.w4(32'hbbdf5cd2),
	.w5(32'hbc362a8e),
	.w6(32'hbc87bff3),
	.w7(32'hbc696657),
	.w8(32'hbc8cf834),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c32e),
	.w1(32'hb8e05b8f),
	.w2(32'hbbaa99f3),
	.w3(32'hbb1c21f2),
	.w4(32'h3b5e5ead),
	.w5(32'hbb0e70eb),
	.w6(32'hba17c7e9),
	.w7(32'h3b24cfce),
	.w8(32'hbac47942),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8512c),
	.w1(32'hbb218d0f),
	.w2(32'hbbbd244d),
	.w3(32'h3b9fd61e),
	.w4(32'hbb04ff4c),
	.w5(32'hbb75b1dc),
	.w6(32'h3afe4cbc),
	.w7(32'hbab41a4a),
	.w8(32'hbbc0b611),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75decb),
	.w1(32'hbb257572),
	.w2(32'hbc04e67b),
	.w3(32'hb8fd39d8),
	.w4(32'h3b08d5aa),
	.w5(32'hbb93a3de),
	.w6(32'hb90a7c9a),
	.w7(32'h3b827a1f),
	.w8(32'hbb569fe4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6bb63),
	.w1(32'hbc515bb9),
	.w2(32'hbc73022c),
	.w3(32'hbc22000d),
	.w4(32'hbc6e69eb),
	.w5(32'hbc76f8b1),
	.w6(32'hbc5c97fa),
	.w7(32'hbc83d481),
	.w8(32'hbc822ecb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8995a),
	.w1(32'h3b48902d),
	.w2(32'h3aa3d74e),
	.w3(32'hbbf92c43),
	.w4(32'h3b23698e),
	.w5(32'h3ac7ff2f),
	.w6(32'h3b913ae7),
	.w7(32'h3b45708b),
	.w8(32'h3b5f14fc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dcaf0),
	.w1(32'hbb4308ef),
	.w2(32'hbb4b8931),
	.w3(32'h3ad8d18c),
	.w4(32'hbb3265b2),
	.w5(32'hbb3807b5),
	.w6(32'hbb70dd26),
	.w7(32'hbb481a00),
	.w8(32'hbb798ba1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40beb8),
	.w1(32'hba8ed780),
	.w2(32'hba4dbdb4),
	.w3(32'hbb845342),
	.w4(32'hb9c1a9a9),
	.w5(32'hba908dc7),
	.w6(32'hbad1287a),
	.w7(32'hbb1847a0),
	.w8(32'hb94012db),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0434e),
	.w1(32'hbaa6211b),
	.w2(32'hbac95568),
	.w3(32'hba02aa8f),
	.w4(32'hbac35df8),
	.w5(32'hbaed4a04),
	.w6(32'hbb1dd97e),
	.w7(32'hba52844c),
	.w8(32'h39044496),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a033),
	.w1(32'h3be051c0),
	.w2(32'hbacac61f),
	.w3(32'hbc0ae275),
	.w4(32'h3c5f4a84),
	.w5(32'h3b7ba6af),
	.w6(32'hbb9ca9d8),
	.w7(32'h3c15a3bd),
	.w8(32'h3b58d28e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04d80c),
	.w1(32'h3b83840c),
	.w2(32'hba7a42ea),
	.w3(32'hbade0625),
	.w4(32'h3b864968),
	.w5(32'hba86b4b3),
	.w6(32'hba3dd9eb),
	.w7(32'h3b4f7e72),
	.w8(32'hbaa9b880),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8fd3),
	.w1(32'h3b3ce7b0),
	.w2(32'h392044f5),
	.w3(32'h3a40916c),
	.w4(32'h3bb3089a),
	.w5(32'h3b071dda),
	.w6(32'h3ac7290c),
	.w7(32'h3bc8adb2),
	.w8(32'hbb01fc7d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba82af),
	.w1(32'hbbeda078),
	.w2(32'hbc2c33b5),
	.w3(32'hbc004ba9),
	.w4(32'hbc1ca322),
	.w5(32'hbc0f65f1),
	.w6(32'hbc8e6dc7),
	.w7(32'hbc7d2957),
	.w8(32'hbc84b924),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985c20f),
	.w1(32'h3c107efd),
	.w2(32'hbbe52efd),
	.w3(32'hb9ba8b40),
	.w4(32'h3c1e5934),
	.w5(32'hbb47d8c5),
	.w6(32'hbba5ba10),
	.w7(32'h3bd3baa1),
	.w8(32'hbb8dd4bb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf3b5),
	.w1(32'hbbe3129c),
	.w2(32'hbc39cf24),
	.w3(32'hbb3e4311),
	.w4(32'hb9d6e9ec),
	.w5(32'hbbc1a634),
	.w6(32'hba48a3d3),
	.w7(32'hbaab4f1f),
	.w8(32'hbc5c08e7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bcfbe),
	.w1(32'h3c003a45),
	.w2(32'hbaeffa63),
	.w3(32'hba8d5f07),
	.w4(32'h3c0f63a5),
	.w5(32'h398a0efc),
	.w6(32'hbab2ae69),
	.w7(32'h3c10e5c5),
	.w8(32'hb8f35ab4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b8cec),
	.w1(32'hbb73d41a),
	.w2(32'hbc369a0d),
	.w3(32'h3b127634),
	.w4(32'h3ba5daea),
	.w5(32'hbbb4f95c),
	.w6(32'h384fb594),
	.w7(32'h3b85a9ce),
	.w8(32'hbc386128),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e7154),
	.w1(32'hb848d8c4),
	.w2(32'hbb82f728),
	.w3(32'hbb476c6c),
	.w4(32'h3b5f845e),
	.w5(32'hba4c7cd6),
	.w6(32'h3ad179ea),
	.w7(32'h3a07108b),
	.w8(32'hbbbec2fd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d8ac),
	.w1(32'h3b3d9df3),
	.w2(32'hbbf288c7),
	.w3(32'hbbe30951),
	.w4(32'h3c1069f8),
	.w5(32'hbb81e69a),
	.w6(32'hbc4a98c3),
	.w7(32'h39d06e54),
	.w8(32'hbc16988d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6af9d7),
	.w1(32'h3b66b68a),
	.w2(32'h3b39c576),
	.w3(32'h3b80cad9),
	.w4(32'h3b98b0e4),
	.w5(32'h3b89eb97),
	.w6(32'h3b9e8363),
	.w7(32'h3b76a60d),
	.w8(32'h3b04051f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691418),
	.w1(32'h3ae2d84d),
	.w2(32'hbc7536af),
	.w3(32'h3a2fb56d),
	.w4(32'h3c130c74),
	.w5(32'hbc345bf9),
	.w6(32'h3b86479c),
	.w7(32'hbb0f9e5c),
	.w8(32'hbcc25161),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da5a9),
	.w1(32'hbb692fef),
	.w2(32'hbc75ddd3),
	.w3(32'hbb93e9d4),
	.w4(32'hbb4e3071),
	.w5(32'hbc12272a),
	.w6(32'hbc20fcd9),
	.w7(32'hbc1e3dbd),
	.w8(32'hbcc05647),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82bcce),
	.w1(32'h3befe275),
	.w2(32'hbc050ee9),
	.w3(32'hbc9f43da),
	.w4(32'h3acfa857),
	.w5(32'hbc22db50),
	.w6(32'hbb948d1b),
	.w7(32'hbb8f63e8),
	.w8(32'hbc7497a6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f64e2),
	.w1(32'h3ca5f5c3),
	.w2(32'hbba35f25),
	.w3(32'h3ba1bf12),
	.w4(32'h3d0cbfc4),
	.w5(32'h3c2b3a3a),
	.w6(32'hbbb675cf),
	.w7(32'h3d04404b),
	.w8(32'h3bcd958b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02dd9c),
	.w1(32'hbadb0ef5),
	.w2(32'hbc8e7fa0),
	.w3(32'hbb81b26a),
	.w4(32'hba356719),
	.w5(32'hbc890aa9),
	.w6(32'hbb9ec6ee),
	.w7(32'hbb4af886),
	.w8(32'hbcaf8c86),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3830ba),
	.w1(32'hbb981d45),
	.w2(32'hbc830104),
	.w3(32'h3ad92b08),
	.w4(32'h3ae6350e),
	.w5(32'hbc056d81),
	.w6(32'h3ad49351),
	.w7(32'h3b37fe13),
	.w8(32'hbc42a6a6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c179),
	.w1(32'h3a538c07),
	.w2(32'h3ace998b),
	.w3(32'h3aae092e),
	.w4(32'h3afc4810),
	.w5(32'h3a9aa4c7),
	.w6(32'h3aa9d217),
	.w7(32'h39a0fbab),
	.w8(32'hba66678b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96c4d9),
	.w1(32'hbb5cbb57),
	.w2(32'hbc65b1e6),
	.w3(32'hbc87bb1b),
	.w4(32'hbb5c6bba),
	.w5(32'hbc2ad00d),
	.w6(32'hbbe4eb9f),
	.w7(32'hbb443abd),
	.w8(32'hbc298684),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41e264),
	.w1(32'hbb42e00b),
	.w2(32'hbc2fcf55),
	.w3(32'hbc0a3226),
	.w4(32'hbc02d59e),
	.w5(32'hbc861d10),
	.w6(32'hba525b46),
	.w7(32'hbb74b4e5),
	.w8(32'hbc6fc09a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba584ddd),
	.w1(32'hba4ea5ed),
	.w2(32'hb9ebaf6e),
	.w3(32'hb97079d1),
	.w4(32'hbaa6661e),
	.w5(32'hbafb3ca1),
	.w6(32'hbb0e57fe),
	.w7(32'hbaca75df),
	.w8(32'hbb3f277e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3986fd),
	.w1(32'hbae2089f),
	.w2(32'hbb17c721),
	.w3(32'hbb62de44),
	.w4(32'hb9ea5b59),
	.w5(32'hba9b2c0a),
	.w6(32'hbb33b1db),
	.w7(32'hbad6d804),
	.w8(32'hbac48d95),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9016c2),
	.w1(32'hbc03f47d),
	.w2(32'hbc5d77b9),
	.w3(32'hbc049af8),
	.w4(32'hbc336ee7),
	.w5(32'hbc7996ee),
	.w6(32'hbbfb33f4),
	.w7(32'hbc836b99),
	.w8(32'hbcbfe5fb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05123),
	.w1(32'hbb023a03),
	.w2(32'hbc8d4f6d),
	.w3(32'h391694d4),
	.w4(32'h39bc2ca8),
	.w5(32'hbc7bf178),
	.w6(32'hbab70d8a),
	.w7(32'hbb3ddd3b),
	.w8(32'hbc975e37),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54b13a),
	.w1(32'hbbb04cd8),
	.w2(32'hbc4ba49d),
	.w3(32'hbc96a20e),
	.w4(32'hbb6b9487),
	.w5(32'hbc0346ba),
	.w6(32'hbc705ac8),
	.w7(32'hbc22b953),
	.w8(32'hbc5b0976),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85217c),
	.w1(32'h3b272bc6),
	.w2(32'hbbd85d6f),
	.w3(32'hbb0d6304),
	.w4(32'h3c204a8b),
	.w5(32'hbb04b562),
	.w6(32'h3ad0d42d),
	.w7(32'h3b7c6b7a),
	.w8(32'hbb8e477b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185d8c),
	.w1(32'h3b232f8d),
	.w2(32'hbbce4331),
	.w3(32'hb9824d0a),
	.w4(32'h3b853b4b),
	.w5(32'hbb86bc1a),
	.w6(32'hbbd06563),
	.w7(32'h39a302b4),
	.w8(32'hbbd07e20),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cad87),
	.w1(32'hbbd88c3a),
	.w2(32'hbc18c9b0),
	.w3(32'hbbcefc06),
	.w4(32'hba51726b),
	.w5(32'hbb7350ed),
	.w6(32'hbae66ef2),
	.w7(32'h3a5e56ce),
	.w8(32'hbbb030e2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a20ab),
	.w1(32'h3a0b51fc),
	.w2(32'hbbc07257),
	.w3(32'hbbabf54f),
	.w4(32'h3b3df305),
	.w5(32'hbba1afc9),
	.w6(32'hba2021b5),
	.w7(32'h3a4e64dc),
	.w8(32'hbbda8ff9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a697436),
	.w1(32'hbb2e250a),
	.w2(32'hbb863cf4),
	.w3(32'h3a3fc692),
	.w4(32'hbaf04272),
	.w5(32'hbb6b8047),
	.w6(32'hbb008b97),
	.w7(32'hbb5857c6),
	.w8(32'hbaf94397),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d6df),
	.w1(32'hbadd1a38),
	.w2(32'hbb0ce3a0),
	.w3(32'hbb0a0ab9),
	.w4(32'hbace86aa),
	.w5(32'hbaf71408),
	.w6(32'hbae9d6ae),
	.w7(32'hbadf118e),
	.w8(32'hbacfd087),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae73ed0),
	.w1(32'hbac3ddb8),
	.w2(32'hbb163449),
	.w3(32'hbad6745a),
	.w4(32'hbb03a8c3),
	.w5(32'hbb19eb47),
	.w6(32'hbad38fa2),
	.w7(32'hbb1a0a48),
	.w8(32'hbb03ca46),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ce96),
	.w1(32'h3afe8647),
	.w2(32'hbaa42683),
	.w3(32'hbabcff3b),
	.w4(32'h3b7d0b1e),
	.w5(32'h39bc50d9),
	.w6(32'h3b0e4cb2),
	.w7(32'hb9e9232d),
	.w8(32'h3a894b7b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba899ed),
	.w1(32'h3b3310ca),
	.w2(32'hbb481518),
	.w3(32'h3b605ac2),
	.w4(32'h3bd1649a),
	.w5(32'hba66e43b),
	.w6(32'h3b7582ff),
	.w7(32'h3c4989a6),
	.w8(32'hbb1a31b1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2da5),
	.w1(32'hbbe4ae45),
	.w2(32'hbbe4e88d),
	.w3(32'hba1a7b25),
	.w4(32'hbbcfbeea),
	.w5(32'hbbcdc0f0),
	.w6(32'hbbda3bec),
	.w7(32'hbbc69d2a),
	.w8(32'hbbbc9fa7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34136a),
	.w1(32'hbc2ea16c),
	.w2(32'hbc33a7e5),
	.w3(32'hbc37d95d),
	.w4(32'hbc511eb0),
	.w5(32'hbc3d421c),
	.w6(32'hbbfb118a),
	.w7(32'hbc35dd65),
	.w8(32'hbc71aa18),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40e71f),
	.w1(32'h3a90bbed),
	.w2(32'hbbf0b9f3),
	.w3(32'hbc33a2b7),
	.w4(32'h3b4ceb9c),
	.w5(32'hbbdd8763),
	.w6(32'hbc310d70),
	.w7(32'hbb13a2e5),
	.w8(32'hbc430962),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05ba1f),
	.w1(32'h3b2c5011),
	.w2(32'hbb2f03e9),
	.w3(32'hbaff3163),
	.w4(32'h3bcff27d),
	.w5(32'hb96984d0),
	.w6(32'h3ac6a35d),
	.w7(32'h3a0eed4a),
	.w8(32'h3ad255d2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b908d),
	.w1(32'h3b595ca1),
	.w2(32'h3aa25704),
	.w3(32'h3b61c32f),
	.w4(32'h3b287727),
	.w5(32'h3b0d4fcd),
	.w6(32'h3b0442fd),
	.w7(32'h3b0cfc05),
	.w8(32'h3a00d2c6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accc8fc),
	.w1(32'h3a30f1d9),
	.w2(32'hb9c1e9de),
	.w3(32'h3af78a7b),
	.w4(32'h3a4df9f2),
	.w5(32'hb9d9a52d),
	.w6(32'h3a814ed9),
	.w7(32'hb96c4977),
	.w8(32'hb97a34e0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f452),
	.w1(32'h3aefa5ae),
	.w2(32'h3ba3b3e6),
	.w3(32'hbb0b6436),
	.w4(32'hbb6c325a),
	.w5(32'hbc0471a1),
	.w6(32'h381fa38f),
	.w7(32'h3ae633f7),
	.w8(32'h3add852a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad54529),
	.w1(32'hbbe8bf0f),
	.w2(32'hbb61cd92),
	.w3(32'hb8b99ead),
	.w4(32'hbb082881),
	.w5(32'hbb416672),
	.w6(32'h3afd78c0),
	.w7(32'hbc1c5daa),
	.w8(32'hbc5fdf28),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5abc6b),
	.w1(32'hbc244099),
	.w2(32'hbd31151e),
	.w3(32'h3b2af313),
	.w4(32'h3b6830cc),
	.w5(32'h3bc50b82),
	.w6(32'hbb9280b6),
	.w7(32'hbbe78cc9),
	.w8(32'hbc3b3ab6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95042),
	.w1(32'h3b6f1118),
	.w2(32'h3b20ba3f),
	.w3(32'hbb028a72),
	.w4(32'h3b9bca9f),
	.w5(32'h3c001172),
	.w6(32'h3b5ba0d8),
	.w7(32'hbb734b09),
	.w8(32'hba1a8ac3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e6675),
	.w1(32'h3aa15741),
	.w2(32'hbae812b9),
	.w3(32'h3b1f2ee0),
	.w4(32'hba3cb3d0),
	.w5(32'hbb93be25),
	.w6(32'hbbaea107),
	.w7(32'h3a1c7dc1),
	.w8(32'hba6550e3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b830),
	.w1(32'hbccc5839),
	.w2(32'hbc316092),
	.w3(32'hbb159805),
	.w4(32'h3c97d528),
	.w5(32'h3c6c7a55),
	.w6(32'hbc0ed1bd),
	.w7(32'hbb3a04f8),
	.w8(32'hbba17824),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8bdb3),
	.w1(32'h3b88c0a3),
	.w2(32'hb9cb8fcb),
	.w3(32'h3c0d86fc),
	.w4(32'h3af3dd5e),
	.w5(32'h3a510661),
	.w6(32'h3b03fb47),
	.w7(32'hbc83d733),
	.w8(32'hbc96da84),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21b22c),
	.w1(32'hbae90fe4),
	.w2(32'hbb0f22de),
	.w3(32'h3b328250),
	.w4(32'h3c10a179),
	.w5(32'h3c81fac7),
	.w6(32'hbc1a6177),
	.w7(32'hbc790464),
	.w8(32'hbc7cbdb4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb864),
	.w1(32'hb9eba04c),
	.w2(32'hbc4c1ce5),
	.w3(32'hb9ae65bf),
	.w4(32'hbad881f1),
	.w5(32'hbb9ade76),
	.w6(32'hb942fad4),
	.w7(32'hbbfc5676),
	.w8(32'hbc823584),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06a81a),
	.w1(32'h3b60056b),
	.w2(32'hb8e37089),
	.w3(32'h3c1bf9c9),
	.w4(32'h3bb79f5c),
	.w5(32'hbbf91930),
	.w6(32'h3b87f106),
	.w7(32'h3c3125ad),
	.w8(32'hbbb65f34),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756e0e),
	.w1(32'h3b2eb45e),
	.w2(32'h3afae82f),
	.w3(32'hbb43b79a),
	.w4(32'h3be9ba5f),
	.w5(32'h3b11151a),
	.w6(32'hb812cbfc),
	.w7(32'h3a877aed),
	.w8(32'hbbeecc9a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac022e2),
	.w1(32'hbc04b97d),
	.w2(32'hbc60cdc8),
	.w3(32'hbaaff7a6),
	.w4(32'h3b29ccd5),
	.w5(32'h3af98251),
	.w6(32'h3ab0e530),
	.w7(32'hbb261a9d),
	.w8(32'hbc353cd7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc796bc5),
	.w1(32'h3999350d),
	.w2(32'hbb93a66b),
	.w3(32'hbb6eeb85),
	.w4(32'h3b3c12cf),
	.w5(32'hbc30fb5f),
	.w6(32'hbc010e0d),
	.w7(32'hbbe36822),
	.w8(32'hbbc7694f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b7d1),
	.w1(32'hbc01631a),
	.w2(32'hbba73fbe),
	.w3(32'hbb15a695),
	.w4(32'h3c2d1679),
	.w5(32'h3b12ef88),
	.w6(32'h3c0b7700),
	.w7(32'h3c54d7e6),
	.w8(32'hbb108881),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bed4f),
	.w1(32'h3ad0c027),
	.w2(32'hb9ba67e6),
	.w3(32'h3acbec13),
	.w4(32'hbb87f4ff),
	.w5(32'hbbe77bd0),
	.w6(32'hbaaae44d),
	.w7(32'h3a9554e2),
	.w8(32'hbb08c5d7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c13b),
	.w1(32'h3c3f4f2d),
	.w2(32'h3bb06791),
	.w3(32'hbc201fe0),
	.w4(32'hbb5a5fe2),
	.w5(32'hbd0fcaf4),
	.w6(32'h3c5c34b2),
	.w7(32'h3d314795),
	.w8(32'h3c005358),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a33e),
	.w1(32'hbc60b9e9),
	.w2(32'h3be0d079),
	.w3(32'hbc88f91e),
	.w4(32'h3bdf0ae4),
	.w5(32'hbc0c384f),
	.w6(32'hbca67a20),
	.w7(32'hbcd46691),
	.w8(32'hbb9ea92f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd044323),
	.w1(32'h38d0037a),
	.w2(32'h3c023ea2),
	.w3(32'hbc006ae9),
	.w4(32'h3a0de53c),
	.w5(32'h3bb5bb52),
	.w6(32'hbafe704b),
	.w7(32'hbb839433),
	.w8(32'hbb44ea64),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a958134),
	.w1(32'h3c10c6c9),
	.w2(32'h3b9918f9),
	.w3(32'h3a63639f),
	.w4(32'hb9376bb9),
	.w5(32'hbbc104b1),
	.w6(32'h3a272f21),
	.w7(32'hbaa2c1c8),
	.w8(32'hba078dd2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a50a1),
	.w1(32'h397869e6),
	.w2(32'hbbc5a5c0),
	.w3(32'hbbad1210),
	.w4(32'h3b19c59e),
	.w5(32'h3b841d25),
	.w6(32'h38c2d55d),
	.w7(32'hbb66e28f),
	.w8(32'hbb15ca6e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55f923),
	.w1(32'h3ba44afb),
	.w2(32'hbb9c76cb),
	.w3(32'hba65fff6),
	.w4(32'h3bf146cb),
	.w5(32'hb920224c),
	.w6(32'hbb9464b9),
	.w7(32'h3b804e56),
	.w8(32'hbb912f32),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46a3b9),
	.w1(32'h3b4a0be7),
	.w2(32'h39bb36be),
	.w3(32'hbcd6fbc1),
	.w4(32'hbc01eccb),
	.w5(32'hbb5d7df1),
	.w6(32'hbc63b562),
	.w7(32'hbc4b382b),
	.w8(32'hbc83aaa7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b6cc0),
	.w1(32'hbb5a01f6),
	.w2(32'h3b17c944),
	.w3(32'h3b3cad5e),
	.w4(32'hbbac061f),
	.w5(32'hbbf4bb98),
	.w6(32'h3b5bc686),
	.w7(32'h3b8c49df),
	.w8(32'h3bac59ab),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25cc6),
	.w1(32'h3b9ae9be),
	.w2(32'hbc5f6e49),
	.w3(32'hbbf54860),
	.w4(32'hbc8a24ea),
	.w5(32'hbcb113f6),
	.w6(32'hbcbff155),
	.w7(32'hbc39c608),
	.w8(32'hbcd2becc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb753bc),
	.w1(32'hbb6adadb),
	.w2(32'hbc40f8b6),
	.w3(32'hbad84f24),
	.w4(32'hbb3dc9e4),
	.w5(32'hbc05347d),
	.w6(32'h3ae5300a),
	.w7(32'hbbcd011c),
	.w8(32'hbc013783),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b4d2),
	.w1(32'hbbde3d68),
	.w2(32'hbc06a355),
	.w3(32'hbc6c9cc1),
	.w4(32'hbbee89b4),
	.w5(32'hbc57e300),
	.w6(32'hb9e21d92),
	.w7(32'hbbc00ff5),
	.w8(32'hbc504cc8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d63634),
	.w1(32'h3ac4ced0),
	.w2(32'hbbebe8f5),
	.w3(32'hbba23a9f),
	.w4(32'h3c2b45a2),
	.w5(32'hbb113aa2),
	.w6(32'hbc0abfd7),
	.w7(32'hba818c04),
	.w8(32'hbc4bfd0c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059e1c),
	.w1(32'hbbf3f6c0),
	.w2(32'hbcabe73a),
	.w3(32'hbbc0840f),
	.w4(32'h3a803b28),
	.w5(32'hbc211ec1),
	.w6(32'hbb5a5eb7),
	.w7(32'h39219a8e),
	.w8(32'hbb30ddf3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108afc),
	.w1(32'h3c0cf8b7),
	.w2(32'h3be5117a),
	.w3(32'hbc25049c),
	.w4(32'h3bbcd54a),
	.w5(32'h3b34f49e),
	.w6(32'h3c237b92),
	.w7(32'h3bf3995c),
	.w8(32'h3b753705),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc780d0),
	.w1(32'h3a546fc9),
	.w2(32'hbc1030b9),
	.w3(32'hb8595bbe),
	.w4(32'h3c8a5ee3),
	.w5(32'h3b92f851),
	.w6(32'h3b9e5bee),
	.w7(32'h3a4551f4),
	.w8(32'hbc6ef558),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b332),
	.w1(32'h3c10c1fb),
	.w2(32'h3b5088e6),
	.w3(32'hbbbbe967),
	.w4(32'h3bbcd04a),
	.w5(32'hbb651e5d),
	.w6(32'hbbe01e30),
	.w7(32'h3bed52fd),
	.w8(32'hb9152c66),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b647760),
	.w1(32'h3c149836),
	.w2(32'h3aa29eab),
	.w3(32'hbb4b7ced),
	.w4(32'h3bfedc41),
	.w5(32'hbae5b996),
	.w6(32'hbb6bfab2),
	.w7(32'h3b09ec6d),
	.w8(32'hbb459091),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ac540),
	.w1(32'hbb6f7694),
	.w2(32'hbb16cc35),
	.w3(32'hbb403bfc),
	.w4(32'hbbde3775),
	.w5(32'hbbeb4a09),
	.w6(32'hb9f3a9e2),
	.w7(32'hba9dc2b4),
	.w8(32'h3a1c0202),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b4931),
	.w1(32'hbaff2ddc),
	.w2(32'hb9518016),
	.w3(32'hbb6472d8),
	.w4(32'hbb778383),
	.w5(32'hbad50604),
	.w6(32'hbb3a3223),
	.w7(32'hbb6444e7),
	.w8(32'hba2daea2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c69a),
	.w1(32'h3b984903),
	.w2(32'hbba78bff),
	.w3(32'hbb814631),
	.w4(32'hbb9a083f),
	.w5(32'hbc693d74),
	.w6(32'h3c4694a1),
	.w7(32'h3c2e00f1),
	.w8(32'h39dcfaef),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38c51b),
	.w1(32'h3b857887),
	.w2(32'hbc012293),
	.w3(32'hbae2778d),
	.w4(32'h3aa049bf),
	.w5(32'hbc2436b0),
	.w6(32'h3ae4edb6),
	.w7(32'h3854fcbb),
	.w8(32'hbb61f6ea),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ca630),
	.w1(32'hbb8814df),
	.w2(32'hbc49a820),
	.w3(32'h3b2f8fd8),
	.w4(32'h3c3da193),
	.w5(32'h3b946d95),
	.w6(32'hbb888840),
	.w7(32'hbc2803e1),
	.w8(32'hbc3eca8e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8071c4),
	.w1(32'h3ace8b4e),
	.w2(32'h3a8411fd),
	.w3(32'hbc0163e2),
	.w4(32'hba231905),
	.w5(32'hbb420018),
	.w6(32'h3b88010e),
	.w7(32'h3b95892b),
	.w8(32'h3bafb2bf),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93df75),
	.w1(32'hbba5968b),
	.w2(32'hbc95365f),
	.w3(32'hbad00ab3),
	.w4(32'hbb4d5495),
	.w5(32'hbc5c7735),
	.w6(32'hbba0c7aa),
	.w7(32'hbcbe7b07),
	.w8(32'hbccf2691),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1396e6),
	.w1(32'h3b0b5895),
	.w2(32'hbb0f8b33),
	.w3(32'h3a614d89),
	.w4(32'h39c9c7ba),
	.w5(32'h3b414951),
	.w6(32'h3b3d0556),
	.w7(32'h3a74155b),
	.w8(32'h3a6aa371),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c0a38),
	.w1(32'h3af88663),
	.w2(32'h3ba7ae40),
	.w3(32'h3bee8486),
	.w4(32'h3b219259),
	.w5(32'h3b00dd86),
	.w6(32'h3a328354),
	.w7(32'hbb26ec39),
	.w8(32'hbb966367),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d21c),
	.w1(32'h3b4a3149),
	.w2(32'hbb7aaaca),
	.w3(32'h3b292dab),
	.w4(32'h3c0f7f4a),
	.w5(32'h3aeebc2f),
	.w6(32'h3be2e7f8),
	.w7(32'h3b8537f3),
	.w8(32'hbb12e38a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8a04),
	.w1(32'hbc01ed29),
	.w2(32'hbc9a69c8),
	.w3(32'hba9d4085),
	.w4(32'hbb817103),
	.w5(32'hbcb5d0d8),
	.w6(32'h3a181a34),
	.w7(32'h3ae83847),
	.w8(32'hbc822b89),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076b64),
	.w1(32'h37fe1454),
	.w2(32'hbc54a980),
	.w3(32'h3b9918d5),
	.w4(32'h3b8ba83e),
	.w5(32'hbc3a9288),
	.w6(32'h3b30896e),
	.w7(32'h3acea43a),
	.w8(32'hbb55cb27),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b4cd7),
	.w1(32'h3be3d1b3),
	.w2(32'hbbc65484),
	.w3(32'hbb6e7268),
	.w4(32'h3a39a701),
	.w5(32'hbc335127),
	.w6(32'h3b4f58f9),
	.w7(32'h3bff22e1),
	.w8(32'hbba8bee5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dbf02),
	.w1(32'hba896e5c),
	.w2(32'hbc3f813f),
	.w3(32'hbb953bb4),
	.w4(32'h3c3b47fe),
	.w5(32'h3c4b3035),
	.w6(32'hba896a7f),
	.w7(32'h3b6396d0),
	.w8(32'hb9f6830a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2da6b),
	.w1(32'hbb56452a),
	.w2(32'hbcfe4bf9),
	.w3(32'h3aa2bcf5),
	.w4(32'hbc39f9b1),
	.w5(32'hbcf4512b),
	.w6(32'hbb0b50ce),
	.w7(32'h3d1135a9),
	.w8(32'h3bd34f46),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c99a2),
	.w1(32'h39214450),
	.w2(32'hbcdb44e6),
	.w3(32'hbc24fc8b),
	.w4(32'hbc0e5816),
	.w5(32'hbcd012f7),
	.w6(32'h3ba77112),
	.w7(32'h3ce06c1d),
	.w8(32'h3ad3b86b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6da798),
	.w1(32'hbc8ad8bf),
	.w2(32'h3c82dd2d),
	.w3(32'hbc227774),
	.w4(32'hb9d23a40),
	.w5(32'hbb81719c),
	.w6(32'hbc2fe30d),
	.w7(32'hbc866356),
	.w8(32'hbca8eef3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7097d7),
	.w1(32'h3c091e37),
	.w2(32'h3bb755cc),
	.w3(32'h3b6cb062),
	.w4(32'h3b387a7b),
	.w5(32'h3b0016fc),
	.w6(32'h3b190e5c),
	.w7(32'h3ad47021),
	.w8(32'h3b8929f8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a257d),
	.w1(32'hb9aedd12),
	.w2(32'hbb009148),
	.w3(32'hbbc298ae),
	.w4(32'h3b21322d),
	.w5(32'h39cf72bd),
	.w6(32'h3b381d7f),
	.w7(32'h3b16d2fd),
	.w8(32'hbaf33dbe),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7d201),
	.w1(32'h3b32f5b9),
	.w2(32'h3bdd1ac2),
	.w3(32'h3a469cf4),
	.w4(32'hbb6339ef),
	.w5(32'hbc03f448),
	.w6(32'h3c13cd2c),
	.w7(32'h3c5ad9ad),
	.w8(32'h3bb0d856),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f74f1d),
	.w1(32'hbb435efc),
	.w2(32'h3a545b90),
	.w3(32'hbbb82600),
	.w4(32'hbc86a5de),
	.w5(32'hbcdd1a8d),
	.w6(32'h3c6758a9),
	.w7(32'h3cfe3a15),
	.w8(32'h3c487018),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d0bb),
	.w1(32'h3b5a9ee5),
	.w2(32'h3c31e409),
	.w3(32'hbb308334),
	.w4(32'h3c6ff825),
	.w5(32'h3c40eb42),
	.w6(32'hbb926562),
	.w7(32'hbc3676d2),
	.w8(32'hbbacbfa7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc762b9),
	.w1(32'hbbe78ea5),
	.w2(32'h3b0f255e),
	.w3(32'hbc2bb222),
	.w4(32'hbbbdd982),
	.w5(32'h3bf474f3),
	.w6(32'hbc76c22f),
	.w7(32'hbc522c7b),
	.w8(32'hbc0eb87f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5c74),
	.w1(32'hba3d6c1d),
	.w2(32'hbbfbf627),
	.w3(32'h3bec27be),
	.w4(32'h3ba82125),
	.w5(32'h3b98f9c9),
	.w6(32'hbb9bea74),
	.w7(32'hbc9431c1),
	.w8(32'hbc2b2493),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944a3b),
	.w1(32'hb8e277d5),
	.w2(32'hba263cf5),
	.w3(32'hba0a64d8),
	.w4(32'h3bcf45fc),
	.w5(32'h3c0155ef),
	.w6(32'hbb2c8ddc),
	.w7(32'hbbfa2d33),
	.w8(32'hbb8990b8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834d6f),
	.w1(32'hbbc473d0),
	.w2(32'hbb6117c7),
	.w3(32'h3af1eff7),
	.w4(32'hbb5b35cd),
	.w5(32'hbb376aac),
	.w6(32'hb91b0a52),
	.w7(32'hbb36776b),
	.w8(32'h3b59ac6d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafaa79),
	.w1(32'hbb6e7863),
	.w2(32'hbc963165),
	.w3(32'h3b66603b),
	.w4(32'hbc17a071),
	.w5(32'hbd0267bf),
	.w6(32'h3c38f799),
	.w7(32'h3cf6e05e),
	.w8(32'h3be6aea3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6779db),
	.w1(32'h3bb6c26a),
	.w2(32'h39bc7861),
	.w3(32'hbc2a5edb),
	.w4(32'hbc50f676),
	.w5(32'hbc9db782),
	.w6(32'h3c06886b),
	.w7(32'h3c9ae834),
	.w8(32'hba7eb77f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb781d21),
	.w1(32'h3adcd176),
	.w2(32'hb9afa8e6),
	.w3(32'hbbf667a9),
	.w4(32'h3b21700e),
	.w5(32'h3b9ad13a),
	.w6(32'h3b13a5ba),
	.w7(32'h39322dbd),
	.w8(32'h3a956948),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d09d5),
	.w1(32'h38a6ea77),
	.w2(32'hbc16090d),
	.w3(32'h3c195eae),
	.w4(32'h3c3d759f),
	.w5(32'hbaff1912),
	.w6(32'h3c7c17fc),
	.w7(32'h3ca6c615),
	.w8(32'hbc28cecd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8731e4),
	.w1(32'h3b6641c6),
	.w2(32'hbc5f4854),
	.w3(32'hbc4957c6),
	.w4(32'h3c39eb33),
	.w5(32'hbaddebda),
	.w6(32'hbc5a8515),
	.w7(32'h3b503520),
	.w8(32'hbb7b1faa),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acabfe),
	.w1(32'hbb9ca908),
	.w2(32'hbc85275e),
	.w3(32'hbb60eb06),
	.w4(32'hbc14a551),
	.w5(32'hbc749539),
	.w6(32'h3b26ccb2),
	.w7(32'h3c051949),
	.w8(32'hb9e64c29),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a90d86),
	.w1(32'h3c0e43eb),
	.w2(32'h3bd15a22),
	.w3(32'hbbf42630),
	.w4(32'hbbab6c4b),
	.w5(32'hbb4d7bb8),
	.w6(32'h3c23f4ea),
	.w7(32'h3c720687),
	.w8(32'hbb65fc1a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f7810),
	.w1(32'hbadaf02d),
	.w2(32'hbbf16efb),
	.w3(32'h3b2ca8f7),
	.w4(32'h3c087d86),
	.w5(32'h3c1d73b2),
	.w6(32'hba941214),
	.w7(32'hbade52ac),
	.w8(32'hbb5ff17a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914047),
	.w1(32'h3bc56f7a),
	.w2(32'h3b1bf779),
	.w3(32'h3bf5a5e8),
	.w4(32'h3afbd119),
	.w5(32'h3bcdde5d),
	.w6(32'h3bc9fd3f),
	.w7(32'h3b32ca04),
	.w8(32'h3b150512),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa04c4e),
	.w1(32'h3b38328a),
	.w2(32'hba265141),
	.w3(32'h3aa50bad),
	.w4(32'hbb675b22),
	.w5(32'hbc85b78d),
	.w6(32'h3c219300),
	.w7(32'h3cab551e),
	.w8(32'h3ac826e0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab807b0),
	.w1(32'hbc0cfd56),
	.w2(32'hbc056709),
	.w3(32'h3b056c75),
	.w4(32'hbbb12ec1),
	.w5(32'hbbefc9b7),
	.w6(32'hbc4959b5),
	.w7(32'hbc1eee11),
	.w8(32'hbc1bd058),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f65da),
	.w1(32'hbb903deb),
	.w2(32'hbc4315e0),
	.w3(32'hbc57e45a),
	.w4(32'hbb627eda),
	.w5(32'hbbe78934),
	.w6(32'hbc5619b7),
	.w7(32'hbbe8fa0b),
	.w8(32'hbbaf884a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fea17),
	.w1(32'hbb33b684),
	.w2(32'h3baf8dea),
	.w3(32'hbb8ec289),
	.w4(32'hbb8a6cc2),
	.w5(32'hb9af97c1),
	.w6(32'h3b104a9b),
	.w7(32'h3b57062a),
	.w8(32'hba64c50a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ad9b),
	.w1(32'hbad10d29),
	.w2(32'hbc760df0),
	.w3(32'hbc240eb3),
	.w4(32'hbca8241e),
	.w5(32'hbd47b338),
	.w6(32'h3c0f042e),
	.w7(32'h3cf651b8),
	.w8(32'hbbeb7011),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52a14),
	.w1(32'hbac2d51d),
	.w2(32'hbbcb11e7),
	.w3(32'hbc98f387),
	.w4(32'h39e454b1),
	.w5(32'hba93410f),
	.w6(32'hbb51040a),
	.w7(32'hbc08c3a8),
	.w8(32'hbbab40c1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841a7be),
	.w1(32'h3addc867),
	.w2(32'h3bacbd57),
	.w3(32'h3aebd0d7),
	.w4(32'h39d35a01),
	.w5(32'hbb6fdd86),
	.w6(32'h3b62f64a),
	.w7(32'h3b2fa4eb),
	.w8(32'h3b027670),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5698d4),
	.w1(32'hbab3ccc9),
	.w2(32'h3b70d283),
	.w3(32'hbb292824),
	.w4(32'h3a545d56),
	.w5(32'h3adc4a9d),
	.w6(32'hbaeabece),
	.w7(32'hbb627e0c),
	.w8(32'hbb47e404),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981cf54),
	.w1(32'h37d38237),
	.w2(32'h3a38a60a),
	.w3(32'hb993e77f),
	.w4(32'hbb24348c),
	.w5(32'hbaed8aa0),
	.w6(32'h3b4a93d9),
	.w7(32'h3a920973),
	.w8(32'h3bbcbe7e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3526),
	.w1(32'h3981296e),
	.w2(32'hbc0640a8),
	.w3(32'hbba4e30b),
	.w4(32'h3ba3a55f),
	.w5(32'hbbb80c9b),
	.w6(32'hbb304c89),
	.w7(32'hbbcb554f),
	.w8(32'hbc406428),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37144f),
	.w1(32'hbcbd13c3),
	.w2(32'hbca43cee),
	.w3(32'hbbbddf52),
	.w4(32'h3b5a863e),
	.w5(32'hbce7509b),
	.w6(32'hbb0a7653),
	.w7(32'h3c2f1883),
	.w8(32'hbbc7012f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd43bff),
	.w1(32'h3b0d81cc),
	.w2(32'hbc000f50),
	.w3(32'hbb3d1bc7),
	.w4(32'h3bb00aa3),
	.w5(32'hbc49499f),
	.w6(32'h3bcb2366),
	.w7(32'h3c8737d2),
	.w8(32'hbbf7019d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95247d),
	.w1(32'h3af62409),
	.w2(32'hbba7264b),
	.w3(32'hbb004d36),
	.w4(32'h3b847d72),
	.w5(32'hbb95d077),
	.w6(32'hbb72b291),
	.w7(32'h3b3799c0),
	.w8(32'h3b4fb479),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00b45),
	.w1(32'h3c06a7f5),
	.w2(32'hbba1b11c),
	.w3(32'hbbc8e136),
	.w4(32'h3c927feb),
	.w5(32'h3b7e75d0),
	.w6(32'hbb9db9e5),
	.w7(32'hbbb42802),
	.w8(32'hbc4c5909),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc856b),
	.w1(32'hbb9bf54d),
	.w2(32'hbb390b53),
	.w3(32'hba716d51),
	.w4(32'hbbd21973),
	.w5(32'hbc43411c),
	.w6(32'hbaa031d4),
	.w7(32'h3946011c),
	.w8(32'hbb810b6a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca530df),
	.w1(32'hbb9e2743),
	.w2(32'hbc393e66),
	.w3(32'hbce0a164),
	.w4(32'hbc911e62),
	.w5(32'hbc8bd47a),
	.w6(32'hbcce4b45),
	.w7(32'hbc80b3dd),
	.w8(32'hbc474673),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34059e),
	.w1(32'h3b6b59e2),
	.w2(32'h3af4e1c4),
	.w3(32'hba834555),
	.w4(32'hbae3294a),
	.w5(32'hba8e6bee),
	.w6(32'h3b9a510d),
	.w7(32'h3b3de5bf),
	.w8(32'h3b6109c1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1509),
	.w1(32'hbb510a02),
	.w2(32'h3ab629f9),
	.w3(32'h3a3ecb5f),
	.w4(32'hbb45be0d),
	.w5(32'hbb1fca46),
	.w6(32'hbad60e24),
	.w7(32'hbb031827),
	.w8(32'h3bb1cb15),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083ffe),
	.w1(32'h3b5d7516),
	.w2(32'hbc7f4783),
	.w3(32'hbb807da4),
	.w4(32'h3bcabd26),
	.w5(32'hbbe64a52),
	.w6(32'hbb352cee),
	.w7(32'h39545105),
	.w8(32'hbc300c29),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb651918),
	.w1(32'h3c13eed6),
	.w2(32'hbc215c87),
	.w3(32'h3b953d60),
	.w4(32'h3b528fba),
	.w5(32'hbcc80ae6),
	.w6(32'h3be0c073),
	.w7(32'h3978e90c),
	.w8(32'hbc98b936),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba355dc0),
	.w1(32'hbbea7f59),
	.w2(32'hbc800732),
	.w3(32'hbbb2850c),
	.w4(32'hbb010b85),
	.w5(32'hbc5e49af),
	.w6(32'hbbf25db2),
	.w7(32'h3b6e5e45),
	.w8(32'hbc111943),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4272b),
	.w1(32'hbc770702),
	.w2(32'hbbc45222),
	.w3(32'hbaf01b73),
	.w4(32'hbc9cc95d),
	.w5(32'hbccd44b9),
	.w6(32'h3c0aec55),
	.w7(32'h3c63f508),
	.w8(32'h3b78d59b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bfb90),
	.w1(32'hbb7449a4),
	.w2(32'hb9d1b499),
	.w3(32'hbbf06da7),
	.w4(32'hbb974da7),
	.w5(32'hbb8e520b),
	.w6(32'h3a5cb8c2),
	.w7(32'h3a4d97ee),
	.w8(32'h3b49cf3e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae21983),
	.w1(32'hbadd697a),
	.w2(32'hbaa669e2),
	.w3(32'hbb511612),
	.w4(32'h3b31815a),
	.w5(32'h3bc65383),
	.w6(32'hbb969977),
	.w7(32'hbc1ddd8d),
	.w8(32'hbba22792),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5646),
	.w1(32'hbbc0043a),
	.w2(32'hbc310de8),
	.w3(32'hbb6dbab6),
	.w4(32'hbc8b1bc4),
	.w5(32'hbcb96c4f),
	.w6(32'hba90bf49),
	.w7(32'hbb977182),
	.w8(32'hbc4b69a3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e9dc4),
	.w1(32'hbc4798e8),
	.w2(32'hbc6a78b1),
	.w3(32'hbca20aae),
	.w4(32'hbc82ffe1),
	.w5(32'hbc837b68),
	.w6(32'hbc0f694a),
	.w7(32'hbc135da7),
	.w8(32'hbc649699),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad806),
	.w1(32'hbbc309bd),
	.w2(32'hbc2d4b6d),
	.w3(32'hbc6b7ac4),
	.w4(32'hbc6b4c02),
	.w5(32'hbc5ea23c),
	.w6(32'hbaeacab2),
	.w7(32'hbb370dbd),
	.w8(32'hbbdcc07d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bde9b),
	.w1(32'h3c0a6ce1),
	.w2(32'hbb1b88b9),
	.w3(32'h3a8df5ad),
	.w4(32'h3c520491),
	.w5(32'h3c55a620),
	.w6(32'hbc84b9b7),
	.w7(32'hbc59582d),
	.w8(32'hbc3c0711),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1b27),
	.w1(32'hbb15c21a),
	.w2(32'hbc516d06),
	.w3(32'hbb45645b),
	.w4(32'h3b846c85),
	.w5(32'hbbe4366e),
	.w6(32'hbb70a0b6),
	.w7(32'h3b81a446),
	.w8(32'hbb1eb5a6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8512),
	.w1(32'hba74437c),
	.w2(32'hbb0e957f),
	.w3(32'hbb3636ac),
	.w4(32'hba87bf88),
	.w5(32'hbb2cc472),
	.w6(32'hbb998f44),
	.w7(32'hbb9ae043),
	.w8(32'hbaf4bd0e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29b31d),
	.w1(32'h3c1598fd),
	.w2(32'hbbb07849),
	.w3(32'hbb43a798),
	.w4(32'hba8c07bb),
	.w5(32'h3c8d95d5),
	.w6(32'hbbe52e62),
	.w7(32'hbb7f9744),
	.w8(32'hbc23fb86),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fbc38),
	.w1(32'hba2e93e8),
	.w2(32'hbb0d2c5d),
	.w3(32'h3b2d9f3c),
	.w4(32'h3b85e090),
	.w5(32'h3b1649c2),
	.w6(32'h3b9bd15b),
	.w7(32'hbafca945),
	.w8(32'h3b4ec6fd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a156a15),
	.w1(32'h3ac0eac1),
	.w2(32'hba977795),
	.w3(32'h3b67755e),
	.w4(32'h3c4071a9),
	.w5(32'h3c95ace4),
	.w6(32'hbb87e76b),
	.w7(32'hbc4dccfd),
	.w8(32'hbc157d6a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9daba8),
	.w1(32'h3aaf0695),
	.w2(32'hbb4f5e9f),
	.w3(32'h3b3268e3),
	.w4(32'hbae36a75),
	.w5(32'hbb01e962),
	.w6(32'h3b95b42c),
	.w7(32'hbb441292),
	.w8(32'hbb954d4e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99d3cc),
	.w1(32'hbc31533f),
	.w2(32'hbc447f7b),
	.w3(32'h3b225652),
	.w4(32'h3c1eb2b0),
	.w5(32'h3bf08051),
	.w6(32'hbc269ae9),
	.w7(32'hbc890e91),
	.w8(32'hbca7ce71),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38dfd1),
	.w1(32'h3bac32cf),
	.w2(32'hbc8cbc90),
	.w3(32'h3a0065ff),
	.w4(32'h3990b3d5),
	.w5(32'hbcfd5d72),
	.w6(32'h3bbc7d82),
	.w7(32'h3cd2d235),
	.w8(32'h3c03addd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab05d27),
	.w1(32'h3b3ce868),
	.w2(32'hbcda32f3),
	.w3(32'hbc1caeda),
	.w4(32'hbb331c5b),
	.w5(32'h3ad503cd),
	.w6(32'hba14f464),
	.w7(32'hbab2bfe8),
	.w8(32'hbc2236d0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7458),
	.w1(32'hbbb1d50d),
	.w2(32'hbc4826d4),
	.w3(32'hbbceaef7),
	.w4(32'hbbdf2242),
	.w5(32'hbcb7bc8b),
	.w6(32'h3bafc016),
	.w7(32'h3bfa0a7f),
	.w8(32'hbc8ae7bf),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c825),
	.w1(32'hbba1c039),
	.w2(32'h3a929c64),
	.w3(32'hbbbd9ea0),
	.w4(32'hbb81d3f9),
	.w5(32'hbc0bea85),
	.w6(32'h3b3afe54),
	.w7(32'hb9cffc75),
	.w8(32'hbb548244),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7934c0b),
	.w1(32'h3a70a263),
	.w2(32'h3b2929fd),
	.w3(32'hbb3be08b),
	.w4(32'h387cd3a0),
	.w5(32'hbb35cba5),
	.w6(32'h3b8eb578),
	.w7(32'h3bde8cc6),
	.w8(32'h397deae1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359c10),
	.w1(32'h3b6d2a7a),
	.w2(32'hba388947),
	.w3(32'hbb8da2cc),
	.w4(32'hbb063e17),
	.w5(32'hbbbe6350),
	.w6(32'h3b76d356),
	.w7(32'h3ac9f5e9),
	.w8(32'hbaf867ac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7848),
	.w1(32'h3b934dda),
	.w2(32'hb8aa4fe8),
	.w3(32'h3a92ad45),
	.w4(32'hbadc3c69),
	.w5(32'hbb7b953e),
	.w6(32'h3a968114),
	.w7(32'hba955d28),
	.w8(32'hbb382ea2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23c57a),
	.w1(32'hbba7c80b),
	.w2(32'hba611358),
	.w3(32'hbb4110c1),
	.w4(32'hbbefedad),
	.w5(32'hbbe82e2d),
	.w6(32'h3a9c95b3),
	.w7(32'h39caa48f),
	.w8(32'h3b1e7e1f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd46a5),
	.w1(32'h3af8d3c1),
	.w2(32'h3b07ad11),
	.w3(32'hbb8f8433),
	.w4(32'hba76168f),
	.w5(32'hbba9358d),
	.w6(32'h3bd52214),
	.w7(32'h3c3e40c7),
	.w8(32'h3b311307),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bc58d),
	.w1(32'hbbd7f964),
	.w2(32'hbc291803),
	.w3(32'hbb1180ba),
	.w4(32'hbc58c78f),
	.w5(32'hbcb7dfd6),
	.w6(32'h3b8d3216),
	.w7(32'h3ca2e25a),
	.w8(32'h3c540fea),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8afa0f),
	.w1(32'h39dfb97f),
	.w2(32'h3b2fa979),
	.w3(32'hbc2a3f15),
	.w4(32'h3bb861ef),
	.w5(32'h3b99c5ce),
	.w6(32'hbba17fe8),
	.w7(32'hbbbc0757),
	.w8(32'hbc05aff0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba91aed),
	.w1(32'hbc1e39cd),
	.w2(32'hbd19c252),
	.w3(32'hba56bb97),
	.w4(32'h3b167c3f),
	.w5(32'hbcec9415),
	.w6(32'hb9a9c98a),
	.w7(32'h3c135ac4),
	.w8(32'hbb245e71),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c324d),
	.w1(32'hbb20d7b4),
	.w2(32'h3ba63ef6),
	.w3(32'hbc284921),
	.w4(32'h3bedd9f0),
	.w5(32'h3baccbf7),
	.w6(32'h3bd9bd3a),
	.w7(32'h3a33e9f0),
	.w8(32'hbbbca349),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b2ab),
	.w1(32'hbc425515),
	.w2(32'hbc5c1e2a),
	.w3(32'hbbe97eb0),
	.w4(32'hbb9515d8),
	.w5(32'hbc5de665),
	.w6(32'hbc16cc63),
	.w7(32'hbc0de8ec),
	.w8(32'hbc256cdc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5748de),
	.w1(32'hbac776b8),
	.w2(32'hbaec483a),
	.w3(32'h3a9cb905),
	.w4(32'hbc5bcf26),
	.w5(32'hbcc502db),
	.w6(32'h3c46317b),
	.w7(32'h3ca06813),
	.w8(32'h3bf122ca),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba61de4),
	.w1(32'h3ac22e82),
	.w2(32'h3b3f5211),
	.w3(32'hbc44115a),
	.w4(32'hba6057df),
	.w5(32'hbbc3adc2),
	.w6(32'h3c08e64e),
	.w7(32'h3c6470a7),
	.w8(32'h3b1c9c62),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1aee4),
	.w1(32'h3b5a5930),
	.w2(32'h3b6c10c4),
	.w3(32'hbb460dd4),
	.w4(32'h3abbcfdd),
	.w5(32'hba06e4b1),
	.w6(32'h3aa1d046),
	.w7(32'hba6df232),
	.w8(32'hbb587540),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba283ab6),
	.w1(32'h3b1bd5b5),
	.w2(32'h3b8506bd),
	.w3(32'hba68f297),
	.w4(32'h3b687a8b),
	.w5(32'h3b95d5b9),
	.w6(32'hb97f7499),
	.w7(32'hbba45ef8),
	.w8(32'hbbcc39c4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd448),
	.w1(32'hbb9b2a7c),
	.w2(32'hbce3f02a),
	.w3(32'h39daef47),
	.w4(32'hbc333729),
	.w5(32'hbcc206b2),
	.w6(32'hbc79cc9e),
	.w7(32'hbb9e7257),
	.w8(32'hbc36d023),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f3cb4),
	.w1(32'h3bb553d2),
	.w2(32'hbb077818),
	.w3(32'hbc3728a5),
	.w4(32'hbad5a206),
	.w5(32'hbb9950b8),
	.w6(32'h3c019de7),
	.w7(32'h3c41b832),
	.w8(32'h3baaec61),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0a810),
	.w1(32'h3ad7db83),
	.w2(32'h39d2a661),
	.w3(32'h3bc844aa),
	.w4(32'h3b36d2ae),
	.w5(32'h393ae528),
	.w6(32'h3b0d391d),
	.w7(32'h3bddb375),
	.w8(32'h3a56e357),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1564f),
	.w1(32'h3a706013),
	.w2(32'h3bcd1a04),
	.w3(32'hba9ca2ce),
	.w4(32'h3b0782fc),
	.w5(32'h3c197944),
	.w6(32'hbb2b9579),
	.w7(32'hbaaa4a5f),
	.w8(32'hbb3818fe),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9274c3),
	.w1(32'h3b6b5210),
	.w2(32'h3b8623da),
	.w3(32'h3bd4f648),
	.w4(32'h3aadedbb),
	.w5(32'hbac12688),
	.w6(32'h3b3e540c),
	.w7(32'h3b63c0fd),
	.w8(32'hba96ad95),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c40fb),
	.w1(32'hbc459b59),
	.w2(32'hbd405ce3),
	.w3(32'hbb8f52e2),
	.w4(32'hbc1cddb1),
	.w5(32'hbc50f6c2),
	.w6(32'hbc863e04),
	.w7(32'hbbe15ee9),
	.w8(32'hbc9038f7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93cf1c),
	.w1(32'hbc0a48bf),
	.w2(32'h3b0cf7fc),
	.w3(32'hbbfde5c7),
	.w4(32'hbb300329),
	.w5(32'h3c945590),
	.w6(32'hbc49f924),
	.w7(32'hbc9ce849),
	.w8(32'hbc19865d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8114c),
	.w1(32'hbc1f3fb1),
	.w2(32'hbc004225),
	.w3(32'h3b8d6169),
	.w4(32'hbb94937e),
	.w5(32'hbb473268),
	.w6(32'hbbbf08da),
	.w7(32'hbb9298a5),
	.w8(32'h394be58e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b70e3),
	.w1(32'h3a95e191),
	.w2(32'h3b11dda2),
	.w3(32'hbaef3bcf),
	.w4(32'h3a0440e7),
	.w5(32'h3b18d734),
	.w6(32'h39c72e52),
	.w7(32'h3b628070),
	.w8(32'h3a4ad274),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ed38d),
	.w1(32'h3c1f5172),
	.w2(32'h3bcf8d49),
	.w3(32'h3b58543d),
	.w4(32'h3c6ac9ab),
	.w5(32'h3c2abe7d),
	.w6(32'hbbd54dbd),
	.w7(32'h3b8b9f78),
	.w8(32'h3b4d5e97),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule