module layer_10_featuremap_155(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bf378),
	.w1(32'hbb00d8d4),
	.w2(32'hbaa934a6),
	.w3(32'hbaa134fb),
	.w4(32'hbb28ca07),
	.w5(32'hbb2aab33),
	.w6(32'hba78a6d9),
	.w7(32'hbacee023),
	.w8(32'hbaaff2b3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c3a04),
	.w1(32'hb9b35267),
	.w2(32'h39e70761),
	.w3(32'hbb17ba60),
	.w4(32'hbab35f57),
	.w5(32'h399ba6a2),
	.w6(32'hb9c5a2f8),
	.w7(32'h3990fc8e),
	.w8(32'h3a05e898),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a522438),
	.w1(32'hbabca0c2),
	.w2(32'hbad10dc0),
	.w3(32'h391e70a9),
	.w4(32'hb8d0e124),
	.w5(32'h37ffbbca),
	.w6(32'hbade57a1),
	.w7(32'hbb104057),
	.w8(32'hba183236),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91053b0),
	.w1(32'h3b946bb4),
	.w2(32'h3a487afa),
	.w3(32'hb92b5fb3),
	.w4(32'hbb1a1c9b),
	.w5(32'hbae3239d),
	.w6(32'hbb23cb57),
	.w7(32'hbb0e4de1),
	.w8(32'hbabab3c4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396546),
	.w1(32'hbad3a05c),
	.w2(32'hbadb3004),
	.w3(32'h39802650),
	.w4(32'h396231a8),
	.w5(32'hba200218),
	.w6(32'hba5a496f),
	.w7(32'hbb322a82),
	.w8(32'hba784e85),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad0472),
	.w1(32'h3a8d9a43),
	.w2(32'hbb0a2779),
	.w3(32'h3afd87f2),
	.w4(32'h3a387a66),
	.w5(32'hbadc9c2f),
	.w6(32'h3a68ffff),
	.w7(32'hba38e021),
	.w8(32'hbab13c72),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22f606),
	.w1(32'hbb0ee50e),
	.w2(32'hba4ea23c),
	.w3(32'hbb31d1f9),
	.w4(32'hbadcf921),
	.w5(32'hb8fba6d4),
	.w6(32'hbae69fdf),
	.w7(32'hbafc0bcb),
	.w8(32'hba7a1ac5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39a2c7),
	.w1(32'h39a11743),
	.w2(32'hba851c18),
	.w3(32'hba7a91c8),
	.w4(32'h3a81b9eb),
	.w5(32'hb9472167),
	.w6(32'h39d44edb),
	.w7(32'hba0ac5a0),
	.w8(32'hb9d3ffa0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fcb94),
	.w1(32'hba778935),
	.w2(32'hbac59164),
	.w3(32'hba86e993),
	.w4(32'hb9fbfe0f),
	.w5(32'hb9b1cd16),
	.w6(32'hbac01d8a),
	.w7(32'hba89e6e6),
	.w8(32'hba008cb9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f794a),
	.w1(32'h3aec4e2d),
	.w2(32'h39296ca9),
	.w3(32'h3941eaed),
	.w4(32'h393b38e4),
	.w5(32'hb9ec91c0),
	.w6(32'h3abe68aa),
	.w7(32'h3a152489),
	.w8(32'hba98222d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e06e5),
	.w1(32'hbb6f8e2d),
	.w2(32'hbaa3528d),
	.w3(32'hbaf66be7),
	.w4(32'h3b1360c8),
	.w5(32'h3b291efb),
	.w6(32'hbb8445a5),
	.w7(32'hbb3f683c),
	.w8(32'hbb035718),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee474f),
	.w1(32'hba50dfdd),
	.w2(32'hba5d478f),
	.w3(32'h3b46faa9),
	.w4(32'h390ce99a),
	.w5(32'hba53dbc1),
	.w6(32'h3a86509f),
	.w7(32'hba026d45),
	.w8(32'hba13f17c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8891c3),
	.w1(32'h3a508c4a),
	.w2(32'h38cb2e8e),
	.w3(32'h3aa9859b),
	.w4(32'hb977efd9),
	.w5(32'hb97c62e9),
	.w6(32'h3a525790),
	.w7(32'h3a7bf465),
	.w8(32'h3a007e09),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392da56f),
	.w1(32'h397b042b),
	.w2(32'hbb4ab6a4),
	.w3(32'hb785c669),
	.w4(32'h3ad30a21),
	.w5(32'hbb04dfbf),
	.w6(32'h3a8fcf0e),
	.w7(32'hbaad4382),
	.w8(32'hbb26e471),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5802b9),
	.w1(32'hbaaacf6b),
	.w2(32'h3a7e4533),
	.w3(32'hbb6f460b),
	.w4(32'hbb47ee05),
	.w5(32'hb96b76e9),
	.w6(32'hbabfdb33),
	.w7(32'hba947745),
	.w8(32'h3a4b6f4e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad74b24),
	.w1(32'hbaad946b),
	.w2(32'hba5a4b68),
	.w3(32'h3ae4162f),
	.w4(32'hba05dacd),
	.w5(32'hb8a49532),
	.w6(32'hba825790),
	.w7(32'hb9ff71da),
	.w8(32'hba62f6a5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba540606),
	.w1(32'hbb3312fe),
	.w2(32'hbb7714af),
	.w3(32'hba985452),
	.w4(32'h3b31fb73),
	.w5(32'h3b4b0b3b),
	.w6(32'hbb689682),
	.w7(32'hbb822766),
	.w8(32'h3a82f383),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae116cf),
	.w1(32'hbaa295f6),
	.w2(32'hba36256c),
	.w3(32'h3b93463c),
	.w4(32'hbb24635d),
	.w5(32'hba830959),
	.w6(32'hbaab18b4),
	.w7(32'hbabcb9af),
	.w8(32'hb867c8b9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872050),
	.w1(32'hba11c81b),
	.w2(32'hb858e337),
	.w3(32'h36e718b4),
	.w4(32'h39c86e41),
	.w5(32'h3abd243d),
	.w6(32'hb90ae6e4),
	.w7(32'hb95a409e),
	.w8(32'h3a9c3114),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacdf21),
	.w1(32'hba868aeb),
	.w2(32'hb90f0121),
	.w3(32'h3a6a1b67),
	.w4(32'hb9caf703),
	.w5(32'h3a37dc82),
	.w6(32'hba7876fa),
	.w7(32'hb9195a51),
	.w8(32'hba189125),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb44eed60),
	.w1(32'h3b4e1cab),
	.w2(32'hbb452f0e),
	.w3(32'hba11ee1a),
	.w4(32'h3a3f01de),
	.w5(32'hbacb3350),
	.w6(32'h3b2210f0),
	.w7(32'h39a0a21c),
	.w8(32'hb89c4645),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92996d3),
	.w1(32'h3ac7fa44),
	.w2(32'h3b8bf9bc),
	.w3(32'hba31d790),
	.w4(32'h3b2c231a),
	.w5(32'h3b6e75cf),
	.w6(32'h39d4872b),
	.w7(32'hb8f8583f),
	.w8(32'hb93a9d58),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9033c),
	.w1(32'h3b82eb0e),
	.w2(32'h3bcd3510),
	.w3(32'h3b405f92),
	.w4(32'h3af3284a),
	.w5(32'h3c1091a7),
	.w6(32'hbb48947e),
	.w7(32'h3b41fc88),
	.w8(32'h3b53130d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e837f),
	.w1(32'hb9dec3f6),
	.w2(32'hba9bd827),
	.w3(32'h3c219110),
	.w4(32'h3a2b81b1),
	.w5(32'hb9220791),
	.w6(32'h3a13c6b7),
	.w7(32'hb78efbf6),
	.w8(32'h38acab34),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804624),
	.w1(32'hb916a453),
	.w2(32'h3946eb77),
	.w3(32'hba823203),
	.w4(32'hb99b7666),
	.w5(32'h38319060),
	.w6(32'hbab7c6ba),
	.w7(32'hb98ef903),
	.w8(32'h3a165755),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99a422),
	.w1(32'hbb69ed8a),
	.w2(32'hbb474b6e),
	.w3(32'h3a4e5edc),
	.w4(32'h3abc27f0),
	.w5(32'h3b3081bd),
	.w6(32'hbb689d97),
	.w7(32'hbae8694d),
	.w8(32'hbb5c1f63),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a355),
	.w1(32'h39b49477),
	.w2(32'h3a28e04c),
	.w3(32'h3a987e5e),
	.w4(32'h3a4f0bcf),
	.w5(32'h3af94d57),
	.w6(32'h3923d1e3),
	.w7(32'h3a383dc1),
	.w8(32'hb915054a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4a4a7),
	.w1(32'h39aadc37),
	.w2(32'h3b46f2a6),
	.w3(32'h39b0c55b),
	.w4(32'h3ae90b05),
	.w5(32'h3aa8ae73),
	.w6(32'hb9300531),
	.w7(32'h3a5e3824),
	.w8(32'h3ab10849),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af41c03),
	.w1(32'hb9426468),
	.w2(32'hbb97ac85),
	.w3(32'h39087a1f),
	.w4(32'h3b5c5d5c),
	.w5(32'h3b4fbf5c),
	.w6(32'hb914a5eb),
	.w7(32'hbb3677b4),
	.w8(32'h3b2b1d2f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b631393),
	.w1(32'h3bc18326),
	.w2(32'hba09679e),
	.w3(32'h3c051a14),
	.w4(32'h3baa3752),
	.w5(32'hbacde664),
	.w6(32'h3b5dfb17),
	.w7(32'hbb58d0eb),
	.w8(32'h3b0ed3da),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01179),
	.w1(32'h3b18194a),
	.w2(32'hba3587bb),
	.w3(32'h3ac6086f),
	.w4(32'h3ac68cbc),
	.w5(32'h39f3edcf),
	.w6(32'h3b0458d7),
	.w7(32'h3aa8e176),
	.w8(32'h3a329b62),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bdfef),
	.w1(32'h3a438008),
	.w2(32'hb945ec5a),
	.w3(32'h39eeb223),
	.w4(32'h38bdd997),
	.w5(32'h3a10f81f),
	.w6(32'h3a29a8a4),
	.w7(32'h3aaa4d70),
	.w8(32'h39c8fa2a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b71164),
	.w1(32'hba3b1102),
	.w2(32'h3a2e7f62),
	.w3(32'hb91c817a),
	.w4(32'h3a710ab8),
	.w5(32'h3b2ec9ee),
	.w6(32'hba5bdc54),
	.w7(32'h39e9a56b),
	.w8(32'h381da245),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d9edb),
	.w1(32'hbaa3d917),
	.w2(32'h3bc507c7),
	.w3(32'h3aa66fbe),
	.w4(32'hbaaab883),
	.w5(32'h3c0dad02),
	.w6(32'hbb2ef6f6),
	.w7(32'h3b5ebbab),
	.w8(32'h3958d9ac),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54ff67),
	.w1(32'hb90c3cfb),
	.w2(32'hba0d8481),
	.w3(32'h3aa61e92),
	.w4(32'hba7e9b7f),
	.w5(32'hb97c6e54),
	.w6(32'hba61f0ad),
	.w7(32'hbab73f9b),
	.w8(32'hbada9d3e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6c7a1),
	.w1(32'h3a050de9),
	.w2(32'hb97c9d1b),
	.w3(32'hbac512d9),
	.w4(32'h3a632107),
	.w5(32'h3ab64af0),
	.w6(32'h3a18eb33),
	.w7(32'h3aa6b095),
	.w8(32'h3a517ca7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f343e),
	.w1(32'hb9c01700),
	.w2(32'hb8be98b6),
	.w3(32'h38ba1a43),
	.w4(32'hbad30a14),
	.w5(32'hb9feec4d),
	.w6(32'hb9adf350),
	.w7(32'h399577ff),
	.w8(32'h3a1efe6b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fe517),
	.w1(32'hb9e789d2),
	.w2(32'h39000d34),
	.w3(32'hb89ef13d),
	.w4(32'hba95bbfa),
	.w5(32'h39a4a8dd),
	.w6(32'hba3729b6),
	.w7(32'hba4a5e94),
	.w8(32'h3962f805),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52187d),
	.w1(32'hba7a903e),
	.w2(32'hba923201),
	.w3(32'h3712eabf),
	.w4(32'hba1a43f6),
	.w5(32'hb9fc062f),
	.w6(32'hb9efae8d),
	.w7(32'hbaa076b1),
	.w8(32'hba69f58d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fd211),
	.w1(32'hbab64a51),
	.w2(32'hba5c3164),
	.w3(32'hbabb2d57),
	.w4(32'hba668274),
	.w5(32'hb8da1bee),
	.w6(32'hba869956),
	.w7(32'hbab3e0a5),
	.w8(32'hba151e59),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1295a),
	.w1(32'h3c02a2de),
	.w2(32'h3bc327a6),
	.w3(32'hb932ee8a),
	.w4(32'h3b9d575b),
	.w5(32'h3b9c820e),
	.w6(32'h3bad2fb8),
	.w7(32'h3b6c0aa8),
	.w8(32'h3b9e952a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8c93),
	.w1(32'hbb13ab68),
	.w2(32'hbaaec3a4),
	.w3(32'h3b763073),
	.w4(32'hba9b81a1),
	.w5(32'hb9f4527a),
	.w6(32'hba6f7b8f),
	.w7(32'hba6bd747),
	.w8(32'hba293cfa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a85fb),
	.w1(32'h393acaf0),
	.w2(32'hba615606),
	.w3(32'hba92840d),
	.w4(32'hba3ee4ba),
	.w5(32'hb9e07c9c),
	.w6(32'h3756f3d4),
	.w7(32'h39fc1702),
	.w8(32'hba0593c0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac674),
	.w1(32'h3b0236fe),
	.w2(32'h3adf830b),
	.w3(32'hba44e9ef),
	.w4(32'h3a96d234),
	.w5(32'h3a84ced3),
	.w6(32'h3b256a35),
	.w7(32'h3ab4398c),
	.w8(32'hba9ee447),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1c99),
	.w1(32'hbaca793b),
	.w2(32'hbac6061b),
	.w3(32'hbb3318ef),
	.w4(32'hba86e687),
	.w5(32'hba7e45c2),
	.w6(32'hbb0ab3af),
	.w7(32'hbb316af2),
	.w8(32'hba664b19),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5872d),
	.w1(32'hba7f57ef),
	.w2(32'h399cec9b),
	.w3(32'hba2fe020),
	.w4(32'h393f5f7f),
	.w5(32'hb94b79f2),
	.w6(32'hbab371d1),
	.w7(32'hba7a0c6c),
	.w8(32'hba7edfd9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fd864),
	.w1(32'hb95cc203),
	.w2(32'h3a973083),
	.w3(32'hbace20d9),
	.w4(32'hb8104721),
	.w5(32'h3ae453dc),
	.w6(32'h3a2ad7dd),
	.w7(32'hbb03dc88),
	.w8(32'hba8afc54),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa54550),
	.w1(32'hba86827d),
	.w2(32'h3aa4966e),
	.w3(32'h3b166cce),
	.w4(32'h3b96a718),
	.w5(32'h3c1fcffc),
	.w6(32'hbb14ca01),
	.w7(32'h3a7f27e7),
	.w8(32'h3b5b604d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4adf),
	.w1(32'h3806ad0a),
	.w2(32'hba06dbcb),
	.w3(32'h3c255c83),
	.w4(32'hb9bba16b),
	.w5(32'h3a24330f),
	.w6(32'hb955abc3),
	.w7(32'h396e05be),
	.w8(32'hba89ff5f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5894c),
	.w1(32'h38addba6),
	.w2(32'hba1181b2),
	.w3(32'hbac60d48),
	.w4(32'h3a22c189),
	.w5(32'hb98dc716),
	.w6(32'h39bf285d),
	.w7(32'hb932f239),
	.w8(32'hb942d71b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba874024),
	.w1(32'hba97652d),
	.w2(32'h3a997f82),
	.w3(32'hba6532c3),
	.w4(32'hba56ad08),
	.w5(32'h3a6551cf),
	.w6(32'h39b63dfc),
	.w7(32'h3adef2c1),
	.w8(32'hb9ed7713),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17be2f),
	.w1(32'hbaa8f4fe),
	.w2(32'h3b76d7ae),
	.w3(32'hba8d41ee),
	.w4(32'h3b7c19ba),
	.w5(32'h3af49a66),
	.w6(32'hbaf28c74),
	.w7(32'h385f5ee7),
	.w8(32'hbabeb551),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887546),
	.w1(32'h3b39285b),
	.w2(32'h3ad276e2),
	.w3(32'h388a4ff0),
	.w4(32'h3b1aa998),
	.w5(32'h3aca5a48),
	.w6(32'h3b333a97),
	.w7(32'h3b48f208),
	.w8(32'h3aaf39db),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab83312),
	.w1(32'hb9429432),
	.w2(32'hbb00c9fe),
	.w3(32'hba80f59e),
	.w4(32'hb9f1b14d),
	.w5(32'hba24bfa8),
	.w6(32'h37f4ad13),
	.w7(32'hbaaeab3d),
	.w8(32'hbac67f79),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a7040),
	.w1(32'h3a401a91),
	.w2(32'h39b45c0e),
	.w3(32'h39cdcb1c),
	.w4(32'hba286d6d),
	.w5(32'h3a344254),
	.w6(32'h3a18c679),
	.w7(32'h3b008bfa),
	.w8(32'h3a27e0a1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399309fa),
	.w1(32'h3c25cdbe),
	.w2(32'h3ab4adc8),
	.w3(32'hba2dcfb2),
	.w4(32'h3bbfb7d8),
	.w5(32'hbac895f0),
	.w6(32'h3c246084),
	.w7(32'h3b080627),
	.w8(32'h3c35bec2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3dff44),
	.w1(32'h3b13419c),
	.w2(32'h3b6a2ee6),
	.w3(32'h3bce3bbf),
	.w4(32'h39051a40),
	.w5(32'h3b073edd),
	.w6(32'h3b2a6178),
	.w7(32'h3b961d02),
	.w8(32'h3b21c506),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b794),
	.w1(32'hb813d1f0),
	.w2(32'h3ab28861),
	.w3(32'h3a007f5a),
	.w4(32'h39d67e0a),
	.w5(32'h39ec8913),
	.w6(32'h3a5ed061),
	.w7(32'h3ab106e6),
	.w8(32'h3a96f80d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa71b45),
	.w1(32'hba674b0c),
	.w2(32'hba02da77),
	.w3(32'h3a9011d9),
	.w4(32'hba73b08c),
	.w5(32'hb8c6713b),
	.w6(32'hba935f60),
	.w7(32'hba98a0f1),
	.w8(32'hba15601c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcc11c),
	.w1(32'hb921009e),
	.w2(32'hba5996ec),
	.w3(32'hb9c18166),
	.w4(32'h39325da7),
	.w5(32'hb996272e),
	.w6(32'h38af0a10),
	.w7(32'hb965b8d5),
	.w8(32'h38d6d2b1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8f88d),
	.w1(32'hbaa2df8a),
	.w2(32'hbaa60765),
	.w3(32'hba38b8cb),
	.w4(32'hba01d6e9),
	.w5(32'h3a1a2069),
	.w6(32'hb8f12f9e),
	.w7(32'hbaa46bf2),
	.w8(32'hb9de6b2f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37596b6b),
	.w1(32'h39f3facd),
	.w2(32'hba1bb2b1),
	.w3(32'h39a3545f),
	.w4(32'h3a28ae00),
	.w5(32'h37e9b29b),
	.w6(32'h3a68451b),
	.w7(32'h38585193),
	.w8(32'h387b16b1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba724e5c),
	.w1(32'hbb1031d1),
	.w2(32'h3a3898c7),
	.w3(32'hb9ef62be),
	.w4(32'hbac1a29f),
	.w5(32'h3b2a7d1a),
	.w6(32'hb9c6f4bb),
	.w7(32'h3a55fb53),
	.w8(32'h3a86da8d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a276467),
	.w1(32'h3a84733e),
	.w2(32'h3a4d6b29),
	.w3(32'h3b0f932c),
	.w4(32'h3974df97),
	.w5(32'h39a3196f),
	.w6(32'h3a9b2fae),
	.w7(32'h39e5b5f1),
	.w8(32'hbaa3e4bf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e864),
	.w1(32'hbaefd41b),
	.w2(32'hbb05db50),
	.w3(32'hbb0032ed),
	.w4(32'hbb255c73),
	.w5(32'hbab5a0f7),
	.w6(32'hbb15e57a),
	.w7(32'hbb1ee480),
	.w8(32'hba6da802),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db30ca),
	.w1(32'h3a9d9ebe),
	.w2(32'h3b4d320b),
	.w3(32'hb97847f3),
	.w4(32'h3a60feb4),
	.w5(32'h39f448cb),
	.w6(32'h398ee49b),
	.w7(32'h3b1c2976),
	.w8(32'h3aa477b8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b0ea5),
	.w1(32'h3b9380ad),
	.w2(32'h3baa3b97),
	.w3(32'hba379449),
	.w4(32'h3b4de1dc),
	.w5(32'h3b85e321),
	.w6(32'h3b4927da),
	.w7(32'h3b4dc19a),
	.w8(32'h3b9227d3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf515a7),
	.w1(32'h3bed07ee),
	.w2(32'h3bfc407a),
	.w3(32'h3b0372a2),
	.w4(32'h3aa55206),
	.w5(32'h3c045ce9),
	.w6(32'hb9f38df3),
	.w7(32'h3b8c0011),
	.w8(32'h3b1f8bd7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1043ba),
	.w1(32'hba4deff3),
	.w2(32'hba69b033),
	.w3(32'h3b9c9b38),
	.w4(32'hb9a77b7f),
	.w5(32'hb692f7e9),
	.w6(32'hb9c7d365),
	.w7(32'hb80db300),
	.w8(32'hba193e43),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba937b1c),
	.w1(32'hbaa79368),
	.w2(32'hb80d7c29),
	.w3(32'hba4f4074),
	.w4(32'h3876f694),
	.w5(32'hba48c3f1),
	.w6(32'hbab9d5a3),
	.w7(32'hba361c73),
	.w8(32'hbb06cb54),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bdf4b),
	.w1(32'hb9c4a3c8),
	.w2(32'hb8cb17bd),
	.w3(32'hbacfbab9),
	.w4(32'hba848317),
	.w5(32'h395ff0fb),
	.w6(32'hba132f89),
	.w7(32'h35baf5e6),
	.w8(32'h3a4041c7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949916),
	.w1(32'hba0bf80f),
	.w2(32'hba4852fc),
	.w3(32'h39309d85),
	.w4(32'hba0f22d8),
	.w5(32'hb813ddb4),
	.w6(32'hb9719e8f),
	.w7(32'hb983b393),
	.w8(32'h3986ffd1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39904354),
	.w1(32'hb9ea9945),
	.w2(32'hba67d0b4),
	.w3(32'hb92894ed),
	.w4(32'hb88a3b1d),
	.w5(32'hb9ae8d7d),
	.w6(32'hb8e67c06),
	.w7(32'hb9c80e3e),
	.w8(32'hb68a8c21),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986e4bb),
	.w1(32'h3a756465),
	.w2(32'hba224357),
	.w3(32'hba28b825),
	.w4(32'h3a28a365),
	.w5(32'h3a97b6fc),
	.w6(32'h3aaec2d6),
	.w7(32'h3ad084da),
	.w8(32'h3a3341dc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c13ab0),
	.w1(32'hba8b3ffa),
	.w2(32'hb9f0c6ed),
	.w3(32'hb9549939),
	.w4(32'hb9f53079),
	.w5(32'hb9701abd),
	.w6(32'hba4bef46),
	.w7(32'hba7a982d),
	.w8(32'hba05de6e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c76bc3),
	.w1(32'hb89372b7),
	.w2(32'h3b0509b2),
	.w3(32'hba0589ff),
	.w4(32'h39e6b59a),
	.w5(32'h3b26911c),
	.w6(32'h3b345081),
	.w7(32'h3b9dd8e5),
	.w8(32'h38eb06f7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadff93b),
	.w1(32'h3ac0cce0),
	.w2(32'hba411791),
	.w3(32'h3b0447e9),
	.w4(32'h3b1aae24),
	.w5(32'hb91d1c42),
	.w6(32'h3abfd1d8),
	.w7(32'hb9319e7e),
	.w8(32'hba2a2741),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3501),
	.w1(32'hb9363196),
	.w2(32'hb9b0f2f5),
	.w3(32'hbab179b6),
	.w4(32'h39254580),
	.w5(32'h3a7f72ac),
	.w6(32'h3a8072b7),
	.w7(32'h3a4283ae),
	.w8(32'h3ac78396),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7965e),
	.w1(32'hbad01c00),
	.w2(32'hbaea7146),
	.w3(32'h3ab526d0),
	.w4(32'hbaef9ef1),
	.w5(32'h3ab5ba98),
	.w6(32'hba8aef14),
	.w7(32'h3b0e2f88),
	.w8(32'hbaa7984e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeed635),
	.w1(32'h3b2fcc01),
	.w2(32'hbae7130e),
	.w3(32'h3a49b1c7),
	.w4(32'h3aefb8ac),
	.w5(32'h392cfa37),
	.w6(32'h3b05b9d3),
	.w7(32'h3a8584ca),
	.w8(32'h39998037),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990a4cb),
	.w1(32'h3bb3cea0),
	.w2(32'h3c0cefcb),
	.w3(32'h3a14e4c6),
	.w4(32'h3b865ab3),
	.w5(32'h3c3cbadc),
	.w6(32'h3b4061a2),
	.w7(32'h3bf312ff),
	.w8(32'h3bd37b20),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38f45f),
	.w1(32'hbab2a8ab),
	.w2(32'hba6783ee),
	.w3(32'h3c2c1b7f),
	.w4(32'hbabc5389),
	.w5(32'hba8e6130),
	.w6(32'hb95d7af9),
	.w7(32'hba3a9665),
	.w8(32'hba921715),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4204),
	.w1(32'h3a8ef576),
	.w2(32'h3a649087),
	.w3(32'hbaf1d764),
	.w4(32'h3b21b19a),
	.w5(32'h3b3c4cd3),
	.w6(32'h3a6f7027),
	.w7(32'h3a98feee),
	.w8(32'h3b24a3c5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2effa9),
	.w1(32'hbaa7ec65),
	.w2(32'hba826ad1),
	.w3(32'h3b15aa40),
	.w4(32'hba928c6c),
	.w5(32'hb9849926),
	.w6(32'hba97ef87),
	.w7(32'hbaef9b36),
	.w8(32'hba897225),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3cb6b),
	.w1(32'hbb03b8b9),
	.w2(32'h39387678),
	.w3(32'hb9dc9f6f),
	.w4(32'h3c137049),
	.w5(32'h3c510919),
	.w6(32'hba7d5090),
	.w7(32'h39f2a132),
	.w8(32'hb9a9d9b2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace4ae3),
	.w1(32'h399bd599),
	.w2(32'h3a9faf38),
	.w3(32'h3c594874),
	.w4(32'hba1fffc0),
	.w5(32'hb9f38d12),
	.w6(32'h38de13b1),
	.w7(32'h3a9114e1),
	.w8(32'h3b691eba),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8905af),
	.w1(32'h39bd8515),
	.w2(32'hba33127d),
	.w3(32'h3a51eacd),
	.w4(32'h399b854b),
	.w5(32'h3a02abb9),
	.w6(32'h39ccc08c),
	.w7(32'hb9ed476f),
	.w8(32'h3b01b413),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ba1c),
	.w1(32'h3ad3805b),
	.w2(32'hba8f09df),
	.w3(32'h3aa36996),
	.w4(32'h3a89d79d),
	.w5(32'h38d43389),
	.w6(32'h3afa65b2),
	.w7(32'h3a86c6be),
	.w8(32'h3a0b9ba9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d647e),
	.w1(32'h39ec0658),
	.w2(32'h39d1027a),
	.w3(32'hb800636d),
	.w4(32'hb8e122d8),
	.w5(32'h3a1bab42),
	.w6(32'h38c90fd7),
	.w7(32'h3a0a1fe2),
	.w8(32'hb85f02a0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8c9fc),
	.w1(32'h3aebb8d1),
	.w2(32'hbaa51729),
	.w3(32'hba90128f),
	.w4(32'h3a301337),
	.w5(32'h394c155e),
	.w6(32'h3a9cccc2),
	.w7(32'h3a9656ca),
	.w8(32'h38e9bf41),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c09938),
	.w1(32'h3abd1c57),
	.w2(32'hba8617a6),
	.w3(32'hba0f7576),
	.w4(32'h39e75a45),
	.w5(32'hb9422525),
	.w6(32'h3adcb2a7),
	.w7(32'h3a804fcd),
	.w8(32'h3a015190),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ec64f),
	.w1(32'h3ab7164e),
	.w2(32'h3a49df09),
	.w3(32'h390c6fbb),
	.w4(32'hb9369c85),
	.w5(32'hb8e41485),
	.w6(32'h3a8f4292),
	.w7(32'h3a2bb085),
	.w8(32'hba3f12ce),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e1a0ee),
	.w1(32'h3b1afefa),
	.w2(32'h3b0b4002),
	.w3(32'hba94814d),
	.w4(32'h3ac15990),
	.w5(32'h3afcaa0d),
	.w6(32'h3ae9b0ee),
	.w7(32'h3b170dda),
	.w8(32'h3abe37e0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e6d89),
	.w1(32'h3bcd5398),
	.w2(32'h3ba54d84),
	.w3(32'h3aa85ce7),
	.w4(32'h3b855ae2),
	.w5(32'h3be1f897),
	.w6(32'h3b4b3c59),
	.w7(32'h3b4e4acb),
	.w8(32'h3bd80741),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b933d),
	.w1(32'hbaf8649f),
	.w2(32'hbac69121),
	.w3(32'h3c1aa878),
	.w4(32'hbaadb29d),
	.w5(32'hba1c8b3d),
	.w6(32'hbb433e63),
	.w7(32'hbb502208),
	.w8(32'hba9d6715),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9fdc2),
	.w1(32'h3a048c1b),
	.w2(32'hba614cf1),
	.w3(32'hba2d902e),
	.w4(32'hba21bea5),
	.w5(32'hb9adb21a),
	.w6(32'hba4e48f4),
	.w7(32'hb96a2dfd),
	.w8(32'hba7e63d7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab243b6),
	.w1(32'h3b071b20),
	.w2(32'h3c57f709),
	.w3(32'hb90e9c93),
	.w4(32'hbab78989),
	.w5(32'h3c6dff0d),
	.w6(32'hbb2214dc),
	.w7(32'h3c46a259),
	.w8(32'h3badfee3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085586),
	.w1(32'hbaaa30e5),
	.w2(32'h3b97e231),
	.w3(32'h3c098638),
	.w4(32'h39ab2e01),
	.w5(32'h3ba56864),
	.w6(32'hbaa9965a),
	.w7(32'h3b6e106d),
	.w8(32'h3b1019dc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10abfe),
	.w1(32'hbafad8c9),
	.w2(32'hba3ac23c),
	.w3(32'h3b6223c6),
	.w4(32'hbac2926d),
	.w5(32'h39c09485),
	.w6(32'hbae8689f),
	.w7(32'hbaef8d08),
	.w8(32'hba59a37c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12c800),
	.w1(32'h3b8c459b),
	.w2(32'h3b2b5218),
	.w3(32'hbaa1ef1c),
	.w4(32'h3b4afd4e),
	.w5(32'h3af170bd),
	.w6(32'h3b67c3cd),
	.w7(32'h3b620875),
	.w8(32'h3b7f98ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92ce81),
	.w1(32'h3b011895),
	.w2(32'h3bad560f),
	.w3(32'h3a8e79bb),
	.w4(32'hba413d18),
	.w5(32'h3b7b978c),
	.w6(32'h3b3a54df),
	.w7(32'h3b67562a),
	.w8(32'h3b85eae0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c3a7),
	.w1(32'h3a251f7e),
	.w2(32'h39ce03e2),
	.w3(32'h3b7244de),
	.w4(32'h3ae9d406),
	.w5(32'hba14caca),
	.w6(32'hba1f0c2d),
	.w7(32'h3a5a81da),
	.w8(32'h3aec4839),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26074),
	.w1(32'h3b0ffb71),
	.w2(32'hba9b4148),
	.w3(32'h3ada58c7),
	.w4(32'h3b380542),
	.w5(32'hba50cfc9),
	.w6(32'h3af2fdd3),
	.w7(32'hb9f68eb4),
	.w8(32'hba8a727b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1ca8),
	.w1(32'h3a079109),
	.w2(32'hb96d83a7),
	.w3(32'hbb2343e8),
	.w4(32'h39c2c0a1),
	.w5(32'h3a4cd489),
	.w6(32'h396f008c),
	.w7(32'h3a2345ea),
	.w8(32'h39df7d01),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef522b),
	.w1(32'h3ac1e5b7),
	.w2(32'hba09ab9e),
	.w3(32'h399995cd),
	.w4(32'h3ad831ab),
	.w5(32'hb9b11ca4),
	.w6(32'h3a51ead0),
	.w7(32'hb99945cb),
	.w8(32'hba14131b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813f36),
	.w1(32'hb9a089fc),
	.w2(32'hb998508a),
	.w3(32'hba951057),
	.w4(32'h3a1538ae),
	.w5(32'h3aa1ab08),
	.w6(32'hb993a465),
	.w7(32'hb93a15db),
	.w8(32'hb81278c2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396126dd),
	.w1(32'hbae26827),
	.w2(32'hbae602a4),
	.w3(32'hb788921a),
	.w4(32'hb9868105),
	.w5(32'hb99b52f3),
	.w6(32'hbb2e5cfa),
	.w7(32'hbb3e415d),
	.w8(32'hbac4aa6b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27343b),
	.w1(32'h3b6de4dd),
	.w2(32'hbac66b6f),
	.w3(32'hb880620c),
	.w4(32'h3ab52fd7),
	.w5(32'hba1b617d),
	.w6(32'h3b69a6dd),
	.w7(32'h3ac7bbbf),
	.w8(32'h3aaa815e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41b712),
	.w1(32'h3a8c13c4),
	.w2(32'hba388bd2),
	.w3(32'h3a0e3d43),
	.w4(32'h3ae01619),
	.w5(32'hb9f001d5),
	.w6(32'h3ab63fa1),
	.w7(32'h38578a84),
	.w8(32'hba0bb951),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabeb4c9),
	.w1(32'hbb1fb999),
	.w2(32'hbb6aeb2a),
	.w3(32'hbadf8bb8),
	.w4(32'hbb095437),
	.w5(32'hbad687ab),
	.w6(32'hbac85a30),
	.w7(32'hbad70393),
	.w8(32'hb8776d1e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba387ca6),
	.w1(32'hbac60c22),
	.w2(32'hba772e2a),
	.w3(32'h38e30dc4),
	.w4(32'hb93defb0),
	.w5(32'hb9d06761),
	.w6(32'hbac63ff8),
	.w7(32'hba8b818c),
	.w8(32'hba76f6c1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66e8b),
	.w1(32'hba8da7cd),
	.w2(32'hbb3d864c),
	.w3(32'hbadb6ec6),
	.w4(32'hba84282e),
	.w5(32'hbb0d7bbe),
	.w6(32'hb97c7c88),
	.w7(32'hbb6e3f9c),
	.w8(32'hbb553143),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87750c),
	.w1(32'hbaa9ae24),
	.w2(32'hba907d8e),
	.w3(32'hbb1a703b),
	.w4(32'hb942fa83),
	.w5(32'hb9bcb227),
	.w6(32'hba8e2393),
	.w7(32'hba2d7faf),
	.w8(32'hba5a0b94),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a19f9),
	.w1(32'hbb116135),
	.w2(32'hbb2614f0),
	.w3(32'hba467b43),
	.w4(32'hbadb3e50),
	.w5(32'hbab7fd68),
	.w6(32'hba6b414c),
	.w7(32'hba99d9be),
	.w8(32'h3a086d80),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87a79d),
	.w1(32'hbb2884d1),
	.w2(32'hba7249df),
	.w3(32'hba9c2a7c),
	.w4(32'hbb17591f),
	.w5(32'hb8f06c97),
	.w6(32'hbb2deab5),
	.w7(32'h3a3b8477),
	.w8(32'hba89d34b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf4a1),
	.w1(32'h3ad245b9),
	.w2(32'hba88347b),
	.w3(32'hbae66441),
	.w4(32'h3b0bf496),
	.w5(32'hba47a9da),
	.w6(32'h3ab4b08e),
	.w7(32'hb99e80b5),
	.w8(32'hba7097b9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6e6a0),
	.w1(32'h390cbdd8),
	.w2(32'hba82372d),
	.w3(32'hbb0053a2),
	.w4(32'h3a272a72),
	.w5(32'hb9eafd62),
	.w6(32'h3a1a8831),
	.w7(32'hb9a189fa),
	.w8(32'h384ea851),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc2383),
	.w1(32'h3a63e52d),
	.w2(32'hba90d251),
	.w3(32'hba253dfc),
	.w4(32'h3a8a12f8),
	.w5(32'hba5bf00a),
	.w6(32'h3a5c5bf4),
	.w7(32'hb9dd88e9),
	.w8(32'h38166c75),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9912ed8),
	.w1(32'h3b38bfd0),
	.w2(32'h3a8e3ab4),
	.w3(32'hba272244),
	.w4(32'h3b05f9f8),
	.w5(32'hb9281688),
	.w6(32'h3a9e349f),
	.w7(32'h39e35443),
	.w8(32'hb7b9abcd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0c92e),
	.w1(32'hbb18579f),
	.w2(32'h3b179766),
	.w3(32'hb99975a8),
	.w4(32'hbaa64ae5),
	.w5(32'h3b5ed15c),
	.w6(32'hbab8dc07),
	.w7(32'h3b09102b),
	.w8(32'h3bb493e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01737),
	.w1(32'hb9757c70),
	.w2(32'h39ebde0d),
	.w3(32'h3b9558f7),
	.w4(32'hba29a8a4),
	.w5(32'h3ab12726),
	.w6(32'hbac5a159),
	.w7(32'h384b990d),
	.w8(32'hba1e4e06),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a853e03),
	.w1(32'h387a7246),
	.w2(32'h393594d2),
	.w3(32'h39aa984a),
	.w4(32'h3817b6d7),
	.w5(32'h3958bf3a),
	.w6(32'hb9e7c7be),
	.w7(32'hb9cf4071),
	.w8(32'hba1c38ff),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03dcd2),
	.w1(32'h36c5f806),
	.w2(32'hba6332da),
	.w3(32'hb9beab50),
	.w4(32'h39e6beac),
	.w5(32'hb96a6990),
	.w6(32'h391ab2b5),
	.w7(32'hb9c75449),
	.w8(32'hb9496eba),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a2b57),
	.w1(32'h3a42bb3e),
	.w2(32'h39819780),
	.w3(32'hba96b2dd),
	.w4(32'h3a987bf7),
	.w5(32'hb8efc610),
	.w6(32'hb89ee018),
	.w7(32'hbaf3da79),
	.w8(32'hba7a4944),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72cf9e),
	.w1(32'h3b9e29eb),
	.w2(32'h3b21285d),
	.w3(32'hbaeb34d6),
	.w4(32'h3b5742d0),
	.w5(32'h3b0eb570),
	.w6(32'h3b78b66c),
	.w7(32'h3ba11b7c),
	.w8(32'h3b5d145c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeea58),
	.w1(32'h3b5b3073),
	.w2(32'hba5390e1),
	.w3(32'h3a1d5a5a),
	.w4(32'h3af19717),
	.w5(32'h3a29b75e),
	.w6(32'h3b591880),
	.w7(32'h3b0c0717),
	.w8(32'h3ab0ab81),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c92dd),
	.w1(32'h38b923ce),
	.w2(32'h37d39e4f),
	.w3(32'h39d8e0a7),
	.w4(32'hb84aca36),
	.w5(32'hb723e822),
	.w6(32'hb88c1ef7),
	.w7(32'hb9326008),
	.w8(32'hb8b3e5ac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879e584),
	.w1(32'hb963b0f5),
	.w2(32'hb8a4dca4),
	.w3(32'hb87028f3),
	.w4(32'hb8853e16),
	.w5(32'hb90dcc10),
	.w6(32'h37e77e9f),
	.w7(32'hb823a72a),
	.w8(32'hb90a8f9b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9abb9),
	.w1(32'h3761ed42),
	.w2(32'hb8aa72b6),
	.w3(32'hb8c253a0),
	.w4(32'hb912befb),
	.w5(32'hb8ad9056),
	.w6(32'h39af78c1),
	.w7(32'h38f5063e),
	.w8(32'h3930cd3d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c2b71c),
	.w1(32'h35ef01ce),
	.w2(32'h363dbeac),
	.w3(32'hb622b4bf),
	.w4(32'h352a2d3c),
	.w5(32'h348b958b),
	.w6(32'hb57b83ad),
	.w7(32'hb64fbb48),
	.w8(32'h355b3ec1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858dc50),
	.w1(32'h37c06d99),
	.w2(32'h37c8d657),
	.w3(32'h38b1a3b2),
	.w4(32'h38795cff),
	.w5(32'h389414e8),
	.w6(32'hb83236c7),
	.w7(32'hb84275ff),
	.w8(32'h362a502c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a2296),
	.w1(32'h38a98a5a),
	.w2(32'h386f6776),
	.w3(32'hb7556033),
	.w4(32'h36859895),
	.w5(32'h37c24134),
	.w6(32'hb84f0f0c),
	.w7(32'hb78cb068),
	.w8(32'h376b7018),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8213b3e),
	.w1(32'hb91a4a52),
	.w2(32'hb91de9e1),
	.w3(32'hb66cc5f9),
	.w4(32'hb890f73d),
	.w5(32'hb87b08ee),
	.w6(32'h37af0660),
	.w7(32'hb80889c2),
	.w8(32'hb7c7afd6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a48f3),
	.w1(32'hb90cd741),
	.w2(32'hb902d1e6),
	.w3(32'hb991903a),
	.w4(32'hb9612d27),
	.w5(32'hb8dec3ee),
	.w6(32'hb9e6e2c6),
	.w7(32'hb9acc17f),
	.w8(32'h37c5dcce),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7e428),
	.w1(32'h38bedb8e),
	.w2(32'h39011216),
	.w3(32'h383b2a9f),
	.w4(32'h3876da38),
	.w5(32'h393025d7),
	.w6(32'h38fcc88b),
	.w7(32'h3911ec17),
	.w8(32'h398752bd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3839c717),
	.w1(32'hb90a0275),
	.w2(32'hb9167190),
	.w3(32'h38cbab6e),
	.w4(32'hb64b42d7),
	.w5(32'hb78b2bcd),
	.w6(32'hb8101f78),
	.w7(32'h377593a4),
	.w8(32'hb7b62b03),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39094de4),
	.w1(32'h396ec378),
	.w2(32'h392758f8),
	.w3(32'hb9b9a81c),
	.w4(32'hb97c64ac),
	.w5(32'h38b96654),
	.w6(32'hb9e19f85),
	.w7(32'hb9da172f),
	.w8(32'hb8251134),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8180d),
	.w1(32'hb8a76e79),
	.w2(32'hb8aafd78),
	.w3(32'hb88fd8c6),
	.w4(32'hb8d7a0f1),
	.w5(32'hb8b9dbaf),
	.w6(32'hb93c8f5e),
	.w7(32'hb9099667),
	.w8(32'hb8599920),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea2dcd),
	.w1(32'hb8a39668),
	.w2(32'hb8ae0ac4),
	.w3(32'hb783f74e),
	.w4(32'hb860679d),
	.w5(32'hb84d75a5),
	.w6(32'hb6fa86a1),
	.w7(32'hb8330198),
	.w8(32'hb879e914),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a0269),
	.w1(32'h39142972),
	.w2(32'hb675c356),
	.w3(32'h38d907c5),
	.w4(32'h38eb6ccd),
	.w5(32'h390fe7ed),
	.w6(32'h39809514),
	.w7(32'h397d2ef1),
	.w8(32'h399812c1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a80e4),
	.w1(32'hb864f2bf),
	.w2(32'hb8770d74),
	.w3(32'h384f5e37),
	.w4(32'h37ea0261),
	.w5(32'hb7438f80),
	.w6(32'h38a74afb),
	.w7(32'h386efb98),
	.w8(32'h38037482),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38803c62),
	.w1(32'h37baf0ba),
	.w2(32'hb79b853e),
	.w3(32'h38b5e851),
	.w4(32'h367579ca),
	.w5(32'h38d672d2),
	.w6(32'h376e3ec1),
	.w7(32'h38a10086),
	.w8(32'h3940b514),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9864d19),
	.w1(32'hb870f0e7),
	.w2(32'h3860e4ea),
	.w3(32'hb9d4898f),
	.w4(32'hb940c1cc),
	.w5(32'h3886982e),
	.w6(32'hba1b6de2),
	.w7(32'hb99f5164),
	.w8(32'hb7ddc03b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363832e2),
	.w1(32'h37287170),
	.w2(32'h365344d8),
	.w3(32'h366f0388),
	.w4(32'h37261b41),
	.w5(32'h3686426c),
	.w6(32'hb598eac3),
	.w7(32'h365f5008),
	.w8(32'h358d4091),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c7a50d),
	.w1(32'h3696a08e),
	.w2(32'hb62918d9),
	.w3(32'h357dace8),
	.w4(32'h36c33f9e),
	.w5(32'h3621d370),
	.w6(32'hb5976071),
	.w7(32'h36726251),
	.w8(32'h35db1bea),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35650810),
	.w1(32'h37560b05),
	.w2(32'h36d21652),
	.w3(32'hb3b7f67f),
	.w4(32'h374fcbfb),
	.w5(32'h37d5047b),
	.w6(32'h369ffa94),
	.w7(32'h37630115),
	.w8(32'h37f1c054),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d947c),
	.w1(32'hb7b2e8df),
	.w2(32'h38d20427),
	.w3(32'hb99c7755),
	.w4(32'hb9267b2e),
	.w5(32'h380ce2a1),
	.w6(32'hb9d38d82),
	.w7(32'hb99ed802),
	.w8(32'hb9185720),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c4767),
	.w1(32'h3922a49a),
	.w2(32'hb904c8ad),
	.w3(32'h3a171a6b),
	.w4(32'h39a38f71),
	.w5(32'hb8b269af),
	.w6(32'h39fb01fd),
	.w7(32'h39e14eb6),
	.w8(32'h39301980),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360084f4),
	.w1(32'h362bcc4b),
	.w2(32'h35d035d5),
	.w3(32'h361b8d76),
	.w4(32'h3697088f),
	.w5(32'h359fbb95),
	.w6(32'h35ad8c97),
	.w7(32'h358a703a),
	.w8(32'h35cdd375),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928aeea),
	.w1(32'h37d5fcd7),
	.w2(32'h37d82f59),
	.w3(32'h39a7e905),
	.w4(32'h39288cfc),
	.w5(32'h39103718),
	.w6(32'h39b979a5),
	.w7(32'h398d4846),
	.w8(32'h3983d386),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851f7eb),
	.w1(32'hb88a1bbd),
	.w2(32'hb8f35f82),
	.w3(32'hb8280882),
	.w4(32'hb90f485c),
	.w5(32'hb7e92d82),
	.w6(32'h38f490dd),
	.w7(32'hb8b4d0e5),
	.w8(32'h371987ed),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b9ef5),
	.w1(32'h39dc5794),
	.w2(32'h3983651c),
	.w3(32'h39f25322),
	.w4(32'h39871dd2),
	.w5(32'h37ae4739),
	.w6(32'h39fb95e2),
	.w7(32'h382b772a),
	.w8(32'h38263959),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928bae6),
	.w1(32'h38c1460b),
	.w2(32'h397cc232),
	.w3(32'h3915f5fc),
	.w4(32'h386d54db),
	.w5(32'h3971d3c7),
	.w6(32'h392d9981),
	.w7(32'h38ac6dc7),
	.w8(32'h39122e8d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da7aa0),
	.w1(32'hb94d1f9c),
	.w2(32'hb8d68dc8),
	.w3(32'hb9b31406),
	.w4(32'hb9978726),
	.w5(32'hb902cb3a),
	.w6(32'hb9d4fbfe),
	.w7(32'hb9e9ee2e),
	.w8(32'hb98606f9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9460dcf),
	.w1(32'hb8487392),
	.w2(32'h383adfde),
	.w3(32'h38824c6e),
	.w4(32'h392aed7a),
	.w5(32'h393b762a),
	.w6(32'h39464f08),
	.w7(32'h390f30ea),
	.w8(32'h39566d68),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393084c0),
	.w1(32'h36ef864f),
	.w2(32'h38d5d56b),
	.w3(32'h39b4d607),
	.w4(32'h39830513),
	.w5(32'h39bada5e),
	.w6(32'h39adfcab),
	.w7(32'h399b4d0b),
	.w8(32'h39adb9aa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa2c27),
	.w1(32'h38995b8c),
	.w2(32'h397d2130),
	.w3(32'hba5314c2),
	.w4(32'hb9ec9ed7),
	.w5(32'h37a232a2),
	.w6(32'hba5cbf6a),
	.w7(32'hba3fe72f),
	.w8(32'hb8a70202),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d931c2),
	.w1(32'hb856eb30),
	.w2(32'h3798a4d8),
	.w3(32'hb7c2a6d4),
	.w4(32'hb87bf368),
	.w5(32'h3615a7a7),
	.w6(32'hb7b6ffa4),
	.w7(32'hb8b33965),
	.w8(32'hb9000348),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a42155),
	.w1(32'h380b3c53),
	.w2(32'h37c2ca7f),
	.w3(32'h371d1d9d),
	.w4(32'h37b076f3),
	.w5(32'h37b7075f),
	.w6(32'h34e9de45),
	.w7(32'h37142ef4),
	.w8(32'h375b3197),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53da9db),
	.w1(32'h366324d1),
	.w2(32'h367af4ca),
	.w3(32'hb5a34ecc),
	.w4(32'h366263f2),
	.w5(32'h36901998),
	.w6(32'h3630cd76),
	.w7(32'h36241af9),
	.w8(32'h36657247),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397455d8),
	.w1(32'h391c1b7a),
	.w2(32'h394fcd01),
	.w3(32'h382d8045),
	.w4(32'hb8c08dfa),
	.w5(32'h37cbc48d),
	.w6(32'hb715a578),
	.w7(32'hb93af003),
	.w8(32'h390a5bc2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e72b5),
	.w1(32'hb5c60176),
	.w2(32'hb67d8f26),
	.w3(32'hb715d439),
	.w4(32'hb5b12788),
	.w5(32'h35f74129),
	.w6(32'hb7885758),
	.w7(32'hb681003a),
	.w8(32'h36e0cf1a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38754e61),
	.w1(32'hb8a3a33f),
	.w2(32'hb9061605),
	.w3(32'h38a854ff),
	.w4(32'h37e1225c),
	.w5(32'h37d81f4b),
	.w6(32'h39395998),
	.w7(32'h395cdd28),
	.w8(32'h393553c3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903570e),
	.w1(32'h3899169d),
	.w2(32'h36dd8deb),
	.w3(32'h3902c885),
	.w4(32'h3885131e),
	.w5(32'h37b554ee),
	.w6(32'h37db9e4e),
	.w7(32'h38ba3cb8),
	.w8(32'hb6eb3f85),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3758e8fd),
	.w1(32'hb967438e),
	.w2(32'hb8e0aa47),
	.w3(32'h38fd9c38),
	.w4(32'hb97d45cf),
	.w5(32'hb90dfbef),
	.w6(32'h394b30aa),
	.w7(32'hb9235386),
	.w8(32'hb97c0c10),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a42db4),
	.w1(32'hb7f5bef3),
	.w2(32'h37887e31),
	.w3(32'hb872308c),
	.w4(32'hb7e4387a),
	.w5(32'h366b102b),
	.w6(32'hb75b9f33),
	.w7(32'hb786f2c0),
	.w8(32'h36acdbf8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812e751),
	.w1(32'h37e1fa74),
	.w2(32'hb740df17),
	.w3(32'h3888d7dc),
	.w4(32'h38a9977e),
	.w5(32'h38489547),
	.w6(32'h36fa0ce1),
	.w7(32'h380aadc3),
	.w8(32'h37c62f87),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901faab),
	.w1(32'h36683d5c),
	.w2(32'h3774b0c6),
	.w3(32'h36d4e242),
	.w4(32'hb81fcb89),
	.w5(32'hb7e96d5a),
	.w6(32'hb898f26b),
	.w7(32'hb8ff08d6),
	.w8(32'hb7645de9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abc6db),
	.w1(32'h386000e2),
	.w2(32'h392cee24),
	.w3(32'h39749077),
	.w4(32'h38945a18),
	.w5(32'h3995196c),
	.w6(32'h394bb46f),
	.w7(32'h3926f44c),
	.w8(32'h39d72859),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936b785),
	.w1(32'hb99ebb09),
	.w2(32'hb9d92b36),
	.w3(32'hb8bd93a2),
	.w4(32'hb9a2bd79),
	.w5(32'hb9cef6b8),
	.w6(32'hb8d3ca14),
	.w7(32'hb963c9c5),
	.w8(32'hb9ba4037),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbac87),
	.w1(32'hb8b3155d),
	.w2(32'hb9666561),
	.w3(32'h39e6f2ab),
	.w4(32'h392ea637),
	.w5(32'hb8e2c6d4),
	.w6(32'h398331a4),
	.w7(32'h39752885),
	.w8(32'h3930c3f9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c2630),
	.w1(32'h38960760),
	.w2(32'h3883fb3f),
	.w3(32'h38802a72),
	.w4(32'h387651de),
	.w5(32'h3876924c),
	.w6(32'hb712c919),
	.w7(32'hb62762fe),
	.w8(32'h38614b2c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39763531),
	.w1(32'h38b6c9a3),
	.w2(32'h3988ef3e),
	.w3(32'h39831662),
	.w4(32'h388ce885),
	.w5(32'h393e7066),
	.w6(32'h39896e7c),
	.w7(32'h39002a62),
	.w8(32'h390327b5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdd08f),
	.w1(32'hb8721dd2),
	.w2(32'hb9451293),
	.w3(32'h38b234f7),
	.w4(32'h38b38898),
	.w5(32'hb8ca3aef),
	.w6(32'h37b167b8),
	.w7(32'hb89b3cb4),
	.w8(32'hb94b847d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d71bbf),
	.w1(32'hb9659fee),
	.w2(32'hb91546f1),
	.w3(32'h38579b7f),
	.w4(32'h3851d2de),
	.w5(32'h38a7e08b),
	.w6(32'h397b8b16),
	.w7(32'h39965db8),
	.w8(32'h39a23424),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812150d),
	.w1(32'hb89d7849),
	.w2(32'hb81571ee),
	.w3(32'hb86e7ac7),
	.w4(32'hb8b21225),
	.w5(32'hb7c7dc6e),
	.w6(32'hb8a2a764),
	.w7(32'hb84dcf09),
	.w8(32'hb80c8328),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ebb44),
	.w1(32'h38688c39),
	.w2(32'h38ac47a5),
	.w3(32'hb93501e2),
	.w4(32'hb8fac8ed),
	.w5(32'h38236e33),
	.w6(32'hb9c0c681),
	.w7(32'hb96b9eff),
	.w8(32'h371f0960),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3683d4cf),
	.w1(32'hb620fdb9),
	.w2(32'hb58d9466),
	.w3(32'hb5706e0b),
	.w4(32'hb6b186cc),
	.w5(32'hb63ad757),
	.w6(32'hb681d25d),
	.w7(32'hb65f8400),
	.w8(32'hb5ab495d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da3511),
	.w1(32'hb7363d07),
	.w2(32'hb8250ac1),
	.w3(32'h390d8868),
	.w4(32'hb5899b37),
	.w5(32'hb7b6c153),
	.w6(32'h38ab54a9),
	.w7(32'h3819bfac),
	.w8(32'hb6912613),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83bd7ae),
	.w1(32'hb81f7b39),
	.w2(32'hb83d2e1a),
	.w3(32'hb76b4019),
	.w4(32'hb7915585),
	.w5(32'hb7c447f4),
	.w6(32'hb8074e25),
	.w7(32'hb7842b8b),
	.w8(32'hb777f5b6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a4057),
	.w1(32'h384e8a84),
	.w2(32'hb6c07147),
	.w3(32'hb7575b3f),
	.w4(32'h3872f32f),
	.w5(32'h3784520a),
	.w6(32'h380aea64),
	.w7(32'h38bad9c9),
	.w8(32'h389ca267),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fb6cfa),
	.w1(32'hb608cb06),
	.w2(32'hb5212f6b),
	.w3(32'hb41ab805),
	.w4(32'hb636cabb),
	.w5(32'hb549fbf5),
	.w6(32'hb4aefeba),
	.w7(32'hb601d4ed),
	.w8(32'hb5b51d9c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec3b9d),
	.w1(32'hb78e9406),
	.w2(32'hb74af8dd),
	.w3(32'hb7b6a67b),
	.w4(32'hb7212e84),
	.w5(32'h360904c7),
	.w6(32'hb7752f5b),
	.w7(32'hb5240ac1),
	.w8(32'h35e72fab),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb795984d),
	.w1(32'hb8c6265c),
	.w2(32'hb8c5984e),
	.w3(32'hb7461b24),
	.w4(32'hb8918f2a),
	.w5(32'hb8c02d35),
	.w6(32'h387bcff4),
	.w7(32'hb74a9d2e),
	.w8(32'hb8596858),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91032a9),
	.w1(32'hb9190f92),
	.w2(32'hb961e335),
	.w3(32'hb9247bff),
	.w4(32'hb9446ed0),
	.w5(32'hb972b972),
	.w6(32'hb907eda8),
	.w7(32'hb99892d6),
	.w8(32'hb97fe587),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fa2c4b),
	.w1(32'hb816bf23),
	.w2(32'hb815cb1b),
	.w3(32'hb71f017e),
	.w4(32'h37b39079),
	.w5(32'hb8276097),
	.w6(32'hb7d9a562),
	.w7(32'hb6e4c390),
	.w8(32'hb8a0dd76),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37880e4d),
	.w1(32'hb784fbb7),
	.w2(32'hb7c55f99),
	.w3(32'h374c8c34),
	.w4(32'hb8045c13),
	.w5(32'hb7abdca7),
	.w6(32'h378e68ff),
	.w7(32'hb81e609d),
	.w8(32'hb88b5acb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16f093),
	.w1(32'hb95026b5),
	.w2(32'hb811b4d3),
	.w3(32'h3a8ce0fa),
	.w4(32'h39a7ae28),
	.w5(32'h39a7c69f),
	.w6(32'h3abd915e),
	.w7(32'h3a6b9902),
	.w8(32'h3a830d32),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886ff4e),
	.w1(32'h39d192c1),
	.w2(32'h3a44e627),
	.w3(32'hb9af26a1),
	.w4(32'h386f08f1),
	.w5(32'h3a078a78),
	.w6(32'hb9fe9b21),
	.w7(32'h3899426d),
	.w8(32'h3a031321),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb850855d),
	.w1(32'hb799a04d),
	.w2(32'h37d05081),
	.w3(32'h37039c61),
	.w4(32'h372ee049),
	.w5(32'h38718fa9),
	.w6(32'hb77b385b),
	.w7(32'h37be0d52),
	.w8(32'h38656810),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c04309),
	.w1(32'h3540df1f),
	.w2(32'h362733d9),
	.w3(32'hb5888e21),
	.w4(32'h36813419),
	.w5(32'h36d851d1),
	.w6(32'h36acb4ae),
	.w7(32'h370058ba),
	.w8(32'h36abcb7d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d65787),
	.w1(32'hb906d068),
	.w2(32'hb912ddd4),
	.w3(32'hb8647a0f),
	.w4(32'hb8772f7e),
	.w5(32'hb86f7d7a),
	.w6(32'hb862d3ad),
	.w7(32'hb8876156),
	.w8(32'hb8b85859),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a48057),
	.w1(32'h36842eff),
	.w2(32'hb61bcba9),
	.w3(32'h3743af55),
	.w4(32'h37252fc6),
	.w5(32'hb62404d2),
	.w6(32'h365ccdb8),
	.w7(32'h35a164f5),
	.w8(32'hb52a6c03),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a9f672),
	.w1(32'h38d15009),
	.w2(32'h389dff4e),
	.w3(32'h38bf751a),
	.w4(32'h38db4cb7),
	.w5(32'h3901f6eb),
	.w6(32'hb77509e8),
	.w7(32'h37440a7b),
	.w8(32'h38762be7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934acbb),
	.w1(32'h3806757f),
	.w2(32'hb8fca542),
	.w3(32'hba154575),
	.w4(32'hb9df17a3),
	.w5(32'hb9154de2),
	.w6(32'hb9d99a79),
	.w7(32'hba2695d0),
	.w8(32'hb9ace6cc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f095f),
	.w1(32'h388d2c6a),
	.w2(32'hb86e03f2),
	.w3(32'h394cd27e),
	.w4(32'hb6ec0a65),
	.w5(32'hb8d4609f),
	.w6(32'h3920daee),
	.w7(32'h379ca5cd),
	.w8(32'h3941ac35),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394cbaba),
	.w1(32'h38fb3efd),
	.w2(32'hb8cccbd1),
	.w3(32'h39036f04),
	.w4(32'h38d78fdf),
	.w5(32'hb858be7a),
	.w6(32'h38826478),
	.w7(32'hb875ee90),
	.w8(32'hb921b16a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9b001),
	.w1(32'h38eb734e),
	.w2(32'hb855bb69),
	.w3(32'h3a13eb2a),
	.w4(32'h39947640),
	.w5(32'h390b3ef8),
	.w6(32'h3a352a38),
	.w7(32'h39d6b6cd),
	.w8(32'h39909beb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3719bb5e),
	.w1(32'h381d1569),
	.w2(32'hb8fb4e4f),
	.w3(32'hb7c6c1f4),
	.w4(32'hb644d96c),
	.w5(32'hb8fd631c),
	.w6(32'h384ef195),
	.w7(32'h37cb9a3d),
	.w8(32'hb81bc68f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d1b5ba),
	.w1(32'h36c78032),
	.w2(32'h372a3b02),
	.w3(32'h340c56fd),
	.w4(32'h3567f264),
	.w5(32'h36af1442),
	.w6(32'hb5bcb9c6),
	.w7(32'h354e33c6),
	.w8(32'h36a95357),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3709a805),
	.w1(32'h36214706),
	.w2(32'h37645d70),
	.w3(32'hb7a88571),
	.w4(32'hb7775dbd),
	.w5(32'hb7b05c96),
	.w6(32'hb78cb587),
	.w7(32'hb7d4cf28),
	.w8(32'hb700eb1d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3786053f),
	.w1(32'h376459ef),
	.w2(32'h37a23816),
	.w3(32'h34402bf4),
	.w4(32'hb60b1da4),
	.w5(32'h36a0149f),
	.w6(32'h34f8f439),
	.w7(32'hb5c00576),
	.w8(32'h36ef6051),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391030f2),
	.w1(32'hb8495549),
	.w2(32'hb8e589d9),
	.w3(32'h390fc871),
	.w4(32'hb7f68016),
	.w5(32'hb887deb9),
	.w6(32'h38087000),
	.w7(32'h381f0f9d),
	.w8(32'h387efd04),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c241d5),
	.w1(32'hb9886845),
	.w2(32'h38366f0e),
	.w3(32'hba0d2ce1),
	.w4(32'hb9ea404e),
	.w5(32'hb6f65c82),
	.w6(32'hba2e1a80),
	.w7(32'hba281b64),
	.w8(32'hb9c6a1ac),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38995f03),
	.w1(32'hb8ab8f86),
	.w2(32'hb90bf7f9),
	.w3(32'h3935b35d),
	.w4(32'h388086e4),
	.w5(32'hb705425f),
	.w6(32'h392a8b39),
	.w7(32'h387e6905),
	.w8(32'hb7d9f9a2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8495c45),
	.w1(32'hb80fcd1e),
	.w2(32'hb70fba72),
	.w3(32'hb820e525),
	.w4(32'hb893ec40),
	.w5(32'hb7c2ac2a),
	.w6(32'hb8389ec6),
	.w7(32'hb8cd16c6),
	.w8(32'hb89b9763),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c2bc0),
	.w1(32'h3954859e),
	.w2(32'h39bd0eef),
	.w3(32'h395553a1),
	.w4(32'h390044b0),
	.w5(32'h3956e88f),
	.w6(32'h38797aab),
	.w7(32'h38950efa),
	.w8(32'h394a166a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39516462),
	.w1(32'h3821d5b3),
	.w2(32'hb8926cd5),
	.w3(32'h391f9d54),
	.w4(32'h3854b52f),
	.w5(32'hb8b3be07),
	.w6(32'h39053cf6),
	.w7(32'hb68683b6),
	.w8(32'hb7bbce54),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398037a7),
	.w1(32'h39041e62),
	.w2(32'hb90b6570),
	.w3(32'h39bb60a2),
	.w4(32'h39317ea7),
	.w5(32'hb8844d96),
	.w6(32'h3a228235),
	.w7(32'h39b68d30),
	.w8(32'h39706768),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b02bf5),
	.w1(32'hb78e74d3),
	.w2(32'hb84b1b19),
	.w3(32'hb72977cd),
	.w4(32'hb747393f),
	.w5(32'hb858da1a),
	.w6(32'hb6b675ad),
	.w7(32'hb5a3df97),
	.w8(32'hb82db855),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357af8c3),
	.w1(32'h35939b9e),
	.w2(32'hb4a28b72),
	.w3(32'hb5cc5c11),
	.w4(32'h340609e5),
	.w5(32'hb40d97a5),
	.w6(32'h3667b71a),
	.w7(32'h34723050),
	.w8(32'h362949e4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af96d0),
	.w1(32'h37947835),
	.w2(32'h371d0a82),
	.w3(32'hb8a71e3c),
	.w4(32'hb82081cb),
	.w5(32'hb702fb54),
	.w6(32'hb977c2f6),
	.w7(32'hb91c52b4),
	.w8(32'hb896feb1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926e735),
	.w1(32'hb92b2a66),
	.w2(32'hb9649a8b),
	.w3(32'h38b59bbb),
	.w4(32'hb8e9f3a5),
	.w5(32'hb8c8161b),
	.w6(32'h38f224f7),
	.w7(32'h38363835),
	.w8(32'h392304b8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b3850),
	.w1(32'h391697de),
	.w2(32'h37a7dbfc),
	.w3(32'h399ffc1b),
	.w4(32'h39702e96),
	.w5(32'h39334b22),
	.w6(32'h3923bb0c),
	.w7(32'h3948cb22),
	.w8(32'h3979e967),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71ad958),
	.w1(32'hb641ea6f),
	.w2(32'h378fb046),
	.w3(32'hb733ac65),
	.w4(32'h369ff525),
	.w5(32'hb6fca8b2),
	.w6(32'h38261cc9),
	.w7(32'h37c44ba6),
	.w8(32'h38a8f593),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d3617),
	.w1(32'h374a0577),
	.w2(32'h3748400d),
	.w3(32'hb60f4ea7),
	.w4(32'h369abef8),
	.w5(32'h37152691),
	.w6(32'h352fda12),
	.w7(32'h36523fa1),
	.w8(32'h378d35a1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63ed7cb),
	.w1(32'h37ea32a6),
	.w2(32'h382f2ae6),
	.w3(32'h36d405bc),
	.w4(32'h381982d7),
	.w5(32'h382d0ad0),
	.w6(32'h37339bef),
	.w7(32'h379c0a48),
	.w8(32'h37be738f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37313c93),
	.w1(32'h3878f02d),
	.w2(32'h38fcec3d),
	.w3(32'h38f89226),
	.w4(32'h38a87bbe),
	.w5(32'h391a1ed2),
	.w6(32'h391aca3f),
	.w7(32'h38e4f3b9),
	.w8(32'h393889e3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec8ec9),
	.w1(32'h39aed73e),
	.w2(32'h38e7e3bc),
	.w3(32'h3a3f54b1),
	.w4(32'h39a9d170),
	.w5(32'hb9368553),
	.w6(32'h3a4e8359),
	.w7(32'h3997098e),
	.w8(32'h397720be),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb814a4c3),
	.w1(32'h3999930e),
	.w2(32'h3a022507),
	.w3(32'hb7ab500f),
	.w4(32'h393574b5),
	.w5(32'h39baa42e),
	.w6(32'hb96fc92e),
	.w7(32'h38292bdc),
	.w8(32'h39992fcb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f62054),
	.w1(32'hb8721625),
	.w2(32'hb88c0803),
	.w3(32'hb9408a51),
	.w4(32'hb8a3b3e6),
	.w5(32'h3702dfcf),
	.w6(32'hb9c8e13e),
	.w7(32'hb9966477),
	.w8(32'hb8aea60d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398255e1),
	.w1(32'h383cd60f),
	.w2(32'hb820c7f5),
	.w3(32'h3931970e),
	.w4(32'h38006083),
	.w5(32'h3703ac56),
	.w6(32'h38e5b7ef),
	.w7(32'hb6768e26),
	.w8(32'h38bf3b25),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36415f35),
	.w1(32'h36a4cf8c),
	.w2(32'h36088ff4),
	.w3(32'h3576c480),
	.w4(32'h361f2c1f),
	.w5(32'h34b2425f),
	.w6(32'h358b7f3e),
	.w7(32'hb47ac33a),
	.w8(32'hb40ce657),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3667041b),
	.w1(32'h36a0cc49),
	.w2(32'h36afec67),
	.w3(32'h359e18ac),
	.w4(32'h362dec3c),
	.w5(32'h366d48e9),
	.w6(32'h3539a926),
	.w7(32'h3584c313),
	.w8(32'h36713088),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371f043c),
	.w1(32'h362992d7),
	.w2(32'hb79f8dc2),
	.w3(32'hb6edd3ad),
	.w4(32'h34a16b52),
	.w5(32'h372dd64f),
	.w6(32'hb630e1ae),
	.w7(32'h36ba22db),
	.w8(32'h37ea2eaf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b554a),
	.w1(32'h36fd54cf),
	.w2(32'h3698489e),
	.w3(32'h3614acdd),
	.w4(32'h361f2a29),
	.w5(32'h3679f93f),
	.w6(32'h3696e46a),
	.w7(32'h368d5dcd),
	.w8(32'hb48df5bb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849ee82),
	.w1(32'hb6f80066),
	.w2(32'hb81d69fb),
	.w3(32'hb85b3f5f),
	.w4(32'hb8462930),
	.w5(32'hb7229d5b),
	.w6(32'hb77825c9),
	.w7(32'hb8141c6b),
	.w8(32'hb7d18aab),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999c9af),
	.w1(32'hb7945c30),
	.w2(32'hb86942cc),
	.w3(32'h38ceb8dd),
	.w4(32'h375d4c29),
	.w5(32'hb770e1cd),
	.w6(32'h388d6ef9),
	.w7(32'h3844e69c),
	.w8(32'h3916750c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961c9a3),
	.w1(32'h391dfa2b),
	.w2(32'h3934fa78),
	.w3(32'h393e81d5),
	.w4(32'h390c898a),
	.w5(32'h38fedadc),
	.w6(32'h38aada22),
	.w7(32'hb7f41cdc),
	.w8(32'h386531e9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6253907),
	.w1(32'h35425acc),
	.w2(32'h36130887),
	.w3(32'hb5a120d3),
	.w4(32'hb6c96df6),
	.w5(32'hb3d53702),
	.w6(32'h364762a7),
	.w7(32'h340d4f00),
	.w8(32'hb61fe27d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c89403),
	.w1(32'h39940fd2),
	.w2(32'h390d9973),
	.w3(32'h39647b4c),
	.w4(32'h39541fe4),
	.w5(32'h38d30bb0),
	.w6(32'h39ae8076),
	.w7(32'h39806a6c),
	.w8(32'h3949783b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd6189),
	.w1(32'hb915fdf5),
	.w2(32'hb91dbb1f),
	.w3(32'hb79fe9bd),
	.w4(32'hb8654e65),
	.w5(32'hb892cdd0),
	.w6(32'hb77ed902),
	.w7(32'h37b0683f),
	.w8(32'h3856974c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3826e9c8),
	.w1(32'hb7b422ae),
	.w2(32'hb8bdb0c8),
	.w3(32'hb816fd45),
	.w4(32'hb8eb61cb),
	.w5(32'hb92a44a0),
	.w6(32'hb890dc10),
	.w7(32'hb90d96a9),
	.w8(32'hb8cee1d2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae77c7),
	.w1(32'hb6316732),
	.w2(32'hb89f9c4d),
	.w3(32'h389b8dc3),
	.w4(32'h389e13eb),
	.w5(32'hb75817aa),
	.w6(32'h39079fec),
	.w7(32'h391cca43),
	.w8(32'h3894923b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73779bd),
	.w1(32'h3650c49c),
	.w2(32'hb66dcf4e),
	.w3(32'h382250d9),
	.w4(32'h388c0ed7),
	.w5(32'h38157f0d),
	.w6(32'h37e90976),
	.w7(32'h3884788e),
	.w8(32'h37cd8b5f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7431b46),
	.w1(32'h38691865),
	.w2(32'h38aec1f4),
	.w3(32'h343e29ea),
	.w4(32'h38a95c15),
	.w5(32'h38ba4e48),
	.w6(32'h3841c0ab),
	.w7(32'h38749cdd),
	.w8(32'h382d5253),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb564039b),
	.w1(32'hb61fbc60),
	.w2(32'h370d02ab),
	.w3(32'hb54ca39b),
	.w4(32'hb645ad50),
	.w5(32'h3735a207),
	.w6(32'hb661f9c5),
	.w7(32'hb6a962f3),
	.w8(32'h3688d8d5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792e39d),
	.w1(32'h3807da4a),
	.w2(32'h37767010),
	.w3(32'h378a74b3),
	.w4(32'h380312c9),
	.w5(32'h375f1db4),
	.w6(32'h36bf94a5),
	.w7(32'h3775da7c),
	.w8(32'hb57c6b73),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394789f3),
	.w1(32'h391bc9df),
	.w2(32'h38eaccce),
	.w3(32'h3941a917),
	.w4(32'h3963b5b2),
	.w5(32'h391bf86f),
	.w6(32'hb82f1e2f),
	.w7(32'h388663e0),
	.w8(32'h390551df),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39544612),
	.w1(32'hb88a8f9b),
	.w2(32'hb942f672),
	.w3(32'h39a9d57b),
	.w4(32'h38518089),
	.w5(32'hb8467b4b),
	.w6(32'h39a256f7),
	.w7(32'h3919bdb0),
	.w8(32'h39301e1f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390effce),
	.w1(32'hb92af2df),
	.w2(32'hb9b50a19),
	.w3(32'h3822996e),
	.w4(32'hb91144f2),
	.w5(32'hb9964a06),
	.w6(32'hb713b7ae),
	.w7(32'hb784d198),
	.w8(32'hb91e2f27),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4a41b),
	.w1(32'h39831d0f),
	.w2(32'h393a2e9f),
	.w3(32'h3996f135),
	.w4(32'h3900c077),
	.w5(32'h38daff84),
	.w6(32'h39b19e2d),
	.w7(32'h39839bb7),
	.w8(32'h39c03272),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ca9b35),
	.w1(32'h373c8cc0),
	.w2(32'hb7b83de9),
	.w3(32'h37982715),
	.w4(32'h36db4647),
	.w5(32'hb7c7ec45),
	.w6(32'hb6e787a1),
	.w7(32'hb749a723),
	.w8(32'hb8165b9e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e532d3),
	.w1(32'hb6d5d54f),
	.w2(32'hb6d0c398),
	.w3(32'hb69082a2),
	.w4(32'hb6ea3dce),
	.w5(32'hb7080358),
	.w6(32'hb7028a69),
	.w7(32'hb7199ab8),
	.w8(32'hb70517ca),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e88c8d),
	.w1(32'hb7ba0a90),
	.w2(32'hb7890270),
	.w3(32'hb71508f3),
	.w4(32'hb792bfcc),
	.w5(32'h3670cb4b),
	.w6(32'h354a7c4c),
	.w7(32'hb5eaf0c3),
	.w8(32'h3702bd71),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36804223),
	.w1(32'h36e10664),
	.w2(32'h365d4beb),
	.w3(32'h36fb4596),
	.w4(32'h36dd158c),
	.w5(32'hb696ddd2),
	.w6(32'hb694641b),
	.w7(32'hb6cea670),
	.w8(32'hb72c98de),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d38f0d),
	.w1(32'h3870ca51),
	.w2(32'h398526a1),
	.w3(32'h36e458ac),
	.w4(32'h39770d95),
	.w5(32'h39a95e1f),
	.w6(32'hb83e9a89),
	.w7(32'h39675268),
	.w8(32'h39a9af46),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86e84e5),
	.w1(32'hb885791d),
	.w2(32'hb816e5b2),
	.w3(32'hb85de275),
	.w4(32'hb7d82e29),
	.w5(32'h3665fba2),
	.w6(32'hb84a1f71),
	.w7(32'hb837796e),
	.w8(32'h36b4528a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88685df),
	.w1(32'hb7f4f31a),
	.w2(32'hb8e6a128),
	.w3(32'hb87cc1da),
	.w4(32'hb880fcff),
	.w5(32'hb9132e31),
	.w6(32'hb80b6264),
	.w7(32'hb88e5bd0),
	.w8(32'hb953b2d5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a39e7f),
	.w1(32'hb7bbc877),
	.w2(32'hb7257987),
	.w3(32'h35a810a1),
	.w4(32'hb81367ef),
	.w5(32'hb82205b1),
	.w6(32'h37a3ae95),
	.w7(32'hb8293d1f),
	.w8(32'hb86f4ac0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8934ce0),
	.w1(32'hb8a5efbb),
	.w2(32'hb882f462),
	.w3(32'hb82b8530),
	.w4(32'hb85465e9),
	.w5(32'hb82a7425),
	.w6(32'hb7579032),
	.w7(32'hb7ca038b),
	.w8(32'hb79cf731),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea1556),
	.w1(32'h38ccd58f),
	.w2(32'h393905d9),
	.w3(32'h38d1039a),
	.w4(32'h38a43b6e),
	.w5(32'h3913c1d7),
	.w6(32'h38bfb044),
	.w7(32'h389f3520),
	.w8(32'h391b5c8e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773d2aa),
	.w1(32'hb6b50708),
	.w2(32'hb6b705a1),
	.w3(32'hb6ecdb53),
	.w4(32'h360c5a83),
	.w5(32'hb59d07f2),
	.w6(32'h368330c0),
	.w7(32'h36ca34f5),
	.w8(32'hb5565759),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af75f8),
	.w1(32'h39c4ba3b),
	.w2(32'h399a1e52),
	.w3(32'h39523c88),
	.w4(32'h390b29fe),
	.w5(32'h389c3ba8),
	.w6(32'h36de57ee),
	.w7(32'hb922f72e),
	.w8(32'hb7979ed1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365a2c75),
	.w1(32'hb68897a2),
	.w2(32'hb68314c2),
	.w3(32'h378e06f4),
	.w4(32'h372749bd),
	.w5(32'h36ef7b80),
	.w6(32'h370596b0),
	.w7(32'h372c197a),
	.w8(32'hb668b7aa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886f789),
	.w1(32'h3913bfc0),
	.w2(32'h3957a652),
	.w3(32'hb90cd48f),
	.w4(32'hb90ac22c),
	.w5(32'h398521ff),
	.w6(32'hb9f11cbe),
	.w7(32'hb9be59ba),
	.w8(32'hb96a8429),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule