module layer_8_featuremap_138(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b06bd),
	.w1(32'hbb9a3a49),
	.w2(32'hbaca58ce),
	.w3(32'h3aac250e),
	.w4(32'hbae9b43b),
	.w5(32'hba4f2dc0),
	.w6(32'h3adec3c4),
	.w7(32'h3a2deddc),
	.w8(32'h3a82aa97),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d30898),
	.w1(32'h3940345b),
	.w2(32'h3a7546db),
	.w3(32'hb9d3f412),
	.w4(32'h3a1d02b2),
	.w5(32'h3a463342),
	.w6(32'hba3b2b6a),
	.w7(32'h38440c0b),
	.w8(32'h39ccd507),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074ec9),
	.w1(32'hbaba8302),
	.w2(32'hba5fb12c),
	.w3(32'hbb1fe332),
	.w4(32'hba8ca5b2),
	.w5(32'hb999cb98),
	.w6(32'hbb42a791),
	.w7(32'hbb0be1ca),
	.w8(32'hba825dcf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cca50),
	.w1(32'hbb664753),
	.w2(32'hb9491e64),
	.w3(32'hbbc81fed),
	.w4(32'hbb4d8711),
	.w5(32'h3a908511),
	.w6(32'hbaddf294),
	.w7(32'hbb816c89),
	.w8(32'h3a998811),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31b139),
	.w1(32'h3b10b780),
	.w2(32'h3ad419ba),
	.w3(32'h3b17ddb6),
	.w4(32'h3b0eaacd),
	.w5(32'h3af3307f),
	.w6(32'h3b16a6bb),
	.w7(32'h3b1f5078),
	.w8(32'h3b3ea5f0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a283),
	.w1(32'h3bd02f3d),
	.w2(32'h3baec013),
	.w3(32'h39b30f09),
	.w4(32'h3aeb4fa4),
	.w5(32'h3b2e9e2d),
	.w6(32'h390ddf1e),
	.w7(32'hba959464),
	.w8(32'h3ae4d0e2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8824511),
	.w1(32'hb83f2779),
	.w2(32'hb8559203),
	.w3(32'hb7b5f062),
	.w4(32'hb6a685c4),
	.w5(32'hb7c0aa6e),
	.w6(32'hb82a7f30),
	.w7(32'hb7b56c5d),
	.w8(32'hb8481980),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba963191),
	.w1(32'hb98c5312),
	.w2(32'h3a4d9fd2),
	.w3(32'hbae79570),
	.w4(32'hbab8959b),
	.w5(32'h388d18eb),
	.w6(32'h39704484),
	.w7(32'h3a50947c),
	.w8(32'h3adffaa3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e93960),
	.w1(32'h3a8d3eec),
	.w2(32'h3a6ab3e1),
	.w3(32'hb9a29736),
	.w4(32'h3944db72),
	.w5(32'h38c94041),
	.w6(32'h3a4ac64c),
	.w7(32'h3a4034e1),
	.w8(32'h3ae30902),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56f821),
	.w1(32'hbb9c02e0),
	.w2(32'hba8029b5),
	.w3(32'hbb517f8a),
	.w4(32'hbb1a6f1f),
	.w5(32'hba22012b),
	.w6(32'hbb289ddb),
	.w7(32'hba8139ea),
	.w8(32'hb98ddf1e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc969),
	.w1(32'hbb47e637),
	.w2(32'h3aabfd8e),
	.w3(32'hb99a3ae7),
	.w4(32'hbb1a8723),
	.w5(32'h3a8bb9b0),
	.w6(32'h3aa5e36a),
	.w7(32'hb8082090),
	.w8(32'h3b037564),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa611a),
	.w1(32'hbb4cdf6c),
	.w2(32'hba8a0724),
	.w3(32'hba65063a),
	.w4(32'hba990991),
	.w5(32'hb9e24300),
	.w6(32'h3af0bd03),
	.w7(32'hba7b30d7),
	.w8(32'hba06f8cc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ddb2),
	.w1(32'h398e1280),
	.w2(32'h3ac6b74a),
	.w3(32'hbaf0f864),
	.w4(32'h39130e58),
	.w5(32'hbac29b96),
	.w6(32'hbb1c9316),
	.w7(32'h3c3e2fbc),
	.w8(32'h3ccbd9d8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054360),
	.w1(32'h3b395eab),
	.w2(32'h39307358),
	.w3(32'hb9dcb59b),
	.w4(32'hba7b2a9c),
	.w5(32'hbaf66c75),
	.w6(32'h3c49b344),
	.w7(32'hbaaef89c),
	.w8(32'hbb16a0d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa88813),
	.w1(32'h3906c1ba),
	.w2(32'hba3c150a),
	.w3(32'h3a0a6b73),
	.w4(32'h3aa32787),
	.w5(32'hb7f4c150),
	.w6(32'hb9ad78ea),
	.w7(32'hba57a045),
	.w8(32'hbafabb00),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeba740),
	.w1(32'hb9e82b78),
	.w2(32'h3b1e2a5a),
	.w3(32'h3b063e11),
	.w4(32'hbbacb6c5),
	.w5(32'hbb625d9d),
	.w6(32'hbaa43d31),
	.w7(32'h3bc1e6fa),
	.w8(32'h3c278564),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93c35f),
	.w1(32'h3ba6bfd9),
	.w2(32'hbb8fd92d),
	.w3(32'hbba576b4),
	.w4(32'h3ab0211d),
	.w5(32'h3b598940),
	.w6(32'h3c20fc1f),
	.w7(32'h3bde6455),
	.w8(32'h3b8a757a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeba331),
	.w1(32'hbc113042),
	.w2(32'h3b305402),
	.w3(32'hbab3d64b),
	.w4(32'hbaedec9c),
	.w5(32'hba63989f),
	.w6(32'h3ab5fff6),
	.w7(32'h3914a223),
	.w8(32'hbb81b318),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e99b3),
	.w1(32'hbc8fdfcd),
	.w2(32'h3ba65c17),
	.w3(32'h3af3adcc),
	.w4(32'hbbb462d3),
	.w5(32'h3c0355c8),
	.w6(32'hbba61989),
	.w7(32'h3a7537a0),
	.w8(32'h3c196933),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c269b1d),
	.w1(32'h3b8b2f57),
	.w2(32'hbaa3544f),
	.w3(32'h3b828201),
	.w4(32'h3b2be103),
	.w5(32'h3bda3408),
	.w6(32'h3c08ddac),
	.w7(32'hbba6c0e0),
	.w8(32'hbc2acad7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6cff),
	.w1(32'hbb82b986),
	.w2(32'h3989fa6f),
	.w3(32'h3b18a34a),
	.w4(32'hbc21b715),
	.w5(32'hba14e210),
	.w6(32'hbbf95a1a),
	.w7(32'hb91153d1),
	.w8(32'h3c22448d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a81cbc),
	.w1(32'hbab9ad87),
	.w2(32'hbb3ee67b),
	.w3(32'hbb6f8def),
	.w4(32'hbb35253d),
	.w5(32'hbb59145a),
	.w6(32'h3c3ebbbc),
	.w7(32'hba432fe5),
	.w8(32'hbb0c2eb8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65472c),
	.w1(32'hbbf207ea),
	.w2(32'hbb7dc629),
	.w3(32'hba36ae4c),
	.w4(32'hbba698f7),
	.w5(32'h3b6dd469),
	.w6(32'hba309d86),
	.w7(32'hb96015af),
	.w8(32'h3b94d911),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8235ac),
	.w1(32'h3b54d002),
	.w2(32'hbb3bfc7f),
	.w3(32'h3a66a851),
	.w4(32'h3b82fd42),
	.w5(32'h3bbbc317),
	.w6(32'h3bb4be94),
	.w7(32'h3b241b78),
	.w8(32'h3ac3ecc0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed5265),
	.w1(32'h3a9b028d),
	.w2(32'hb980b151),
	.w3(32'hb92b2d39),
	.w4(32'hbb3b0e60),
	.w5(32'hbb07f777),
	.w6(32'hb93421d4),
	.w7(32'hbbb69de7),
	.w8(32'hbbd70d91),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50cb91),
	.w1(32'hbb83a09e),
	.w2(32'hbba6d24f),
	.w3(32'h3bd882c6),
	.w4(32'hbc03def4),
	.w5(32'hbbeedb31),
	.w6(32'h3a85861a),
	.w7(32'hbba86201),
	.w8(32'hbc155138),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6c57),
	.w1(32'hbc086201),
	.w2(32'h3bb6c141),
	.w3(32'hbbbfebc1),
	.w4(32'h3ac19e8c),
	.w5(32'hbb017f9f),
	.w6(32'hbc1e1b8b),
	.w7(32'h3b08a6ef),
	.w8(32'h3a381be5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc667c0),
	.w1(32'hbd6be5f6),
	.w2(32'hbd16cc2a),
	.w3(32'h3c0c2d86),
	.w4(32'hbd4ede9d),
	.w5(32'hbd3d65cd),
	.w6(32'h3d69577f),
	.w7(32'h3c624ef9),
	.w8(32'hbc93152a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7858ad),
	.w1(32'hbc03fb2b),
	.w2(32'h3a986470),
	.w3(32'hbc4fca8d),
	.w4(32'h38e32623),
	.w5(32'hbb41b017),
	.w6(32'h3c2090f2),
	.w7(32'hbab9d4f7),
	.w8(32'hbab772b4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f710e),
	.w1(32'h38b8d4a7),
	.w2(32'hbbf8ea22),
	.w3(32'hbb566d20),
	.w4(32'hba9c72e4),
	.w5(32'h3ab7d37c),
	.w6(32'hbafc6023),
	.w7(32'h3ac07bb9),
	.w8(32'h3bc0d054),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9450d6),
	.w1(32'hbbcc0ee1),
	.w2(32'h3a29ccc2),
	.w3(32'hb85bcbb8),
	.w4(32'h3b96e05e),
	.w5(32'h3b366f90),
	.w6(32'h3c1e4b81),
	.w7(32'h3ab014b4),
	.w8(32'h3aa097f4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a8d59),
	.w1(32'h3723d306),
	.w2(32'hbbba62fc),
	.w3(32'h3b8d1bf3),
	.w4(32'hbc0ac89d),
	.w5(32'hbb93673b),
	.w6(32'hb9a58a82),
	.w7(32'hbba57fb8),
	.w8(32'h3c412144),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc66499),
	.w1(32'hbbd40031),
	.w2(32'hbb8616ee),
	.w3(32'hbc1f6442),
	.w4(32'h3be4871c),
	.w5(32'h3c9b483f),
	.w6(32'h3b1432fc),
	.w7(32'hbc8d9bc5),
	.w8(32'h3a81f4cc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a19f),
	.w1(32'h3b42a4c6),
	.w2(32'h3ad699c8),
	.w3(32'h384cc360),
	.w4(32'hbb7e29d3),
	.w5(32'hbbc74adc),
	.w6(32'hbc32479c),
	.w7(32'h3b03309f),
	.w8(32'hbbdcfa4f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be72567),
	.w1(32'h3b56fb64),
	.w2(32'h3b397c02),
	.w3(32'h369ac224),
	.w4(32'h3bb7d12a),
	.w5(32'h3b947850),
	.w6(32'hbbd7b009),
	.w7(32'hba33c8c5),
	.w8(32'h3ae32cd0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03bc22),
	.w1(32'hbbdf5251),
	.w2(32'hbc0f86a8),
	.w3(32'h3b4c6470),
	.w4(32'hbb1e0481),
	.w5(32'hbae425c7),
	.w6(32'h3b104ef7),
	.w7(32'hbbf836fc),
	.w8(32'hbbb4f3f5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae3cb0),
	.w1(32'hbaf7eb15),
	.w2(32'hbc35af62),
	.w3(32'hbb4e7c00),
	.w4(32'hbbbaf6f0),
	.w5(32'hba82eb40),
	.w6(32'hbbc3381a),
	.w7(32'hbc69f592),
	.w8(32'hba853c8d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f37c8),
	.w1(32'hbbf3402a),
	.w2(32'hbaea8f31),
	.w3(32'hbb6cffdc),
	.w4(32'hbb2b6afd),
	.w5(32'hbb2ca666),
	.w6(32'hbc76b18c),
	.w7(32'hbb48dbb1),
	.w8(32'hbb9a4142),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4a14),
	.w1(32'hbadc4bf0),
	.w2(32'hbb0177a1),
	.w3(32'hb90be792),
	.w4(32'h3a24e3ed),
	.w5(32'hba6f55dc),
	.w6(32'hbabc6bd6),
	.w7(32'h3c2611ce),
	.w8(32'h3c4764c1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390942dd),
	.w1(32'hbb55c5fc),
	.w2(32'h3ab161bb),
	.w3(32'hba5ae498),
	.w4(32'h3c20931c),
	.w5(32'h3c12773d),
	.w6(32'h3c10e89f),
	.w7(32'h3caab9e7),
	.w8(32'h3d0191b5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0bb27),
	.w1(32'h3c3b5535),
	.w2(32'h3b58173c),
	.w3(32'h3aa380c6),
	.w4(32'hbc2b82d1),
	.w5(32'hbb5e9417),
	.w6(32'h3cf79b92),
	.w7(32'hbba00766),
	.w8(32'hbb691c0a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181201),
	.w1(32'hb9c69433),
	.w2(32'hbbc0c99b),
	.w3(32'hbbd09581),
	.w4(32'hbbc8da7f),
	.w5(32'hbc369471),
	.w6(32'h3b684f60),
	.w7(32'hbbb004be),
	.w8(32'hbadf24fe),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd921c7),
	.w1(32'hba3b5724),
	.w2(32'hbae3b14f),
	.w3(32'hbbd57ec8),
	.w4(32'h3bb2eed3),
	.w5(32'h3c37581f),
	.w6(32'h3bc4cf3e),
	.w7(32'h3c8eb2ee),
	.w8(32'h3ced7cd9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ec82b),
	.w1(32'h3b27f7f0),
	.w2(32'hba349502),
	.w3(32'h3bc76a69),
	.w4(32'hb9aa38f8),
	.w5(32'hbbef5d93),
	.w6(32'h3caad587),
	.w7(32'h3bccecfd),
	.w8(32'h3c73c44c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c343927),
	.w1(32'h39daf918),
	.w2(32'hba6fbf1c),
	.w3(32'hbb0d2360),
	.w4(32'hbb2a67dc),
	.w5(32'h3b313c8c),
	.w6(32'h3bdb12d3),
	.w7(32'h39c50213),
	.w8(32'h3ac34e21),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc691c44),
	.w1(32'hbc1def1d),
	.w2(32'hbb844aa1),
	.w3(32'hbade9cda),
	.w4(32'hbafca752),
	.w5(32'hbb506e8f),
	.w6(32'hbb30c554),
	.w7(32'h3badc20c),
	.w8(32'h3c45570e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64800),
	.w1(32'h3c023c05),
	.w2(32'hbc413b3a),
	.w3(32'hbbee0341),
	.w4(32'h3a03412f),
	.w5(32'hbb621f01),
	.w6(32'h3b9a0476),
	.w7(32'h3bdcfb76),
	.w8(32'h3bfaf146),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfba671),
	.w1(32'hbbce625b),
	.w2(32'hba5742a8),
	.w3(32'hbb924b90),
	.w4(32'hbb8b3375),
	.w5(32'h3baf02ec),
	.w6(32'h3baa10e5),
	.w7(32'hbbebf71d),
	.w8(32'hba99e54a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c9c0b),
	.w1(32'hbb20c37d),
	.w2(32'hbb97a599),
	.w3(32'hba85c218),
	.w4(32'hbb409a95),
	.w5(32'hbb60acbb),
	.w6(32'hba0b5b4c),
	.w7(32'h39b16fd9),
	.w8(32'h3b242fd2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037b7a),
	.w1(32'hbb9e9fa2),
	.w2(32'hbb12af34),
	.w3(32'hbc024537),
	.w4(32'hbc0334d5),
	.w5(32'hbc005bca),
	.w6(32'h3aaf5772),
	.w7(32'h3992b055),
	.w8(32'h3b4411fb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1401),
	.w1(32'hb9f4bbb6),
	.w2(32'hbb702ebb),
	.w3(32'hbc80be17),
	.w4(32'hbc3f4b8f),
	.w5(32'hbc5c39e2),
	.w6(32'hbbde96ab),
	.w7(32'hbc6c35a9),
	.w8(32'hbc1ca2e7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a4ee),
	.w1(32'hbbe7e128),
	.w2(32'h3a5c70cb),
	.w3(32'hbc5a68c7),
	.w4(32'hbbaf8998),
	.w5(32'hbb8e44d9),
	.w6(32'hbad4b1eb),
	.w7(32'hb918d5bb),
	.w8(32'h39c787d0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d42b2),
	.w1(32'hbc09f84b),
	.w2(32'h3b657c6a),
	.w3(32'h3b3cef0f),
	.w4(32'hbad865b0),
	.w5(32'hba24ccfc),
	.w6(32'h3b2b91f9),
	.w7(32'h3ad9ea74),
	.w8(32'h3b8e5d02),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b5a75),
	.w1(32'hbbaba3c7),
	.w2(32'hbb20926c),
	.w3(32'h3a8b438a),
	.w4(32'h3b07e9d3),
	.w5(32'hbb6225ee),
	.w6(32'hba13ed22),
	.w7(32'h3ba21d28),
	.w8(32'h3b9efd7c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b998053),
	.w1(32'h3b2f8aa0),
	.w2(32'hba2b45be),
	.w3(32'hbac1ce0c),
	.w4(32'hbae2fbff),
	.w5(32'hbacb82a5),
	.w6(32'h3a8c5fda),
	.w7(32'hbbd7515c),
	.w8(32'hbba39243),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ea90e),
	.w1(32'hbbaffc7f),
	.w2(32'hba3d184e),
	.w3(32'hbbbff44e),
	.w4(32'hbb3f2cf8),
	.w5(32'h3b642255),
	.w6(32'hbb94e894),
	.w7(32'h3a76aa4e),
	.w8(32'h3b8828c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae3328),
	.w1(32'h3b27d4d6),
	.w2(32'h3c382786),
	.w3(32'hbbac2dd5),
	.w4(32'h3bfb3ed2),
	.w5(32'h3be8c659),
	.w6(32'h3ab135b6),
	.w7(32'h3c918499),
	.w8(32'h3cbb850e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be193a5),
	.w1(32'h3b3e9457),
	.w2(32'hbc0668ba),
	.w3(32'h3c2ba83c),
	.w4(32'hbc719f8d),
	.w5(32'hbc17ec14),
	.w6(32'h3cbfe4d8),
	.w7(32'h3c237114),
	.w8(32'h3c1e5654),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39da62),
	.w1(32'hbbc1eb84),
	.w2(32'hb9db5446),
	.w3(32'h3b09d9cb),
	.w4(32'hbae09984),
	.w5(32'hbbbccf76),
	.w6(32'h3c710081),
	.w7(32'h3b7a280e),
	.w8(32'h3c1b4e2f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9a0be),
	.w1(32'h3b264dec),
	.w2(32'h3aede2dd),
	.w3(32'hbb5bd4cc),
	.w4(32'hbba2e219),
	.w5(32'hbc17bdcc),
	.w6(32'hba039b82),
	.w7(32'h3b341b62),
	.w8(32'h3bfb4734),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6e476),
	.w1(32'h3b93b3ae),
	.w2(32'h3aad41db),
	.w3(32'hbb355627),
	.w4(32'hbba726d5),
	.w5(32'hbc5f7a77),
	.w6(32'h3bb1f469),
	.w7(32'h3c67a657),
	.w8(32'h3bdcf07b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fb921),
	.w1(32'h3b8c951f),
	.w2(32'hba716df1),
	.w3(32'hbc0739a8),
	.w4(32'h3a123b07),
	.w5(32'hbaf3b775),
	.w6(32'h3c449594),
	.w7(32'hbbf9c45d),
	.w8(32'hbc2b28ba),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8845fa),
	.w1(32'hbb37cce3),
	.w2(32'h3bd20223),
	.w3(32'hbafb8879),
	.w4(32'hbbf084cc),
	.w5(32'hbb59af5d),
	.w6(32'hbbe26da3),
	.w7(32'hbb2ba898),
	.w8(32'hbb5641d8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3d0a),
	.w1(32'h3acdcf79),
	.w2(32'hbb093ad4),
	.w3(32'hb98d649c),
	.w4(32'hbb82c60c),
	.w5(32'h3bda6f34),
	.w6(32'hbb3c3a63),
	.w7(32'h3c8097f4),
	.w8(32'h3d1c44e5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e21a1),
	.w1(32'hba0a7351),
	.w2(32'h3bc553ff),
	.w3(32'h3a754420),
	.w4(32'hba43e8f5),
	.w5(32'hbb32de39),
	.w6(32'h3cd4204d),
	.w7(32'h3ac12e6f),
	.w8(32'h3bfbaf50),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd47e80),
	.w1(32'h3c336b69),
	.w2(32'h3a7c7f3d),
	.w3(32'hba8beb23),
	.w4(32'hb9214903),
	.w5(32'hb8e03898),
	.w6(32'h3c1b864f),
	.w7(32'hbbe4b40f),
	.w8(32'hbbe9f2a6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27fe0),
	.w1(32'h3b8819f1),
	.w2(32'h3b705ef4),
	.w3(32'h3b275dfd),
	.w4(32'hbada79a0),
	.w5(32'hbab5303f),
	.w6(32'hbb69e437),
	.w7(32'h3bcf4558),
	.w8(32'h3becff93),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72a228),
	.w1(32'hbb58d317),
	.w2(32'hbb737091),
	.w3(32'h39bee1ae),
	.w4(32'h3a9f261c),
	.w5(32'h3b790178),
	.w6(32'h3b9a23ac),
	.w7(32'hbbb16c6c),
	.w8(32'h3b9018e0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5355),
	.w1(32'hbc0ce4a6),
	.w2(32'hba03a218),
	.w3(32'hbba4f3bb),
	.w4(32'hbbd238ce),
	.w5(32'hbc212cea),
	.w6(32'hbc436b70),
	.w7(32'hbbb7d86a),
	.w8(32'hbb9008bc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b959e),
	.w1(32'h3b0bd2ad),
	.w2(32'h3b0fc879),
	.w3(32'hbb7a93d8),
	.w4(32'hbb194282),
	.w5(32'h3b4832f7),
	.w6(32'h3a8aa467),
	.w7(32'h3a089827),
	.w8(32'h3bc5f5f0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64f796),
	.w1(32'hbbc6cc99),
	.w2(32'h3b285d5e),
	.w3(32'h3b0bcf8c),
	.w4(32'h3a0f3697),
	.w5(32'hbb46225e),
	.w6(32'h3a6224bb),
	.w7(32'h3a8ee95a),
	.w8(32'h3b3ade39),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5532cb),
	.w1(32'h3b295826),
	.w2(32'hbba77174),
	.w3(32'h3af82ca5),
	.w4(32'hbb24c510),
	.w5(32'hbac233c5),
	.w6(32'h3bc355f6),
	.w7(32'h3a28470f),
	.w8(32'h39a20609),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7384),
	.w1(32'hbaa7ad5b),
	.w2(32'hbba06246),
	.w3(32'h3afc2d53),
	.w4(32'h3a40c942),
	.w5(32'h3abf841f),
	.w6(32'hbb04fbda),
	.w7(32'hbc774c23),
	.w8(32'hbc2cbd98),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b3da),
	.w1(32'hbb81ff41),
	.w2(32'hbb2e737f),
	.w3(32'hbb8f8198),
	.w4(32'hbad729a1),
	.w5(32'h3bb0e649),
	.w6(32'hbc50e44d),
	.w7(32'h3c017825),
	.w8(32'h3c88f4ea),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7dcf),
	.w1(32'hbc343d73),
	.w2(32'hbbb8438e),
	.w3(32'hba7a9d1d),
	.w4(32'h3ab3d3c1),
	.w5(32'hb80f0364),
	.w6(32'h3c1701a2),
	.w7(32'hbb31961e),
	.w8(32'hbac03029),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d977),
	.w1(32'h3b1193fc),
	.w2(32'h3af39537),
	.w3(32'hbae79cf0),
	.w4(32'h3b3a5d34),
	.w5(32'h3b23acbc),
	.w6(32'h3acd73e0),
	.w7(32'h3b820648),
	.w8(32'h3add5817),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6488b2),
	.w1(32'h3b2d74fe),
	.w2(32'hb8b15736),
	.w3(32'hbafd5ede),
	.w4(32'hb902229d),
	.w5(32'hbbeeeb56),
	.w6(32'h3b37deb2),
	.w7(32'hbb9a1a2c),
	.w8(32'h3a6f88db),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf249bc),
	.w1(32'hba911fe0),
	.w2(32'hbbfb9416),
	.w3(32'h3b45deba),
	.w4(32'hb9e36f86),
	.w5(32'hbb43de89),
	.w6(32'h3c3d7150),
	.w7(32'hbb3349f0),
	.w8(32'h39d5228a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006ac4),
	.w1(32'hbbc048dc),
	.w2(32'hba64f6c0),
	.w3(32'hbb43a39f),
	.w4(32'hbaf1d900),
	.w5(32'h3b1b8a25),
	.w6(32'h3b25fd66),
	.w7(32'h398824a4),
	.w8(32'h3b4c6c8c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8614e2),
	.w1(32'hbb063674),
	.w2(32'hba3e4a85),
	.w3(32'hb9d6829e),
	.w4(32'h3c883790),
	.w5(32'h3c95f8bb),
	.w6(32'h3a98bdcb),
	.w7(32'hbc3bcfb7),
	.w8(32'hbc09684e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3f35),
	.w1(32'hbc880a79),
	.w2(32'hb9cbc6d5),
	.w3(32'h3afd623f),
	.w4(32'hbb9be983),
	.w5(32'h3b223dea),
	.w6(32'hbbd14a14),
	.w7(32'h3b0d0038),
	.w8(32'h3b73ac01),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc50a1),
	.w1(32'hbc00451b),
	.w2(32'h3bf14b8d),
	.w3(32'h3bdeccfa),
	.w4(32'hbb5f7781),
	.w5(32'hbc5d0918),
	.w6(32'hbab46421),
	.w7(32'hbb5e7452),
	.w8(32'h3b3d591c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa44d2),
	.w1(32'h3c7ad4a7),
	.w2(32'h3a02eb2d),
	.w3(32'h3af1067e),
	.w4(32'h3b813721),
	.w5(32'h3c97e392),
	.w6(32'hbb9015b2),
	.w7(32'hbb8b0480),
	.w8(32'hbcdaa039),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b93d9),
	.w1(32'h3b855ec8),
	.w2(32'hbc62498d),
	.w3(32'hbbb9bbee),
	.w4(32'hbc129432),
	.w5(32'hbc97a978),
	.w6(32'hbc1acb82),
	.w7(32'hbb51f0eb),
	.w8(32'h3d08226b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be73c12),
	.w1(32'hbc5e9efa),
	.w2(32'hba56be79),
	.w3(32'h3b314a90),
	.w4(32'h3c8691c7),
	.w5(32'h3c1e52a2),
	.w6(32'h3d003e70),
	.w7(32'hbd186424),
	.w8(32'hba7b6c7b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2a28),
	.w1(32'hbba8668b),
	.w2(32'hba993616),
	.w3(32'h3c21d711),
	.w4(32'h3b439219),
	.w5(32'h398856dc),
	.w6(32'h3cee1e13),
	.w7(32'h3b09a0fe),
	.w8(32'hbc85ce10),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94e289),
	.w1(32'h3ac8ab80),
	.w2(32'hbb8af1bc),
	.w3(32'h3aa039a3),
	.w4(32'h3a9454c2),
	.w5(32'hbb4bca84),
	.w6(32'hbb0a55e8),
	.w7(32'h3c35d0a7),
	.w8(32'h3c41429c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc263e25),
	.w1(32'hbc7b15ed),
	.w2(32'h3959b35c),
	.w3(32'hbc50ae31),
	.w4(32'hbc048366),
	.w5(32'h3b5f0c3c),
	.w6(32'hbc9eab6f),
	.w7(32'hbb46c05b),
	.w8(32'h3b947918),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6370c5),
	.w1(32'h3bc0abe9),
	.w2(32'hbbf25948),
	.w3(32'h3aaaedb8),
	.w4(32'h3c24fe97),
	.w5(32'h3b85f8b5),
	.w6(32'hba696b04),
	.w7(32'hbb661218),
	.w8(32'h3b8ef7b1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f37b5),
	.w1(32'h3b9a8bb6),
	.w2(32'hbc25905c),
	.w3(32'hbb87fda5),
	.w4(32'h3c9859f8),
	.w5(32'h3c923f65),
	.w6(32'hbbcf942e),
	.w7(32'h3bb68673),
	.w8(32'hbc503a6e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd079033),
	.w1(32'hbbe98561),
	.w2(32'hbbaa71de),
	.w3(32'hbc433c6a),
	.w4(32'hbc7d3521),
	.w5(32'hbc8cb24d),
	.w6(32'hbcc4f88f),
	.w7(32'hbb92129d),
	.w8(32'h3a1facfa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badd795),
	.w1(32'h3c60e866),
	.w2(32'hbcce5c51),
	.w3(32'h3ac9af63),
	.w4(32'hba31ef5f),
	.w5(32'h3d04e178),
	.w6(32'h3b21371e),
	.w7(32'h3ce9cca4),
	.w8(32'h3d88f80e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4e44ac),
	.w1(32'hbd490d9f),
	.w2(32'h3c141351),
	.w3(32'h3b515d7b),
	.w4(32'h3bf4383a),
	.w5(32'h3c043f90),
	.w6(32'hbb60b0c0),
	.w7(32'hbc04e8df),
	.w8(32'hbcde3011),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd6e3d),
	.w1(32'h3b935518),
	.w2(32'h3bebe4fc),
	.w3(32'h3c0525c2),
	.w4(32'hbc591501),
	.w5(32'hbc76e146),
	.w6(32'hbc616696),
	.w7(32'h3bba7bd1),
	.w8(32'h3d552bec),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a708),
	.w1(32'hbc7cefb8),
	.w2(32'h3a1737a4),
	.w3(32'h3a8cb70c),
	.w4(32'h3ace4020),
	.w5(32'h3bb35bf3),
	.w6(32'h3cdb7a92),
	.w7(32'h3b7c3ce2),
	.w8(32'h3bc0fddb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914cd8),
	.w1(32'hbb8ac80d),
	.w2(32'hbc05bc86),
	.w3(32'h3b0afb31),
	.w4(32'h3b04b100),
	.w5(32'hbc2edbbb),
	.w6(32'h3b1d056b),
	.w7(32'hbcbb7ec8),
	.w8(32'h3c86503d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05e95c),
	.w1(32'hbcb4b415),
	.w2(32'h3cbfed0b),
	.w3(32'hbc215ff8),
	.w4(32'hbd235d4c),
	.w5(32'hbd31c713),
	.w6(32'h3c269997),
	.w7(32'hba3d4f8a),
	.w8(32'h3c9d1552),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2fece3),
	.w1(32'h3c313bb5),
	.w2(32'hbc0834d0),
	.w3(32'hbb72d080),
	.w4(32'h3c5f29d2),
	.w5(32'h3ad2d2cc),
	.w6(32'h3c959e6f),
	.w7(32'hbbd65f70),
	.w8(32'hbd087f0f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c836d),
	.w1(32'h3c240f7e),
	.w2(32'h3bd93bf9),
	.w3(32'h3bd0b9b8),
	.w4(32'h3b3c1bfe),
	.w5(32'hb9a3d0bd),
	.w6(32'hbcd17017),
	.w7(32'h3ba057eb),
	.w8(32'h3b0a60a7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad94d7e),
	.w1(32'h3b918b9a),
	.w2(32'h3cb0a2ce),
	.w3(32'h3b9069ec),
	.w4(32'hbccfb510),
	.w5(32'hbcbd4d80),
	.w6(32'h3c00c778),
	.w7(32'h3ca429d7),
	.w8(32'hbbc485bb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2165c),
	.w1(32'h3cac8c71),
	.w2(32'hbc9d1ca3),
	.w3(32'hbc37a648),
	.w4(32'hbbb47c11),
	.w5(32'hbba512ec),
	.w6(32'hbc9cf67f),
	.w7(32'hbc8d5424),
	.w8(32'hbb7835a5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96b3d5),
	.w1(32'h3c2b5cf0),
	.w2(32'h3b3b2e17),
	.w3(32'hbc1cbf20),
	.w4(32'h3ca09b98),
	.w5(32'h3bef554b),
	.w6(32'h3bd4c933),
	.w7(32'hbc720362),
	.w8(32'hbc8d3961),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e470),
	.w1(32'hb9297cf9),
	.w2(32'hbaf83f3d),
	.w3(32'h3b5e9a3b),
	.w4(32'h3b1c3717),
	.w5(32'h3cabedc8),
	.w6(32'h3b1dc362),
	.w7(32'hbb1bf2b5),
	.w8(32'hbd125209),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03fac),
	.w1(32'h3c826a86),
	.w2(32'hbbd19fe6),
	.w3(32'h3bfa3d14),
	.w4(32'h3b6378dd),
	.w5(32'hbadd2b5a),
	.w6(32'hbc2e250e),
	.w7(32'hbbff643c),
	.w8(32'hbb62dd7d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9e063),
	.w1(32'hbbfe07ec),
	.w2(32'hbbd1811f),
	.w3(32'hbc117f14),
	.w4(32'h3c7ae128),
	.w5(32'hb8b51173),
	.w6(32'hbc4c197c),
	.w7(32'hbb6ad30c),
	.w8(32'h3c069422),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5794ec),
	.w1(32'hbab78289),
	.w2(32'hba7c92f4),
	.w3(32'h3b93a9d0),
	.w4(32'hbbf3d5a8),
	.w5(32'hb9cc68ad),
	.w6(32'hbb8786f5),
	.w7(32'h3ca4013e),
	.w8(32'h3d4e226e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5154bf),
	.w1(32'hbc9c3085),
	.w2(32'h3bff44b9),
	.w3(32'hbbebc579),
	.w4(32'hbc1c7307),
	.w5(32'hbc8fc3a7),
	.w6(32'hbbecbf31),
	.w7(32'hbc682f66),
	.w8(32'hbc4576f9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7984d1),
	.w1(32'h3d161b4e),
	.w2(32'h3ab2aef3),
	.w3(32'hbae0d1d5),
	.w4(32'hbab2bd7d),
	.w5(32'hbbfd6a31),
	.w6(32'h3c153e65),
	.w7(32'hba67de59),
	.w8(32'hba18ef2c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0263a6),
	.w1(32'h3b95dc6d),
	.w2(32'h3c66fef0),
	.w3(32'hba92c869),
	.w4(32'h3a9a334c),
	.w5(32'h3c9568c2),
	.w6(32'h3bfbb076),
	.w7(32'h3cd29914),
	.w8(32'hbba44cb8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29432a),
	.w1(32'hba3d5bd6),
	.w2(32'h3c9b4c8a),
	.w3(32'h3b036fa1),
	.w4(32'hbc9ed73b),
	.w5(32'hbba75f92),
	.w6(32'hbc81534a),
	.w7(32'h3ac3d4df),
	.w8(32'h3b9327fc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae8473),
	.w1(32'h3ce0aa67),
	.w2(32'h3c2614ea),
	.w3(32'h3b2b3bfd),
	.w4(32'hbb0c0f6d),
	.w5(32'h3ba6f0bd),
	.w6(32'hbc4de539),
	.w7(32'h3b40966b),
	.w8(32'h3b7815e4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a16ac),
	.w1(32'h3b7f2745),
	.w2(32'h3b76755d),
	.w3(32'h3ab4ee68),
	.w4(32'h3c00c84e),
	.w5(32'h3acc3466),
	.w6(32'h3b4f88ee),
	.w7(32'hbca60afa),
	.w8(32'hbbf83b74),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11fe0b),
	.w1(32'h3c49b6a0),
	.w2(32'hbc0ec49e),
	.w3(32'h3b4be0a0),
	.w4(32'hbc24fba0),
	.w5(32'hbc28954d),
	.w6(32'h3c1d9be1),
	.w7(32'h3b7d2f61),
	.w8(32'h3d672d10),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc886fc6),
	.w1(32'h3c495479),
	.w2(32'hbc9f2bac),
	.w3(32'hbb683a0c),
	.w4(32'hbc91e6e5),
	.w5(32'hbc0a5d73),
	.w6(32'h3b5a481d),
	.w7(32'hbcbdbaa3),
	.w8(32'hbc9e45b0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9054),
	.w1(32'h3b8ddae0),
	.w2(32'hbc8b6c31),
	.w3(32'hbcd0abee),
	.w4(32'h3c3e611a),
	.w5(32'h3c3d87ab),
	.w6(32'hbcb591e7),
	.w7(32'h3bbe27ad),
	.w8(32'h3bf1b2f0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4d3e5),
	.w1(32'hbc1aac27),
	.w2(32'hbcd8d933),
	.w3(32'h3aacead1),
	.w4(32'h3ce90ce4),
	.w5(32'h3c62db50),
	.w6(32'hbb86e832),
	.w7(32'hbc525133),
	.w8(32'h3c2c6084),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3bc18),
	.w1(32'hbc85ec7e),
	.w2(32'hbbcc9610),
	.w3(32'h3c3cd300),
	.w4(32'h3c82b250),
	.w5(32'h391ff2de),
	.w6(32'h3cf925c5),
	.w7(32'h3bb32f76),
	.w8(32'hbbe71f8b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4dca3),
	.w1(32'hbc853b3c),
	.w2(32'hbb4fd4ef),
	.w3(32'h3b4e8a9b),
	.w4(32'hbbace036),
	.w5(32'hbba7cff6),
	.w6(32'hbc509623),
	.w7(32'hb947aa3a),
	.w8(32'h3a9a0c3a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22e35b),
	.w1(32'hbad9f85a),
	.w2(32'h3afc2c8a),
	.w3(32'hbb663efc),
	.w4(32'hbb94cd3a),
	.w5(32'hbc4ab1b1),
	.w6(32'h3b832bc9),
	.w7(32'h3b68e40f),
	.w8(32'h3bb9ee33),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2343),
	.w1(32'hbb13357a),
	.w2(32'h3bea0aed),
	.w3(32'hbc0768f2),
	.w4(32'h3b958580),
	.w5(32'h3bbfcd31),
	.w6(32'h3c4d8d2e),
	.w7(32'hba953734),
	.w8(32'hbcdca04b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c603bd3),
	.w1(32'h3c906a25),
	.w2(32'hbbf8d54c),
	.w3(32'h3c24ef7c),
	.w4(32'hbcaa4e31),
	.w5(32'hbc4171cf),
	.w6(32'hbb939069),
	.w7(32'hbc9750b4),
	.w8(32'h3c9a391c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3300ac),
	.w1(32'h3a8412d0),
	.w2(32'hbbe90853),
	.w3(32'hbb774bf2),
	.w4(32'h3b2fe098),
	.w5(32'h3cd62917),
	.w6(32'h3bd5ef30),
	.w7(32'h3d33b0bf),
	.w8(32'h3cc932a9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2a013a),
	.w1(32'hbcae9f26),
	.w2(32'hb9152f64),
	.w3(32'h3c4546e2),
	.w4(32'hb9d895b8),
	.w5(32'hbbaf393e),
	.w6(32'h3be3ca4b),
	.w7(32'h3b3241ce),
	.w8(32'h3a5b57f9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b093c),
	.w1(32'hba114b6f),
	.w2(32'hbaf6d5fc),
	.w3(32'hbb4c26ec),
	.w4(32'h3c6177c1),
	.w5(32'h3d001060),
	.w6(32'h3b8d1c05),
	.w7(32'hbcd6b2b9),
	.w8(32'hbdc4f490),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16d27b),
	.w1(32'h3cd16a5b),
	.w2(32'hba70d08a),
	.w3(32'h3c05fbf7),
	.w4(32'h3cb97c94),
	.w5(32'h3bcb7679),
	.w6(32'hbd2e0e7a),
	.w7(32'h38be8338),
	.w8(32'hbd27d173),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84942f0),
	.w1(32'hbc8bd136),
	.w2(32'hbad07b63),
	.w3(32'h3aa36a38),
	.w4(32'h3b02dedf),
	.w5(32'h3bf2fb9b),
	.w6(32'hbcf4a103),
	.w7(32'hbabb0314),
	.w8(32'hbb1cc75a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad12b97),
	.w1(32'hbbe112a8),
	.w2(32'h39ce202e),
	.w3(32'hba908ada),
	.w4(32'h3c3fdd2e),
	.w5(32'hbc0d0363),
	.w6(32'hbb9f36ae),
	.w7(32'hbc1c8b16),
	.w8(32'hbce34fb0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bcba5),
	.w1(32'hbab3f075),
	.w2(32'hbca89c02),
	.w3(32'h3b1084ba),
	.w4(32'hbc032a4c),
	.w5(32'hbc114d91),
	.w6(32'h3ca36ed2),
	.w7(32'hbba6e1ae),
	.w8(32'h3b74caa4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule