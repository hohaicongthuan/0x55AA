module layer_10_featuremap_509(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc116eae),
	.w1(32'h3cc3a026),
	.w2(32'hbb1712ba),
	.w3(32'h3c440b02),
	.w4(32'hbcb92bfd),
	.w5(32'h3c6c4016),
	.w6(32'h3b121924),
	.w7(32'hbc105094),
	.w8(32'hbb24a945),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6c46d),
	.w1(32'h3c2adb0c),
	.w2(32'h3c064a31),
	.w3(32'h3bc623e6),
	.w4(32'h3ce69d0a),
	.w5(32'hbc2c0342),
	.w6(32'hbccb68d5),
	.w7(32'hbc1cde8f),
	.w8(32'h399c3136),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696a12),
	.w1(32'hba9325eb),
	.w2(32'hbb4696d8),
	.w3(32'hb952e77c),
	.w4(32'h3c3ff069),
	.w5(32'hbd181e88),
	.w6(32'h3c3f0de1),
	.w7(32'hbc1aa454),
	.w8(32'hbc44ef8d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e67952),
	.w1(32'hbb5b82d6),
	.w2(32'h3b8b7027),
	.w3(32'h3b81d2f3),
	.w4(32'hbc597858),
	.w5(32'hbc9c9635),
	.w6(32'hbbb5f92c),
	.w7(32'h3bb0b27c),
	.w8(32'hbb6c2edf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1200ea),
	.w1(32'hbb5472da),
	.w2(32'h3c015366),
	.w3(32'hbb46e5c2),
	.w4(32'h3ba58fe3),
	.w5(32'h3746612f),
	.w6(32'h3c0e325d),
	.w7(32'hbb9da37b),
	.w8(32'h3b2fe780),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3fea9),
	.w1(32'h39ef2ea7),
	.w2(32'h3caee871),
	.w3(32'h3b8ea2ab),
	.w4(32'hbc1b3a20),
	.w5(32'hbb9634b1),
	.w6(32'hbae64f7f),
	.w7(32'hbbbac7e5),
	.w8(32'h3bbc7416),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c403d35),
	.w1(32'hbc28f41a),
	.w2(32'hbb840593),
	.w3(32'h3c17cb78),
	.w4(32'hbc2ab86d),
	.w5(32'hbc078688),
	.w6(32'h3b5e881d),
	.w7(32'hbd5923ec),
	.w8(32'hbc97178d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00a52c),
	.w1(32'hbcc1a9c7),
	.w2(32'hbba4f101),
	.w3(32'h3b8e02ee),
	.w4(32'hbcf2b603),
	.w5(32'hba3ad839),
	.w6(32'h3c1ae88c),
	.w7(32'hbc1940f3),
	.w8(32'h3bd0ed42),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91463e0),
	.w1(32'hbaa67e2a),
	.w2(32'hba076af5),
	.w3(32'hbcbb236f),
	.w4(32'h3c1a04f0),
	.w5(32'hbbf4d696),
	.w6(32'hbbdebd6a),
	.w7(32'hbbdb1a6c),
	.w8(32'hbb4b58a5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2775be),
	.w1(32'hbc4c6f46),
	.w2(32'hbbe15b44),
	.w3(32'hbb8eace5),
	.w4(32'hbca031fa),
	.w5(32'h3c92f641),
	.w6(32'h3b5178cb),
	.w7(32'h3af0ebbe),
	.w8(32'h3a8b82a0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc950e14),
	.w1(32'hba654cf6),
	.w2(32'hb78152f0),
	.w3(32'h3bcd6722),
	.w4(32'h3aa118bc),
	.w5(32'hbbaef7ea),
	.w6(32'h3914a3f1),
	.w7(32'h3bf90f37),
	.w8(32'h3b2f00af),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dcc38),
	.w1(32'hba942cce),
	.w2(32'h3bcee670),
	.w3(32'hbc30fb94),
	.w4(32'h3c236cb5),
	.w5(32'h3a8f5c11),
	.w6(32'h3c122254),
	.w7(32'h3b73e344),
	.w8(32'hbc323849),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb09600),
	.w1(32'hba3cba17),
	.w2(32'hbc851203),
	.w3(32'hbc303d6e),
	.w4(32'hbcfde0cc),
	.w5(32'h3b552214),
	.w6(32'h3c3ae57e),
	.w7(32'hbc28325e),
	.w8(32'h3c69cd49),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1eacc),
	.w1(32'hbb02f115),
	.w2(32'hbc4438ec),
	.w3(32'h3ac24884),
	.w4(32'hbc8621e7),
	.w5(32'hbbf7cbd7),
	.w6(32'hb78c5cbf),
	.w7(32'h3b91b811),
	.w8(32'h3cc610e7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9380e7),
	.w1(32'h3c449008),
	.w2(32'hbb92cb7a),
	.w3(32'h3ad5f6a8),
	.w4(32'h3c814242),
	.w5(32'h3be2f4d4),
	.w6(32'hbc8989c6),
	.w7(32'h3c8331b9),
	.w8(32'hbad9f6f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcacf330),
	.w1(32'hbc829311),
	.w2(32'hbc253957),
	.w3(32'hbc560289),
	.w4(32'hbb81a63c),
	.w5(32'hbc9fcb89),
	.w6(32'hbbf03529),
	.w7(32'h3b38aa91),
	.w8(32'h3bc79bc7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5e5e9),
	.w1(32'h3b83adf0),
	.w2(32'h3b3d664b),
	.w3(32'hbc3d9a00),
	.w4(32'h3a4ddf72),
	.w5(32'hbb28c354),
	.w6(32'h3c0f0fca),
	.w7(32'h3c119347),
	.w8(32'hbc03f171),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20abcb),
	.w1(32'hbc79e9a2),
	.w2(32'hbbebcb64),
	.w3(32'hbc646aab),
	.w4(32'hbca639c9),
	.w5(32'h3c16423d),
	.w6(32'h3ca06c4c),
	.w7(32'h39a8c986),
	.w8(32'h3ac7d113),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2e3cf),
	.w1(32'hbc7fcc49),
	.w2(32'hbbb08bb1),
	.w3(32'hbaaaa157),
	.w4(32'h3b984d73),
	.w5(32'h39a53eb5),
	.w6(32'h3c378674),
	.w7(32'hbb92c1fa),
	.w8(32'h3d2bcbf1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9543c24),
	.w1(32'h3a980f44),
	.w2(32'h39f3653e),
	.w3(32'hbb2b4cad),
	.w4(32'h3b5ac7bc),
	.w5(32'h3bc92208),
	.w6(32'hbc99c275),
	.w7(32'hbccad58b),
	.w8(32'h3bb75b80),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4970d0),
	.w1(32'h3d1aa0a5),
	.w2(32'hbc4018c3),
	.w3(32'hbbdedb73),
	.w4(32'h3b9300c9),
	.w5(32'h3bd2be41),
	.w6(32'hba4e408a),
	.w7(32'hbb1898d3),
	.w8(32'hbc2c5cf0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b81f4),
	.w1(32'h3b822bfd),
	.w2(32'hbbba1424),
	.w3(32'h3c11dcfd),
	.w4(32'hbc3c296b),
	.w5(32'hbc6c46d2),
	.w6(32'h3ba16804),
	.w7(32'h3b9bdd60),
	.w8(32'h3b5dda98),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf907e1),
	.w1(32'hbb28c402),
	.w2(32'hbc96e48d),
	.w3(32'hbc26eea1),
	.w4(32'h3cbffb9a),
	.w5(32'hbbcbd10a),
	.w6(32'h3cf51441),
	.w7(32'h3c3ac2e4),
	.w8(32'h390bec97),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cbdab),
	.w1(32'hbd150b38),
	.w2(32'hbb428b17),
	.w3(32'hbc878a7d),
	.w4(32'hbc2b899a),
	.w5(32'h3c706963),
	.w6(32'h3c9132ee),
	.w7(32'hbbd2b87b),
	.w8(32'h3add8e5d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a215586),
	.w1(32'h3cd636e4),
	.w2(32'h3c030b69),
	.w3(32'hbbb3a0d3),
	.w4(32'h3cbebbf4),
	.w5(32'h3c4eba3c),
	.w6(32'hbca24422),
	.w7(32'hbc9ab48d),
	.w8(32'hbc01b487),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bdd4d),
	.w1(32'h3b41c006),
	.w2(32'hbba176ab),
	.w3(32'h3c31fa05),
	.w4(32'h3b986286),
	.w5(32'h3d26ed7f),
	.w6(32'h3c009542),
	.w7(32'hbba7e56c),
	.w8(32'hbb3b365d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2de4fc),
	.w1(32'h3ad93172),
	.w2(32'h3cc05867),
	.w3(32'hbb4b65e4),
	.w4(32'hbc2628e5),
	.w5(32'hbb2e8b93),
	.w6(32'h3a8951b7),
	.w7(32'hbbe6bd3d),
	.w8(32'hbb99f8ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77b447),
	.w1(32'h3c2f9df2),
	.w2(32'hbc3649af),
	.w3(32'hbc2e03c4),
	.w4(32'hbcd82f87),
	.w5(32'hbc453294),
	.w6(32'hbc8e134c),
	.w7(32'hbc9f72f4),
	.w8(32'h3b738e6d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279667),
	.w1(32'h3c71fd82),
	.w2(32'h3b8ca52a),
	.w3(32'h39cadcb7),
	.w4(32'h3b6738b0),
	.w5(32'h3b03043d),
	.w6(32'h3b4bab4a),
	.w7(32'hbb90f687),
	.w8(32'h3b7f417e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b086),
	.w1(32'h3cee38a8),
	.w2(32'h3c62f89f),
	.w3(32'hbc7703ed),
	.w4(32'h394934a1),
	.w5(32'hbc40e93a),
	.w6(32'hbbe78030),
	.w7(32'hbce2f83d),
	.w8(32'hbc332df7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d932c),
	.w1(32'h39a8ffac),
	.w2(32'h3c4125c9),
	.w3(32'h3b821a3e),
	.w4(32'h3bb5469c),
	.w5(32'h3b28801b),
	.w6(32'h3c2cf2cd),
	.w7(32'h3b1ce3c0),
	.w8(32'h3c341516),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1784c),
	.w1(32'hbbade0d0),
	.w2(32'h3b9944ea),
	.w3(32'h3b3b2799),
	.w4(32'hbc05c1b2),
	.w5(32'h3cae0121),
	.w6(32'h3bee4c6f),
	.w7(32'hbd86e8c2),
	.w8(32'hbd12f4f6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831cb9),
	.w1(32'hbbd283af),
	.w2(32'hbc0667da),
	.w3(32'h3b0ef367),
	.w4(32'h3bb131a5),
	.w5(32'h3c16db7c),
	.w6(32'h3ca8d222),
	.w7(32'h3b1d15e9),
	.w8(32'h3b8d1b62),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c456055),
	.w1(32'h3b8ef65a),
	.w2(32'hbb0d62b6),
	.w3(32'hbc1cdc22),
	.w4(32'hbc6bb93e),
	.w5(32'h3aa8b710),
	.w6(32'hbb8467ed),
	.w7(32'hbba0a514),
	.w8(32'hbb0292ce),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b4a5),
	.w1(32'hbbf2abc3),
	.w2(32'h3bd87c3d),
	.w3(32'hbb8aa818),
	.w4(32'hbc05ecea),
	.w5(32'h3929b0ab),
	.w6(32'hba5736e1),
	.w7(32'h3b15b691),
	.w8(32'h3c16f604),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8713),
	.w1(32'hbbd66419),
	.w2(32'hbca76a5d),
	.w3(32'h3c18a4af),
	.w4(32'h3b0ffc8e),
	.w5(32'h3c3edd70),
	.w6(32'h3b93de43),
	.w7(32'h3c0041f5),
	.w8(32'hbb2f4702),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88acf0),
	.w1(32'hbc705652),
	.w2(32'hbd269220),
	.w3(32'h3c299f25),
	.w4(32'h3c5fdd43),
	.w5(32'hbb988e87),
	.w6(32'h3c70f79f),
	.w7(32'h3c6ff74c),
	.w8(32'h3c6c6f59),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8924f3),
	.w1(32'h3cf419c3),
	.w2(32'h3cce0711),
	.w3(32'hbbea9c4c),
	.w4(32'h3cfbc835),
	.w5(32'h3c5548c1),
	.w6(32'hbcae2730),
	.w7(32'hbc41d044),
	.w8(32'hbb38459b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051a05),
	.w1(32'h3cbddc12),
	.w2(32'h3ccc46ae),
	.w3(32'hbb098717),
	.w4(32'hbc550389),
	.w5(32'hbc5480ad),
	.w6(32'h399fdacb),
	.w7(32'hbc6de606),
	.w8(32'hbce7c37c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c588213),
	.w1(32'h3c6eec17),
	.w2(32'hbb7d9707),
	.w3(32'h3b94eb85),
	.w4(32'hba4f97f1),
	.w5(32'hbb08eca5),
	.w6(32'hbbe66a23),
	.w7(32'h3aef2055),
	.w8(32'hbb8d1db0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba006048),
	.w1(32'h3b875717),
	.w2(32'h3bf8a71f),
	.w3(32'hbbf00689),
	.w4(32'hbc84aee8),
	.w5(32'h3b5a16f0),
	.w6(32'h3b041f40),
	.w7(32'hbb8b8c9a),
	.w8(32'h3bd118e7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54b5f4),
	.w1(32'hbc135b86),
	.w2(32'hbc8315b0),
	.w3(32'hbc669558),
	.w4(32'h39aba1ae),
	.w5(32'h3bc8ce27),
	.w6(32'h3cd81e8f),
	.w7(32'h3c0fe0b6),
	.w8(32'hbc18a893),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78c02f),
	.w1(32'h3c3c94d1),
	.w2(32'hbca9971d),
	.w3(32'h3c28d073),
	.w4(32'h3b908ca0),
	.w5(32'hba9531da),
	.w6(32'hbad26c26),
	.w7(32'h3c3f5145),
	.w8(32'h3bd898be),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa1674),
	.w1(32'hbbd446a9),
	.w2(32'h3af13508),
	.w3(32'hbc5f742e),
	.w4(32'hbc63c670),
	.w5(32'hba3c2f58),
	.w6(32'h3b458056),
	.w7(32'hbb216dfc),
	.w8(32'h3c475447),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a62f1),
	.w1(32'h3bbcac42),
	.w2(32'hbb0adc33),
	.w3(32'hba58b0c5),
	.w4(32'h3c5d6d61),
	.w5(32'h391673a9),
	.w6(32'hb893701c),
	.w7(32'hbbe30a45),
	.w8(32'h3bccded8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce28ac),
	.w1(32'hbb1d8c1b),
	.w2(32'hbba27a7f),
	.w3(32'hba8bc88a),
	.w4(32'h3c6191af),
	.w5(32'hbbaeaac9),
	.w6(32'h3b2a2dbb),
	.w7(32'hbbbeec7c),
	.w8(32'h3b22c99e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d18e0),
	.w1(32'h3ad59f16),
	.w2(32'hbc666600),
	.w3(32'hbbb0bbd1),
	.w4(32'hbb7aa453),
	.w5(32'h3b5686c3),
	.w6(32'hbbaa07da),
	.w7(32'h3b8a62a8),
	.w8(32'h3bbf57aa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdca3d0),
	.w1(32'hbc71dcba),
	.w2(32'h3cff6d7a),
	.w3(32'hbb1aa8a4),
	.w4(32'hbcb67086),
	.w5(32'hbc822109),
	.w6(32'h3d411b7e),
	.w7(32'h3c39e627),
	.w8(32'h3c1c177e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a53a),
	.w1(32'hbbfee2bb),
	.w2(32'hbb1fbcba),
	.w3(32'hbbe36f95),
	.w4(32'hbb3b762d),
	.w5(32'hbb88f93e),
	.w6(32'hbae6c233),
	.w7(32'hbbd43769),
	.w8(32'h39ca81aa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb86f99),
	.w1(32'h3afde34c),
	.w2(32'hbb553647),
	.w3(32'hbbd990be),
	.w4(32'hbb77296f),
	.w5(32'hbd13b13b),
	.w6(32'h3c3cc45b),
	.w7(32'h3b18735a),
	.w8(32'hbbc91d03),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8cef),
	.w1(32'h3bcda1ba),
	.w2(32'h3b0d1355),
	.w3(32'h3aa82e48),
	.w4(32'hbbfc2d44),
	.w5(32'h3a50eaf8),
	.w6(32'hbb0c3d42),
	.w7(32'hbbae0677),
	.w8(32'hba7f5b83),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18288b),
	.w1(32'hba9a0f0f),
	.w2(32'h3c54aa08),
	.w3(32'hbb2112bf),
	.w4(32'h3ae49849),
	.w5(32'hbbc4fff8),
	.w6(32'hbc4e0ee5),
	.w7(32'h3b8732d2),
	.w8(32'hbac25f93),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b851d),
	.w1(32'h3c139c2f),
	.w2(32'hba757d93),
	.w3(32'hbc15590a),
	.w4(32'hbb9f73e8),
	.w5(32'h3a253157),
	.w6(32'hbc1c13e9),
	.w7(32'hbb557496),
	.w8(32'h3c33ddb0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a2099),
	.w1(32'hbc9890c4),
	.w2(32'hbbcfe25c),
	.w3(32'hbccd086a),
	.w4(32'hbce34cfe),
	.w5(32'hbb577007),
	.w6(32'h3c84de4d),
	.w7(32'hbad9d2f0),
	.w8(32'h3bd58555),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b2ec),
	.w1(32'hbb013be9),
	.w2(32'hbb935e0c),
	.w3(32'hbaf77b1e),
	.w4(32'h3a827001),
	.w5(32'h3b4262f4),
	.w6(32'h3c54eaf0),
	.w7(32'h3c3b25f0),
	.w8(32'hbc32f7f0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7f0e2),
	.w1(32'h3b68b708),
	.w2(32'h3b590d60),
	.w3(32'h3aa21969),
	.w4(32'hbc09eb39),
	.w5(32'hbc556538),
	.w6(32'h3b810132),
	.w7(32'hba8ae33d),
	.w8(32'h3b3e1104),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a710),
	.w1(32'h3b792fb2),
	.w2(32'h3b193fbd),
	.w3(32'hbb333084),
	.w4(32'h3bf258f2),
	.w5(32'h37babe1b),
	.w6(32'h3b3ae0cb),
	.w7(32'h3c955988),
	.w8(32'hbc3d24c2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815b98),
	.w1(32'h3b596d14),
	.w2(32'hbba02688),
	.w3(32'hbbc2923f),
	.w4(32'h3bdf3b95),
	.w5(32'h3c26322d),
	.w6(32'hbc072ea2),
	.w7(32'h3ce0bf87),
	.w8(32'h3b8f0e5d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b9c80),
	.w1(32'h3b637bd2),
	.w2(32'hbc1474f3),
	.w3(32'h3c5d5d74),
	.w4(32'h3c1eab8a),
	.w5(32'hba71b849),
	.w6(32'h3b5945fd),
	.w7(32'h3ae59118),
	.w8(32'hbc294fae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0089fe),
	.w1(32'hbb969bc0),
	.w2(32'hbb42e339),
	.w3(32'h3afb8532),
	.w4(32'h3c44a70a),
	.w5(32'hbc51220b),
	.w6(32'h3c031232),
	.w7(32'h3a664810),
	.w8(32'h39614e70),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd161488),
	.w1(32'hbc92aedc),
	.w2(32'hbc17a55a),
	.w3(32'hbc367644),
	.w4(32'hba142c23),
	.w5(32'h3c58e3d0),
	.w6(32'h3c83341a),
	.w7(32'h39328e57),
	.w8(32'h3c625a07),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aa042),
	.w1(32'hbbfee7d0),
	.w2(32'h3a2845fd),
	.w3(32'h3c0484d5),
	.w4(32'hbc3206d1),
	.w5(32'hbc2b6af3),
	.w6(32'hbb53addb),
	.w7(32'hbc7d7e23),
	.w8(32'h3c23b714),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb216f3f),
	.w1(32'h3b3e0542),
	.w2(32'h3bc61215),
	.w3(32'hba3e1d3d),
	.w4(32'h3c82705c),
	.w5(32'hbc5c1c3c),
	.w6(32'h393f8ebc),
	.w7(32'h3b56fc41),
	.w8(32'hbcb84362),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5250ed),
	.w1(32'hbbb2b6d9),
	.w2(32'hb8e12766),
	.w3(32'h3bb22b6b),
	.w4(32'hbc15b8e8),
	.w5(32'h39c0165c),
	.w6(32'hbbab8d2b),
	.w7(32'h3b1625a4),
	.w8(32'hbaf9ed14),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc51b5),
	.w1(32'h3b5cecc3),
	.w2(32'hb9f6ceb0),
	.w3(32'h3aed353f),
	.w4(32'hbc503cdb),
	.w5(32'hbc182961),
	.w6(32'hbba3548f),
	.w7(32'h3bc59937),
	.w8(32'h3a78c3d8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc125bf8),
	.w1(32'h3b4fa17d),
	.w2(32'h3c03faca),
	.w3(32'h3aa6f52b),
	.w4(32'h3b1b00bd),
	.w5(32'hbc7892f1),
	.w6(32'hba85eaef),
	.w7(32'h3c1c5c52),
	.w8(32'h3c21e314),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc3a61),
	.w1(32'hbb202d1a),
	.w2(32'h3b376ad0),
	.w3(32'h3aeadd0b),
	.w4(32'hbc85c487),
	.w5(32'h3c04de24),
	.w6(32'hbb8b1374),
	.w7(32'hbbd12a11),
	.w8(32'h3c9b8026),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c209dbe),
	.w1(32'h3a897d79),
	.w2(32'hbc8c00b7),
	.w3(32'h3c348dce),
	.w4(32'hbbce1439),
	.w5(32'hbbf68198),
	.w6(32'h3c509ce8),
	.w7(32'h3bb880b1),
	.w8(32'h3c85c632),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc513698),
	.w1(32'hbb8a4347),
	.w2(32'hba54b4e1),
	.w3(32'hbbc458f2),
	.w4(32'h3a7d019d),
	.w5(32'hbc018495),
	.w6(32'h3c67d4f4),
	.w7(32'hbc180ae5),
	.w8(32'hbb8a25dd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f020b),
	.w1(32'h3cd52414),
	.w2(32'hba578d02),
	.w3(32'h3b5075bf),
	.w4(32'h3ca1710a),
	.w5(32'h3b8a01ca),
	.w6(32'hbc80eec0),
	.w7(32'hbc78dbf5),
	.w8(32'h3b1f9cc3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981a64f),
	.w1(32'hbc8e9e25),
	.w2(32'hbbab7f08),
	.w3(32'h3b5db251),
	.w4(32'h3a411598),
	.w5(32'hba726a53),
	.w6(32'h3b3848a9),
	.w7(32'h3c2d2846),
	.w8(32'hbc2b1deb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafafd86),
	.w1(32'hbb869e49),
	.w2(32'hb9d45a2b),
	.w3(32'h3c87951a),
	.w4(32'h3b9e2349),
	.w5(32'h3b8c7a91),
	.w6(32'h3b1af5be),
	.w7(32'h3ba4db48),
	.w8(32'hbb9a51b3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17b00c),
	.w1(32'hba334db3),
	.w2(32'h3c507e19),
	.w3(32'h3b9e6f45),
	.w4(32'hb8e3144b),
	.w5(32'hbac3097a),
	.w6(32'hbad535d1),
	.w7(32'h3b07871c),
	.w8(32'hbc18db2c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc142a76),
	.w1(32'hbb699ba0),
	.w2(32'hbc086ca8),
	.w3(32'hbc519d00),
	.w4(32'hbc06bcd1),
	.w5(32'hb9d32051),
	.w6(32'hbb4fc314),
	.w7(32'h3bc56b24),
	.w8(32'h3c268cfe),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9204af),
	.w1(32'h3ae6e566),
	.w2(32'h3b6427ca),
	.w3(32'h3c884e60),
	.w4(32'h3a04c35d),
	.w5(32'h38e95ffe),
	.w6(32'h3b7f3977),
	.w7(32'h3b81bdc0),
	.w8(32'hbadb520c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24831e),
	.w1(32'hbc8cc7e1),
	.w2(32'h3b8475b8),
	.w3(32'h3b24d1c6),
	.w4(32'hbc506c8f),
	.w5(32'h39fa64db),
	.w6(32'h3bf8a88a),
	.w7(32'hbbde155c),
	.w8(32'hba35ae10),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceab8cb),
	.w1(32'hbc3026f4),
	.w2(32'hbc055599),
	.w3(32'h3af4fb04),
	.w4(32'hbc99b45a),
	.w5(32'h3b185e07),
	.w6(32'h3c546a41),
	.w7(32'h3c2c75fd),
	.w8(32'hbba77e5b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5819d9),
	.w1(32'hbc79bf2e),
	.w2(32'h3becf099),
	.w3(32'hbc316f51),
	.w4(32'h3ae1577c),
	.w5(32'h3b3fa812),
	.w6(32'hbbf6014f),
	.w7(32'h3b00ccbf),
	.w8(32'hb8caf418),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4c22f),
	.w1(32'h39a63642),
	.w2(32'hbc6a230d),
	.w3(32'hbbb18d02),
	.w4(32'hbb00e548),
	.w5(32'hba13df05),
	.w6(32'h3ae94e1c),
	.w7(32'hbb0069f5),
	.w8(32'h3a04dcb7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac73f8),
	.w1(32'hbc8c333b),
	.w2(32'h3ba0cf4d),
	.w3(32'h3bb90883),
	.w4(32'hbbca1f9b),
	.w5(32'hbb94cc70),
	.w6(32'h3c0ce5f9),
	.w7(32'hbc09db49),
	.w8(32'h3b0f1ddb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb7d1),
	.w1(32'hbc8b9467),
	.w2(32'hbc161018),
	.w3(32'hbbb1a1ce),
	.w4(32'h3a175bd9),
	.w5(32'h3ab8e871),
	.w6(32'hbc453f03),
	.w7(32'hbb7da8db),
	.w8(32'h3b516213),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71a1dc),
	.w1(32'h3bc80ede),
	.w2(32'hbb6f2027),
	.w3(32'h3b1869bc),
	.w4(32'hbbbad2b4),
	.w5(32'h3b9e3599),
	.w6(32'hbcb7e4cd),
	.w7(32'hbb9e27a3),
	.w8(32'h3cb6b95b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8aeec),
	.w1(32'hbba6689d),
	.w2(32'hbc1b42bd),
	.w3(32'hbc4f5b19),
	.w4(32'h3b586710),
	.w5(32'hbc13fc90),
	.w6(32'h3c5236fa),
	.w7(32'hbc856b73),
	.w8(32'h3be20192),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8671e9),
	.w1(32'hb9a57e1f),
	.w2(32'hbaf54fcb),
	.w3(32'h3c25a9c8),
	.w4(32'hbc4d6f06),
	.w5(32'h3b5c4df7),
	.w6(32'h3a98d01e),
	.w7(32'h3acf8e1e),
	.w8(32'h3cce6eac),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e92c5),
	.w1(32'h3c5628e9),
	.w2(32'hbb151ac2),
	.w3(32'h3c220bda),
	.w4(32'h3bc6235c),
	.w5(32'hbc09db9c),
	.w6(32'hbab42812),
	.w7(32'hbb2e5b60),
	.w8(32'hbc0d1114),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1e0da),
	.w1(32'h3bea1ed0),
	.w2(32'h3ca9a89d),
	.w3(32'hbc89118d),
	.w4(32'h3b7bd3d3),
	.w5(32'h3c755bd3),
	.w6(32'h3d2dfb5d),
	.w7(32'h3b3041a4),
	.w8(32'h3c3340dc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87cbce),
	.w1(32'h3c4cb0a4),
	.w2(32'h3cadfdfa),
	.w3(32'h3cba326d),
	.w4(32'h3cae5dc8),
	.w5(32'h3d07b4bf),
	.w6(32'hbb3b3421),
	.w7(32'h39d47948),
	.w8(32'h3b625aaa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc561991),
	.w1(32'h3b210de3),
	.w2(32'hbbd45e7e),
	.w3(32'h3c12d9d1),
	.w4(32'hbb07ff7c),
	.w5(32'hbc178ed4),
	.w6(32'h3bb2832a),
	.w7(32'h3aa4b321),
	.w8(32'hbb6f3aaa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74307f),
	.w1(32'hbc057f62),
	.w2(32'hbbe86df7),
	.w3(32'h3d1724f8),
	.w4(32'h3beeb1bf),
	.w5(32'hbc7f5421),
	.w6(32'h3c0e75b7),
	.w7(32'h3c3174d3),
	.w8(32'h3c61bd3f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02dca),
	.w1(32'hbc1f3480),
	.w2(32'hbbe739be),
	.w3(32'hbc23ed82),
	.w4(32'hbcc3490c),
	.w5(32'hbb28afe6),
	.w6(32'h3d371151),
	.w7(32'hbbc185c5),
	.w8(32'hbbdea3cf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e159),
	.w1(32'h3cab279c),
	.w2(32'hbc743a9a),
	.w3(32'hbbd1cc5f),
	.w4(32'hbbb99f86),
	.w5(32'hbc07a1ba),
	.w6(32'hbc5ecd26),
	.w7(32'hbb2f74f8),
	.w8(32'hbbd76464),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8f5c5),
	.w1(32'hbcb1ac76),
	.w2(32'hbd0c25a6),
	.w3(32'h3c0aca1d),
	.w4(32'h3cd1bb08),
	.w5(32'hbc2f734f),
	.w6(32'h3bafe352),
	.w7(32'h3b1dc01c),
	.w8(32'h3c8d0511),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f655f),
	.w1(32'h3cd44ac5),
	.w2(32'h3d0115de),
	.w3(32'h3bedb88e),
	.w4(32'hbae100eb),
	.w5(32'hbc676882),
	.w6(32'hb9040d78),
	.w7(32'hbc9f2d0f),
	.w8(32'h3d04d320),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0429e0),
	.w1(32'hbc7952e0),
	.w2(32'hbc7d53d2),
	.w3(32'h3a7a86e5),
	.w4(32'h3d022ea6),
	.w5(32'h3d255190),
	.w6(32'hbc0292df),
	.w7(32'hbb9c4cd2),
	.w8(32'hbb0fafb8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f5049),
	.w1(32'h3c0693af),
	.w2(32'h3afed2b5),
	.w3(32'hbd106c1f),
	.w4(32'hbc4fc001),
	.w5(32'h3ad0cb51),
	.w6(32'h3c248b66),
	.w7(32'hbc0fa196),
	.w8(32'h3c67d1d0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f1921),
	.w1(32'h3d45a272),
	.w2(32'hbbbb7ec8),
	.w3(32'hbc3169de),
	.w4(32'h3cd4ddb5),
	.w5(32'hbbfcba3a),
	.w6(32'h3c39af3d),
	.w7(32'hbaf2d5af),
	.w8(32'h38dcd7ec),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c549b9d),
	.w1(32'h3c2322db),
	.w2(32'h3c4e2ca5),
	.w3(32'h3b9b4d64),
	.w4(32'h3ca97b64),
	.w5(32'h37a2cb58),
	.w6(32'hbafa3d11),
	.w7(32'h3bc4d1d0),
	.w8(32'h3a9d2f49),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35109a),
	.w1(32'hbcb51fdc),
	.w2(32'h3b919638),
	.w3(32'hbacddac6),
	.w4(32'hbb580c56),
	.w5(32'hbc1f9292),
	.w6(32'h3d35804f),
	.w7(32'hbc36a9b8),
	.w8(32'h3c725c3f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd021438),
	.w1(32'hbd001431),
	.w2(32'hbbfb141c),
	.w3(32'h3c109222),
	.w4(32'hbbfd6219),
	.w5(32'hbc0de2b8),
	.w6(32'hbc6733f0),
	.w7(32'h3c86ad38),
	.w8(32'h3c4c77e4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c857c),
	.w1(32'hbd08aeb0),
	.w2(32'hbd123f60),
	.w3(32'h3b122995),
	.w4(32'h3a3f2cbc),
	.w5(32'hbc1034c6),
	.w6(32'h3c8e3f0b),
	.w7(32'hbbc4f5ff),
	.w8(32'h3d44e4c1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36710b),
	.w1(32'h3cffe809),
	.w2(32'hbc0a96c6),
	.w3(32'h3d156648),
	.w4(32'h3ce6cd89),
	.w5(32'h3b9562b8),
	.w6(32'hbbed6b3e),
	.w7(32'h3bc33c1d),
	.w8(32'hbc7db720),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0466),
	.w1(32'h3caf4b64),
	.w2(32'h3c600645),
	.w3(32'h3ba087d6),
	.w4(32'hbad77a0a),
	.w5(32'hbabfc512),
	.w6(32'hbbf63abb),
	.w7(32'hba98e405),
	.w8(32'h3c5562ca),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafac64),
	.w1(32'hbd55361e),
	.w2(32'hbc74d983),
	.w3(32'h3d0422dc),
	.w4(32'h3c3376f0),
	.w5(32'h3c3da2a5),
	.w6(32'h3c233c42),
	.w7(32'h3cb10194),
	.w8(32'h3bdba2bd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0f384),
	.w1(32'h3cab7693),
	.w2(32'h3c7529b8),
	.w3(32'h3bd4e199),
	.w4(32'hbc2402b9),
	.w5(32'hbb708ce6),
	.w6(32'h3c47fe2f),
	.w7(32'h3c524c3d),
	.w8(32'hb9bdded1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd098598),
	.w1(32'hbce48a67),
	.w2(32'hbcac94a6),
	.w3(32'hb8ff3026),
	.w4(32'hbbb05371),
	.w5(32'hbc625683),
	.w6(32'h3d0d4601),
	.w7(32'h3c213b80),
	.w8(32'hbc695f74),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2067),
	.w1(32'h3b358e42),
	.w2(32'hbc352cfd),
	.w3(32'hbc1574a3),
	.w4(32'hbb2902bf),
	.w5(32'hbbe4eb26),
	.w6(32'hbbf064fe),
	.w7(32'h3be6b6f2),
	.w8(32'h3b554a89),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b33eb),
	.w1(32'hb85132a5),
	.w2(32'h3b98d7ff),
	.w3(32'hbd2a56a8),
	.w4(32'hbb6f5489),
	.w5(32'h3b8a4601),
	.w6(32'h3b5d3be6),
	.w7(32'h3adcc8a6),
	.w8(32'hbb993821),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3d85a),
	.w1(32'hbbbad664),
	.w2(32'h3b4451f6),
	.w3(32'h3cdb98cf),
	.w4(32'h3d12f62a),
	.w5(32'h3af1f0a8),
	.w6(32'hbc96ebb4),
	.w7(32'hbbc5e82a),
	.w8(32'hbcedeb4c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3064e7),
	.w1(32'hbc2aab54),
	.w2(32'h3b95290d),
	.w3(32'hbba43242),
	.w4(32'hbc874435),
	.w5(32'hbd080586),
	.w6(32'h3bf835f0),
	.w7(32'hbb02f785),
	.w8(32'hbc0aa864),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c0e46),
	.w1(32'hbd02011d),
	.w2(32'h3cb2f1dc),
	.w3(32'h3c5a3d13),
	.w4(32'h3d072753),
	.w5(32'hbb86b35f),
	.w6(32'hbba230cd),
	.w7(32'hbc00396c),
	.w8(32'h3be03d2a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b305db8),
	.w1(32'hba9b025e),
	.w2(32'h3cba8242),
	.w3(32'hbc47c60e),
	.w4(32'h3c026bb7),
	.w5(32'h37ec108f),
	.w6(32'hbcf091f1),
	.w7(32'h3c287d53),
	.w8(32'h3b527804),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d66221c),
	.w1(32'h3d08fbd6),
	.w2(32'hbc3640fb),
	.w3(32'h3c8b1e0e),
	.w4(32'h3c46e5fa),
	.w5(32'h3c2abaad),
	.w6(32'hbbb146f2),
	.w7(32'h3c04a562),
	.w8(32'h3c65ba62),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3deae4),
	.w1(32'h3d30b92a),
	.w2(32'h3b6dcbac),
	.w3(32'h3b09c371),
	.w4(32'h3ae17a70),
	.w5(32'hbc65cffc),
	.w6(32'hbb310d14),
	.w7(32'h3c3094eb),
	.w8(32'h3c53477d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc967e16),
	.w1(32'hbb5df5bf),
	.w2(32'hbc565c65),
	.w3(32'hbc84b947),
	.w4(32'hbb081508),
	.w5(32'h3cad3e90),
	.w6(32'hbc1d56c7),
	.w7(32'h3a9e3e06),
	.w8(32'h3b3dfb97),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df469),
	.w1(32'hbabc517f),
	.w2(32'h3a92c3d8),
	.w3(32'hbcce0b6d),
	.w4(32'h3b4393b7),
	.w5(32'hbb97d1e9),
	.w6(32'h3c23cc3f),
	.w7(32'h3ccaa776),
	.w8(32'h3c9de9c6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d6df9),
	.w1(32'h3b9b098e),
	.w2(32'h3ae48fa5),
	.w3(32'h3bed6057),
	.w4(32'h3afafa3a),
	.w5(32'h3c15d218),
	.w6(32'h3b561ed6),
	.w7(32'h3ad2909f),
	.w8(32'h3b770d33),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5f35),
	.w1(32'h3c09ccad),
	.w2(32'hbc09d882),
	.w3(32'h3c145927),
	.w4(32'h3c3fc891),
	.w5(32'h3ceabb18),
	.w6(32'h3c6624b4),
	.w7(32'h3c46b890),
	.w8(32'hbb9f2574),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd05be5),
	.w1(32'hb8d3361a),
	.w2(32'h3ca6bacd),
	.w3(32'h3ad36dbf),
	.w4(32'h3b68ca90),
	.w5(32'h3af00e3e),
	.w6(32'hbae57e16),
	.w7(32'h3a3b4a4e),
	.w8(32'h3b2fdc30),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81251d),
	.w1(32'hbc04fb99),
	.w2(32'h3bb3fd57),
	.w3(32'hbbc88a1a),
	.w4(32'h3c38213b),
	.w5(32'h3c25a7d1),
	.w6(32'hbafd2158),
	.w7(32'h3b5710aa),
	.w8(32'h3cf2840c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950b15c),
	.w1(32'h3a7b3d5c),
	.w2(32'h3c4d79e3),
	.w3(32'hbc6958f1),
	.w4(32'h397179d1),
	.w5(32'hbc1518fa),
	.w6(32'h38a69781),
	.w7(32'h3c99aed7),
	.w8(32'h3c477167),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49ef14),
	.w1(32'h3a3d0d0d),
	.w2(32'hbb886d22),
	.w3(32'h3b0720d8),
	.w4(32'hbb8ac4d9),
	.w5(32'hbc983e7a),
	.w6(32'hb91fd23b),
	.w7(32'hbc0296ce),
	.w8(32'h3b1dfe8d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd245a16),
	.w1(32'hbabac851),
	.w2(32'h3c7e4244),
	.w3(32'h3ca84832),
	.w4(32'hbbb4ce8c),
	.w5(32'h3ba1c567),
	.w6(32'h3c6a764d),
	.w7(32'h3be9535c),
	.w8(32'h3b0288ca),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57bc94),
	.w1(32'h3cb26f13),
	.w2(32'h3c1a31cc),
	.w3(32'hbaec0d11),
	.w4(32'h3c143f6e),
	.w5(32'hbb472978),
	.w6(32'hbb68f438),
	.w7(32'hbcf64390),
	.w8(32'hbc598484),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81e1f8),
	.w1(32'hbb4bc203),
	.w2(32'h3bdbad4c),
	.w3(32'hb98eb549),
	.w4(32'hbc799278),
	.w5(32'h3bc1d998),
	.w6(32'hba98b5c4),
	.w7(32'hbb2c50c8),
	.w8(32'h3b810f46),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036a6f),
	.w1(32'hbb479c26),
	.w2(32'h39636c4b),
	.w3(32'h3ac9ba53),
	.w4(32'h3c814834),
	.w5(32'h39d33277),
	.w6(32'hbb693701),
	.w7(32'h3c47fd20),
	.w8(32'h3b030efd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2937f2),
	.w1(32'hb9096455),
	.w2(32'hbb33392b),
	.w3(32'hbaf37d57),
	.w4(32'h3b231c0d),
	.w5(32'hbcbdce91),
	.w6(32'h3b8bfa1c),
	.w7(32'hbabf0c4c),
	.w8(32'h388f9a01),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e5ce1),
	.w1(32'h3a4a3e66),
	.w2(32'h3a3ee438),
	.w3(32'h3b21c713),
	.w4(32'h3b32f2e5),
	.w5(32'hbbf43adc),
	.w6(32'hbb9dfc5c),
	.w7(32'hbc448ef2),
	.w8(32'h3bc07e3d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05877f),
	.w1(32'hbba907ed),
	.w2(32'hbc2412d9),
	.w3(32'h3bb81a69),
	.w4(32'hbb5a5a78),
	.w5(32'hbcd7e254),
	.w6(32'h3a8d95db),
	.w7(32'h39f847d2),
	.w8(32'hbb1f524e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd006342),
	.w1(32'h3ca6b5f8),
	.w2(32'h3b36f805),
	.w3(32'hbc5f73bb),
	.w4(32'hbcc99e7a),
	.w5(32'hba6b809e),
	.w6(32'h3c056686),
	.w7(32'h3bf1014f),
	.w8(32'h3b84527d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb187a22),
	.w1(32'hbb8b086e),
	.w2(32'hba9a945c),
	.w3(32'h3b4d3d93),
	.w4(32'hbbe9b500),
	.w5(32'hbb89f0e4),
	.w6(32'h3aeb9b84),
	.w7(32'h3c2b0980),
	.w8(32'hbb35e013),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb645dd1),
	.w1(32'hba89526b),
	.w2(32'h3ba46ace),
	.w3(32'h3aaeaa56),
	.w4(32'h3c79b01e),
	.w5(32'hbc21c957),
	.w6(32'hba73e2bf),
	.w7(32'h3b50b3b6),
	.w8(32'h3badefac),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc69bf2),
	.w1(32'hba38d659),
	.w2(32'h3c5cc2a1),
	.w3(32'hbb7a3b73),
	.w4(32'hbbf06895),
	.w5(32'h3af92577),
	.w6(32'hbb780d5b),
	.w7(32'h3aebb23b),
	.w8(32'hbc86c7a0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba79069),
	.w1(32'hbba08c59),
	.w2(32'h3b0fe772),
	.w3(32'h3bad9dde),
	.w4(32'h396eb185),
	.w5(32'h3bfe52cf),
	.w6(32'hbac8015d),
	.w7(32'h3b940dee),
	.w8(32'hbc090476),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9113c5),
	.w1(32'hbcabe8bd),
	.w2(32'hbbb53b39),
	.w3(32'hbb476c55),
	.w4(32'h3c6dc494),
	.w5(32'h3c8bd39d),
	.w6(32'hbb9be04f),
	.w7(32'h3c0c0cb3),
	.w8(32'h3a4a3625),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9faa2),
	.w1(32'hbc82ffe9),
	.w2(32'hbacc8681),
	.w3(32'hbb2e3d68),
	.w4(32'hbc143d03),
	.w5(32'hbc1b6f8b),
	.w6(32'h3a3decae),
	.w7(32'hbb61f370),
	.w8(32'h3b15ecff),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170b7c),
	.w1(32'h3c04a669),
	.w2(32'hbba0b51d),
	.w3(32'h3c2df8c5),
	.w4(32'hbbb035a6),
	.w5(32'hbc1db2d9),
	.w6(32'hbbe0fc22),
	.w7(32'h3b9d56a0),
	.w8(32'hbad21e1f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3dd7a),
	.w1(32'hbc416cb7),
	.w2(32'h3b4bf5d8),
	.w3(32'hbc3b8ed1),
	.w4(32'hbc185e1a),
	.w5(32'hba24e619),
	.w6(32'h3ba510f7),
	.w7(32'h3b8d463c),
	.w8(32'hbb9aa17d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd095ec),
	.w1(32'hbc6135e2),
	.w2(32'hbc4f87d6),
	.w3(32'h3b940049),
	.w4(32'h3c3731a1),
	.w5(32'hbc4665c9),
	.w6(32'h3c07ce06),
	.w7(32'h3c12469f),
	.w8(32'h3c466fa8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba73a0),
	.w1(32'h3c9a2059),
	.w2(32'hbc0610f2),
	.w3(32'h3b804cc1),
	.w4(32'h3bee3f32),
	.w5(32'h3b203424),
	.w6(32'h3aa5f223),
	.w7(32'h3b26941b),
	.w8(32'hbc048445),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79a364),
	.w1(32'hbbce9923),
	.w2(32'hbac40a21),
	.w3(32'hbc06706f),
	.w4(32'h3cd31912),
	.w5(32'hbc3e8353),
	.w6(32'hb8d4869e),
	.w7(32'h38ba9679),
	.w8(32'hbaade908),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce928c9),
	.w1(32'hbada6165),
	.w2(32'h3b2067a0),
	.w3(32'hbbf9e7b9),
	.w4(32'h3b824aa4),
	.w5(32'h3a4d6c5c),
	.w6(32'hbc25cff8),
	.w7(32'h3abef0bc),
	.w8(32'hbc6edc25),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e32ad),
	.w1(32'h3cb0aaa6),
	.w2(32'h3c84571f),
	.w3(32'hbc5f444a),
	.w4(32'h3c72ea09),
	.w5(32'hbb6294fb),
	.w6(32'h3b8bda65),
	.w7(32'hbba2fd46),
	.w8(32'hbc874fd2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3309),
	.w1(32'hbbd8e65d),
	.w2(32'hbc99dfa0),
	.w3(32'h3c01bcdb),
	.w4(32'hbb6255d5),
	.w5(32'hba5727d9),
	.w6(32'hbb613c83),
	.w7(32'h3bbbd0ac),
	.w8(32'h3bb7d738),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4391),
	.w1(32'hbb4f6109),
	.w2(32'hba689b04),
	.w3(32'hba8c1c0a),
	.w4(32'hb9a6dedf),
	.w5(32'hbbf65250),
	.w6(32'h3b655eb4),
	.w7(32'hbb27d814),
	.w8(32'h3bb12c1c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69b0d4),
	.w1(32'hba62984e),
	.w2(32'hbc5dac79),
	.w3(32'h3c93ada0),
	.w4(32'h3bfa5e9c),
	.w5(32'h3c193442),
	.w6(32'hbc5dcf98),
	.w7(32'hbbc65d11),
	.w8(32'hbc717c60),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a851),
	.w1(32'hbccff3bc),
	.w2(32'hb9fbc2b5),
	.w3(32'hbc2371ce),
	.w4(32'hbb5f04ae),
	.w5(32'hbbcac3eb),
	.w6(32'hbb186c72),
	.w7(32'hbc3c136a),
	.w8(32'hbb3b2f68),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1bf0),
	.w1(32'hbabfc9ea),
	.w2(32'h3b679a1a),
	.w3(32'hba23d365),
	.w4(32'h3bc0f0ef),
	.w5(32'hb9f728d6),
	.w6(32'h3bbb50cb),
	.w7(32'hbb832aee),
	.w8(32'h3a58c79f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4389b3),
	.w1(32'hbc24ddc3),
	.w2(32'hbb776717),
	.w3(32'hbcbdc79e),
	.w4(32'hbc74e537),
	.w5(32'hbb67f3c1),
	.w6(32'h3b884c97),
	.w7(32'h3bcca5ad),
	.w8(32'h3c43da57),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf07a50),
	.w1(32'h3c6ce0b0),
	.w2(32'hbc7b6f32),
	.w3(32'hbb01263b),
	.w4(32'hba2c9ef7),
	.w5(32'hbd009e77),
	.w6(32'hbb81fe56),
	.w7(32'h3ba60ad5),
	.w8(32'hba44e6b7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1605e6),
	.w1(32'hbc5b5b37),
	.w2(32'hbb19f561),
	.w3(32'hbb7d5422),
	.w4(32'hbcdc5ffa),
	.w5(32'h3bdfddca),
	.w6(32'h3c62f007),
	.w7(32'hbc749f7e),
	.w8(32'hbb20986b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5e9c3),
	.w1(32'h3d06ff21),
	.w2(32'hbbda208e),
	.w3(32'h3ca8ebf4),
	.w4(32'hbc241f7e),
	.w5(32'hbb448d3b),
	.w6(32'h3a7c7056),
	.w7(32'hbae79312),
	.w8(32'hb903e3c4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3460ca),
	.w1(32'hbc441abf),
	.w2(32'h3b2b2f82),
	.w3(32'h3c3c2380),
	.w4(32'hbcae9c82),
	.w5(32'h3a052914),
	.w6(32'h3c982ec9),
	.w7(32'h3c3b4ffe),
	.w8(32'h3ae0fc96),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc49b7c),
	.w1(32'h3bec03ca),
	.w2(32'h3aab5a4f),
	.w3(32'hbafa08d9),
	.w4(32'hbc4f3476),
	.w5(32'h39f468a8),
	.w6(32'h3b77063f),
	.w7(32'hbc8de31b),
	.w8(32'hbbe2f061),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2345f4),
	.w1(32'h3c1da017),
	.w2(32'h3b205f87),
	.w3(32'hbaa37d01),
	.w4(32'h3bcbd67d),
	.w5(32'hba0fcccc),
	.w6(32'hbc03eb04),
	.w7(32'hbc32bd1c),
	.w8(32'hbb5c00ac),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b410241),
	.w1(32'hba8dd514),
	.w2(32'hbc48fa4a),
	.w3(32'h3c0c9b63),
	.w4(32'h3c226402),
	.w5(32'hbb933ff0),
	.w6(32'h3be6c1da),
	.w7(32'hbb5647fc),
	.w8(32'hbbb22825),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8385c),
	.w1(32'hbb587d4a),
	.w2(32'h3c01d602),
	.w3(32'hbb31beb9),
	.w4(32'hbc23b737),
	.w5(32'h3b394b2b),
	.w6(32'h3b1dc761),
	.w7(32'h3aac5fbe),
	.w8(32'h3cc05874),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bf6fb),
	.w1(32'hbab15642),
	.w2(32'h3b92e381),
	.w3(32'h3b0d4c52),
	.w4(32'h3a6df22b),
	.w5(32'h3abb76fa),
	.w6(32'h3c2fd0f0),
	.w7(32'h3b95ea22),
	.w8(32'h3bf42a3d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca27f28),
	.w1(32'h3c704f9a),
	.w2(32'h3a35f15f),
	.w3(32'h3af2db34),
	.w4(32'h3c650440),
	.w5(32'h3b98d70a),
	.w6(32'h3a199373),
	.w7(32'hbb060d15),
	.w8(32'hb824d685),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0609b),
	.w1(32'hba263bf3),
	.w2(32'hba5f287f),
	.w3(32'h3b14642c),
	.w4(32'hbbba191b),
	.w5(32'hbb01669b),
	.w6(32'h3be8a9fa),
	.w7(32'h3b025935),
	.w8(32'hbb8ba5e6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb71afb),
	.w1(32'hbb001af0),
	.w2(32'h3b947e16),
	.w3(32'h3b1aa715),
	.w4(32'hbc167271),
	.w5(32'h3c3ed964),
	.w6(32'h3bde4513),
	.w7(32'h3af3e037),
	.w8(32'hbb6aa35f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaced02),
	.w1(32'hbbeb4e84),
	.w2(32'hbc408fde),
	.w3(32'hbc0c9639),
	.w4(32'hbb4f6586),
	.w5(32'hbb1fafa9),
	.w6(32'h3c229dda),
	.w7(32'h3934ef19),
	.w8(32'h3b864852),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c104099),
	.w1(32'h3c66e93b),
	.w2(32'h3b5b4174),
	.w3(32'h3c074533),
	.w4(32'hbb182917),
	.w5(32'h3892a153),
	.w6(32'h3ba17662),
	.w7(32'h3aae6c65),
	.w8(32'h3bec91c2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd66471),
	.w1(32'hbb176cad),
	.w2(32'h3b60e615),
	.w3(32'hbb9caa4c),
	.w4(32'h3b4c0613),
	.w5(32'hbb086e41),
	.w6(32'hbab19f08),
	.w7(32'hbaed7fb5),
	.w8(32'h3c69f04b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed72f1),
	.w1(32'hbb8cee0c),
	.w2(32'h3b405beb),
	.w3(32'h3a42b562),
	.w4(32'hbc5e9701),
	.w5(32'hbb35866e),
	.w6(32'hbbacfa43),
	.w7(32'hbaf0fbc0),
	.w8(32'hbb781e46),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c991a05),
	.w1(32'h3c00a583),
	.w2(32'hbbec53bb),
	.w3(32'h3b56cbec),
	.w4(32'hbad52098),
	.w5(32'hbbcf51cb),
	.w6(32'h3c8c381e),
	.w7(32'h3bb0b26d),
	.w8(32'h3b0cc462),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbbe1),
	.w1(32'h3bd0e7b1),
	.w2(32'h3a6917b7),
	.w3(32'hbcbecb5e),
	.w4(32'hbbd27844),
	.w5(32'h3a36b0ae),
	.w6(32'hbbc3119d),
	.w7(32'h3b6e0491),
	.w8(32'h3c5789ab),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa13c57),
	.w1(32'h3c75d1a6),
	.w2(32'h3cd58f92),
	.w3(32'hbc1488a2),
	.w4(32'hbbbcfced),
	.w5(32'hbc2dc925),
	.w6(32'hbb602a57),
	.w7(32'hbd293347),
	.w8(32'h3bc9832b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a916a),
	.w1(32'h3c912f10),
	.w2(32'hbb850777),
	.w3(32'h3c15ac72),
	.w4(32'h3ba90fbf),
	.w5(32'hbba58355),
	.w6(32'hbc2af068),
	.w7(32'h3c516529),
	.w8(32'hbc2c3625),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c782ac9),
	.w1(32'hbc48256b),
	.w2(32'hbbdc2dcb),
	.w3(32'hbb0902e1),
	.w4(32'hbba10373),
	.w5(32'hbc3a718c),
	.w6(32'hbb41d0cd),
	.w7(32'h3c1621d6),
	.w8(32'h394514a8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e66a0),
	.w1(32'hbc1ec278),
	.w2(32'h3d54aed7),
	.w3(32'h3c093f09),
	.w4(32'hbcdf73a0),
	.w5(32'hbc466ae3),
	.w6(32'hbbf8fffe),
	.w7(32'h3b892399),
	.w8(32'hbb16250d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf6fdf),
	.w1(32'h3c80bf63),
	.w2(32'h3ba2dc5a),
	.w3(32'hbbfdbdb8),
	.w4(32'hbb7fa52a),
	.w5(32'hbb9304cb),
	.w6(32'hbc30b5e9),
	.w7(32'h3c3d7d3f),
	.w8(32'hbb8e219d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b482bc7),
	.w1(32'hb9f576b4),
	.w2(32'hbad115db),
	.w3(32'hbc62763c),
	.w4(32'h3b095a8b),
	.w5(32'hbb9a5fa5),
	.w6(32'hbbe90320),
	.w7(32'h3cad33e8),
	.w8(32'hbc3e4750),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1aab89),
	.w1(32'hbbaf71a0),
	.w2(32'hbb2323c2),
	.w3(32'hbcfc8031),
	.w4(32'hbc80635f),
	.w5(32'hbb64a56b),
	.w6(32'h3c0495fe),
	.w7(32'h3c163dc9),
	.w8(32'h3c39fef1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8072c2),
	.w1(32'hbcc92386),
	.w2(32'hbc988ae6),
	.w3(32'h3c39794f),
	.w4(32'hbd34dec6),
	.w5(32'hbbeedc13),
	.w6(32'h3c616a7e),
	.w7(32'h3c0d46f5),
	.w8(32'hbafb538c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51a66b),
	.w1(32'h3c4e4804),
	.w2(32'hbca1ba16),
	.w3(32'hbc4ab33d),
	.w4(32'hbc8edbfe),
	.w5(32'hbb6788f1),
	.w6(32'h3c06c96c),
	.w7(32'h3d09cc3a),
	.w8(32'h3c202aeb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf575c8),
	.w1(32'hbadd288e),
	.w2(32'h3c359335),
	.w3(32'h3c2cd525),
	.w4(32'h3b3fe24b),
	.w5(32'h3ac12511),
	.w6(32'hbbec076a),
	.w7(32'hb9df73cd),
	.w8(32'hbc43bac2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950d4ad),
	.w1(32'hbbeb7b15),
	.w2(32'hbc0751c5),
	.w3(32'h3c059c5d),
	.w4(32'hbc035863),
	.w5(32'hbbff383f),
	.w6(32'hbacc12e8),
	.w7(32'hbc3bc92e),
	.w8(32'hba800ae4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57174a),
	.w1(32'h3a2ef41e),
	.w2(32'h3c38e5ed),
	.w3(32'hbb497155),
	.w4(32'h3bcb6d09),
	.w5(32'h3a6f0d77),
	.w6(32'hbc9155ee),
	.w7(32'hbb4cdd06),
	.w8(32'hbbb93f3a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3ed5a),
	.w1(32'h3a8999df),
	.w2(32'hbafd794a),
	.w3(32'hbbe0b831),
	.w4(32'hbabc7f0f),
	.w5(32'h3cdfc57e),
	.w6(32'hbbb7d3cf),
	.w7(32'h3c13c3c1),
	.w8(32'hbc3d7319),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f56b4),
	.w1(32'h3c0762ea),
	.w2(32'h3aac8bc5),
	.w3(32'hbcc517dd),
	.w4(32'h3c1fc475),
	.w5(32'h3b02b254),
	.w6(32'h3cbe5345),
	.w7(32'h3a278312),
	.w8(32'hbbc95c15),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83221a),
	.w1(32'hbc405dc7),
	.w2(32'h3c6bacd4),
	.w3(32'hbca2e4c1),
	.w4(32'hbbcbb106),
	.w5(32'hbac3f2a4),
	.w6(32'hbb01b9b7),
	.w7(32'h3c6c3dec),
	.w8(32'h39fe0b0d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7c99),
	.w1(32'hbb2d0dfb),
	.w2(32'h3c304f49),
	.w3(32'hbaf9ef99),
	.w4(32'h3acc3505),
	.w5(32'hbc11a912),
	.w6(32'h3c2462ba),
	.w7(32'h3c378c02),
	.w8(32'h3a2fb6ad),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95edc),
	.w1(32'hbb5546c0),
	.w2(32'hbbe0a197),
	.w3(32'hbbd01e28),
	.w4(32'h3b875864),
	.w5(32'hbb1f2fa8),
	.w6(32'h3904cb49),
	.w7(32'hbd0b8e3b),
	.w8(32'h3b51c6b7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaaa7b),
	.w1(32'hbc48f147),
	.w2(32'h3b4d2aa1),
	.w3(32'h3a711963),
	.w4(32'hbbfa8115),
	.w5(32'h3b8fff29),
	.w6(32'hbc656ddc),
	.w7(32'hb9a5e970),
	.w8(32'h3be1697f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f3d0),
	.w1(32'hba884689),
	.w2(32'hbc374c8c),
	.w3(32'hbb632633),
	.w4(32'hb9852e74),
	.w5(32'h3a818ce1),
	.w6(32'h3ba339f6),
	.w7(32'hbb5297fd),
	.w8(32'hb923e5a9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc5a4),
	.w1(32'hbc200027),
	.w2(32'hbc9e29db),
	.w3(32'hbbcb1c40),
	.w4(32'hbbdc6072),
	.w5(32'hbbcb1456),
	.w6(32'hbb4da771),
	.w7(32'h3b85dc53),
	.w8(32'h3c59763d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098385),
	.w1(32'h3c54e2ae),
	.w2(32'h3a4cb909),
	.w3(32'hbbeadac5),
	.w4(32'hbc982850),
	.w5(32'hbc8d6e81),
	.w6(32'hbb885436),
	.w7(32'hbbdde230),
	.w8(32'h3d83adf0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01ca93),
	.w1(32'hbc259815),
	.w2(32'h3c026e48),
	.w3(32'hbba7ba10),
	.w4(32'hba98750c),
	.w5(32'hbbd18c09),
	.w6(32'h3d0526f8),
	.w7(32'h3cc6675d),
	.w8(32'h3afe7c61),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced6cdb),
	.w1(32'hba05d9a1),
	.w2(32'h3c8fa49e),
	.w3(32'hbbce72c5),
	.w4(32'h3b657161),
	.w5(32'hbb90b5c4),
	.w6(32'hbb36d2c0),
	.w7(32'hbc30ee8f),
	.w8(32'hbb6c9b05),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a362a),
	.w1(32'hbb987119),
	.w2(32'hbba579f9),
	.w3(32'h3ccac985),
	.w4(32'hbbc9bfd4),
	.w5(32'h3c4bf5da),
	.w6(32'h3c9e3b6b),
	.w7(32'h3c1f85a5),
	.w8(32'h3a9a73da),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a28d0),
	.w1(32'hbbbb6dbd),
	.w2(32'h3c08175d),
	.w3(32'hbb899ddc),
	.w4(32'hba328a11),
	.w5(32'hba046b81),
	.w6(32'h3ba7ff08),
	.w7(32'hbb21891d),
	.w8(32'h3aebb724),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e50c),
	.w1(32'h3c3f7508),
	.w2(32'hbb875af7),
	.w3(32'h3b5648f5),
	.w4(32'h3ab8e556),
	.w5(32'hba328d3e),
	.w6(32'hbc1f7a0c),
	.w7(32'h3be43283),
	.w8(32'hbc7217f2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164c16),
	.w1(32'hbc047161),
	.w2(32'hbbc9e0c9),
	.w3(32'hb9b49710),
	.w4(32'hbc288fef),
	.w5(32'h3a89c182),
	.w6(32'h3bd907a3),
	.w7(32'hbc1a0b4f),
	.w8(32'h3b188a35),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25c6b0),
	.w1(32'h3a96bbb0),
	.w2(32'h3bc67e35),
	.w3(32'h3b2aeee3),
	.w4(32'hbbf60cc6),
	.w5(32'h39bed9ce),
	.w6(32'h3accd039),
	.w7(32'h3b5eb7ec),
	.w8(32'hbc6e56a8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c883167),
	.w1(32'h3b6748bb),
	.w2(32'hba73ed8a),
	.w3(32'hbbd36c98),
	.w4(32'h3c012c3a),
	.w5(32'h3cb7a826),
	.w6(32'h3b9e424f),
	.w7(32'h3cbb16e9),
	.w8(32'h3b5587f9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896a1c),
	.w1(32'h3cb88b92),
	.w2(32'hba52014c),
	.w3(32'hbc3b2749),
	.w4(32'h3ae06bf8),
	.w5(32'h3bd68d89),
	.w6(32'hbcb7a0b0),
	.w7(32'hbc8517bd),
	.w8(32'h3c0afea7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58edd6),
	.w1(32'hbc51ec53),
	.w2(32'hbc2e2a92),
	.w3(32'h3bd76414),
	.w4(32'h3d2ac79b),
	.w5(32'hbbe16c82),
	.w6(32'hbc5f4dec),
	.w7(32'h3ca79bab),
	.w8(32'h3c290770),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc225548),
	.w1(32'hba207f83),
	.w2(32'h3a5fcf72),
	.w3(32'hbc6242be),
	.w4(32'hbaec6212),
	.w5(32'hbc687feb),
	.w6(32'h3c6c4511),
	.w7(32'h3b99ac6e),
	.w8(32'h3ad1c8a6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3aea),
	.w1(32'h3be628aa),
	.w2(32'hbc035175),
	.w3(32'hb99765d9),
	.w4(32'h3b82b4cf),
	.w5(32'hb9dc806d),
	.w6(32'h3a17579e),
	.w7(32'h3b0365d6),
	.w8(32'h3c17996d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4b751),
	.w1(32'h3b43476f),
	.w2(32'h3ca7baa7),
	.w3(32'h3ada4d1d),
	.w4(32'h3c052020),
	.w5(32'hbb2a3184),
	.w6(32'hbc5d8576),
	.w7(32'h3b330201),
	.w8(32'h3c831ef7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7520b8),
	.w1(32'h3bc409e6),
	.w2(32'h3ba9fb3d),
	.w3(32'hbbc64dfb),
	.w4(32'hbacbdfeb),
	.w5(32'h3a465b7b),
	.w6(32'h3b3b7939),
	.w7(32'h3c32ba41),
	.w8(32'h3bfaa465),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7fdd2),
	.w1(32'h3c5ce64f),
	.w2(32'hbbbdf23c),
	.w3(32'h3d0b8a42),
	.w4(32'hbb13da33),
	.w5(32'hbc885327),
	.w6(32'h3be7c201),
	.w7(32'h3b0cf8d9),
	.w8(32'h39588e69),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7464f),
	.w1(32'h3bd21b67),
	.w2(32'h3c3a36ef),
	.w3(32'hbc0a52bf),
	.w4(32'hbc0a64f7),
	.w5(32'h3b696d22),
	.w6(32'hbd493eb1),
	.w7(32'h39b23dcc),
	.w8(32'hbc01a40a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951053),
	.w1(32'h3c2abfdf),
	.w2(32'hbbbdcfa0),
	.w3(32'hbcad93e9),
	.w4(32'h3c0506bc),
	.w5(32'h3c304ccd),
	.w6(32'hbc2f8a26),
	.w7(32'hbadb3c0c),
	.w8(32'h3b18086f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab86e3d),
	.w1(32'h3b80be84),
	.w2(32'hbb65eb94),
	.w3(32'h3c8352cd),
	.w4(32'h3bfbed9b),
	.w5(32'h3bdd2c20),
	.w6(32'h3b24cd6c),
	.w7(32'h3bebce13),
	.w8(32'hbb7d7a7a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976d4a1),
	.w1(32'hbb1df36b),
	.w2(32'hbb268d96),
	.w3(32'hbca867e2),
	.w4(32'h3ba93a27),
	.w5(32'h3c1fd0f8),
	.w6(32'h3c0d116e),
	.w7(32'h3b88202b),
	.w8(32'h3acbaae8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d045),
	.w1(32'hbc02ac0f),
	.w2(32'hba865f5b),
	.w3(32'hba25beba),
	.w4(32'h3ac51583),
	.w5(32'hbb966e4b),
	.w6(32'h3bbc7b83),
	.w7(32'h3902efa7),
	.w8(32'hb9c0433e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082661),
	.w1(32'hbbecf662),
	.w2(32'h3b299c9d),
	.w3(32'hbc006ccc),
	.w4(32'hbc6c2f05),
	.w5(32'h3ab9ebff),
	.w6(32'h3bd687ab),
	.w7(32'h3c523e86),
	.w8(32'hbcd50af9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff68b),
	.w1(32'hbc5fe3e2),
	.w2(32'hbaf016dc),
	.w3(32'hbb551e9a),
	.w4(32'hbc805efe),
	.w5(32'hbc4ee0d9),
	.w6(32'h3beaba9f),
	.w7(32'hbbfd8b80),
	.w8(32'hbbbf8094),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b502295),
	.w1(32'h39b871e8),
	.w2(32'h3bd18ff9),
	.w3(32'h3be5d807),
	.w4(32'hbb2a463d),
	.w5(32'h3b0722db),
	.w6(32'h3b957941),
	.w7(32'hbc71c1ea),
	.w8(32'hbbfa3083),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4df7bf),
	.w1(32'hba9b2ad2),
	.w2(32'hb8350066),
	.w3(32'hbb9ce5ae),
	.w4(32'h3c01c8e4),
	.w5(32'hbc0500e4),
	.w6(32'h3c43cb8c),
	.w7(32'hbc13a09a),
	.w8(32'h3ab01537),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95cd69),
	.w1(32'hbb3b2637),
	.w2(32'h3a7f7c4f),
	.w3(32'h3b40c1d9),
	.w4(32'h3b0287ed),
	.w5(32'hbbf51b84),
	.w6(32'hbc294432),
	.w7(32'h3c1aba1e),
	.w8(32'h3c8ea502),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4613ab),
	.w1(32'hbd0a20da),
	.w2(32'hbbd20750),
	.w3(32'h3bab592e),
	.w4(32'hbc1277b2),
	.w5(32'hb9ddd5b8),
	.w6(32'h3b75ae84),
	.w7(32'h3c111a5a),
	.w8(32'hbb9dd039),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c74b),
	.w1(32'hbbf1009d),
	.w2(32'h3c09986a),
	.w3(32'hba052415),
	.w4(32'h3a9711f0),
	.w5(32'hbb8c93e3),
	.w6(32'hbb19c019),
	.w7(32'h3b8532c1),
	.w8(32'h3c576c00),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc849da2),
	.w1(32'hbc1baad5),
	.w2(32'hbbeddf78),
	.w3(32'h3b00d9c2),
	.w4(32'hbb4bafdc),
	.w5(32'h3b8220a4),
	.w6(32'h3aa09078),
	.w7(32'h3b9a9f74),
	.w8(32'h3c095f2b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8015a3),
	.w1(32'h3c18ab91),
	.w2(32'h3c383a25),
	.w3(32'h3bdebb8f),
	.w4(32'h3c6e3dbf),
	.w5(32'h3c9c02fb),
	.w6(32'hbb87027c),
	.w7(32'hbabb0fc4),
	.w8(32'hbc346e56),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24323f),
	.w1(32'hbca2e34a),
	.w2(32'hb9f19a87),
	.w3(32'h3c3c111d),
	.w4(32'h3bb1740a),
	.w5(32'hbc2e0d73),
	.w6(32'hbaad6952),
	.w7(32'hbbdc900b),
	.w8(32'hbb54ce6a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77e4c5),
	.w1(32'h3b322ba8),
	.w2(32'hbbb86e76),
	.w3(32'h3b8df445),
	.w4(32'hbb9abdaf),
	.w5(32'hbc85332f),
	.w6(32'h3c94096c),
	.w7(32'hba081e3a),
	.w8(32'h3cc20e56),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd40b2),
	.w1(32'hbd64b4a1),
	.w2(32'h3b140454),
	.w3(32'hbc275d5d),
	.w4(32'hbcdf82c7),
	.w5(32'h3b5bd0b3),
	.w6(32'h3cf27fec),
	.w7(32'h3c87c080),
	.w8(32'h3c9d4950),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d32f5),
	.w1(32'hbc800bcb),
	.w2(32'hbba0a260),
	.w3(32'h3ad569df),
	.w4(32'hba7669a9),
	.w5(32'hbb0d93c2),
	.w6(32'h3bf47a2b),
	.w7(32'h3c08682d),
	.w8(32'hbb3677a9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca5f01),
	.w1(32'h3c03b864),
	.w2(32'h3c22d403),
	.w3(32'hbbb2572a),
	.w4(32'hbb5dc67a),
	.w5(32'hbb00643d),
	.w6(32'hbc1cf3cb),
	.w7(32'h392de83f),
	.w8(32'hbc128267),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22199c),
	.w1(32'h3c4cf0e1),
	.w2(32'h3cb9dc53),
	.w3(32'hbbba25f7),
	.w4(32'hbb45d867),
	.w5(32'h3c409633),
	.w6(32'hbbf5c2f3),
	.w7(32'hbc6b5850),
	.w8(32'h3bf348b5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb17420),
	.w1(32'h3b836e26),
	.w2(32'h3b61320a),
	.w3(32'hbc1af6d6),
	.w4(32'h3a94c9d5),
	.w5(32'h3ba2a33e),
	.w6(32'hbb6a4649),
	.w7(32'hbbf687d8),
	.w8(32'hbaab33e9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e9f9),
	.w1(32'hbc51694c),
	.w2(32'hba9d38f1),
	.w3(32'hba192f21),
	.w4(32'hbbcd9ab8),
	.w5(32'hbbb7fc70),
	.w6(32'hbbb9d91a),
	.w7(32'h3d07b1dc),
	.w8(32'h3c36b8b3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29db71),
	.w1(32'h3bc1d9e3),
	.w2(32'h3c0a37b2),
	.w3(32'hbc9444d2),
	.w4(32'hbb149c53),
	.w5(32'hbc88e91a),
	.w6(32'hbbb502d6),
	.w7(32'hbc114669),
	.w8(32'hbabe5c9f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19ae8b),
	.w1(32'h3beccae7),
	.w2(32'h3b3149a3),
	.w3(32'h3c240211),
	.w4(32'h3baa3f03),
	.w5(32'hbca0c212),
	.w6(32'hbc129691),
	.w7(32'h3c084f15),
	.w8(32'hbb42920c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40bf32),
	.w1(32'h3cc06475),
	.w2(32'hbaa8d80b),
	.w3(32'h3c1e272c),
	.w4(32'h3aa7e40e),
	.w5(32'hbb6cb617),
	.w6(32'hbc180313),
	.w7(32'hbd197f77),
	.w8(32'hbbf7af85),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ad455),
	.w1(32'hbc7667c5),
	.w2(32'h3bd0271c),
	.w3(32'h3cafaae5),
	.w4(32'hbc46a0b5),
	.w5(32'hbbce6700),
	.w6(32'hbc199b95),
	.w7(32'hbc414934),
	.w8(32'hbca76fcb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e8f5),
	.w1(32'h3c86276d),
	.w2(32'h3c075e88),
	.w3(32'h3a47b268),
	.w4(32'hbc03837a),
	.w5(32'hbcb1b3d1),
	.w6(32'h3b3991e9),
	.w7(32'hbb2b5543),
	.w8(32'h3c4570c0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e40aa),
	.w1(32'h3b07db94),
	.w2(32'h3c6183a0),
	.w3(32'h3a827557),
	.w4(32'h3c0aa5f0),
	.w5(32'hbc0bc6b4),
	.w6(32'hbc0dd9b5),
	.w7(32'h3c8db887),
	.w8(32'h3cd5f1c8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6717b),
	.w1(32'hbd0997dd),
	.w2(32'hbc27ff9c),
	.w3(32'hbb3c8f64),
	.w4(32'hbc7b234a),
	.w5(32'h3c34793c),
	.w6(32'h3cca990f),
	.w7(32'hbc1e1824),
	.w8(32'h3b88eb69),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56bf87),
	.w1(32'hbc880ffd),
	.w2(32'hbbee3657),
	.w3(32'h3b3292c1),
	.w4(32'h38a33eb5),
	.w5(32'hbbb37324),
	.w6(32'h3c299321),
	.w7(32'h3b0b8ad5),
	.w8(32'h3ad83512),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba568f3),
	.w1(32'hbabf65b2),
	.w2(32'h3c8e2635),
	.w3(32'hbb3c422f),
	.w4(32'h3aee5485),
	.w5(32'h3baca610),
	.w6(32'hbb565f07),
	.w7(32'hbc8e6675),
	.w8(32'h3ad71566),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229194),
	.w1(32'hbc868a4e),
	.w2(32'h3b4b96ee),
	.w3(32'hbc594bb7),
	.w4(32'hbc10d1b2),
	.w5(32'hbc64a9ce),
	.w6(32'h3c5267da),
	.w7(32'h3b9a5764),
	.w8(32'hbc242c84),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae598e2),
	.w1(32'h3b6dc0dd),
	.w2(32'hbc490e29),
	.w3(32'h3cac82d9),
	.w4(32'hb9cb9b0c),
	.w5(32'h3b75782c),
	.w6(32'hbbb028f6),
	.w7(32'h3a0d7eb9),
	.w8(32'h3c75b9ab),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9af29f),
	.w1(32'hbbba95aa),
	.w2(32'hbbc94c1e),
	.w3(32'hbc3cbb6c),
	.w4(32'h3b329c6a),
	.w5(32'hbb2efd84),
	.w6(32'h3c4eb79f),
	.w7(32'h3c18ddbe),
	.w8(32'hb9fce5d8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5f79),
	.w1(32'h3984d2d3),
	.w2(32'h3b2b391a),
	.w3(32'hbc8188fb),
	.w4(32'h3ac6a8af),
	.w5(32'hbb39699c),
	.w6(32'hbc0649a8),
	.w7(32'hba9fe24d),
	.w8(32'h3b7e1bdd),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72cfa6),
	.w1(32'h3c0e0128),
	.w2(32'h3c9d6855),
	.w3(32'h3ad951c5),
	.w4(32'h3ae06806),
	.w5(32'hbc5e834c),
	.w6(32'hbc7ca146),
	.w7(32'hbb5ada60),
	.w8(32'hbaa95f15),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0f9f),
	.w1(32'hb7a30d9c),
	.w2(32'hbc0195cf),
	.w3(32'hbca332c9),
	.w4(32'h3c2a48ce),
	.w5(32'hbb0ad571),
	.w6(32'h3a443be0),
	.w7(32'h3c0f1557),
	.w8(32'hbb37958f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc45971),
	.w1(32'hbb667bcb),
	.w2(32'h3952ad7c),
	.w3(32'hbb9f39db),
	.w4(32'hbcb7ec61),
	.w5(32'hbc5f9aec),
	.w6(32'hbc51719b),
	.w7(32'hbc41bc8a),
	.w8(32'h3c6b3f7c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63af7f),
	.w1(32'hbc4af7ad),
	.w2(32'h3960a185),
	.w3(32'hbc81d7c7),
	.w4(32'hbb8b3a3f),
	.w5(32'h3b58ee03),
	.w6(32'hbd4118c6),
	.w7(32'h3b0f64a7),
	.w8(32'h3c8620ec),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb16211),
	.w1(32'h3c10a87a),
	.w2(32'hbcfe4143),
	.w3(32'hbb06bb2d),
	.w4(32'hbc4a6813),
	.w5(32'hbb97699f),
	.w6(32'hbb8c17ec),
	.w7(32'h3b53f9fa),
	.w8(32'hbc819d56),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ea9a1),
	.w1(32'hbcde1bae),
	.w2(32'h3ac2c77a),
	.w3(32'h3b89ef6b),
	.w4(32'hbb8f7ed9),
	.w5(32'hba6a0721),
	.w6(32'h3894c5ea),
	.w7(32'hbba327a1),
	.w8(32'h3ac1a864),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c179c7f),
	.w1(32'hbcae3080),
	.w2(32'hbd02de69),
	.w3(32'h3b9fadac),
	.w4(32'hbb845ad2),
	.w5(32'h3be773da),
	.w6(32'h3a7f1bd7),
	.w7(32'hbb4a7404),
	.w8(32'hbc03929d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c285),
	.w1(32'hbb46eb5d),
	.w2(32'hbbd598be),
	.w3(32'hbb371c2e),
	.w4(32'h3b89c9b4),
	.w5(32'hbca6e8fe),
	.w6(32'h3c2f4b4d),
	.w7(32'h3c08dbe9),
	.w8(32'h3a726818),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c661bf3),
	.w1(32'h3bf4b0ea),
	.w2(32'h3c39555b),
	.w3(32'h3afced2c),
	.w4(32'hbc85030f),
	.w5(32'h3c0f9bcb),
	.w6(32'hbb6a6838),
	.w7(32'h3c3b5e56),
	.w8(32'h3b1a66fd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57b999),
	.w1(32'hbbe99d8f),
	.w2(32'hbc771d0b),
	.w3(32'hbbc85c46),
	.w4(32'hbb89879d),
	.w5(32'h3c00fb04),
	.w6(32'h3c967999),
	.w7(32'hbae6b616),
	.w8(32'hbc1d7e43),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1fe07),
	.w1(32'h3c12e9bb),
	.w2(32'h39d2c3aa),
	.w3(32'h3c524505),
	.w4(32'h3c0ccb51),
	.w5(32'h3c60f5b3),
	.w6(32'hbbaaaa3f),
	.w7(32'h3c911850),
	.w8(32'h3d7f391a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba685782),
	.w1(32'hbae7cc05),
	.w2(32'h3c016222),
	.w3(32'hba0477fc),
	.w4(32'h3b861608),
	.w5(32'hbbb21237),
	.w6(32'h3b6cc712),
	.w7(32'h3bc3025a),
	.w8(32'hbbac1c49),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a8db),
	.w1(32'hbcc07879),
	.w2(32'h3bc60c43),
	.w3(32'hbb92bd90),
	.w4(32'hbc0f4e4c),
	.w5(32'h3c1340a8),
	.w6(32'hbc5dcaad),
	.w7(32'h3c5018f2),
	.w8(32'hbb2b7bb0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c252ddd),
	.w1(32'hbc25b814),
	.w2(32'h3d26966d),
	.w3(32'h3cc4be2b),
	.w4(32'h3c21e523),
	.w5(32'hbc4239a5),
	.w6(32'h3b63b8ea),
	.w7(32'hbbd6d714),
	.w8(32'hbd1c70de),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7ba4),
	.w1(32'hbc9585f2),
	.w2(32'h3d2ee7bb),
	.w3(32'hbbd321a1),
	.w4(32'h3c722547),
	.w5(32'hbc637aa0),
	.w6(32'h3b46c5b9),
	.w7(32'hbc317c9c),
	.w8(32'h3c6c4939),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058a3e),
	.w1(32'h3c238696),
	.w2(32'h3bf6458e),
	.w3(32'h3b87c5a4),
	.w4(32'hbb67f58f),
	.w5(32'hbab3aee2),
	.w6(32'h3a27a607),
	.w7(32'hbba73746),
	.w8(32'h3c6bf1e7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7a149),
	.w1(32'hbd2629c0),
	.w2(32'hb794554a),
	.w3(32'hbc73771a),
	.w4(32'hb95d0e15),
	.w5(32'h3a45910a),
	.w6(32'h3b97835f),
	.w7(32'hbc7876af),
	.w8(32'h3c7b2b71),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab2756),
	.w1(32'h3c59c466),
	.w2(32'hbbc7e78d),
	.w3(32'hbbc4880b),
	.w4(32'h3bde0718),
	.w5(32'h3c6bbe6d),
	.w6(32'hbb366313),
	.w7(32'h3bb37e6a),
	.w8(32'hbb7bae5a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5cdc),
	.w1(32'h3bf94c7b),
	.w2(32'h3c53c8a7),
	.w3(32'hbc58be18),
	.w4(32'h3b12ac7c),
	.w5(32'h3c82d35c),
	.w6(32'hbc63e41c),
	.w7(32'h3c880b2f),
	.w8(32'h3ba902c5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule