module layer_8_featuremap_152(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45d2f9),
	.w1(32'h3c17ff0f),
	.w2(32'h3ba582b0),
	.w3(32'hbc0c703f),
	.w4(32'hbb5929e4),
	.w5(32'hbb12593d),
	.w6(32'hbc3ef733),
	.w7(32'hbbadc178),
	.w8(32'h3a8b33cd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba338a5),
	.w1(32'hba5a68ab),
	.w2(32'hbb090ad1),
	.w3(32'hbb828731),
	.w4(32'hbadc3d5b),
	.w5(32'hbb0d9431),
	.w6(32'hbb0f30d5),
	.w7(32'h3963e4e3),
	.w8(32'hba429f47),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10011e),
	.w1(32'h3b407339),
	.w2(32'h3b3cdbba),
	.w3(32'hbb3c23ec),
	.w4(32'h3abcb072),
	.w5(32'h399d2b72),
	.w6(32'hbb24c1eb),
	.w7(32'h3b1395e3),
	.w8(32'h3a028887),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3066f3),
	.w1(32'hbbc6ccc8),
	.w2(32'hbcb17d07),
	.w3(32'hbc6229fa),
	.w4(32'hbc2bc507),
	.w5(32'hbcd2f52d),
	.w6(32'hbc889e9f),
	.w7(32'hbc334e08),
	.w8(32'hbc67d8d6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc224f80),
	.w1(32'hbb769fe3),
	.w2(32'hbb87e7e0),
	.w3(32'hbc0b30c9),
	.w4(32'hbad5ef87),
	.w5(32'hbb0afe0e),
	.w6(32'hbbe46e80),
	.w7(32'hbabd2cfc),
	.w8(32'hbb53c308),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb849c),
	.w1(32'h3c2567a2),
	.w2(32'h3c19733f),
	.w3(32'hbc1f98d7),
	.w4(32'h3cb6056a),
	.w5(32'h3c56a10f),
	.w6(32'hbbfadff2),
	.w7(32'h3c69497b),
	.w8(32'h3b8acf92),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b8c4d),
	.w1(32'h37cdf206),
	.w2(32'h38ccee25),
	.w3(32'h3997071d),
	.w4(32'hb7c2aed8),
	.w5(32'h38234440),
	.w6(32'h399793b0),
	.w7(32'h37fadc34),
	.w8(32'h38555411),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f42b50),
	.w1(32'h3bc3098e),
	.w2(32'h3bc11726),
	.w3(32'hbc28c3df),
	.w4(32'hbb59f428),
	.w5(32'hbb547ace),
	.w6(32'hbab512dd),
	.w7(32'h3bd25069),
	.w8(32'h3b428aa7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58ffd2),
	.w1(32'hba369ed8),
	.w2(32'hb99be630),
	.w3(32'hbb12ada0),
	.w4(32'hbb14112a),
	.w5(32'hbb3cac6b),
	.w6(32'hbacc99e3),
	.w7(32'h3a08c2f0),
	.w8(32'h39eb3ead),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd1843),
	.w1(32'h3b8993ca),
	.w2(32'h3b659874),
	.w3(32'hbbed3137),
	.w4(32'hb9903084),
	.w5(32'hbb071803),
	.w6(32'hbc8c4670),
	.w7(32'hbbb0d7d7),
	.w8(32'hbbb8c108),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c01d),
	.w1(32'h3bde5689),
	.w2(32'h396206da),
	.w3(32'hbc611434),
	.w4(32'hbbf59be7),
	.w5(32'hbc23bca4),
	.w6(32'hbbe3e7e6),
	.w7(32'h3b4d984b),
	.w8(32'h3b221080),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e50d5),
	.w1(32'hba9a2111),
	.w2(32'hba8f62e9),
	.w3(32'hbc53a984),
	.w4(32'hbb4d2992),
	.w5(32'hb993ed50),
	.w6(32'hbca3848c),
	.w7(32'hb98fa9b9),
	.w8(32'h3abf8e4f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33f257),
	.w1(32'h3a525782),
	.w2(32'h39c873b3),
	.w3(32'hbc19519d),
	.w4(32'h3afc022f),
	.w5(32'hb9fe392c),
	.w6(32'hbc25319a),
	.w7(32'h3b219f43),
	.w8(32'hbbb973d1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e2f8c),
	.w1(32'h3aa596cf),
	.w2(32'h3bad534c),
	.w3(32'h3b57f8e8),
	.w4(32'h3b21a7e5),
	.w5(32'h3b32d45f),
	.w6(32'hba333bb6),
	.w7(32'h3b942723),
	.w8(32'h3b62ccbd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6a3c1),
	.w1(32'h3bdd533b),
	.w2(32'h3bcc3206),
	.w3(32'h3bc49a24),
	.w4(32'h3a8b8d77),
	.w5(32'h3b91dc8f),
	.w6(32'h3bc2d5c9),
	.w7(32'h3b77dcbb),
	.w8(32'h3bd48e5f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc138f),
	.w1(32'h3bc324f5),
	.w2(32'hbb8d4fae),
	.w3(32'h3bd2c3b5),
	.w4(32'hbbc7a9fa),
	.w5(32'hbba25a0b),
	.w6(32'h3bb79cce),
	.w7(32'hbb98ea08),
	.w8(32'hbc3bb4d8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4ce94),
	.w1(32'hbb99c1ea),
	.w2(32'h3bf09719),
	.w3(32'hbb9339bc),
	.w4(32'h3b53e4b1),
	.w5(32'h3c0f6f8c),
	.w6(32'hbbbf2a79),
	.w7(32'h3ae88dba),
	.w8(32'h3c00b3a4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc552e2e),
	.w1(32'hbb5e1f1b),
	.w2(32'hbb9549ae),
	.w3(32'hbc4812b0),
	.w4(32'hbbd66d14),
	.w5(32'hbc53a4b3),
	.w6(32'hbc7e7c39),
	.w7(32'hbbf6caec),
	.w8(32'h3b38faa8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77d8c8),
	.w1(32'h3cc5a5c2),
	.w2(32'h3c6605da),
	.w3(32'hbd287b29),
	.w4(32'hbc44f2e6),
	.w5(32'hbc982cf6),
	.w6(32'hbd071f9f),
	.w7(32'hbab0af9c),
	.w8(32'h3b9b2e32),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2a73a7),
	.w1(32'hbb6e17ba),
	.w2(32'h3af4420d),
	.w3(32'hbd27d31d),
	.w4(32'hbbe487d0),
	.w5(32'hbc974053),
	.w6(32'hbd473fef),
	.w7(32'hbc1730d9),
	.w8(32'hbcc2b698),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6930c9),
	.w1(32'h3b58f99b),
	.w2(32'h3a56409c),
	.w3(32'hbcae0c29),
	.w4(32'h3c0d92b2),
	.w5(32'h3c7ecdee),
	.w6(32'hbcb6e73b),
	.w7(32'h3bda7943),
	.w8(32'h3c85e9c5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe0d8d),
	.w1(32'hbb31d585),
	.w2(32'hbbdf8c5f),
	.w3(32'hba2cbbda),
	.w4(32'h3bbf4e40),
	.w5(32'h3bc3451f),
	.w6(32'h3b81c029),
	.w7(32'hba6d45d9),
	.w8(32'h39a16119),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8edc1f),
	.w1(32'h3c509875),
	.w2(32'h3cc04176),
	.w3(32'hbc461282),
	.w4(32'hbc1ca885),
	.w5(32'hbc13986c),
	.w6(32'hbbcff884),
	.w7(32'h3a5823fd),
	.w8(32'h3c3a0077),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0da99b),
	.w1(32'hbaaaf5f5),
	.w2(32'h3c14187d),
	.w3(32'hbc2c9418),
	.w4(32'h3c1b343f),
	.w5(32'hbad190fb),
	.w6(32'hbc89d19e),
	.w7(32'h3c3d62d1),
	.w8(32'h3a867480),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483965),
	.w1(32'hbaad8c09),
	.w2(32'h3b15b366),
	.w3(32'h39574881),
	.w4(32'h3c16e799),
	.w5(32'hbac31464),
	.w6(32'h3a276508),
	.w7(32'h3bab983e),
	.w8(32'hbb5c0e9c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50d4b2),
	.w1(32'h3c6d4917),
	.w2(32'h3c63283c),
	.w3(32'hbca0b2ef),
	.w4(32'h3c36932b),
	.w5(32'h3cfa6700),
	.w6(32'hbc3d0b34),
	.w7(32'h3cf8b4ef),
	.w8(32'h3d354265),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9aee),
	.w1(32'hbc7f27f1),
	.w2(32'h3b6289d2),
	.w3(32'h3aeccd38),
	.w4(32'hbc15b753),
	.w5(32'hbc2af0d7),
	.w6(32'h3c1d2423),
	.w7(32'h3c1be5e3),
	.w8(32'h3c2cb6ff),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6334f),
	.w1(32'h3d739ee7),
	.w2(32'h3d912710),
	.w3(32'hbd86c4f4),
	.w4(32'h3c97f48e),
	.w5(32'h3c51b3b7),
	.w6(32'hbd94e9a4),
	.w7(32'h3d073353),
	.w8(32'h3d484739),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73fbbf),
	.w1(32'h3bf84d79),
	.w2(32'h3afe1f51),
	.w3(32'hbcd24323),
	.w4(32'hbbac9d07),
	.w5(32'h3c0b8b73),
	.w6(32'hbc4865b9),
	.w7(32'hbbe07b80),
	.w8(32'h3bb7f68f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd84741),
	.w1(32'hbb871588),
	.w2(32'hbb0205ed),
	.w3(32'hbb3cd0a8),
	.w4(32'hbd0fccc7),
	.w5(32'hbcc742c0),
	.w6(32'hba680a42),
	.w7(32'hba2ef89e),
	.w8(32'hbb23ff5e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c795835),
	.w1(32'h3c37f5bd),
	.w2(32'h3bc4ad3f),
	.w3(32'hbc050a53),
	.w4(32'hbb4ae0e4),
	.w5(32'h3b3681c5),
	.w6(32'h3b69a0e3),
	.w7(32'h3b24ba5b),
	.w8(32'h3bdd4289),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55c29a),
	.w1(32'h3c493412),
	.w2(32'hba141a61),
	.w3(32'hbb252361),
	.w4(32'h3c00ecf8),
	.w5(32'hbbb69cb4),
	.w6(32'h3b47c271),
	.w7(32'hbb753a8f),
	.w8(32'hbc6804f1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfda3cb),
	.w1(32'hbbd35a51),
	.w2(32'hbca7fa03),
	.w3(32'hbbcffaaf),
	.w4(32'hbd02c143),
	.w5(32'hbc83419d),
	.w6(32'hbc6314c6),
	.w7(32'hbc848ba9),
	.w8(32'hbc2e705d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb701d0),
	.w1(32'hbbbb4d80),
	.w2(32'hb848715f),
	.w3(32'h3c280886),
	.w4(32'h3c161662),
	.w5(32'h3c2fc799),
	.w6(32'h3a94df7a),
	.w7(32'h3a8a7611),
	.w8(32'h3b7bf461),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba6858),
	.w1(32'hbc35e610),
	.w2(32'h3b03cfbc),
	.w3(32'hb96e44f3),
	.w4(32'h3c568b69),
	.w5(32'h3a787343),
	.w6(32'hbbf7d0a6),
	.w7(32'h3c466119),
	.w8(32'hbb39a74d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1cd65),
	.w1(32'h3c5a47a0),
	.w2(32'hb9af0222),
	.w3(32'hbbe330ed),
	.w4(32'hbd115d63),
	.w5(32'hbc370008),
	.w6(32'hbabc2723),
	.w7(32'hbcb0301f),
	.w8(32'hbc128254),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc06ca8),
	.w1(32'h3a9ddf6a),
	.w2(32'hbb31fb45),
	.w3(32'h3bec17e5),
	.w4(32'hbbf74068),
	.w5(32'hbc77485c),
	.w6(32'h3b872ac7),
	.w7(32'h3b10ce61),
	.w8(32'hba2b185f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412b06),
	.w1(32'hbbe7b6d7),
	.w2(32'hbbc1bb2f),
	.w3(32'hbc6ff733),
	.w4(32'hbb3700b8),
	.w5(32'hbb8b2d4b),
	.w6(32'hbb3fc4ae),
	.w7(32'hbb921bb5),
	.w8(32'hbbab99d5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0eed4),
	.w1(32'h3c290618),
	.w2(32'hbadd77f7),
	.w3(32'h3b5bc9c4),
	.w4(32'hbafc35b3),
	.w5(32'h3b42d108),
	.w6(32'h3c23ac12),
	.w7(32'hbc1e31b1),
	.w8(32'hbc26999f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4274),
	.w1(32'hbc3ed303),
	.w2(32'hbace576e),
	.w3(32'h3b242778),
	.w4(32'hbbca5eec),
	.w5(32'hbbb59b23),
	.w6(32'hbb741914),
	.w7(32'hbc612ac2),
	.w8(32'hbc7fe90f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9ae4fe),
	.w1(32'h3b38d67b),
	.w2(32'hbb8513b4),
	.w3(32'hbdbf4fb4),
	.w4(32'hbc9bf17e),
	.w5(32'hbc8f629d),
	.w6(32'hbdd2506e),
	.w7(32'hbb971a48),
	.w8(32'h3bd6c80c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb087110),
	.w1(32'h3c4728a9),
	.w2(32'h3bd584de),
	.w3(32'hbc224e15),
	.w4(32'hbb9b7f9e),
	.w5(32'h3a94437e),
	.w6(32'hbbb52bf6),
	.w7(32'h3c4bd9ea),
	.w8(32'h3c6c7367),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accbbc4),
	.w1(32'hbacc4d8f),
	.w2(32'h3ba0600e),
	.w3(32'hbcac25e3),
	.w4(32'hbc036e86),
	.w5(32'hbc12f1be),
	.w6(32'hbc047b65),
	.w7(32'hbc0a2c09),
	.w8(32'hbc24f30c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc881a06),
	.w1(32'h3c249007),
	.w2(32'h3c55045b),
	.w3(32'hbc060ef3),
	.w4(32'hba8ec555),
	.w5(32'h3a13e64b),
	.w6(32'hba9c47a8),
	.w7(32'h3bf69cb8),
	.w8(32'h3b5acecf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e89a9),
	.w1(32'h3c8db9c2),
	.w2(32'h3c9ab391),
	.w3(32'hbca447ab),
	.w4(32'hbc5c9fc3),
	.w5(32'hbbbaafe2),
	.w6(32'hbc1b4edf),
	.w7(32'h3af045a6),
	.w8(32'h3c27156d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c312cfe),
	.w1(32'h3cb977b5),
	.w2(32'h3c00498c),
	.w3(32'hbacb2e55),
	.w4(32'hbbadb208),
	.w5(32'hbaba27ae),
	.w6(32'h3b44280f),
	.w7(32'h3b8dc762),
	.w8(32'h3c3ade63),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80ce40),
	.w1(32'h3a8595aa),
	.w2(32'h3c1ca211),
	.w3(32'hbb9da56f),
	.w4(32'hbb26a5e4),
	.w5(32'h3bca5acd),
	.w6(32'h3a669612),
	.w7(32'h3b74080e),
	.w8(32'h3c5aa714),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf5bac4),
	.w1(32'h3ca19f4a),
	.w2(32'h3c7d84b4),
	.w3(32'hbbb5a9fb),
	.w4(32'hbc485c88),
	.w5(32'hbc088076),
	.w6(32'h3c0c504b),
	.w7(32'h3b6df7e7),
	.w8(32'h3c2ee351),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd516a),
	.w1(32'h3c8c4c9f),
	.w2(32'hbb8d3027),
	.w3(32'hba12b428),
	.w4(32'h3a0f7952),
	.w5(32'h3a39bbfc),
	.w6(32'hbb3bef5c),
	.w7(32'h3b934e0c),
	.w8(32'h3b9eacc6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8de884),
	.w1(32'hbc8bc9ca),
	.w2(32'hbc130868),
	.w3(32'hbca6af14),
	.w4(32'hbc89f252),
	.w5(32'hbcfefb3c),
	.w6(32'hbce2be81),
	.w7(32'hbc6fb7e9),
	.w8(32'hbcb5822e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d07d8),
	.w1(32'hbc7ae661),
	.w2(32'hbc4751fa),
	.w3(32'hbca4c8cf),
	.w4(32'h3c2c7998),
	.w5(32'h3ba454a4),
	.w6(32'hbce15cd0),
	.w7(32'h3c99233d),
	.w8(32'h3c407094),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd5906),
	.w1(32'h3d1a046e),
	.w2(32'h3ce1646a),
	.w3(32'hbd865577),
	.w4(32'h3c60ee2e),
	.w5(32'h3c6065e6),
	.w6(32'hbd1f7516),
	.w7(32'h3cc16da3),
	.w8(32'h3d3f2f4a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa31668),
	.w1(32'h3c039532),
	.w2(32'h3b71c2a1),
	.w3(32'hbb2678ef),
	.w4(32'hba4807b4),
	.w5(32'hbbc2207d),
	.w6(32'h3bea809c),
	.w7(32'hbaba1df8),
	.w8(32'hbc449177),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba482294),
	.w1(32'h3c14e420),
	.w2(32'h3c0c908f),
	.w3(32'hbc5dbe1f),
	.w4(32'hbb9b8ea8),
	.w5(32'h3ae06d5e),
	.w6(32'hbcd8d827),
	.w7(32'hbc638682),
	.w8(32'hbbd9fd7b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99234f),
	.w1(32'h3b0b68c7),
	.w2(32'hbb875e64),
	.w3(32'h3b259d94),
	.w4(32'hbbaf9d26),
	.w5(32'hba5f7aad),
	.w6(32'h3a0a9317),
	.w7(32'h3bec1119),
	.w8(32'h3bfb2611),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03466e),
	.w1(32'h3cbbb993),
	.w2(32'h3bc68093),
	.w3(32'hbc89c3fb),
	.w4(32'hbb8e660e),
	.w5(32'hbbac76d6),
	.w6(32'h3a70bd47),
	.w7(32'h3bdf7da8),
	.w8(32'hbb934072),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc845993),
	.w1(32'hbb3a21db),
	.w2(32'hb9c40b51),
	.w3(32'hbbd2bfca),
	.w4(32'h3a536d22),
	.w5(32'hbb904113),
	.w6(32'hbc34df3a),
	.w7(32'hbc47018d),
	.w8(32'hbc4fd46a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc387cd7),
	.w1(32'h3c390ed6),
	.w2(32'h3cbbcc33),
	.w3(32'hbcd9d826),
	.w4(32'h3c317583),
	.w5(32'h3c684de3),
	.w6(32'hbce4418d),
	.w7(32'h3c21a601),
	.w8(32'h3d03a7bf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e6504),
	.w1(32'h3d0cc079),
	.w2(32'h3c828dec),
	.w3(32'hbb2b8721),
	.w4(32'hbb3865a1),
	.w5(32'hbb11d37b),
	.w6(32'h3c901985),
	.w7(32'h3bfa7d41),
	.w8(32'h3bab4d50),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54b93b),
	.w1(32'hbaef5b00),
	.w2(32'hbbcdf4a2),
	.w3(32'hbc712b80),
	.w4(32'h3b464bb4),
	.w5(32'hbb983e9c),
	.w6(32'hbc74d882),
	.w7(32'hbba204de),
	.w8(32'hba0fbb75),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7000f2),
	.w1(32'hbcaf5122),
	.w2(32'hbb38207a),
	.w3(32'hbba81152),
	.w4(32'hbbdffca9),
	.w5(32'hbc19f614),
	.w6(32'hbbb9af8d),
	.w7(32'hbbff82eb),
	.w8(32'hbb97e338),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba118c69),
	.w1(32'h3a993bbb),
	.w2(32'h3bf69931),
	.w3(32'hbb7b6ef9),
	.w4(32'h3aceadbe),
	.w5(32'hbbd263c2),
	.w6(32'h3b0c25fe),
	.w7(32'h3a436b0d),
	.w8(32'hbbf7ab6c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd240afa),
	.w1(32'h3c750112),
	.w2(32'hbc267dda),
	.w3(32'hbd1bba0f),
	.w4(32'hbb156029),
	.w5(32'h3b8ddde1),
	.w6(32'hbd2211bc),
	.w7(32'h3bfbe68b),
	.w8(32'h3c95eb72),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008eb7),
	.w1(32'h3a569ead),
	.w2(32'h3bdad6f0),
	.w3(32'hbbe465c7),
	.w4(32'hbb395360),
	.w5(32'hbbb5ec21),
	.w6(32'hbbf143bb),
	.w7(32'hbbff5800),
	.w8(32'hbc189ec8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62d257),
	.w1(32'hba4547e6),
	.w2(32'h3bfbeaa1),
	.w3(32'h3b133a62),
	.w4(32'h3ba51d0b),
	.w5(32'h3bbfbc61),
	.w6(32'hbbae9e43),
	.w7(32'h3b61c6fb),
	.w8(32'h3c1252b5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7992),
	.w1(32'h3c3c94a4),
	.w2(32'h3c3c79c3),
	.w3(32'hbc005b4f),
	.w4(32'h3baa08ad),
	.w5(32'hbc0e19d3),
	.w6(32'hbb77af20),
	.w7(32'h3b8a8ff5),
	.w8(32'hbbddae23),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf98f6),
	.w1(32'h3c0c4937),
	.w2(32'hbabb3ec1),
	.w3(32'hbbbd0595),
	.w4(32'h3bdd978c),
	.w5(32'hbbad5c89),
	.w6(32'hbb638355),
	.w7(32'h3c552278),
	.w8(32'hba06d76e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c0deb),
	.w1(32'hb97e4f16),
	.w2(32'hbae2bfec),
	.w3(32'hbc7ef96e),
	.w4(32'h3bd943a5),
	.w5(32'h3b360012),
	.w6(32'hbc9cf3ae),
	.w7(32'h3c024712),
	.w8(32'h3b3a3eb0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8782dc),
	.w1(32'hbc2ba1cb),
	.w2(32'hbc7398ad),
	.w3(32'h3ae29f97),
	.w4(32'hbb9e6af5),
	.w5(32'hbb9b5d3b),
	.w6(32'h3b78bf7a),
	.w7(32'hbb030475),
	.w8(32'hbc3585e7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad2def),
	.w1(32'h3b4985b7),
	.w2(32'h3c972049),
	.w3(32'hbd655832),
	.w4(32'hbcae45e2),
	.w5(32'hbca80394),
	.w6(32'hbcbfc88e),
	.w7(32'h3c1d8211),
	.w8(32'h3c9fd6be),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9222f3),
	.w1(32'h3bb99119),
	.w2(32'hbbb0622f),
	.w3(32'hbbbc7e0c),
	.w4(32'h3bd0e55a),
	.w5(32'h3a5e28ee),
	.w6(32'h3ab34aad),
	.w7(32'hbbc45e83),
	.w8(32'hbc296f27),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bdd18),
	.w1(32'hbb80daa9),
	.w2(32'hbb0f11c8),
	.w3(32'hbcf70567),
	.w4(32'hbc5d09cb),
	.w5(32'hbc11b59f),
	.w6(32'hbcf50d8f),
	.w7(32'hbbaaf7f2),
	.w8(32'h3bf8ced3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d52c3),
	.w1(32'h3b280b79),
	.w2(32'h3a5cd6e6),
	.w3(32'h3bc1fa83),
	.w4(32'hbb97e161),
	.w5(32'hbbc22e50),
	.w6(32'h3bbb8477),
	.w7(32'h3a834526),
	.w8(32'h3a139b72),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52b0b),
	.w1(32'h3b197416),
	.w2(32'hbcac8e79),
	.w3(32'hbc85e39c),
	.w4(32'hbc58559d),
	.w5(32'hbb7437f1),
	.w6(32'hbc8ba0c7),
	.w7(32'hbc3524a8),
	.w8(32'hbc00037e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45ff4b),
	.w1(32'h3c58168f),
	.w2(32'h3c090d7c),
	.w3(32'hbb551751),
	.w4(32'hbc4db28f),
	.w5(32'hbc7a9344),
	.w6(32'hbb274dad),
	.w7(32'h3bd6d6de),
	.w8(32'h3b958fe2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22ba89),
	.w1(32'h3b151f3a),
	.w2(32'hbbf21667),
	.w3(32'hbc890065),
	.w4(32'hbbfc42b4),
	.w5(32'hbba311a5),
	.w6(32'hbbac6e8e),
	.w7(32'hbbb1c4e6),
	.w8(32'hbad17c90),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc209ffd),
	.w1(32'hbc25338d),
	.w2(32'h3af40fb0),
	.w3(32'hbb7a58cd),
	.w4(32'h3aa9ff86),
	.w5(32'h3b202828),
	.w6(32'hbc26bf71),
	.w7(32'h3ae42a7d),
	.w8(32'h3b7de371),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0ab8),
	.w1(32'h3c34b205),
	.w2(32'h3b6c6273),
	.w3(32'hbce06a10),
	.w4(32'hbbdbb6d5),
	.w5(32'hbb51b46a),
	.w6(32'hbc36ae87),
	.w7(32'h3bf708d1),
	.w8(32'h3c44f79f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d87c),
	.w1(32'h3b17215e),
	.w2(32'h3b309c39),
	.w3(32'hbc4e4b63),
	.w4(32'hbb5f3388),
	.w5(32'hbc034a7a),
	.w6(32'hbc59ffca),
	.w7(32'hbc2d5484),
	.w8(32'hbc69b7a6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ee22),
	.w1(32'hbc63c1f5),
	.w2(32'h3aa20d62),
	.w3(32'hbc6d69b2),
	.w4(32'h3b900777),
	.w5(32'hbb656c1b),
	.w6(32'hbc7f6898),
	.w7(32'h3ba1bd07),
	.w8(32'hbb479f4d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02030a),
	.w1(32'h3ac59a27),
	.w2(32'hba52e665),
	.w3(32'hba85cd61),
	.w4(32'hbc1772d0),
	.w5(32'hbb824587),
	.w6(32'hba52ab8d),
	.w7(32'hbb9eae91),
	.w8(32'hbb877998),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1898e2),
	.w1(32'h3c2951d0),
	.w2(32'h3c96b79a),
	.w3(32'hbb996d89),
	.w4(32'h3bf444b7),
	.w5(32'hbae3e0a0),
	.w6(32'hbc003949),
	.w7(32'h3bec6c2a),
	.w8(32'h391ac3b0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1e9ee),
	.w1(32'h3be1990a),
	.w2(32'h3bcc7420),
	.w3(32'hbd1f5375),
	.w4(32'hbc07e3f4),
	.w5(32'hbc108165),
	.w6(32'hbcff9ef3),
	.w7(32'h3be449c9),
	.w8(32'h3bf79966),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd95780),
	.w1(32'hbcb5926b),
	.w2(32'hbcc8178a),
	.w3(32'hbdbea9b6),
	.w4(32'hbc17ea48),
	.w5(32'hbca19f1a),
	.w6(32'hbdbe9dfe),
	.w7(32'hbcadd676),
	.w8(32'hba87f9fe),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc777570),
	.w1(32'h3cc5d96a),
	.w2(32'h3cb7243c),
	.w3(32'hbd6e7571),
	.w4(32'hbbabd884),
	.w5(32'hbaa9cb9b),
	.w6(32'hbd4af483),
	.w7(32'h3c28161d),
	.w8(32'h3cbe28b9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7f90),
	.w1(32'hbc0b0540),
	.w2(32'h3c009ec8),
	.w3(32'hbc6bd1ab),
	.w4(32'hbc858d47),
	.w5(32'hbc6c9383),
	.w6(32'hbc988a14),
	.w7(32'hbc05f279),
	.w8(32'hba7cb91d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb8d0d),
	.w1(32'h3b3e574c),
	.w2(32'hbcc58f61),
	.w3(32'h3bf09bea),
	.w4(32'hbcf48152),
	.w5(32'hbce585b5),
	.w6(32'h3c026716),
	.w7(32'hbcf04b56),
	.w8(32'hbd08e287),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4b80a),
	.w1(32'hbc9365e9),
	.w2(32'hba2aad2d),
	.w3(32'hbc9067f2),
	.w4(32'hbb3979a7),
	.w5(32'h3b136204),
	.w6(32'hbcb48ca4),
	.w7(32'hba4715b0),
	.w8(32'h3b600b21),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8527e),
	.w1(32'h3c1f8f99),
	.w2(32'hbb48865a),
	.w3(32'h3c1c1169),
	.w4(32'hb9e0b033),
	.w5(32'hbb5473b9),
	.w6(32'h3c1eb46f),
	.w7(32'hba8eb795),
	.w8(32'hbb8af791),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8e283),
	.w1(32'hbae3cda2),
	.w2(32'h3c27e147),
	.w3(32'hbb485936),
	.w4(32'h3a788099),
	.w5(32'h3be57acc),
	.w6(32'h3aeae19a),
	.w7(32'h3c3a2b7a),
	.w8(32'h3c9bb099),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84fedd),
	.w1(32'hbba34d40),
	.w2(32'h3bf22b61),
	.w3(32'hbbd25781),
	.w4(32'h3bba5025),
	.w5(32'hbb00fb3c),
	.w6(32'hbb784e92),
	.w7(32'h3c012811),
	.w8(32'h3b81942e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2d62f),
	.w1(32'h3bbe9a86),
	.w2(32'h3bc433f2),
	.w3(32'h3b2a6d2e),
	.w4(32'h3b5bdffa),
	.w5(32'h3b75f3c0),
	.w6(32'h3b82f8d3),
	.w7(32'h3bfe2340),
	.w8(32'h3c4297f7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf100de),
	.w1(32'h3c336e67),
	.w2(32'hbac3f915),
	.w3(32'hbce26a61),
	.w4(32'hbc1e9429),
	.w5(32'hbc43dd4e),
	.w6(32'hbc784e3b),
	.w7(32'hbb4f9078),
	.w8(32'h3b9714de),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf639be),
	.w1(32'h3a9eb233),
	.w2(32'h3c5512da),
	.w3(32'hbc90f016),
	.w4(32'hbb41cd5c),
	.w5(32'hb949b98d),
	.w6(32'hbc8650f4),
	.w7(32'h3b6ca2bb),
	.w8(32'hba4b7dd7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aea8e),
	.w1(32'h3b958488),
	.w2(32'hbc1c2e52),
	.w3(32'hbc6ef512),
	.w4(32'hbba1d969),
	.w5(32'hbbea0aae),
	.w6(32'hbcc0e5bb),
	.w7(32'hbbb9f3f3),
	.w8(32'hbc0d1ef4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cfbd4),
	.w1(32'h3bdb9242),
	.w2(32'h3becc3cd),
	.w3(32'hbc8e09f7),
	.w4(32'h3c637f60),
	.w5(32'hbb69e764),
	.w6(32'hbc5d43e5),
	.w7(32'h3bbce046),
	.w8(32'hbbd933f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d626c),
	.w1(32'hbc53093f),
	.w2(32'h3bc94fae),
	.w3(32'hbd1ef5ef),
	.w4(32'hba15e53e),
	.w5(32'h3bea90df),
	.w6(32'hbd171276),
	.w7(32'h3c0dc372),
	.w8(32'h3c373489),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac54a8e),
	.w1(32'hbbc7fa3d),
	.w2(32'hbb8793ef),
	.w3(32'h3aa0d550),
	.w4(32'h3b3fe643),
	.w5(32'hbb8a669a),
	.w6(32'hbb214448),
	.w7(32'hbb09a33b),
	.w8(32'hbbaa6a3f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaee5d4),
	.w1(32'hbbce2ee9),
	.w2(32'h3d44705d),
	.w3(32'h3a52e94b),
	.w4(32'h3d5a6b3a),
	.w5(32'h3bd54c5c),
	.w6(32'hbbbd6134),
	.w7(32'h3d486b3c),
	.w8(32'h3b45befa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a500),
	.w1(32'hbb72bdf9),
	.w2(32'h3bd052c2),
	.w3(32'hbb262193),
	.w4(32'hbb054b8d),
	.w5(32'hbb8d6488),
	.w6(32'hbbd087ac),
	.w7(32'hbb45d748),
	.w8(32'hbba0595b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888720),
	.w1(32'hbc69fe9c),
	.w2(32'h38de63d1),
	.w3(32'hbb5ba54f),
	.w4(32'hba84cd78),
	.w5(32'hbabf22bf),
	.w6(32'hbbcaa432),
	.w7(32'h39ea0f5d),
	.w8(32'hbb38e5de),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba724b32),
	.w1(32'hbb978e02),
	.w2(32'hbafa8cd6),
	.w3(32'hbaf2f4cc),
	.w4(32'h3ac01434),
	.w5(32'hbc00eb39),
	.w6(32'hbb90ecb8),
	.w7(32'hba7dde93),
	.w8(32'hbc3ea98c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc04c1),
	.w1(32'h3bc8bd72),
	.w2(32'h3c683b6f),
	.w3(32'h3c06062b),
	.w4(32'h3bb455cf),
	.w5(32'hbc403386),
	.w6(32'h3be1429b),
	.w7(32'h3bd6ed3e),
	.w8(32'hbc1e76d3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f7a12),
	.w1(32'h3bdc3a09),
	.w2(32'h3bd4bb31),
	.w3(32'hbc832e76),
	.w4(32'h3af3fc82),
	.w5(32'hbb12df54),
	.w6(32'hbcb25047),
	.w7(32'hbb5e365b),
	.w8(32'hbb90df43),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8879),
	.w1(32'h39ec6e4c),
	.w2(32'hbb15bb44),
	.w3(32'hb9eace1b),
	.w4(32'h3c0d71d2),
	.w5(32'hbbf09a81),
	.w6(32'hbb9998cf),
	.w7(32'h3bb55b96),
	.w8(32'hbbf85489),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39954288),
	.w1(32'h3c627bfd),
	.w2(32'h3c9e7183),
	.w3(32'hbcf90314),
	.w4(32'h3af19473),
	.w5(32'hbc99dc44),
	.w6(32'hbc6b5b6e),
	.w7(32'h3c8fc683),
	.w8(32'h39628674),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc19c3c),
	.w1(32'hbb3d375d),
	.w2(32'h3c77e890),
	.w3(32'hbc609a59),
	.w4(32'hbc002ba7),
	.w5(32'h3ad99d82),
	.w6(32'hbc8077d0),
	.w7(32'h399e2656),
	.w8(32'hbbcc1285),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c759),
	.w1(32'hbba7f3dc),
	.w2(32'hb8ff3a2e),
	.w3(32'hbb2eea3b),
	.w4(32'h3be7b141),
	.w5(32'h3b09e7e1),
	.w6(32'hbc8292b6),
	.w7(32'h3be091d9),
	.w8(32'h3b55ecc2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af08524),
	.w1(32'h3aa332fe),
	.w2(32'hbc21266b),
	.w3(32'hbb5e4f7c),
	.w4(32'hbbbb5462),
	.w5(32'hbc398537),
	.w6(32'hb8d3c346),
	.w7(32'hbc0f6c59),
	.w8(32'hbc1f1613),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02dde8),
	.w1(32'hbbb8ad81),
	.w2(32'h3c55b25e),
	.w3(32'h3ac60ca7),
	.w4(32'h3bd1a319),
	.w5(32'hbbf1f755),
	.w6(32'hb9b40723),
	.w7(32'h3b143ad9),
	.w8(32'hbb84ad7d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb17047),
	.w1(32'hba1b79ec),
	.w2(32'h3bd96a0f),
	.w3(32'hbcb4b929),
	.w4(32'h3b92b55b),
	.w5(32'h3b2d815c),
	.w6(32'hbcdc6a51),
	.w7(32'h3b615287),
	.w8(32'h3a0234e3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98dd40),
	.w1(32'hbbbd77af),
	.w2(32'hbc5148a0),
	.w3(32'hbcf258b2),
	.w4(32'hbc09a4ee),
	.w5(32'hba71f0c9),
	.w6(32'hbcc76364),
	.w7(32'hbbf023a5),
	.w8(32'h3be4c171),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a4859),
	.w1(32'hbbacbbc9),
	.w2(32'hbc74636e),
	.w3(32'hbbc158fe),
	.w4(32'h3bf6ee56),
	.w5(32'hbc3fd55a),
	.w6(32'hbc00b878),
	.w7(32'h3be8a68b),
	.w8(32'hbc947ae0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0705f4),
	.w1(32'hbbc67c4d),
	.w2(32'hbc96c683),
	.w3(32'hbbb7c264),
	.w4(32'hbc90cae0),
	.w5(32'hbc841766),
	.w6(32'hbba99a1f),
	.w7(32'hbc85bc25),
	.w8(32'hbc4ca126),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc309cb7),
	.w1(32'hbb2a9b58),
	.w2(32'h39ccb3e6),
	.w3(32'hbb9500f2),
	.w4(32'h3bb7c5f8),
	.w5(32'hbb3dd669),
	.w6(32'h39ffede0),
	.w7(32'h3a4a4190),
	.w8(32'hbb47da30),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56f4eb),
	.w1(32'h3c10b5eb),
	.w2(32'hbc241d38),
	.w3(32'h3bf5e356),
	.w4(32'hbc1e0579),
	.w5(32'h3b56a696),
	.w6(32'hbbad3ae2),
	.w7(32'hbc399a3e),
	.w8(32'hbb04ba6c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3758ff),
	.w1(32'h3b524f02),
	.w2(32'hbad71f57),
	.w3(32'hbbd27aed),
	.w4(32'h3baddd63),
	.w5(32'h3b7072db),
	.w6(32'hbbf9c09b),
	.w7(32'h3ba6c1ab),
	.w8(32'h3b557b8f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f3daf),
	.w1(32'h3c4a1009),
	.w2(32'h3bd1682f),
	.w3(32'hbc4e89e3),
	.w4(32'h3b398758),
	.w5(32'h3b19765c),
	.w6(32'hbbcb670c),
	.w7(32'h3c27c0c4),
	.w8(32'h3c01c2c6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b797d),
	.w1(32'h3a00ba0b),
	.w2(32'h3bf7d4c8),
	.w3(32'h3a476aea),
	.w4(32'h3aefea4a),
	.w5(32'h3b2a9b27),
	.w6(32'h3b039473),
	.w7(32'h3b6caeb2),
	.w8(32'hbab323e0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b899e67),
	.w1(32'hbb5b65bf),
	.w2(32'hb72ea0a8),
	.w3(32'hbb9fc52c),
	.w4(32'hbb21b112),
	.w5(32'hbbb2099e),
	.w6(32'hbb75f0a2),
	.w7(32'hbb5d31ef),
	.w8(32'hbbe51da5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26f31),
	.w1(32'h3b8c4e9e),
	.w2(32'hba99c930),
	.w3(32'hbc43c203),
	.w4(32'hbbaa42eb),
	.w5(32'hbc3cc460),
	.w6(32'hbcb08cdb),
	.w7(32'hbc66710b),
	.w8(32'hbbeb457c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257723),
	.w1(32'hbc417a7b),
	.w2(32'h3c2447e1),
	.w3(32'hbc4b4bb3),
	.w4(32'hbc49b147),
	.w5(32'hbb2feafc),
	.w6(32'hbc0f769d),
	.w7(32'hbbb8bfa3),
	.w8(32'hbb4fc834),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04d58a),
	.w1(32'h3b5b4301),
	.w2(32'h3a85fd6d),
	.w3(32'hbb8fd01c),
	.w4(32'h3ae9e7e9),
	.w5(32'h3b4b0031),
	.w6(32'hbc0c6649),
	.w7(32'h39c317b6),
	.w8(32'h3b889da5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd67a3a),
	.w1(32'h3b429618),
	.w2(32'hbb88b287),
	.w3(32'h3b017f52),
	.w4(32'h3c662fb4),
	.w5(32'h3cae7430),
	.w6(32'h3b31e98f),
	.w7(32'hb91d3686),
	.w8(32'h3c4c48eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833192),
	.w1(32'hbbbc69f8),
	.w2(32'h3b996427),
	.w3(32'h3bea60ce),
	.w4(32'h3c04d478),
	.w5(32'hbbe3fa69),
	.w6(32'h3c616dc4),
	.w7(32'hbbc7773b),
	.w8(32'hbc01c613),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b455122),
	.w1(32'h3aa39343),
	.w2(32'hba578fa5),
	.w3(32'h3b785fca),
	.w4(32'hbb3874c8),
	.w5(32'hbb5c6563),
	.w6(32'h3a8d6f9b),
	.w7(32'hbb438853),
	.w8(32'h3b4faa49),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78d6a3),
	.w1(32'h3be545af),
	.w2(32'hbb944e30),
	.w3(32'hb8841797),
	.w4(32'hbba2bb47),
	.w5(32'hbbb76307),
	.w6(32'hbb0f2370),
	.w7(32'hbb4e056f),
	.w8(32'hbc6f5ca6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a87f),
	.w1(32'hba99ad85),
	.w2(32'h3c2941c6),
	.w3(32'hbc848178),
	.w4(32'hba8b6a56),
	.w5(32'h3aa8bd71),
	.w6(32'hbb66b173),
	.w7(32'h3b76f31d),
	.w8(32'h3bc6b42c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule