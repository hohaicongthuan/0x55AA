module layer_6_featuremap_75(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a68e),
	.w1(32'hbadc02c2),
	.w2(32'h3a9ac987),
	.w3(32'hbb83846f),
	.w4(32'h3b0f293c),
	.w5(32'h3b158bda),
	.w6(32'hbb9feb2b),
	.w7(32'h399544c8),
	.w8(32'hb849abec),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c783b),
	.w1(32'h3c9a4807),
	.w2(32'h3c961a91),
	.w3(32'h3c3b86d4),
	.w4(32'h3c1cf555),
	.w5(32'h3c378387),
	.w6(32'h3ced427b),
	.w7(32'h3cedc6b1),
	.w8(32'h3d11d2c9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67c2ea),
	.w1(32'h3cab9e69),
	.w2(32'h3bede444),
	.w3(32'h3cabb36d),
	.w4(32'h3d03f86e),
	.w5(32'h3c93949d),
	.w6(32'h3cf939ec),
	.w7(32'hbab88866),
	.w8(32'hbab1b366),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99ec9f),
	.w1(32'h3ad62b78),
	.w2(32'h38119337),
	.w3(32'h3b95035c),
	.w4(32'h3b5b2e13),
	.w5(32'hba7390b5),
	.w6(32'h3bbaac78),
	.w7(32'h3b199fb8),
	.w8(32'h393eace6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c291),
	.w1(32'hbbd8192c),
	.w2(32'h3aa7654d),
	.w3(32'h3ba92c92),
	.w4(32'h37f19c1f),
	.w5(32'hbbeeec20),
	.w6(32'h3b3b9bb2),
	.w7(32'hbad7a474),
	.w8(32'hbbc68eac),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2a5ca),
	.w1(32'h3b0e3e0f),
	.w2(32'h3c015c00),
	.w3(32'hbbc0aad5),
	.w4(32'h39dcb91e),
	.w5(32'h3aeb51fa),
	.w6(32'hbb2a904a),
	.w7(32'h3b2c1b4f),
	.w8(32'h3b790a13),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83182d),
	.w1(32'hbbe28631),
	.w2(32'hb9e03f79),
	.w3(32'hbc2ce597),
	.w4(32'hbbfd6154),
	.w5(32'hbb9c1002),
	.w6(32'hbb6ce1ef),
	.w7(32'h3ab0d328),
	.w8(32'h3b55ab86),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5193),
	.w1(32'h3ce076d4),
	.w2(32'h3cebfa31),
	.w3(32'hbc5520ee),
	.w4(32'hbc153f35),
	.w5(32'hbb8fa2c8),
	.w6(32'h3c24457c),
	.w7(32'h3c257539),
	.w8(32'h3c6b902a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc073f0),
	.w1(32'hba738be0),
	.w2(32'h3bfe17cf),
	.w3(32'hbb6d00e2),
	.w4(32'h3b196854),
	.w5(32'h3bc9a096),
	.w6(32'h3c1e8c72),
	.w7(32'hbb5b64c2),
	.w8(32'h3b6d7143),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a069),
	.w1(32'h3b82527e),
	.w2(32'h3bc2d533),
	.w3(32'hbb73dd63),
	.w4(32'h3b87698d),
	.w5(32'h39155c98),
	.w6(32'h3b3f93e1),
	.w7(32'h3bcb5760),
	.w8(32'hb7935aff),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1587c5),
	.w1(32'hbcf17d76),
	.w2(32'hbd0b1388),
	.w3(32'hbc9253f6),
	.w4(32'hbca5ac85),
	.w5(32'hbca2eb08),
	.w6(32'hbd2b0c6c),
	.w7(32'hbd6e52b6),
	.w8(32'hbd42c21f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfd62b),
	.w1(32'h3caafdca),
	.w2(32'h3c8e72c1),
	.w3(32'hbbb63456),
	.w4(32'hbc0b1f28),
	.w5(32'hbb15f00b),
	.w6(32'h3c2eef66),
	.w7(32'h3c02b01e),
	.w8(32'h3b99198e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439a0e),
	.w1(32'hbb26008d),
	.w2(32'h3c7884bb),
	.w3(32'hba75c1b6),
	.w4(32'h3c5e949b),
	.w5(32'hbba7dc7a),
	.w6(32'h38f89cd9),
	.w7(32'h3c910de6),
	.w8(32'hb9ef4c32),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0409f5),
	.w1(32'h3c03e1c1),
	.w2(32'h3c9e5c58),
	.w3(32'h3c8aad3e),
	.w4(32'h3ce1c5c6),
	.w5(32'h3c7ec9bb),
	.w6(32'h3c9c290c),
	.w7(32'h3ccdef7c),
	.w8(32'h3c8ce57f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc82226),
	.w1(32'h3c0aecbc),
	.w2(32'h3b2fb233),
	.w3(32'h3b41c1bd),
	.w4(32'h3b7f6405),
	.w5(32'hba133297),
	.w6(32'h3a405630),
	.w7(32'hbb01af22),
	.w8(32'hbba50f17),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babae20),
	.w1(32'h3bc7d2a1),
	.w2(32'h3bc77e81),
	.w3(32'hbb80d364),
	.w4(32'hbabdcff5),
	.w5(32'h3b222cd5),
	.w6(32'h3a213ec6),
	.w7(32'h3bc00e79),
	.w8(32'h3c00ea13),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dfafd),
	.w1(32'hbd28c97a),
	.w2(32'hbd64cde8),
	.w3(32'hbd8124dc),
	.w4(32'hbda71e0d),
	.w5(32'hbd46afed),
	.w6(32'hbdbdedf2),
	.w7(32'hbde0c6ed),
	.w8(32'hbd9e13f3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa44c6),
	.w1(32'hbb9d6510),
	.w2(32'hbb20b31a),
	.w3(32'hbbd1730f),
	.w4(32'hbac9f8be),
	.w5(32'hb9d3c7a0),
	.w6(32'hbb872622),
	.w7(32'h3a7f3690),
	.w8(32'h3a88dbd0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31401),
	.w1(32'h3bafe65c),
	.w2(32'h3b916c3c),
	.w3(32'h3af12fc5),
	.w4(32'hbb33db58),
	.w5(32'hbb976731),
	.w6(32'h3bc9b410),
	.w7(32'h3b57c1c1),
	.w8(32'hbaf0eeb0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ae47e),
	.w1(32'hbc1d1f40),
	.w2(32'hbb9897f6),
	.w3(32'h3ae32cad),
	.w4(32'h3c39175f),
	.w5(32'h3c0bbc69),
	.w6(32'hbc6d13c0),
	.w7(32'hbc0b9cca),
	.w8(32'hbb3b2d28),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe01a31),
	.w1(32'h3b20372f),
	.w2(32'h3ad4cbac),
	.w3(32'h3afea734),
	.w4(32'hba38b25b),
	.w5(32'hbb1d0041),
	.w6(32'h3aca5f5d),
	.w7(32'hba0c331d),
	.w8(32'h38f2b75e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958456),
	.w1(32'h3c873a4b),
	.w2(32'h3b2e1757),
	.w3(32'h3ba2d968),
	.w4(32'h3b7ed059),
	.w5(32'h3958539a),
	.w6(32'h3bcf250d),
	.w7(32'hbc151ae3),
	.w8(32'hbbf81be4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0302),
	.w1(32'hbb750145),
	.w2(32'h3a6248fe),
	.w3(32'h3bdffd5f),
	.w4(32'h3c2b5b95),
	.w5(32'h3c391019),
	.w6(32'h3a4e15c6),
	.w7(32'hbc0daf2c),
	.w8(32'h3c4a779c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d8cd),
	.w1(32'h3bef478d),
	.w2(32'h3b02d4f0),
	.w3(32'h3c4df157),
	.w4(32'h3d05312f),
	.w5(32'h3c38de23),
	.w6(32'h3b3ad4a2),
	.w7(32'hbabd0b5c),
	.w8(32'hb97f18ff),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c694357),
	.w1(32'h3c5d87b4),
	.w2(32'h3cb727cd),
	.w3(32'h3cb5c22b),
	.w4(32'hba39d5de),
	.w5(32'hbad09cd6),
	.w6(32'h3d1fc5b4),
	.w7(32'h3cb49686),
	.w8(32'h3c5e5312),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d255515),
	.w1(32'hbbd2861d),
	.w2(32'hbc501425),
	.w3(32'h3a5d9727),
	.w4(32'h3bdf2c40),
	.w5(32'h3c556f81),
	.w6(32'hbb99829f),
	.w7(32'hbc6f813e),
	.w8(32'hbc409ef8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d69bf),
	.w1(32'h3bf9bd91),
	.w2(32'h3c5c8781),
	.w3(32'hb910713c),
	.w4(32'h3b177b55),
	.w5(32'h3b47fff2),
	.w6(32'h3c98a381),
	.w7(32'h3cbd9fcb),
	.w8(32'h3c954055),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9b298),
	.w1(32'h3a922691),
	.w2(32'h3b9609eb),
	.w3(32'hba3461c7),
	.w4(32'hba51db2b),
	.w5(32'hba45829b),
	.w6(32'h3adbabdd),
	.w7(32'h3b56ef19),
	.w8(32'h38b09f0f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2398e),
	.w1(32'h3b0f7f00),
	.w2(32'hbb5f5a7a),
	.w3(32'hba9fce9a),
	.w4(32'hbbacea51),
	.w5(32'h39e49de6),
	.w6(32'hbb08088e),
	.w7(32'hbbc8d7f0),
	.w8(32'hba7d6690),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34a63b),
	.w1(32'h3be1fbd8),
	.w2(32'h3c670ebf),
	.w3(32'h3cb52983),
	.w4(32'h3c8003e2),
	.w5(32'h3c674582),
	.w6(32'h3c501e3b),
	.w7(32'h3b72d3ce),
	.w8(32'h3ca0806f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d6c7d),
	.w1(32'h3c2e1cc6),
	.w2(32'h3bcdaef1),
	.w3(32'h3bcedf92),
	.w4(32'hbbc29f12),
	.w5(32'hbbcdea13),
	.w6(32'h3c27edbd),
	.w7(32'hba281226),
	.w8(32'hbbe4070a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5368),
	.w1(32'hbc8b6ff8),
	.w2(32'hbc88309a),
	.w3(32'hbbc0a5f2),
	.w4(32'h3c33a325),
	.w5(32'h3b713695),
	.w6(32'hbc2e3601),
	.w7(32'hbc030256),
	.w8(32'hbae3b61e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc824b5),
	.w1(32'hbbfbb82f),
	.w2(32'hbbbc3b94),
	.w3(32'hb9cfe78f),
	.w4(32'h3c14f0e1),
	.w5(32'h3b1f8d10),
	.w6(32'hbca75128),
	.w7(32'hbcda15fe),
	.w8(32'hbbf77f13),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0454a),
	.w1(32'hbcedf083),
	.w2(32'hbd112866),
	.w3(32'hbccce9a8),
	.w4(32'hbc3ee15f),
	.w5(32'hbc0d9df5),
	.w6(32'hbd3b2596),
	.w7(32'hbd43fcd8),
	.w8(32'hbd1b5ad0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9a192),
	.w1(32'h3b5b8daf),
	.w2(32'h3b763ab2),
	.w3(32'h3b10ae47),
	.w4(32'h3b914680),
	.w5(32'h3c01306d),
	.w6(32'hba8ad167),
	.w7(32'h3b03032a),
	.w8(32'h3bbf40cf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a24c6),
	.w1(32'h3c381140),
	.w2(32'h3bd8e3fd),
	.w3(32'h3a7eb692),
	.w4(32'hbb952e72),
	.w5(32'h3a0f1446),
	.w6(32'h3bde09eb),
	.w7(32'h3b48b6c0),
	.w8(32'hbbf6a726),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1599df),
	.w1(32'h3b0b67d8),
	.w2(32'h3b66bcbc),
	.w3(32'h3bb6c15f),
	.w4(32'h3c1da06c),
	.w5(32'h3bb0f39e),
	.w6(32'h3ae1b232),
	.w7(32'h3c043d72),
	.w8(32'h3aa6553e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa3b05),
	.w1(32'hbba3821d),
	.w2(32'hbb95da36),
	.w3(32'hbb716294),
	.w4(32'hbb74875c),
	.w5(32'h3b7d0c07),
	.w6(32'hbbbdcc12),
	.w7(32'hbb939022),
	.w8(32'h3b0b7a12),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf82b1),
	.w1(32'h3cd28f77),
	.w2(32'h3cb65bfa),
	.w3(32'hbc300e61),
	.w4(32'h3c3a2152),
	.w5(32'h3ca3d8c9),
	.w6(32'h3ca821b1),
	.w7(32'h3ce8a932),
	.w8(32'h3ccb3286),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1345df),
	.w1(32'h3cfb67f3),
	.w2(32'h3cde6a3c),
	.w3(32'hbbf72cf9),
	.w4(32'h3b13fa03),
	.w5(32'h3c8b14c6),
	.w6(32'hbbc49ef7),
	.w7(32'h3a5d65d4),
	.w8(32'h3bc76b5e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f9b54),
	.w1(32'h3a8d3037),
	.w2(32'h3bd2194e),
	.w3(32'h3ad99801),
	.w4(32'h3c15c529),
	.w5(32'h3c4e874b),
	.w6(32'hbc3a31c6),
	.w7(32'hba975e1d),
	.w8(32'h3b14ed9d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0db1f0),
	.w1(32'h3b8c88f5),
	.w2(32'h3bd04489),
	.w3(32'h3b30ac7a),
	.w4(32'h3bd944bc),
	.w5(32'h3be25fbf),
	.w6(32'h3a1913e9),
	.w7(32'h3ba70b92),
	.w8(32'h3bd9fb82),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32888f),
	.w1(32'hbbefe7f5),
	.w2(32'hbb4ca70b),
	.w3(32'hbb902597),
	.w4(32'h3b9d4fae),
	.w5(32'h3ae9f61f),
	.w6(32'hbc4618c2),
	.w7(32'hbbce9e0e),
	.w8(32'hbb6f8ef5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a74d18),
	.w1(32'h3cbfe7fd),
	.w2(32'h3c9edf3e),
	.w3(32'h3cbc250f),
	.w4(32'h3ce3062c),
	.w5(32'h3ccd3444),
	.w6(32'h3d1b28bf),
	.w7(32'h3d24751b),
	.w8(32'h3d0b8669),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae3646),
	.w1(32'h3c5c3a77),
	.w2(32'h3c28bf34),
	.w3(32'h3ba0027f),
	.w4(32'h3c1b0232),
	.w5(32'h3c144060),
	.w6(32'h3aaecc5d),
	.w7(32'h3bc0b27b),
	.w8(32'h3bb939d0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc287de),
	.w1(32'h3cc98321),
	.w2(32'h3c331c75),
	.w3(32'h3c05f10d),
	.w4(32'h3cff0274),
	.w5(32'h3d06712b),
	.w6(32'h3b036b87),
	.w7(32'hba2ec946),
	.w8(32'h3c99c03f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f1d02),
	.w1(32'h3c8ebf29),
	.w2(32'h3cbf3fa3),
	.w3(32'h3b879bb5),
	.w4(32'h3b426ceb),
	.w5(32'hbc3176a4),
	.w6(32'h3c3c09a1),
	.w7(32'h3cab3a97),
	.w8(32'h3a9801ce),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb361106),
	.w1(32'hbdb59bac),
	.w2(32'hbdbfafd3),
	.w3(32'hbd45edaa),
	.w4(32'hbd819fcc),
	.w5(32'hbd05b142),
	.w6(32'hbdcdd8f8),
	.w7(32'hbe08caab),
	.w8(32'hbd9304a4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01663c),
	.w1(32'h3c3584d5),
	.w2(32'h3c51ee95),
	.w3(32'h3b5a964c),
	.w4(32'h3b94c61f),
	.w5(32'h3b9e4bdb),
	.w6(32'hbad9805a),
	.w7(32'h3ad42826),
	.w8(32'h3ae1c9a9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb617d),
	.w1(32'hbcd9dcbc),
	.w2(32'hbcb39493),
	.w3(32'hbad4ef6c),
	.w4(32'hbc29c841),
	.w5(32'hbc6db988),
	.w6(32'hbc6ab9e6),
	.w7(32'hbc98109e),
	.w8(32'hbca76eca),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f489),
	.w1(32'hba3f8605),
	.w2(32'h3b1e0711),
	.w3(32'hbad176c4),
	.w4(32'hbab6f8e4),
	.w5(32'hbbed1d8c),
	.w6(32'h3ad0ba5e),
	.w7(32'h3ac8f78f),
	.w8(32'hbb87548e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b9d71),
	.w1(32'h3c33f4fd),
	.w2(32'h3c3663a4),
	.w3(32'h3bf207e6),
	.w4(32'h3c486997),
	.w5(32'h3c3365af),
	.w6(32'h3b50b84f),
	.w7(32'h3c246f4e),
	.w8(32'h3ba5506d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70430e),
	.w1(32'h3c1acdcb),
	.w2(32'h3c22e380),
	.w3(32'hbb1d1504),
	.w4(32'hba94f285),
	.w5(32'hbb75c289),
	.w6(32'hbb012243),
	.w7(32'hbb14ad20),
	.w8(32'hbb831f86),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21f988),
	.w1(32'hb9fe65c4),
	.w2(32'h3c366420),
	.w3(32'hbc93150b),
	.w4(32'hbbdf316b),
	.w5(32'h3b625149),
	.w6(32'hbca5fcd4),
	.w7(32'hbc2169f5),
	.w8(32'h3c0e0a47),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8202b3),
	.w1(32'h3bbe54b8),
	.w2(32'h3c204ad3),
	.w3(32'h3bb583a3),
	.w4(32'h3c3f56c4),
	.w5(32'h3bff8f6a),
	.w6(32'h3c22720b),
	.w7(32'h3c7033c7),
	.w8(32'h3c363167),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ba86a),
	.w1(32'hbc327df1),
	.w2(32'hbc46bab2),
	.w3(32'hb9dd5529),
	.w4(32'hbc0ef246),
	.w5(32'h3a580721),
	.w6(32'hbb04f71c),
	.w7(32'hbc2bade0),
	.w8(32'hbbd603be),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17a7c),
	.w1(32'hbd100ca7),
	.w2(32'hbd1226f0),
	.w3(32'hbd2a3083),
	.w4(32'hbd289f63),
	.w5(32'hbd13e19e),
	.w6(32'hbd3f3d72),
	.w7(32'hbd400fb8),
	.w8(32'hbd23f43d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16761e),
	.w1(32'h3bc60d65),
	.w2(32'h3bb9983b),
	.w3(32'h3ad87288),
	.w4(32'h3ba2cf30),
	.w5(32'hbafdcabd),
	.w6(32'h3bb05a09),
	.w7(32'h3c06086e),
	.w8(32'h3bfbda34),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a304),
	.w1(32'h3c2776d4),
	.w2(32'h3c790280),
	.w3(32'h3c36830f),
	.w4(32'h3c6fecb1),
	.w5(32'h3c41c4e1),
	.w6(32'h3c395faa),
	.w7(32'h3c901ae7),
	.w8(32'h3c81e82c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fbda4),
	.w1(32'h3970df66),
	.w2(32'hbb18141a),
	.w3(32'h3c66553f),
	.w4(32'h3bb4113c),
	.w5(32'h3b4ba410),
	.w6(32'h3c0128dc),
	.w7(32'h3abe3ced),
	.w8(32'hbb60781e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eb94f),
	.w1(32'h3c1ee057),
	.w2(32'h3c9c869a),
	.w3(32'h3c39aee2),
	.w4(32'h3ca22833),
	.w5(32'h3c780d4d),
	.w6(32'h3c83ea8d),
	.w7(32'h3cc14ba5),
	.w8(32'h3ca1d2d6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf9093),
	.w1(32'h3ae3a76b),
	.w2(32'h3b4254e1),
	.w3(32'hbaffc909),
	.w4(32'hbb56c951),
	.w5(32'hbc13af83),
	.w6(32'hbaae3dd3),
	.w7(32'hbbf4a4d5),
	.w8(32'hbbc2a0ce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e144a),
	.w1(32'h3c476130),
	.w2(32'h3c7f4eb9),
	.w3(32'h3d1283c9),
	.w4(32'h3c1acda2),
	.w5(32'h3b9ea696),
	.w6(32'h3ca62dc1),
	.w7(32'h3be37ba7),
	.w8(32'h3c67f972),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ffb4),
	.w1(32'hbd3007e7),
	.w2(32'hbd3c7e4f),
	.w3(32'hbd3a3345),
	.w4(32'hbd368345),
	.w5(32'hbd0bdaa4),
	.w6(32'hbd66a906),
	.w7(32'hbd73341e),
	.w8(32'hbd443fe2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule