module layer_8_featuremap_149(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2d8f),
	.w1(32'h391de8e8),
	.w2(32'h3a83bd08),
	.w3(32'h3bdce339),
	.w4(32'h3ae6e1c7),
	.w5(32'hb9008ab8),
	.w6(32'h3bd1f078),
	.w7(32'h3b75f079),
	.w8(32'h3aa40fe1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac286e5),
	.w1(32'h3b04626a),
	.w2(32'h3a489125),
	.w3(32'h3accb88f),
	.w4(32'h3a05082a),
	.w5(32'h3a5e83d8),
	.w6(32'h3b108ee2),
	.w7(32'h3aa80f0e),
	.w8(32'h3a860eba),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba7807),
	.w1(32'h3b26029d),
	.w2(32'h3b35581e),
	.w3(32'hba4ad4da),
	.w4(32'hba2417f5),
	.w5(32'h3a0b43b0),
	.w6(32'hbb5ae0fb),
	.w7(32'hbabfbba4),
	.w8(32'h39b62d7d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff5aa2),
	.w1(32'h3a6ac19c),
	.w2(32'h3ae43a90),
	.w3(32'hba1c28d7),
	.w4(32'hbaab1d52),
	.w5(32'hbaa1484f),
	.w6(32'h39cf65f3),
	.w7(32'hb96e2a6e),
	.w8(32'hba89cc9c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096b1b),
	.w1(32'h3a63aa80),
	.w2(32'h39fb5941),
	.w3(32'h3ad6ff75),
	.w4(32'h38d7c50e),
	.w5(32'hba48b87d),
	.w6(32'h3b83e576),
	.w7(32'h3b1da0fe),
	.w8(32'h3a15a3f2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a450686),
	.w1(32'h3b63697f),
	.w2(32'h38fb505e),
	.w3(32'hba5679d8),
	.w4(32'h3b473e8c),
	.w5(32'h39ac30ae),
	.w6(32'hbb8cf194),
	.w7(32'hbadca1a5),
	.w8(32'hbb8f90b0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f2350b),
	.w1(32'hb7ba8e2c),
	.w2(32'hb74f771c),
	.w3(32'h379502ea),
	.w4(32'hb7ad4e25),
	.w5(32'hb78a1374),
	.w6(32'h37b7b212),
	.w7(32'hb69a1745),
	.w8(32'hb74fbb3a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913c4d),
	.w1(32'h3a76ff7e),
	.w2(32'h3b26c8bb),
	.w3(32'hbadae6d4),
	.w4(32'hbb9c7176),
	.w5(32'hbaa3252b),
	.w6(32'h3b4f003e),
	.w7(32'hb9d5270f),
	.w8(32'h3ad253f3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfcb86),
	.w1(32'hbab6cbea),
	.w2(32'h3a2f4d46),
	.w3(32'hba4c828d),
	.w4(32'hbb75d1fa),
	.w5(32'hbab11ca1),
	.w6(32'hb9e78a38),
	.w7(32'hba0e2db7),
	.w8(32'h3a7bd5de),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85d983),
	.w1(32'h3b3a733c),
	.w2(32'h3a723706),
	.w3(32'h3bc50c31),
	.w4(32'h3ae63ef2),
	.w5(32'h39915a85),
	.w6(32'h3bd84c0f),
	.w7(32'h3b8781ed),
	.w8(32'h3b9cb202),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a13a5),
	.w1(32'hbae42a42),
	.w2(32'h39e3d0a6),
	.w3(32'h3b7fd67a),
	.w4(32'hbaef03b1),
	.w5(32'hbb02ffba),
	.w6(32'h3bab1020),
	.w7(32'h3a394fc6),
	.w8(32'hba8eeffd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b21e),
	.w1(32'hba71d7f5),
	.w2(32'hbb2309bc),
	.w3(32'h3b22af9e),
	.w4(32'h3a0c70cd),
	.w5(32'hbb56add6),
	.w6(32'h3b6d9cbd),
	.w7(32'h3b77f7cb),
	.w8(32'h3adc913e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c368ac),
	.w1(32'h3b02b398),
	.w2(32'h3b04efc7),
	.w3(32'h39c11259),
	.w4(32'h3a069bf7),
	.w5(32'hb98e3d00),
	.w6(32'hbaa94904),
	.w7(32'hbb1bda31),
	.w8(32'h3c397623),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec6fb2),
	.w1(32'h3b1e43ab),
	.w2(32'hbba114a4),
	.w3(32'h3afb7923),
	.w4(32'h3b240366),
	.w5(32'h3b8b17a8),
	.w6(32'h3c47be69),
	.w7(32'hbb378b69),
	.w8(32'hba83b254),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb575d60),
	.w1(32'h3b090806),
	.w2(32'hbac6113b),
	.w3(32'hb9174ab8),
	.w4(32'h3ab91084),
	.w5(32'h3a39b9dc),
	.w6(32'h3adbaa26),
	.w7(32'hba5d0b76),
	.w8(32'hba9ebd3c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eaeb51),
	.w1(32'h3b56c3f8),
	.w2(32'hbb7bd50c),
	.w3(32'h3a42d960),
	.w4(32'hbc0e9089),
	.w5(32'hba4e913a),
	.w6(32'h3ab44744),
	.w7(32'h3b881780),
	.w8(32'h3c1ce46d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc557760),
	.w1(32'hbc70096f),
	.w2(32'h3b7d161b),
	.w3(32'hba40dd67),
	.w4(32'hbbf39db4),
	.w5(32'hbc78b0e3),
	.w6(32'h3c5f0db3),
	.w7(32'hbbcf28b3),
	.w8(32'hbc1341bb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac16ffd),
	.w1(32'h3be08779),
	.w2(32'h38a2530e),
	.w3(32'h3baa88df),
	.w4(32'hbb2d400b),
	.w5(32'hb9d5def4),
	.w6(32'h3ad2b400),
	.w7(32'h3b9220cd),
	.w8(32'h3c7715f8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499072),
	.w1(32'hbc96645e),
	.w2(32'h3b133897),
	.w3(32'h3c63dbba),
	.w4(32'hbc778cae),
	.w5(32'hbc53383c),
	.w6(32'h3cce2402),
	.w7(32'h3c0eb3d5),
	.w8(32'h3c4b65e4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8397eb),
	.w1(32'hbba6abed),
	.w2(32'hbc0f0988),
	.w3(32'h3bb8b6a8),
	.w4(32'hbaa1e6f2),
	.w5(32'hbce0935d),
	.w6(32'h3c58aa86),
	.w7(32'hbc621a6f),
	.w8(32'hbca6ce71),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc665c8),
	.w1(32'hbba02d1b),
	.w2(32'hbbd09463),
	.w3(32'hbb0ef306),
	.w4(32'h3b907da2),
	.w5(32'hbcb43a8c),
	.w6(32'h3c9bd69b),
	.w7(32'h3bccd21d),
	.w8(32'h3c957bb5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69649a),
	.w1(32'hbc43a687),
	.w2(32'h3ae466c7),
	.w3(32'hbb89f271),
	.w4(32'h3c537305),
	.w5(32'hbb9f090a),
	.w6(32'h3d1f2aeb),
	.w7(32'hbc5e1bc3),
	.w8(32'h3c2022db),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156dfa),
	.w1(32'hbcb2efba),
	.w2(32'h3b0bf4f0),
	.w3(32'h3cc8d521),
	.w4(32'hbc42f4b2),
	.w5(32'hbc0892a1),
	.w6(32'h3d026337),
	.w7(32'hbc10ccdb),
	.w8(32'hbc3f4839),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc011d2),
	.w1(32'hbbcc377f),
	.w2(32'hbad0e0dc),
	.w3(32'h3c230889),
	.w4(32'hba91ec26),
	.w5(32'h3be770f9),
	.w6(32'hbc370f1a),
	.w7(32'hbb18c1bc),
	.w8(32'hbb9d6920),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dd317),
	.w1(32'h3af0bdb4),
	.w2(32'hbb624215),
	.w3(32'h39107886),
	.w4(32'hbb4ae322),
	.w5(32'hba87faa9),
	.w6(32'hbbf7bc83),
	.w7(32'hb982e4d8),
	.w8(32'h3b026d19),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca126e),
	.w1(32'h3b9ea3ae),
	.w2(32'h3ba90a04),
	.w3(32'h3c42e1db),
	.w4(32'hbc06e3b1),
	.w5(32'hba3dd9e6),
	.w6(32'h3c68bf30),
	.w7(32'h3d144b4b),
	.w8(32'hbc1b65cb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0056c2),
	.w1(32'h3bb624f5),
	.w2(32'h3b4eab91),
	.w3(32'h3a8151e9),
	.w4(32'h3bd03ba6),
	.w5(32'h3b614077),
	.w6(32'hbd07482b),
	.w7(32'h3b33691e),
	.w8(32'h3a481649),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd15b948),
	.w1(32'hbda5b1e8),
	.w2(32'hbd51cc73),
	.w3(32'hbc899f54),
	.w4(32'h3bff3dc5),
	.w5(32'hbbf3d8ef),
	.w6(32'h3d37c7cc),
	.w7(32'hbb92931e),
	.w8(32'hbb571b19),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5cb72),
	.w1(32'hbc65d4dc),
	.w2(32'hbc388a10),
	.w3(32'h3bf3725a),
	.w4(32'hbc373807),
	.w5(32'hbb83853f),
	.w6(32'h3c57a668),
	.w7(32'hbcb480b6),
	.w8(32'h3c785642),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae4b84),
	.w1(32'hbcc715a8),
	.w2(32'hbc357418),
	.w3(32'hbbd2bf09),
	.w4(32'h3b11339f),
	.w5(32'hbc44e6eb),
	.w6(32'h3c03b9a0),
	.w7(32'hbcc5b061),
	.w8(32'hbc7c35e1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4f55),
	.w1(32'h3a9d9c5a),
	.w2(32'hbaa7756a),
	.w3(32'hbc85c62b),
	.w4(32'h3b4aaeaa),
	.w5(32'h39d0a4d2),
	.w6(32'h3cc0c78f),
	.w7(32'hba437103),
	.w8(32'hbac4bc7e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3206f),
	.w1(32'h392009d1),
	.w2(32'hbc3fdb0b),
	.w3(32'hbaa9d705),
	.w4(32'hbcd36e7a),
	.w5(32'hbbbb2020),
	.w6(32'h3b3a1acc),
	.w7(32'hbd183fd9),
	.w8(32'h3c8af0c7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c552e4d),
	.w1(32'hbbf6de49),
	.w2(32'h3a7610f3),
	.w3(32'h3ca00817),
	.w4(32'h3c6cb890),
	.w5(32'hb8f5eeb0),
	.w6(32'h3d1156fa),
	.w7(32'h3ad5ab47),
	.w8(32'hbc14a08e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e00b),
	.w1(32'h3bc70f12),
	.w2(32'hbb901404),
	.w3(32'hbb83c0bd),
	.w4(32'hbc4a9f23),
	.w5(32'hbc1f8c99),
	.w6(32'h3b2bfa87),
	.w7(32'h3c820816),
	.w8(32'h3c8c95e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133010),
	.w1(32'hbc125514),
	.w2(32'h3a1a7e0c),
	.w3(32'h3923b89b),
	.w4(32'h3c1a8605),
	.w5(32'h3b2df1f3),
	.w6(32'hbc4a10c5),
	.w7(32'h3ba8a443),
	.w8(32'h3c379a7a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be37879),
	.w1(32'h3af627e8),
	.w2(32'h3aef6eb9),
	.w3(32'h3c23f3c3),
	.w4(32'hba168c9d),
	.w5(32'hbaee5de4),
	.w6(32'h3c58be62),
	.w7(32'hbc981d2f),
	.w8(32'hbba372fd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde2b55),
	.w1(32'hbbd3874d),
	.w2(32'hbc179667),
	.w3(32'h3c3d81ae),
	.w4(32'hbc206821),
	.w5(32'hbc40b65d),
	.w6(32'hbce5fb6f),
	.w7(32'h3c51db8f),
	.w8(32'h3d32944e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e53d),
	.w1(32'hbbcb37e4),
	.w2(32'hbb204111),
	.w3(32'hbc793fb1),
	.w4(32'hba8a6605),
	.w5(32'h3b9e824b),
	.w6(32'h3c30fac1),
	.w7(32'h3c35a6d1),
	.w8(32'h3b89507a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb3d7a),
	.w1(32'h3ba1ec68),
	.w2(32'hbc133e83),
	.w3(32'h3ba9ede0),
	.w4(32'hbcb97518),
	.w5(32'hbc83a8be),
	.w6(32'hbb9fb686),
	.w7(32'hbc554adb),
	.w8(32'h3bcc2435),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974f37e),
	.w1(32'hbcbd261e),
	.w2(32'h3c3b69e4),
	.w3(32'h3bf90879),
	.w4(32'hbbbfbf89),
	.w5(32'hbbf525c2),
	.w6(32'h3a933dc5),
	.w7(32'hbad4702f),
	.w8(32'hba76e880),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb60b2c),
	.w1(32'h378cec22),
	.w2(32'hbbf3cf29),
	.w3(32'h3b7edfa0),
	.w4(32'hbc0d0691),
	.w5(32'hbc4e36dc),
	.w6(32'h3c01ee64),
	.w7(32'h3bf36a1c),
	.w8(32'hbbfeff74),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca60a6),
	.w1(32'hbaf28cf1),
	.w2(32'h3bb2dfe6),
	.w3(32'hbab50e49),
	.w4(32'h3ca7e59e),
	.w5(32'h3c4b68ec),
	.w6(32'hbc2cab40),
	.w7(32'hb956d320),
	.w8(32'hbd306866),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaea21),
	.w1(32'h3be35805),
	.w2(32'h3ba07d1f),
	.w3(32'hb84d13f2),
	.w4(32'hbc38e99e),
	.w5(32'hbc5b0a03),
	.w6(32'hbc891053),
	.w7(32'hbcabfc96),
	.w8(32'h3d03aa80),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14c543),
	.w1(32'hbc61718c),
	.w2(32'hbac4318f),
	.w3(32'h3ca6f475),
	.w4(32'hba46138f),
	.w5(32'hbb8c49d6),
	.w6(32'h3a90a8ef),
	.w7(32'hba945cd3),
	.w8(32'h3b861357),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce945),
	.w1(32'hbb14a060),
	.w2(32'hb90d9d00),
	.w3(32'h3b807da2),
	.w4(32'h3b011d51),
	.w5(32'h3a28c873),
	.w6(32'h3c75863f),
	.w7(32'hbc92d907),
	.w8(32'hbcd041a9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33dca8),
	.w1(32'hbc1ea30b),
	.w2(32'h3c07a426),
	.w3(32'h3be63696),
	.w4(32'h3c126bd4),
	.w5(32'h3caf1f68),
	.w6(32'h3b9f41b5),
	.w7(32'hba9c1ee7),
	.w8(32'hbae92f7a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3abc),
	.w1(32'h3c39d507),
	.w2(32'hbc388246),
	.w3(32'h3bf6d0d4),
	.w4(32'h3c226c46),
	.w5(32'hbcb9ccd9),
	.w6(32'hbc972bb7),
	.w7(32'h3b917b96),
	.w8(32'hbbdddb28),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d09be),
	.w1(32'h3af041fa),
	.w2(32'h3b7c4822),
	.w3(32'hbbda3403),
	.w4(32'hbc1461a3),
	.w5(32'hbc2079af),
	.w6(32'h3ccaa56e),
	.w7(32'hbc33f68c),
	.w8(32'hbb8dad25),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20aedf),
	.w1(32'h3ba90cac),
	.w2(32'hbb160869),
	.w3(32'hbbacb85e),
	.w4(32'hbb8ef831),
	.w5(32'hbc57523b),
	.w6(32'h3b9e3cb7),
	.w7(32'hbc7ded2d),
	.w8(32'hbcd032c5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab460),
	.w1(32'hbbb24ba8),
	.w2(32'hbc459939),
	.w3(32'hbc8b5f93),
	.w4(32'hbc7e5e7d),
	.w5(32'hbc288794),
	.w6(32'hbc53b25f),
	.w7(32'hbbe98ed6),
	.w8(32'hbc600508),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dc0bd),
	.w1(32'hbb8de744),
	.w2(32'hbc539370),
	.w3(32'hbc242e94),
	.w4(32'h3c447bce),
	.w5(32'h3c913972),
	.w6(32'hbc099d25),
	.w7(32'h3ce02276),
	.w8(32'hbd3cfe4b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8182de),
	.w1(32'h3cac4190),
	.w2(32'h3bd89ab8),
	.w3(32'hbbde21a0),
	.w4(32'hbcaab696),
	.w5(32'hbcee3d67),
	.w6(32'hbc598b94),
	.w7(32'h3c0e53db),
	.w8(32'hbaebc1db),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03db24),
	.w1(32'hbb5ca21c),
	.w2(32'hba154743),
	.w3(32'hbc2c5dcf),
	.w4(32'hbc8ba346),
	.w5(32'h3b85cc3b),
	.w6(32'h3c6e762e),
	.w7(32'hbb50aeb8),
	.w8(32'hbc6d9f1f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1992),
	.w1(32'h3c23735c),
	.w2(32'hbb757d28),
	.w3(32'h3c6e755c),
	.w4(32'h3b84bd05),
	.w5(32'h3a85d840),
	.w6(32'hbc9aee7b),
	.w7(32'h3a43f7b8),
	.w8(32'h3bf28e6c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac105e),
	.w1(32'hbb1293f7),
	.w2(32'h3c66986c),
	.w3(32'hba6ca5ea),
	.w4(32'h3c0b8e4a),
	.w5(32'h3cc3dfe0),
	.w6(32'h3b673953),
	.w7(32'h3a97cdbe),
	.w8(32'h3d43800d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb34317),
	.w1(32'hbc50f48d),
	.w2(32'hbc1e7a5a),
	.w3(32'hbccd18d8),
	.w4(32'hbb58c4ef),
	.w5(32'hbbbc34a5),
	.w6(32'hbc0d2877),
	.w7(32'hba80dce2),
	.w8(32'h3a08aeb4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeef1ee),
	.w1(32'hbb47cb7c),
	.w2(32'h3ba9a61a),
	.w3(32'hbbb851ed),
	.w4(32'hbbe74e33),
	.w5(32'hbb768c90),
	.w6(32'hbbd859fc),
	.w7(32'hba7bbe79),
	.w8(32'hbb80c96f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf2f70),
	.w1(32'h3b78c99a),
	.w2(32'h3c2a0cbc),
	.w3(32'hbaf9d1e6),
	.w4(32'h3c6d396a),
	.w5(32'hbc7bc091),
	.w6(32'hbba00e16),
	.w7(32'h3aeabfe7),
	.w8(32'h3c091350),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc667a),
	.w1(32'hbc071a15),
	.w2(32'hbb656c65),
	.w3(32'hbb586c07),
	.w4(32'hbb0b8ba8),
	.w5(32'hbafcd817),
	.w6(32'h3b52799b),
	.w7(32'hbb9318eb),
	.w8(32'h3af9b19d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b8e3),
	.w1(32'hb9ce7990),
	.w2(32'h3a2708d4),
	.w3(32'h3a756ff2),
	.w4(32'hbcf8eb4f),
	.w5(32'h3b89a9f2),
	.w6(32'h3b3b1469),
	.w7(32'h3c821488),
	.w8(32'h3cba88de),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc776f70),
	.w1(32'hba991ad2),
	.w2(32'hbbae42fb),
	.w3(32'h3ce36562),
	.w4(32'h3c2eee88),
	.w5(32'h3ca4e702),
	.w6(32'hbd2bd98d),
	.w7(32'hbbd07ad3),
	.w8(32'hbc753b00),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c204c4f),
	.w1(32'h3bea7275),
	.w2(32'hbaa6dcf8),
	.w3(32'h3c78bcf3),
	.w4(32'h3c0dc773),
	.w5(32'hb9c052b4),
	.w6(32'hbc971a60),
	.w7(32'h3c0cbc5c),
	.w8(32'h3bdd3d25),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9f361),
	.w1(32'h3b880fd9),
	.w2(32'hbc2ea79b),
	.w3(32'h3b1bdd80),
	.w4(32'hbc17eb4a),
	.w5(32'hbc2b0138),
	.w6(32'h3cd6d764),
	.w7(32'hbb16ca70),
	.w8(32'hbbd18450),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a4f28),
	.w1(32'hb924f86c),
	.w2(32'hbb71cedb),
	.w3(32'hbc1d5d23),
	.w4(32'h3b8e0146),
	.w5(32'hbb381b5a),
	.w6(32'hbbc26bcb),
	.w7(32'hbbec77a3),
	.w8(32'hbb7ba348),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe75b6),
	.w1(32'h3a9b625d),
	.w2(32'h3af00cb5),
	.w3(32'hb827e93c),
	.w4(32'hbc16c80b),
	.w5(32'hbb8b3a35),
	.w6(32'h3c77f5fb),
	.w7(32'hbbe93fdf),
	.w8(32'h3c332902),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806710e),
	.w1(32'hbc47f551),
	.w2(32'hbb8326ed),
	.w3(32'hbbc7d343),
	.w4(32'hbb8ed14c),
	.w5(32'hbc618559),
	.w6(32'h3bdf09e8),
	.w7(32'hb96b0ffa),
	.w8(32'hbc180b0c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac05718),
	.w1(32'h3c6fe5ea),
	.w2(32'h3aef1862),
	.w3(32'hbc018080),
	.w4(32'hbc657776),
	.w5(32'hbcab9a8a),
	.w6(32'hbc527051),
	.w7(32'hbb6f2568),
	.w8(32'hbcb53a73),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67474),
	.w1(32'h3b1eb52a),
	.w2(32'h3b2c138e),
	.w3(32'h3c19b2de),
	.w4(32'hbaf3e30c),
	.w5(32'hbbe462a4),
	.w6(32'hba8e3429),
	.w7(32'h3b135a29),
	.w8(32'hbb544ddb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb67dd6),
	.w1(32'hbc503556),
	.w2(32'h3ba9b837),
	.w3(32'hbb07191a),
	.w4(32'h3c2072cd),
	.w5(32'h3cb5a59e),
	.w6(32'h3b9726d5),
	.w7(32'hb9db278a),
	.w8(32'h3b9ff172),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add08a2),
	.w1(32'hbc94fee4),
	.w2(32'hbbc81e4c),
	.w3(32'h3bc142f5),
	.w4(32'h3a5b9ae8),
	.w5(32'hbcce622e),
	.w6(32'h3bfa04a5),
	.w7(32'hbaea1fa7),
	.w8(32'hbc8a75fa),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d5252),
	.w1(32'hbb17721b),
	.w2(32'h3a6fcdc4),
	.w3(32'hbc7fb2c7),
	.w4(32'h3b546bf7),
	.w5(32'hbbbe49f7),
	.w6(32'h3b254aa2),
	.w7(32'hbbcff35a),
	.w8(32'hbcc5ebd4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c63d),
	.w1(32'h3be6763d),
	.w2(32'hbc46a852),
	.w3(32'h3aba8dda),
	.w4(32'hbba1bb51),
	.w5(32'hbbbb5e62),
	.w6(32'hbc59f41d),
	.w7(32'hbb8ea6bd),
	.w8(32'hbb99f15b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56ebee),
	.w1(32'h398e0f16),
	.w2(32'h3bf5725f),
	.w3(32'hbb5f1cad),
	.w4(32'h3a29ae5e),
	.w5(32'hbbad6c27),
	.w6(32'hbc1fc8f0),
	.w7(32'hbc005769),
	.w8(32'h3beff144),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52965c),
	.w1(32'h3b9fcacd),
	.w2(32'hbae9a5ae),
	.w3(32'h3b9d6cb1),
	.w4(32'hbd1acbf0),
	.w5(32'hbbbc4a11),
	.w6(32'h3c652fbf),
	.w7(32'h3d029b14),
	.w8(32'h3d310272),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc825cb6),
	.w1(32'h3c234cc4),
	.w2(32'hbc74d50d),
	.w3(32'h3c7178c5),
	.w4(32'hbc00b2e0),
	.w5(32'hbceafa61),
	.w6(32'hbd03f8e7),
	.w7(32'hbc44424a),
	.w8(32'hbc5040c5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5fd55),
	.w1(32'hbba72fb1),
	.w2(32'hbc0959bb),
	.w3(32'hbbdb5eb4),
	.w4(32'hbb7112e5),
	.w5(32'hbb88f1e9),
	.w6(32'h3c7850ce),
	.w7(32'hbbc0ee46),
	.w8(32'hbc55525d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4f930),
	.w1(32'hbb916dd5),
	.w2(32'h369158b6),
	.w3(32'h3aac05ae),
	.w4(32'hb917fc77),
	.w5(32'hb8b66d46),
	.w6(32'hbbf763f9),
	.w7(32'h38e55433),
	.w8(32'hb86c435f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec174a),
	.w1(32'hbbd529b5),
	.w2(32'hbb8d1349),
	.w3(32'h3b2066ad),
	.w4(32'hbb92d191),
	.w5(32'hbbd31d5a),
	.w6(32'h3bef075a),
	.w7(32'hb8b27973),
	.w8(32'hbb64361d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89c978),
	.w1(32'hbb54c14f),
	.w2(32'hbb583c24),
	.w3(32'h3ad0df82),
	.w4(32'hbac069fc),
	.w5(32'hbb3314ab),
	.w6(32'h3b7bc081),
	.w7(32'h3af9429c),
	.w8(32'h3acb32d4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df417e),
	.w1(32'hba382319),
	.w2(32'hba862041),
	.w3(32'hb9dbdd9f),
	.w4(32'hba26333c),
	.w5(32'hba07bcdf),
	.w6(32'hb9b54e4b),
	.w7(32'hb9798e15),
	.w8(32'hb94eb59e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fcc108),
	.w1(32'h39f68036),
	.w2(32'hb86ef060),
	.w3(32'h39b76e0c),
	.w4(32'h398f05ba),
	.w5(32'h38cc0879),
	.w6(32'h3899f820),
	.w7(32'h38c08ebf),
	.w8(32'hb977ed34),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6a2ae),
	.w1(32'hb9eed383),
	.w2(32'h3a630bfe),
	.w3(32'h3b1c03e7),
	.w4(32'h3aa44863),
	.w5(32'h3acce2ff),
	.w6(32'hbaacce6a),
	.w7(32'hbabb2f05),
	.w8(32'h390dcf92),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954c41),
	.w1(32'hbab85033),
	.w2(32'h3a941b4e),
	.w3(32'h3ba3691a),
	.w4(32'hbad25196),
	.w5(32'hbb3fe1db),
	.w6(32'h3c262f7c),
	.w7(32'h3b863b6e),
	.w8(32'h3aa7f9e0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999ef59),
	.w1(32'hbad0eed5),
	.w2(32'hbc23b635),
	.w3(32'h38b7ab80),
	.w4(32'hbb56374b),
	.w5(32'hbc23b1e9),
	.w6(32'hbae266aa),
	.w7(32'h3b33588a),
	.w8(32'hbb8b6af1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1afd),
	.w1(32'hbb7ebd45),
	.w2(32'hb9bb443b),
	.w3(32'h3c3556b0),
	.w4(32'hba954502),
	.w5(32'hbbf68a5e),
	.w6(32'h3c8dbcc0),
	.w7(32'h3c0b6212),
	.w8(32'h3b9b5d5d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78f46e),
	.w1(32'hbb222431),
	.w2(32'hbaf3d3bd),
	.w3(32'h3bae5073),
	.w4(32'hbb7b9a62),
	.w5(32'hbb9565ee),
	.w6(32'h3b536ca8),
	.w7(32'h39cd3fac),
	.w8(32'hbb59ce6b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b57e4),
	.w1(32'hb9d0bb12),
	.w2(32'hb99c16b5),
	.w3(32'hb9d61537),
	.w4(32'hb85709e2),
	.w5(32'hb8c16ca8),
	.w6(32'h39919296),
	.w7(32'hb9673f27),
	.w8(32'hb80f16e6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f65ce1),
	.w1(32'h391a7de2),
	.w2(32'h378529a5),
	.w3(32'h39515b44),
	.w4(32'hb85c020e),
	.w5(32'hb8b53c69),
	.w6(32'h392b4c2d),
	.w7(32'hb7e892e0),
	.w8(32'hb9482fa4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88377ce),
	.w1(32'h383ff5f6),
	.w2(32'h38c62ead),
	.w3(32'h38a0f27b),
	.w4(32'hb77bf026),
	.w5(32'hb804f1ff),
	.w6(32'h384ac150),
	.w7(32'hb93c7b7f),
	.w8(32'hb8d9fad5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421dd7),
	.w1(32'hb9a5a1f1),
	.w2(32'hb9ca82d3),
	.w3(32'h3afd50b3),
	.w4(32'hb82c7968),
	.w5(32'hbb3a7bcc),
	.w6(32'h3b74da27),
	.w7(32'hb9f82b41),
	.w8(32'hb9f89501),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae030ea),
	.w1(32'hbb0cbfdc),
	.w2(32'hbb21f327),
	.w3(32'hbaa6b888),
	.w4(32'hbab46807),
	.w5(32'hbb152cf2),
	.w6(32'hba0c3797),
	.w7(32'hbaf4c647),
	.w8(32'hbab72207),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f956e),
	.w1(32'hb98d7dba),
	.w2(32'h3a092243),
	.w3(32'h3a6f50cd),
	.w4(32'h3a878848),
	.w5(32'hba017c48),
	.w6(32'h3a71df55),
	.w7(32'hb9d6e2d5),
	.w8(32'hb9c91c5e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13a06f),
	.w1(32'hba3b0195),
	.w2(32'h3a9e1bfd),
	.w3(32'hbab153b8),
	.w4(32'h3a225dd8),
	.w5(32'h3af213ec),
	.w6(32'hba67e9bf),
	.w7(32'hba03d36c),
	.w8(32'h3a15f206),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d504e),
	.w1(32'h3802f5c3),
	.w2(32'hba115261),
	.w3(32'h3b0dd0f1),
	.w4(32'hba3cfda7),
	.w5(32'hbb1c8e6e),
	.w6(32'h3b80ff38),
	.w7(32'h3b0079e3),
	.w8(32'hba07dc50),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad331c6),
	.w1(32'h38eeeb00),
	.w2(32'hb9e0a285),
	.w3(32'h3b653b61),
	.w4(32'h3a8d02a2),
	.w5(32'h38653682),
	.w6(32'h3b4aca36),
	.w7(32'h3a9d202f),
	.w8(32'h3a724d0a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b32af),
	.w1(32'hb963ef7e),
	.w2(32'hb996953a),
	.w3(32'h3bb8d95b),
	.w4(32'h39089a6e),
	.w5(32'hba1da617),
	.w6(32'h3bfbe99b),
	.w7(32'h3b91eca0),
	.w8(32'h3abae6eb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c74b9),
	.w1(32'hbb26284d),
	.w2(32'hba8f922c),
	.w3(32'h3b1e2a7a),
	.w4(32'hbb8ee2c7),
	.w5(32'hbb452be2),
	.w6(32'h3c2e72cb),
	.w7(32'h3b6ef7d8),
	.w8(32'h3ae38774),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38863654),
	.w1(32'h39180985),
	.w2(32'hb9a9c034),
	.w3(32'h37ee2cd1),
	.w4(32'h3a22aa99),
	.w5(32'hb9c889bb),
	.w6(32'h3921e6e5),
	.w7(32'hb81ccffe),
	.w8(32'h39c15cb5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3cd4),
	.w1(32'hb89186d0),
	.w2(32'h39844011),
	.w3(32'h3a8d4e17),
	.w4(32'hb74e2b8a),
	.w5(32'h38f91e21),
	.w6(32'h3a33f814),
	.w7(32'h38488b28),
	.w8(32'h391caece),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39484ad1),
	.w1(32'h37e5568b),
	.w2(32'hb8809e7b),
	.w3(32'h392f7042),
	.w4(32'hb93956c2),
	.w5(32'hb8e87536),
	.w6(32'h388778cc),
	.w7(32'hb89ea486),
	.w8(32'hb90e522f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39356af7),
	.w1(32'h39ae4420),
	.w2(32'hb9ce007a),
	.w3(32'hb9257421),
	.w4(32'hb9ad6258),
	.w5(32'hb974c273),
	.w6(32'h39cb572d),
	.w7(32'h38864b42),
	.w8(32'hba3bf8a7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1a16),
	.w1(32'hb9c7c9c9),
	.w2(32'h37ed2841),
	.w3(32'h3b0cfba3),
	.w4(32'h39b4b3d2),
	.w5(32'h38a42c2b),
	.w6(32'h3aeb8540),
	.w7(32'h3ac58a35),
	.w8(32'h3a8c1bd9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926105),
	.w1(32'h3a80a5e3),
	.w2(32'h3a8c3a34),
	.w3(32'h3a916732),
	.w4(32'h3a67ae87),
	.w5(32'h3a945c02),
	.w6(32'h3aab0958),
	.w7(32'h3ab8d70a),
	.w8(32'h3ab6abb0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9758c9),
	.w1(32'h3a21aedd),
	.w2(32'h3aa68f50),
	.w3(32'h37ea2471),
	.w4(32'h3aa2af87),
	.w5(32'h3b8d0346),
	.w6(32'hba9934b7),
	.w7(32'hb998c7b2),
	.w8(32'h3aadbc1d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba174f7f),
	.w1(32'h397ef203),
	.w2(32'hb99c5796),
	.w3(32'hba9f3d38),
	.w4(32'hba042b5f),
	.w5(32'h3a354e43),
	.w6(32'hbb30af39),
	.w7(32'hbaa44588),
	.w8(32'hbaace754),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05b78e),
	.w1(32'hbaefb2fe),
	.w2(32'h3b033b2a),
	.w3(32'h39d1ead1),
	.w4(32'hb980e0a7),
	.w5(32'hbb82167c),
	.w6(32'h3b42eb6f),
	.w7(32'hbadcf316),
	.w8(32'hba9c79b9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d513a),
	.w1(32'hbb2ecba4),
	.w2(32'hbab851c9),
	.w3(32'h3aa98ffc),
	.w4(32'hbb48dd9f),
	.w5(32'hbb123d31),
	.w6(32'h3b8fe137),
	.w7(32'h3a894295),
	.w8(32'hbb33eedb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bec79),
	.w1(32'h3b17620c),
	.w2(32'h3a78c909),
	.w3(32'hb9f7cf87),
	.w4(32'hb91d5c44),
	.w5(32'h38050819),
	.w6(32'hbb27afbc),
	.w7(32'h38f04460),
	.w8(32'h38ca08b3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39741e99),
	.w1(32'h3acd1fad),
	.w2(32'hba5c6ca8),
	.w3(32'hb95b8abb),
	.w4(32'h3abf3ae7),
	.w5(32'hb8b04a7a),
	.w6(32'hbb1538b9),
	.w7(32'hba6460a6),
	.w8(32'hbac85707),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3cd5a),
	.w1(32'hba6979a6),
	.w2(32'h3b0046a9),
	.w3(32'h3b09fc6b),
	.w4(32'hb9b6256c),
	.w5(32'h3b3bc85e),
	.w6(32'h3b93fac5),
	.w7(32'h3b8a9d9e),
	.w8(32'h3b3f4a41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9f4d5),
	.w1(32'hb902473b),
	.w2(32'hbb32217a),
	.w3(32'h3a7798e5),
	.w4(32'h3b02dcb2),
	.w5(32'hbaa45bc4),
	.w6(32'h3a9d4094),
	.w7(32'h3b5797b7),
	.w8(32'h3b4e3aa2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b41d),
	.w1(32'hbb69130f),
	.w2(32'hbb357262),
	.w3(32'hbb6c3e7b),
	.w4(32'hbaa2e363),
	.w5(32'hbadd2781),
	.w6(32'hbb491409),
	.w7(32'hba0e4583),
	.w8(32'hbaf9f9a1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2681e8),
	.w1(32'h3b623332),
	.w2(32'h3b61dc8a),
	.w3(32'hba1cd530),
	.w4(32'h3b6e51df),
	.w5(32'h3b346f85),
	.w6(32'hbb40e74e),
	.w7(32'hbac0d4b8),
	.w8(32'h3a0125f5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9168335),
	.w1(32'hbaa1c791),
	.w2(32'hba0284d6),
	.w3(32'hb9daae9c),
	.w4(32'hb937ac7f),
	.w5(32'hb92dadb7),
	.w6(32'h3a352a41),
	.w7(32'hb9af40a9),
	.w8(32'hb90cdfb1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f62df),
	.w1(32'h399dc62b),
	.w2(32'h3788e6c1),
	.w3(32'h3a805316),
	.w4(32'h3a1a24fc),
	.w5(32'hba807ca2),
	.w6(32'h3a427aa2),
	.w7(32'hbac0b1d2),
	.w8(32'hbb02f6fa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df730e),
	.w1(32'hba95b48e),
	.w2(32'hb98d4b15),
	.w3(32'hb89ac63a),
	.w4(32'h39d4200a),
	.w5(32'h3903b113),
	.w6(32'h3b29589b),
	.w7(32'h3aba1974),
	.w8(32'h389e3f8c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf909d),
	.w1(32'h3a1ce81f),
	.w2(32'hba35e09a),
	.w3(32'h39d3297b),
	.w4(32'h3aacc535),
	.w5(32'hb90ecfeb),
	.w6(32'h390ab437),
	.w7(32'h3a883fcd),
	.w8(32'hba0c82a4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39393b1a),
	.w1(32'hba8c79a0),
	.w2(32'hbb0c977a),
	.w3(32'hba5343d5),
	.w4(32'hb9e189b4),
	.w5(32'hbb2b57f2),
	.w6(32'h38f6f272),
	.w7(32'hb98d43d3),
	.w8(32'hba9454da),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899a07b),
	.w1(32'h38f42917),
	.w2(32'h398a6271),
	.w3(32'h382f5f09),
	.w4(32'h39ab79b8),
	.w5(32'h39917704),
	.w6(32'h37ec85ae),
	.w7(32'h394cd211),
	.w8(32'hba1a6fbd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abf0ed),
	.w1(32'hba055834),
	.w2(32'h3965516f),
	.w3(32'hb91fb091),
	.w4(32'hb9430e68),
	.w5(32'h3944c8c8),
	.w6(32'h3a759aff),
	.w7(32'h3a1e6f19),
	.w8(32'h3a17564d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d23ab),
	.w1(32'h36e4282c),
	.w2(32'hba9b5759),
	.w3(32'h3b00b89d),
	.w4(32'h3a579473),
	.w5(32'h3a7ca6be),
	.w6(32'hb723bdfa),
	.w7(32'hb9f0c76c),
	.w8(32'h3a8eed65),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eee55e),
	.w1(32'hbb357320),
	.w2(32'hbb53c506),
	.w3(32'h3b922140),
	.w4(32'h39e68f2c),
	.w5(32'hbb0eba7e),
	.w6(32'h3bd489ee),
	.w7(32'h3b96643c),
	.w8(32'h3a12893a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba769fd3),
	.w1(32'hba9efffb),
	.w2(32'hbaab676b),
	.w3(32'hba85b9f3),
	.w4(32'hb9b2419d),
	.w5(32'h37bdb455),
	.w6(32'hba832eff),
	.w7(32'hba12f40c),
	.w8(32'hb9a45460),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f01744),
	.w1(32'h3abb94a7),
	.w2(32'hb699541d),
	.w3(32'h3a2b61c4),
	.w4(32'h3aebb755),
	.w5(32'h3a3581e9),
	.w6(32'hba2a33d5),
	.w7(32'h39a6a2c5),
	.w8(32'hba0b537c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b1648),
	.w1(32'h3abc3520),
	.w2(32'h3aac57f6),
	.w3(32'h3a967074),
	.w4(32'h3a92e73a),
	.w5(32'h3afd466a),
	.w6(32'h3ae64ce2),
	.w7(32'h3b29cb73),
	.w8(32'h3b1c14fa),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4e8c),
	.w1(32'hba9dbe33),
	.w2(32'hba876807),
	.w3(32'hbb3b95f0),
	.w4(32'hbaa8e559),
	.w5(32'hba5a5227),
	.w6(32'hbae1e30c),
	.w7(32'hb95786d6),
	.w8(32'h398bf437),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a082e80),
	.w1(32'hba11e276),
	.w2(32'hba5e6525),
	.w3(32'h3b518d94),
	.w4(32'h3ac4d9fb),
	.w5(32'h3a10f313),
	.w6(32'h3b7c42b4),
	.w7(32'h3b37dfe6),
	.w8(32'h3af907e9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913441),
	.w1(32'hbafa7839),
	.w2(32'hbad0db47),
	.w3(32'h38899f49),
	.w4(32'hb90fe684),
	.w5(32'hbae4879c),
	.w6(32'h3a9b8b45),
	.w7(32'h3a49f96b),
	.w8(32'hbaa6609b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule