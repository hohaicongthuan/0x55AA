module layer_10_featuremap_119(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb973add3),
	.w1(32'h3a66db12),
	.w2(32'h3b2108e5),
	.w3(32'hb8f593ca),
	.w4(32'hba5abc01),
	.w5(32'h3a0c1f44),
	.w6(32'h37d737f2),
	.w7(32'hba41bbc1),
	.w8(32'hb939dafe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a7659),
	.w1(32'h3a253e14),
	.w2(32'h3992d63e),
	.w3(32'h3a1d8b7f),
	.w4(32'h39b3619c),
	.w5(32'h3979f4b8),
	.w6(32'h3a0416f7),
	.w7(32'h3934d4bf),
	.w8(32'hb74da719),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a843b6),
	.w1(32'hb7aeb49c),
	.w2(32'h38fda826),
	.w3(32'h39b94b5d),
	.w4(32'h39a29d0b),
	.w5(32'h397673ed),
	.w6(32'h3950cf20),
	.w7(32'h3907f537),
	.w8(32'hb79b0964),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cdb84),
	.w1(32'hbace3305),
	.w2(32'hba8d70ff),
	.w3(32'h3a0e440f),
	.w4(32'h395623d1),
	.w5(32'h399bd85d),
	.w6(32'hb9cad028),
	.w7(32'hba3ac1ee),
	.w8(32'hba5ac8b3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cc549),
	.w1(32'h39a1f4ce),
	.w2(32'h39733e26),
	.w3(32'h39a5d945),
	.w4(32'h39a2b31d),
	.w5(32'h38adf2cb),
	.w6(32'h394eb7e3),
	.w7(32'h376bceac),
	.w8(32'hb9e11f78),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2b8e5),
	.w1(32'h399d7649),
	.w2(32'hb8c7120b),
	.w3(32'h38e5e89f),
	.w4(32'h39f69717),
	.w5(32'hb715c1b9),
	.w6(32'h3a05a3aa),
	.w7(32'h393a9f2c),
	.w8(32'h3725c252),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378d8a31),
	.w1(32'h3a1e18ff),
	.w2(32'h3a0f530c),
	.w3(32'h39eee58c),
	.w4(32'h3a349cfc),
	.w5(32'h3a2dcfbf),
	.w6(32'h3a5becd0),
	.w7(32'h39ed6068),
	.w8(32'h396fec82),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c8af1),
	.w1(32'hba1704f6),
	.w2(32'hba4b4ecf),
	.w3(32'h3a27c5ce),
	.w4(32'hb9196aaa),
	.w5(32'hb96a108f),
	.w6(32'h38e234d9),
	.w7(32'hb92cc74d),
	.w8(32'hba086efc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946dc5a),
	.w1(32'hb9c2778e),
	.w2(32'hb947f965),
	.w3(32'hb947fe66),
	.w4(32'hb98d65a1),
	.w5(32'h384fecd5),
	.w6(32'hb9e06bae),
	.w7(32'hb99a8c9c),
	.w8(32'hb92b37cb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02df02),
	.w1(32'h3a94a820),
	.w2(32'h39a06b77),
	.w3(32'hb8064308),
	.w4(32'h3a6fb19d),
	.w5(32'h3787d01c),
	.w6(32'h3a39af66),
	.w7(32'h38f6fac0),
	.w8(32'hb82facfd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39864a7b),
	.w1(32'hba446782),
	.w2(32'hba7ab2d5),
	.w3(32'h3a0c1929),
	.w4(32'h3917f0d7),
	.w5(32'h37d4978e),
	.w6(32'hb966aba9),
	.w7(32'hb9c4ea5a),
	.w8(32'hb9fb1816),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf303f3),
	.w1(32'hba829e84),
	.w2(32'hb90c9c07),
	.w3(32'hb8226822),
	.w4(32'h395fc869),
	.w5(32'hb983306d),
	.w6(32'h3a15ca4f),
	.w7(32'h3821c41b),
	.w8(32'hb9bc1f08),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954c024),
	.w1(32'hb8da016b),
	.w2(32'hb98ecbf1),
	.w3(32'hb8ab240f),
	.w4(32'h395ba92b),
	.w5(32'h37040111),
	.w6(32'hb9b4e597),
	.w7(32'hb9f396c5),
	.w8(32'hb96f0115),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db915b),
	.w1(32'hba1610d2),
	.w2(32'hba3b3dde),
	.w3(32'h3993e387),
	.w4(32'hb97e1944),
	.w5(32'hb9de352f),
	.w6(32'hba0269cb),
	.w7(32'hba0463b2),
	.w8(32'hb9f4e5c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f82588),
	.w1(32'hb9bf5cae),
	.w2(32'h3922227e),
	.w3(32'hb978b6d7),
	.w4(32'hba47f588),
	.w5(32'hba59b3d9),
	.w6(32'hba41527a),
	.w7(32'hbaa5e0b9),
	.w8(32'hbaded088),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6a3f7),
	.w1(32'hb985d4d4),
	.w2(32'hb9a5efe1),
	.w3(32'hb952cd65),
	.w4(32'hb9b76f7b),
	.w5(32'hb9aa8a8b),
	.w6(32'hb9a75ea0),
	.w7(32'hb9fc31bb),
	.w8(32'hba1aa797),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b8d08b),
	.w1(32'hb815e2ae),
	.w2(32'hb69e445c),
	.w3(32'h38ce139d),
	.w4(32'h390eb4d0),
	.w5(32'hb99b579d),
	.w6(32'hb9450876),
	.w7(32'h384b6325),
	.w8(32'h38715119),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0bec8),
	.w1(32'hba48ebfd),
	.w2(32'hb9a94b72),
	.w3(32'h3a8df575),
	.w4(32'h3a655d06),
	.w5(32'h3647b000),
	.w6(32'h3a3e3c03),
	.w7(32'h390234b7),
	.w8(32'hb9aebd61),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9209b35),
	.w1(32'hba14a916),
	.w2(32'hb9abaaec),
	.w3(32'h3a2eefdd),
	.w4(32'h39c727f5),
	.w5(32'hb7d8c331),
	.w6(32'h3981acc1),
	.w7(32'h375a9586),
	.w8(32'hb9087726),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907cd1c),
	.w1(32'hb92d2938),
	.w2(32'hb79536e4),
	.w3(32'h38c90e9a),
	.w4(32'hb88a8eca),
	.w5(32'h39542e2c),
	.w6(32'hb8ccd789),
	.w7(32'hb8bcb514),
	.w8(32'hb886076b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373c7e59),
	.w1(32'hba051c5a),
	.w2(32'hb9e328ae),
	.w3(32'h37de07e1),
	.w4(32'h38c14b28),
	.w5(32'hb887ff47),
	.w6(32'hb9a57322),
	.w7(32'hb99d6bd9),
	.w8(32'hb982543b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf587a),
	.w1(32'h3aa11cb9),
	.w2(32'h3a6b9fc3),
	.w3(32'h38ded041),
	.w4(32'h397a055d),
	.w5(32'hb83a0103),
	.w6(32'hba2031a2),
	.w7(32'hbab43bbb),
	.w8(32'hbac98355),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ebb38),
	.w1(32'hba5a7e09),
	.w2(32'hbab3ff05),
	.w3(32'h3a37080b),
	.w4(32'h3989114e),
	.w5(32'hba90856b),
	.w6(32'h38ca7daf),
	.w7(32'hba209774),
	.w8(32'hba695306),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb9950),
	.w1(32'h3a4682ad),
	.w2(32'hb883ae3d),
	.w3(32'h3954b27c),
	.w4(32'h38d152a9),
	.w5(32'hb8e70b70),
	.w6(32'hba2be607),
	.w7(32'hb99769b4),
	.w8(32'hba029930),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974b87a),
	.w1(32'h39dfbb31),
	.w2(32'h38bf2490),
	.w3(32'hba1970e0),
	.w4(32'hb9a397e3),
	.w5(32'hb93a2bf6),
	.w6(32'hba183041),
	.w7(32'hb9381630),
	.w8(32'hb9f2ba1e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e6ebb),
	.w1(32'h3a2034fc),
	.w2(32'h3a6f2c34),
	.w3(32'h391510d7),
	.w4(32'h39c0e41f),
	.w5(32'hba116c2e),
	.w6(32'h39a5fb01),
	.w7(32'hb9b621dd),
	.w8(32'hba05a1bf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f6caa),
	.w1(32'h38b37e82),
	.w2(32'h39098b62),
	.w3(32'hba271e61),
	.w4(32'h393ef8d1),
	.w5(32'h392f5f57),
	.w6(32'h38ce6bbf),
	.w7(32'h37dd42a5),
	.w8(32'hb8a24697),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac0668),
	.w1(32'hb9d9e7d9),
	.w2(32'hb91e765a),
	.w3(32'hb99e771f),
	.w4(32'h3987646f),
	.w5(32'h39b8e975),
	.w6(32'hb993fd66),
	.w7(32'hb98bcaec),
	.w8(32'h38507c70),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2da58),
	.w1(32'hba3eae7c),
	.w2(32'hba38067e),
	.w3(32'hb7d9b244),
	.w4(32'hb9a5dce0),
	.w5(32'hba0a2866),
	.w6(32'hb7c2a46e),
	.w7(32'hb9e5d674),
	.w8(32'h39116d4e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95dee20),
	.w1(32'hb97cf391),
	.w2(32'hb955a945),
	.w3(32'hb9b37f73),
	.w4(32'hba4e4068),
	.w5(32'hba619c55),
	.w6(32'hba946fff),
	.w7(32'hba1098ce),
	.w8(32'hb990b99c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39095dab),
	.w1(32'hb9120b34),
	.w2(32'hb97c6627),
	.w3(32'hb94b9419),
	.w4(32'h38a1c3f6),
	.w5(32'hb8bf8daf),
	.w6(32'hb8ea72a6),
	.w7(32'hb8a5d216),
	.w8(32'hb8f6f86c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d2dd1),
	.w1(32'hb87442df),
	.w2(32'hb82b0e2c),
	.w3(32'hb83f6498),
	.w4(32'h38916ae5),
	.w5(32'h382fa586),
	.w6(32'hb8cf51f4),
	.w7(32'hb92bf705),
	.w8(32'hb99601f8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d15dc),
	.w1(32'hb80935c1),
	.w2(32'hb928db72),
	.w3(32'h399791dc),
	.w4(32'h39bd243b),
	.w5(32'h388f62a7),
	.w6(32'hba259d76),
	.w7(32'hb9a6c1a2),
	.w8(32'hb9884238),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a685f),
	.w1(32'hba0d01cf),
	.w2(32'h3a46ad33),
	.w3(32'hba239951),
	.w4(32'hba8e3336),
	.w5(32'hb7fe4531),
	.w6(32'h378b2d9f),
	.w7(32'h384f3d15),
	.w8(32'h38d404e6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c0114),
	.w1(32'h39c5d7d1),
	.w2(32'h39a08b81),
	.w3(32'h3a3ff56d),
	.w4(32'h3a53f078),
	.w5(32'h39c69d27),
	.w6(32'h3a873df8),
	.w7(32'h3a15c96e),
	.w8(32'h3877c8d6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39333432),
	.w1(32'hb979215b),
	.w2(32'h37a44f29),
	.w3(32'h39e5ff94),
	.w4(32'h39f1449b),
	.w5(32'h39d42e7c),
	.w6(32'h389b0021),
	.w7(32'hb8695a7f),
	.w8(32'hb8a98efd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc239c),
	.w1(32'h39dc16d3),
	.w2(32'h383cf183),
	.w3(32'h39cb711d),
	.w4(32'h3a77d735),
	.w5(32'h39fabe09),
	.w6(32'h3a819481),
	.w7(32'h3925b487),
	.w8(32'h376bb2de),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f6a60),
	.w1(32'h3a19a282),
	.w2(32'h39ab5701),
	.w3(32'hb98d4dad),
	.w4(32'h39155d32),
	.w5(32'h39249ce8),
	.w6(32'hba0fff14),
	.w7(32'hb988692b),
	.w8(32'hb9e93d91),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e483da),
	.w1(32'h36b99d77),
	.w2(32'h39692346),
	.w3(32'hb8d0acbf),
	.w4(32'h37477531),
	.w5(32'h398280e9),
	.w6(32'hba00374a),
	.w7(32'hb90ec1ed),
	.w8(32'hb9a78596),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981e539),
	.w1(32'h3a21e229),
	.w2(32'h39c61b7a),
	.w3(32'hb9308e48),
	.w4(32'h39bd8c56),
	.w5(32'h399beaf9),
	.w6(32'h3a060578),
	.w7(32'h39a20975),
	.w8(32'h36ed4807),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ca14b),
	.w1(32'hba51999d),
	.w2(32'hb9bd67d4),
	.w3(32'h3943d06d),
	.w4(32'hba27539f),
	.w5(32'hb9a769e1),
	.w6(32'hba1b846a),
	.w7(32'hb9679b47),
	.w8(32'hb85bf97f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897dbe5),
	.w1(32'hb99779ef),
	.w2(32'h3918d43b),
	.w3(32'h3707b2f0),
	.w4(32'h3946b05b),
	.w5(32'hb8f89f6c),
	.w6(32'h39e7e7ff),
	.w7(32'h39438d3c),
	.w8(32'h39259137),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c99db6),
	.w1(32'h38e2c8a0),
	.w2(32'h3686162d),
	.w3(32'h37808e52),
	.w4(32'h395595de),
	.w5(32'h398100d2),
	.w6(32'hb89e5fc7),
	.w7(32'hb8ee62bc),
	.w8(32'hb93b6e46),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d9238),
	.w1(32'h3a18c4f4),
	.w2(32'hb94aaa0d),
	.w3(32'h39d983cd),
	.w4(32'h3a49133e),
	.w5(32'h39a74db9),
	.w6(32'h39cc5f0b),
	.w7(32'hb93daa25),
	.w8(32'h38221aba),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a34c7),
	.w1(32'h3a0bb9ea),
	.w2(32'hb986d38a),
	.w3(32'h3a64748a),
	.w4(32'h38a30202),
	.w5(32'h382c65b1),
	.w6(32'hbaeaad59),
	.w7(32'hbac15ffc),
	.w8(32'hbaaa5024),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af5847),
	.w1(32'h39317084),
	.w2(32'hb8d890cc),
	.w3(32'h394e3338),
	.w4(32'hb81f8f17),
	.w5(32'h3927f60c),
	.w6(32'hba7cb2dd),
	.w7(32'hba59a1aa),
	.w8(32'hba60ba58),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d02249),
	.w1(32'hba510151),
	.w2(32'hb9cd681e),
	.w3(32'h3a3cd0aa),
	.w4(32'hba91ba3e),
	.w5(32'hba62dc84),
	.w6(32'hba1f978c),
	.w7(32'hba4326ae),
	.w8(32'hbaa1c23a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf859f),
	.w1(32'hbb09f578),
	.w2(32'hbacd30a2),
	.w3(32'h3a84a700),
	.w4(32'hb9144b20),
	.w5(32'hba6f95ff),
	.w6(32'h3978ec8c),
	.w7(32'hba5a0c38),
	.w8(32'hba341a26),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984b7d0),
	.w1(32'hb90932bc),
	.w2(32'h3924c508),
	.w3(32'hb66659d0),
	.w4(32'hb8bb1f00),
	.w5(32'h3927a496),
	.w6(32'hb8c3634a),
	.w7(32'hb93c9505),
	.w8(32'hb922bd5b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902f89f),
	.w1(32'hb9e91486),
	.w2(32'hba24a0a9),
	.w3(32'h38ea0666),
	.w4(32'hb9a8780a),
	.w5(32'hba003255),
	.w6(32'hb997b6d6),
	.w7(32'hb9c913d6),
	.w8(32'hb9d4ec40),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af19d4),
	.w1(32'hba207741),
	.w2(32'hba12a579),
	.w3(32'hb95048bf),
	.w4(32'hba33bfc6),
	.w5(32'hba2904e0),
	.w6(32'hb9dcd53b),
	.w7(32'hb9f129eb),
	.w8(32'hb9ec5693),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba106031),
	.w1(32'hbadb2374),
	.w2(32'hba95b4d4),
	.w3(32'hba4b0bb9),
	.w4(32'hb67d406b),
	.w5(32'h3aa5b715),
	.w6(32'hba523d6d),
	.w7(32'hb9e8e280),
	.w8(32'h39a0e3a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15041b),
	.w1(32'hb9973fb9),
	.w2(32'hb9efdfce),
	.w3(32'h3a737fd2),
	.w4(32'hb900eb4b),
	.w5(32'hb982a041),
	.w6(32'h360759f8),
	.w7(32'hb9c907f7),
	.w8(32'hb9c5d6c1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e37b70),
	.w1(32'hb9d7d8a7),
	.w2(32'hba1e19a0),
	.w3(32'h3a44748d),
	.w4(32'h3a943da1),
	.w5(32'hb75b87c4),
	.w6(32'h3a81f055),
	.w7(32'h39e9a468),
	.w8(32'hb98ceccf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c19bcd),
	.w1(32'h3911e9d0),
	.w2(32'h38f20246),
	.w3(32'h39135a8c),
	.w4(32'h391d2b3a),
	.w5(32'hb90cff31),
	.w6(32'h38f5fb11),
	.w7(32'h37546c0b),
	.w8(32'hba16029a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b80ec6),
	.w1(32'hba360196),
	.w2(32'hb902533e),
	.w3(32'hb9832af9),
	.w4(32'hb966bda4),
	.w5(32'hb984488d),
	.w6(32'hba238eb4),
	.w7(32'hb91ddfb5),
	.w8(32'h39055ca2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968e2fe),
	.w1(32'hba4021ea),
	.w2(32'hba174d0b),
	.w3(32'hba2fed6c),
	.w4(32'hba151128),
	.w5(32'hba095b0d),
	.w6(32'hba418dfe),
	.w7(32'hb9e548cd),
	.w8(32'hb9a03920),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d46b95),
	.w1(32'hb98a09a5),
	.w2(32'h39cbf8a4),
	.w3(32'hb88a664c),
	.w4(32'hb93ab7db),
	.w5(32'hb88528f6),
	.w6(32'h38732bea),
	.w7(32'h39790072),
	.w8(32'hb928373e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8b577),
	.w1(32'h3a1f160e),
	.w2(32'h39f79336),
	.w3(32'h3835a388),
	.w4(32'h39eeba0e),
	.w5(32'h39450cc4),
	.w6(32'h3a3a0218),
	.w7(32'h39f239a6),
	.w8(32'h397dcef1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f6f2d),
	.w1(32'hb91d992a),
	.w2(32'hb927a180),
	.w3(32'h39833c94),
	.w4(32'hb73c2410),
	.w5(32'h387fac4d),
	.w6(32'hb8f01b7f),
	.w7(32'hb8aef71a),
	.w8(32'hb9169bfc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f9c38),
	.w1(32'h3978570b),
	.w2(32'h38d3a630),
	.w3(32'h390ef8fa),
	.w4(32'h3a192d07),
	.w5(32'h39722590),
	.w6(32'h3a10d5be),
	.w7(32'h3970fe42),
	.w8(32'h39348525),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38891b76),
	.w1(32'h3809398c),
	.w2(32'hb95d9c70),
	.w3(32'h398d983d),
	.w4(32'hb90292b0),
	.w5(32'h3911e204),
	.w6(32'hba0c9b72),
	.w7(32'hba0648c1),
	.w8(32'hb98e66c6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e020b9),
	.w1(32'hba1113b4),
	.w2(32'hb9952694),
	.w3(32'hb90f4664),
	.w4(32'h3909dead),
	.w5(32'h39cbbce7),
	.w6(32'hba94d1c6),
	.w7(32'hbac641f8),
	.w8(32'hbac6724a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bdcb6),
	.w1(32'h3a3ca4a1),
	.w2(32'h39e04eb0),
	.w3(32'h37c001e4),
	.w4(32'h3a548a3a),
	.w5(32'h3a1417ee),
	.w6(32'h3a54b22c),
	.w7(32'h39d59451),
	.w8(32'h39ac16fa),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ba8f3),
	.w1(32'h39d7f075),
	.w2(32'h399a4bcb),
	.w3(32'h3a48821e),
	.w4(32'h394c60e0),
	.w5(32'h38eaa478),
	.w6(32'h39595895),
	.w7(32'hb8eb9dc7),
	.w8(32'hb902cfe0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997d842),
	.w1(32'hba349f73),
	.w2(32'h38ab8758),
	.w3(32'h3927028e),
	.w4(32'hb9a5c744),
	.w5(32'h39ee1ca9),
	.w6(32'hb9a9eb74),
	.w7(32'hb9a2951f),
	.w8(32'h39557acc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39869ba7),
	.w1(32'hba86830f),
	.w2(32'hb85fd26d),
	.w3(32'h3a95d644),
	.w4(32'hba541a6c),
	.w5(32'hb95809c0),
	.w6(32'hba402a9c),
	.w7(32'hba1ad6bf),
	.w8(32'hb9d1826c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b08ad),
	.w1(32'hb9911797),
	.w2(32'hba5a4583),
	.w3(32'h3988e523),
	.w4(32'hb8222103),
	.w5(32'hba07b15a),
	.w6(32'hba24aa74),
	.w7(32'hba0089ed),
	.w8(32'hba18dd99),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f9ea3),
	.w1(32'hb9ae6f7a),
	.w2(32'hba066d4b),
	.w3(32'hb731cf4a),
	.w4(32'hb9070718),
	.w5(32'hb9f30d9b),
	.w6(32'hba21124e),
	.w7(32'hb9bf439f),
	.w8(32'hba23ccd6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a13ef),
	.w1(32'h3a15296a),
	.w2(32'h39b732b4),
	.w3(32'hba228b01),
	.w4(32'hb9df2424),
	.w5(32'hba002acc),
	.w6(32'hba806d19),
	.w7(32'hba108582),
	.w8(32'hba988ae7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c48168),
	.w1(32'h394db2e8),
	.w2(32'h3998f231),
	.w3(32'hb8f8f6ba),
	.w4(32'h39c4472d),
	.w5(32'h39a10d6c),
	.w6(32'h39c4a111),
	.w7(32'h396ffc6d),
	.w8(32'h389cc125),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ff178),
	.w1(32'hba0031c2),
	.w2(32'hb9da8a73),
	.w3(32'h3987fe82),
	.w4(32'hb93bfc7e),
	.w5(32'hb9bf570f),
	.w6(32'hb9cf8aae),
	.w7(32'hb984e9ad),
	.w8(32'hb9bd593a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9937666),
	.w1(32'hb98a4299),
	.w2(32'hb9308c35),
	.w3(32'hb9269683),
	.w4(32'hb881ea7e),
	.w5(32'h37ff70f2),
	.w6(32'hb8e3dcce),
	.w7(32'hb8c7c8dd),
	.w8(32'hb8f18d32),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9898117),
	.w1(32'hba039e1e),
	.w2(32'hb9802a07),
	.w3(32'h37ce8708),
	.w4(32'h389171f9),
	.w5(32'h38c0abe9),
	.w6(32'hb92b6d9a),
	.w7(32'hb98f3f95),
	.w8(32'hb9c042b0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9865a81),
	.w1(32'h39144272),
	.w2(32'h38339ae0),
	.w3(32'h37e7de54),
	.w4(32'h39768a08),
	.w5(32'h3917c91a),
	.w6(32'h3a377aab),
	.w7(32'h394711c3),
	.w8(32'h392cad05),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991a7d8),
	.w1(32'hba94c6d0),
	.w2(32'h39516d9c),
	.w3(32'h3a15f5f5),
	.w4(32'h397abe24),
	.w5(32'h384faea2),
	.w6(32'h3765a71e),
	.w7(32'hb9132cda),
	.w8(32'hb8acf02b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a856833),
	.w1(32'hba66e535),
	.w2(32'hba8ef4ec),
	.w3(32'hb89c02e5),
	.w4(32'h382c0210),
	.w5(32'hb9183c15),
	.w6(32'hb9ac346b),
	.w7(32'hba16102a),
	.w8(32'hb9d22ee4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba424292),
	.w1(32'h38354fd9),
	.w2(32'hb886c50f),
	.w3(32'hba003295),
	.w4(32'h389ae2b9),
	.w5(32'hb902692a),
	.w6(32'hba6599ea),
	.w7(32'hb9b6072c),
	.w8(32'hb9ff609f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85676aa),
	.w1(32'h3a18d40e),
	.w2(32'h38dd0737),
	.w3(32'hb9a3a896),
	.w4(32'h3a225182),
	.w5(32'hb9809b92),
	.w6(32'hb725258a),
	.w7(32'hb91bad80),
	.w8(32'hba8c3e01),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ccd91),
	.w1(32'hb9d4280a),
	.w2(32'hb9ebc536),
	.w3(32'hba6579a5),
	.w4(32'h38ac3f38),
	.w5(32'hb9c9ecca),
	.w6(32'hb96e2748),
	.w7(32'hb919e916),
	.w8(32'hb974b61c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9049867),
	.w1(32'hba19b7c6),
	.w2(32'hba79028b),
	.w3(32'hb95ea359),
	.w4(32'hba052ada),
	.w5(32'hba2a62aa),
	.w6(32'hba509118),
	.w7(32'hba3d052f),
	.w8(32'hba09eefe),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edbc57),
	.w1(32'hb886b946),
	.w2(32'hb8ef2484),
	.w3(32'h396372fc),
	.w4(32'h393f01c5),
	.w5(32'hb65fcb86),
	.w6(32'h3a403be5),
	.w7(32'h3940b1a0),
	.w8(32'h37a29bd2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c5a9c),
	.w1(32'hb9f283e5),
	.w2(32'hb99af868),
	.w3(32'h3915d77d),
	.w4(32'hb9782e96),
	.w5(32'hb95286a0),
	.w6(32'hb82218c5),
	.w7(32'hb90198be),
	.w8(32'h3882e096),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e0d7aa),
	.w1(32'h3a17c3d6),
	.w2(32'h39f2b462),
	.w3(32'hb8dd3e9a),
	.w4(32'h39a31a08),
	.w5(32'h38fbb2e6),
	.w6(32'h39d80eca),
	.w7(32'h393d6652),
	.w8(32'h38f5b95a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e694b4),
	.w1(32'hb92c1e00),
	.w2(32'hb98e6e99),
	.w3(32'h3989fe43),
	.w4(32'hb994ccb3),
	.w5(32'hb98738e2),
	.w6(32'hb9e76ba3),
	.w7(32'hba0f1736),
	.w8(32'hb98aea48),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928b544),
	.w1(32'hb9a97315),
	.w2(32'hb96c76a1),
	.w3(32'hb9f2e339),
	.w4(32'hb9a8b66c),
	.w5(32'hb922f811),
	.w6(32'hb9e0440b),
	.w7(32'hb9be5471),
	.w8(32'hb8e2d78d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a0786),
	.w1(32'hb9dfd3bf),
	.w2(32'hb81ea0b6),
	.w3(32'hb8830469),
	.w4(32'hb9f7a6fd),
	.w5(32'hba59d24b),
	.w6(32'hba35109f),
	.w7(32'hb9cc55fa),
	.w8(32'hba04a3b1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b133f8),
	.w1(32'hb9a4a529),
	.w2(32'hb9af1ad7),
	.w3(32'hba4117dd),
	.w4(32'hb7962d84),
	.w5(32'hb90d9a8d),
	.w6(32'hb9726eb9),
	.w7(32'hb904770c),
	.w8(32'hb949b34e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82dd5e2),
	.w1(32'h399a19e8),
	.w2(32'h3844a7c1),
	.w3(32'hb82783b8),
	.w4(32'hb90539a9),
	.w5(32'hb9b43d08),
	.w6(32'h3978b388),
	.w7(32'hb8abfc12),
	.w8(32'hba3d18ff),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9432aa5),
	.w1(32'hba11fd67),
	.w2(32'hba097cae),
	.w3(32'h39abd610),
	.w4(32'h39cc6798),
	.w5(32'hb94030c1),
	.w6(32'hb8fd7c57),
	.w7(32'hb98dbadc),
	.w8(32'hba1d9f79),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e58a3c),
	.w1(32'hb91c57c0),
	.w2(32'hb8f193e9),
	.w3(32'hb941e2c5),
	.w4(32'h391d11f0),
	.w5(32'h394e9c72),
	.w6(32'hb9cebde6),
	.w7(32'hb92690fa),
	.w8(32'hb99949f7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a42f3),
	.w1(32'h39378f94),
	.w2(32'hb9cda3c5),
	.w3(32'h39fe882e),
	.w4(32'hb9733035),
	.w5(32'hba4d8e43),
	.w6(32'h388bd9b4),
	.w7(32'hba29fca5),
	.w8(32'hb9d6798c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f05c26),
	.w1(32'h3a0fdca0),
	.w2(32'h3a050bab),
	.w3(32'h391d5ade),
	.w4(32'h3a0c74b3),
	.w5(32'h39615083),
	.w6(32'h3a009669),
	.w7(32'h3989625e),
	.w8(32'h37d18e2c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5b6c),
	.w1(32'hba835090),
	.w2(32'hbac45899),
	.w3(32'h38cc3f6c),
	.w4(32'hba5e3c13),
	.w5(32'hbab44e3d),
	.w6(32'hba8dc797),
	.w7(32'hba8f335b),
	.w8(32'hba834f05),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3da8b),
	.w1(32'h3959e365),
	.w2(32'h39b201dc),
	.w3(32'hb98a6bab),
	.w4(32'h39ac733d),
	.w5(32'hb8fe4c51),
	.w6(32'h38c4fcc1),
	.w7(32'h38ecc56d),
	.w8(32'hb98bf1b2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdaf54),
	.w1(32'h3a606deb),
	.w2(32'h39b11882),
	.w3(32'h38e84364),
	.w4(32'h399b1733),
	.w5(32'hb9cf05ef),
	.w6(32'hb7cdec7b),
	.w7(32'h38197735),
	.w8(32'hb9abf869),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a82fdc),
	.w1(32'hb9acfbb9),
	.w2(32'hba086c61),
	.w3(32'h3723b628),
	.w4(32'hb90fc9fc),
	.w5(32'hb9288a73),
	.w6(32'hb9a9f7ca),
	.w7(32'hb9c14cf2),
	.w8(32'hb922c801),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c620f),
	.w1(32'hba90aa60),
	.w2(32'hba09058b),
	.w3(32'h3a0e32ee),
	.w4(32'hb91dbd0f),
	.w5(32'hb94df292),
	.w6(32'hba985b73),
	.w7(32'hba80bd95),
	.w8(32'hba903293),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b0375),
	.w1(32'h3a23a721),
	.w2(32'h3a6c3411),
	.w3(32'h398116d7),
	.w4(32'h3aac846d),
	.w5(32'h3a517753),
	.w6(32'h3a8ceeda),
	.w7(32'h3a77d449),
	.w8(32'h39ad2420),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49c64b),
	.w1(32'hba86c65b),
	.w2(32'hba9459c9),
	.w3(32'h3a8b61bb),
	.w4(32'h39681997),
	.w5(32'hb92c8ee9),
	.w6(32'h3a2e73f0),
	.w7(32'hba649cf0),
	.w8(32'hb9d958c3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980ebae),
	.w1(32'hb9914338),
	.w2(32'h3965dcd0),
	.w3(32'hb9a51176),
	.w4(32'hba678929),
	.w5(32'hba2e588a),
	.w6(32'hb9c60920),
	.w7(32'hb909d175),
	.w8(32'h398a1e02),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f2c67),
	.w1(32'h3a9cf2fc),
	.w2(32'hb9065b43),
	.w3(32'hb9bd036c),
	.w4(32'h3993113c),
	.w5(32'h388666f9),
	.w6(32'hba51bb24),
	.w7(32'hb95d6dd8),
	.w8(32'hba76e709),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a910384),
	.w1(32'hba6f3406),
	.w2(32'hbab447fe),
	.w3(32'h3ae1d8e0),
	.w4(32'h381f5f03),
	.w5(32'hba0acfb5),
	.w6(32'h3a0fe895),
	.w7(32'hb9fae311),
	.w8(32'hb99b20fa),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba216208),
	.w1(32'hba18cc5a),
	.w2(32'hba4961f8),
	.w3(32'hba0625d9),
	.w4(32'h38fcf469),
	.w5(32'hb9e7fa5c),
	.w6(32'hb955737f),
	.w7(32'hb8dc84d1),
	.w8(32'hb9b599be),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab43868),
	.w1(32'h393e8209),
	.w2(32'hba8c1664),
	.w3(32'h3aaca342),
	.w4(32'h3a28b4d1),
	.w5(32'h3a3f96ea),
	.w6(32'h398d3a5e),
	.w7(32'hba0d2a19),
	.w8(32'hba1da69d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36211ed6),
	.w1(32'h39ab4bcc),
	.w2(32'h3a00c5e9),
	.w3(32'h394e088b),
	.w4(32'h39e76107),
	.w5(32'h3a383cf9),
	.w6(32'h3940d472),
	.w7(32'hb89f9217),
	.w8(32'h38aeb8fe),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383067b4),
	.w1(32'h396678e6),
	.w2(32'h3830c9af),
	.w3(32'hb80db40e),
	.w4(32'h39f248ce),
	.w5(32'h39409e1a),
	.w6(32'h3952a969),
	.w7(32'hb8549102),
	.w8(32'hb8c32742),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a17d5b),
	.w1(32'hb99c0d2f),
	.w2(32'hb9b55941),
	.w3(32'h392a6fef),
	.w4(32'h39029406),
	.w5(32'hb88afa95),
	.w6(32'hb9d32f5d),
	.w7(32'hb99cd855),
	.w8(32'hb9ad64d0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913638e),
	.w1(32'hb92bdd86),
	.w2(32'hba4b223c),
	.w3(32'h37b25247),
	.w4(32'hb912c79b),
	.w5(32'hb9dea7ac),
	.w6(32'hba35b43e),
	.w7(32'hba30c2cc),
	.w8(32'hba1fad3c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111790),
	.w1(32'h39a774ae),
	.w2(32'hba628f7f),
	.w3(32'hb9e83177),
	.w4(32'hb9eec308),
	.w5(32'hba742315),
	.w6(32'hba924f99),
	.w7(32'hba9f4ba5),
	.w8(32'hbab19fd2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c54e37),
	.w1(32'h37d8acda),
	.w2(32'hb8e9511b),
	.w3(32'hb9013caf),
	.w4(32'hb894e8e3),
	.w5(32'h3a079aba),
	.w6(32'hb9f3321b),
	.w7(32'hb9b23012),
	.w8(32'hb9a6c9a4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8daca01),
	.w1(32'h39d539ec),
	.w2(32'h3a82fd56),
	.w3(32'hb8ce40ba),
	.w4(32'h39dbd9d8),
	.w5(32'h3ab86885),
	.w6(32'hba762d76),
	.w7(32'hba859570),
	.w8(32'hba1d3128),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21fc16),
	.w1(32'hb9e0b639),
	.w2(32'hb9eb14e4),
	.w3(32'h3a48b761),
	.w4(32'h38a8efc2),
	.w5(32'h3831c63c),
	.w6(32'h38489163),
	.w7(32'hb7498fe2),
	.w8(32'hb9504a02),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39420c8d),
	.w1(32'hb5faa7e2),
	.w2(32'hb9af839d),
	.w3(32'h39a1d031),
	.w4(32'h39e281fa),
	.w5(32'hb9f6aa20),
	.w6(32'h395ccd7b),
	.w7(32'hb7e6a19f),
	.w8(32'hb9da8ae9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371481cf),
	.w1(32'h3a3ecd73),
	.w2(32'h399e34e0),
	.w3(32'hb8b3d158),
	.w4(32'h3a2fc42a),
	.w5(32'h3a3aefcc),
	.w6(32'hb9f28c61),
	.w7(32'hba0c752b),
	.w8(32'hb96a6ef0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a24c2e),
	.w1(32'hb9ca7980),
	.w2(32'hba2853ba),
	.w3(32'h38342992),
	.w4(32'hb89b0c91),
	.w5(32'hb9763799),
	.w6(32'hb9a6f600),
	.w7(32'hb9af59cf),
	.w8(32'hb987f4f1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4f62),
	.w1(32'hb95d30c2),
	.w2(32'hb9c174b1),
	.w3(32'hb99351d5),
	.w4(32'h37b7c2b6),
	.w5(32'hb8e7d8a7),
	.w6(32'hb95d3b8b),
	.w7(32'hb918eb31),
	.w8(32'hb8e2783b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bab600),
	.w1(32'hb9098fc6),
	.w2(32'hb9a690b3),
	.w3(32'hb92d7e92),
	.w4(32'h39558784),
	.w5(32'hb7b97423),
	.w6(32'hb8818bbe),
	.w7(32'hb88146b0),
	.w8(32'hb72ddbda),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4320c),
	.w1(32'h3a3dea8e),
	.w2(32'h39b063fd),
	.w3(32'hb96f71c2),
	.w4(32'h3923d42e),
	.w5(32'h3a5aad55),
	.w6(32'hba3ca3c6),
	.w7(32'hba803f7e),
	.w8(32'hba2934b2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391791dc),
	.w1(32'h39920466),
	.w2(32'h39a9d817),
	.w3(32'h3a284c80),
	.w4(32'hb93334b2),
	.w5(32'h39e3e169),
	.w6(32'hb9692ff0),
	.w7(32'h3811ba26),
	.w8(32'h39297c29),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fea9d2),
	.w1(32'hb89764fd),
	.w2(32'hba237cbb),
	.w3(32'h3a10497d),
	.w4(32'h39d8556e),
	.w5(32'hb9ac3eb6),
	.w6(32'hb842b7b1),
	.w7(32'hb9858318),
	.w8(32'hba2918f9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8bdd4),
	.w1(32'hba4df450),
	.w2(32'hba3dc4b9),
	.w3(32'h39994b84),
	.w4(32'hb94adb23),
	.w5(32'hb9c05119),
	.w6(32'hb914e486),
	.w7(32'hb99f7fa0),
	.w8(32'hb883e738),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97238e8),
	.w1(32'h3891d704),
	.w2(32'hb9342dca),
	.w3(32'hb9bd66c7),
	.w4(32'hb91b976c),
	.w5(32'hb91b9ba5),
	.w6(32'hba167fcb),
	.w7(32'hb9bc8e7c),
	.w8(32'hba1a62f4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d7c47),
	.w1(32'h3aae85e3),
	.w2(32'h3af15f76),
	.w3(32'hb8f9868e),
	.w4(32'hb9d45146),
	.w5(32'h3929bbfa),
	.w6(32'hb962c806),
	.w7(32'hba3607a2),
	.w8(32'hba426236),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5b7bd),
	.w1(32'h39882344),
	.w2(32'hba1ac9a6),
	.w3(32'h3a69437b),
	.w4(32'h39256531),
	.w5(32'hba1d36a3),
	.w6(32'h39c7a921),
	.w7(32'hb9a45920),
	.w8(32'hb9fdc643),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f2a69),
	.w1(32'hb9a9b042),
	.w2(32'hb9ccff65),
	.w3(32'h38d77829),
	.w4(32'h383171a2),
	.w5(32'hb8e751d8),
	.w6(32'hb9873c64),
	.w7(32'hb971dbe4),
	.w8(32'hb958f485),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9970e0c),
	.w1(32'hba79581e),
	.w2(32'h3b9a7e1e),
	.w3(32'hb8b892b5),
	.w4(32'h3ac21d4b),
	.w5(32'h3b102058),
	.w6(32'h3a47b5c3),
	.w7(32'h3ad5d6b7),
	.w8(32'h3ac7752c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38f9b5),
	.w1(32'h3a57d041),
	.w2(32'h3a2e439d),
	.w3(32'h3a9da16f),
	.w4(32'h3a9afb2b),
	.w5(32'h3a51f130),
	.w6(32'h3ac7df4a),
	.w7(32'h39c2aee0),
	.w8(32'h3b040c49),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18f50c),
	.w1(32'hb998a222),
	.w2(32'hbbdfdbd3),
	.w3(32'h3aadbf80),
	.w4(32'hba599054),
	.w5(32'hbc0d0943),
	.w6(32'hbb6629c4),
	.w7(32'h3aa4193e),
	.w8(32'h3bf1decb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa5ae),
	.w1(32'hb8f29d16),
	.w2(32'hbb75e7d4),
	.w3(32'hba5469d3),
	.w4(32'hbb1f0338),
	.w5(32'hbb104e09),
	.w6(32'hba495298),
	.w7(32'hbb1039df),
	.w8(32'h3a721c61),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae01ea2),
	.w1(32'h3b0f9df6),
	.w2(32'h3b7a7414),
	.w3(32'hba45f29b),
	.w4(32'h3b90d9ed),
	.w5(32'h3a6179f4),
	.w6(32'h3ad0760d),
	.w7(32'hba91076f),
	.w8(32'h3b0c5698),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e28b7),
	.w1(32'h3bb5f09b),
	.w2(32'hbb076d7e),
	.w3(32'hbaa0eb0a),
	.w4(32'hbaccbb81),
	.w5(32'hba5f1d95),
	.w6(32'h3b6e0465),
	.w7(32'hbb0a87f8),
	.w8(32'hb9ede27f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617dd7),
	.w1(32'hbb975bd8),
	.w2(32'h3cdf36ff),
	.w3(32'h3ab4086c),
	.w4(32'h39b31a50),
	.w5(32'h3ca60828),
	.w6(32'h3ba3f555),
	.w7(32'h3c833f8c),
	.w8(32'hbb20d67d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb348e),
	.w1(32'h3b0e1175),
	.w2(32'h3b0715fd),
	.w3(32'h3b8ddb28),
	.w4(32'h3b140d7e),
	.w5(32'h3b124e9f),
	.w6(32'h3b414e96),
	.w7(32'h3b6deea0),
	.w8(32'h3b33a02d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33d193),
	.w1(32'hbb423b3d),
	.w2(32'h3b905e2e),
	.w3(32'h3b10527d),
	.w4(32'hba83d7ec),
	.w5(32'h38afc29a),
	.w6(32'hba976406),
	.w7(32'h3b0b6e15),
	.w8(32'h37c7b548),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152274),
	.w1(32'hbab3358b),
	.w2(32'h398c11b3),
	.w3(32'hbb0c731d),
	.w4(32'h38246490),
	.w5(32'hba96edf3),
	.w6(32'hb9cf1d72),
	.w7(32'hba9c7599),
	.w8(32'h3aaefc81),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842ed2),
	.w1(32'hb8ee7e10),
	.w2(32'hb9b4f307),
	.w3(32'h3926c45a),
	.w4(32'h3a37cc1f),
	.w5(32'hba71da51),
	.w6(32'hb84a38a4),
	.w7(32'hbae5095a),
	.w8(32'hba0dbaf6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9957dc5),
	.w1(32'h3b4fef12),
	.w2(32'hb8aa9a3b),
	.w3(32'hb954e3ab),
	.w4(32'hba1e780f),
	.w5(32'hba11d52b),
	.w6(32'h3b0e6b98),
	.w7(32'hb9c9ea7c),
	.w8(32'h3aa40b31),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ab9c4),
	.w1(32'hba327ec1),
	.w2(32'hbad9026b),
	.w3(32'hb89112d5),
	.w4(32'hbad86922),
	.w5(32'hbb3c5627),
	.w6(32'h3ab8d39b),
	.w7(32'hbb29953d),
	.w8(32'hb9abe353),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eb0bef),
	.w1(32'h3aeea1a3),
	.w2(32'hbafc228b),
	.w3(32'h3ae70860),
	.w4(32'hbbb2b6e3),
	.w5(32'hba2f4195),
	.w6(32'h3b5ad496),
	.w7(32'hbaa60ee5),
	.w8(32'h3a581574),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03dbf2),
	.w1(32'hbae2f92a),
	.w2(32'hb9729fdf),
	.w3(32'h3ad6cdc7),
	.w4(32'h3a1dd3f7),
	.w5(32'hba8fe802),
	.w6(32'hb9e0662c),
	.w7(32'hbb0f604a),
	.w8(32'hba54e15c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae143aa),
	.w1(32'hbb576abc),
	.w2(32'hbc044355),
	.w3(32'hbaa0eb57),
	.w4(32'hbb278059),
	.w5(32'hbbbae9a1),
	.w6(32'hbb921d23),
	.w7(32'hbbc10fff),
	.w8(32'h3a466c44),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bac468),
	.w1(32'h3ae38976),
	.w2(32'h3bb85f74),
	.w3(32'hb9a0fa23),
	.w4(32'hbc360fa7),
	.w5(32'h3c149b24),
	.w6(32'h3bf988d4),
	.w7(32'hbb938e4f),
	.w8(32'h3ae0971e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a7b4),
	.w1(32'hba8df950),
	.w2(32'hbaf73b92),
	.w3(32'h3bdf088d),
	.w4(32'h3a5566eb),
	.w5(32'hba23b4d1),
	.w6(32'h394074b3),
	.w7(32'hbaff70b4),
	.w8(32'hba437ef9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c9b35),
	.w1(32'h3a956235),
	.w2(32'h3bf661c8),
	.w3(32'h39adda54),
	.w4(32'h3b235792),
	.w5(32'h3b628d8f),
	.w6(32'h3b72ebee),
	.w7(32'h3bd28db0),
	.w8(32'h3bef4518),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3374),
	.w1(32'h3b39cb55),
	.w2(32'h3b12401d),
	.w3(32'h3ae574b3),
	.w4(32'hba9f96a2),
	.w5(32'h3922756d),
	.w6(32'h39a0ad8d),
	.w7(32'h392650ff),
	.w8(32'h3ade73d6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2ec8),
	.w1(32'hb9f0ddce),
	.w2(32'h3b55852a),
	.w3(32'hb9264d89),
	.w4(32'hb95f15ef),
	.w5(32'h3a92088d),
	.w6(32'hb8ea2948),
	.w7(32'h39eee101),
	.w8(32'h3a3f6d2b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fba4b),
	.w1(32'hba68a42e),
	.w2(32'hbac14832),
	.w3(32'hb8b378f4),
	.w4(32'hba29bd59),
	.w5(32'hba58e2fc),
	.w6(32'hba265d13),
	.w7(32'hbad3bdb7),
	.w8(32'hb958daa0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8af7e),
	.w1(32'h3832daf3),
	.w2(32'h39a16f6e),
	.w3(32'h39306296),
	.w4(32'h38beeb6e),
	.w5(32'h3a409bc4),
	.w6(32'h3a1e7cf4),
	.w7(32'h3a75800a),
	.w8(32'h3a8a80a3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8922f),
	.w1(32'h3ac7d50f),
	.w2(32'h3850cdfb),
	.w3(32'h3a5aef9f),
	.w4(32'h3c72bbf5),
	.w5(32'hbbdb1ee3),
	.w6(32'hba9d8a0e),
	.w7(32'hbbbd2db6),
	.w8(32'hbb9c07f8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0756da),
	.w1(32'h3a55fe24),
	.w2(32'h39d6c85f),
	.w3(32'hbb3dee5f),
	.w4(32'h3a52573c),
	.w5(32'h3b08fa99),
	.w6(32'h3ab312d9),
	.w7(32'h3b253153),
	.w8(32'h3a9a56e0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7536e),
	.w1(32'hbaebd050),
	.w2(32'h39e7278d),
	.w3(32'h3b2211ca),
	.w4(32'hb9ceaf00),
	.w5(32'hba1b0fe7),
	.w6(32'h388ded12),
	.w7(32'hba18bcba),
	.w8(32'h3ad4d979),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0b0d7),
	.w1(32'hbabdde95),
	.w2(32'hbb70e652),
	.w3(32'h38a30bdb),
	.w4(32'hbb5381d9),
	.w5(32'hba7c64ea),
	.w6(32'hbb62d03d),
	.w7(32'hbb4298c3),
	.w8(32'h3a3db819),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264429),
	.w1(32'hbb52b533),
	.w2(32'hbb88fd5b),
	.w3(32'h39ccf50c),
	.w4(32'hbaf075fc),
	.w5(32'hbb691537),
	.w6(32'h3abd09c6),
	.w7(32'hbb01815e),
	.w8(32'hbac1178b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ab14c),
	.w1(32'hb93e41c4),
	.w2(32'hbb1b1807),
	.w3(32'hbb462a95),
	.w4(32'hb96f832e),
	.w5(32'hbad114c5),
	.w6(32'h39419528),
	.w7(32'hbab4e692),
	.w8(32'hba1d45ef),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884ecf8),
	.w1(32'h3b7a6a87),
	.w2(32'hbba46f9f),
	.w3(32'hba683f45),
	.w4(32'hbaf96a9f),
	.w5(32'hba9add0e),
	.w6(32'hbb072aeb),
	.w7(32'hbac6ab3a),
	.w8(32'hbaacbd9d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba808a7),
	.w1(32'h3aa65ae4),
	.w2(32'hba750f59),
	.w3(32'h3ab532aa),
	.w4(32'h3aed0fef),
	.w5(32'hba4cccdb),
	.w6(32'h3b5a35a9),
	.w7(32'hb8e75dd5),
	.w8(32'h3ab14930),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b406ae),
	.w1(32'h3a9e1354),
	.w2(32'h399db6eb),
	.w3(32'h3a77f1a2),
	.w4(32'hb9427bf3),
	.w5(32'h3821715c),
	.w6(32'h3ab95f52),
	.w7(32'h3a3ed2f3),
	.w8(32'h3b0e9856),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17b8a7),
	.w1(32'hba387c60),
	.w2(32'h39bf6395),
	.w3(32'h3accfa7b),
	.w4(32'hb7a746b0),
	.w5(32'hb9ab0a8b),
	.w6(32'h394da558),
	.w7(32'h39602c47),
	.w8(32'h397c28fd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cf731),
	.w1(32'hba881b0b),
	.w2(32'h39aa43ae),
	.w3(32'hba0955c6),
	.w4(32'h39969ed1),
	.w5(32'hba8a58cf),
	.w6(32'hb9072980),
	.w7(32'hba35208e),
	.w8(32'hb89bfd95),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47782a),
	.w1(32'h3b9aea2a),
	.w2(32'h3b45370e),
	.w3(32'hba41719a),
	.w4(32'h3b7caf74),
	.w5(32'h3b2d2bec),
	.w6(32'h3bbddbe1),
	.w7(32'hb9e62e0c),
	.w8(32'hbaa4f542),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389662),
	.w1(32'hbba08b2c),
	.w2(32'hbb3e5a97),
	.w3(32'hbba885b2),
	.w4(32'hbb9828a3),
	.w5(32'hbc011c1f),
	.w6(32'hbb84caee),
	.w7(32'hbb635f95),
	.w8(32'hbb9aec52),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f66e),
	.w1(32'h3ad0b722),
	.w2(32'hbaf90116),
	.w3(32'hbb305e7a),
	.w4(32'hbb348787),
	.w5(32'hbadb8228),
	.w6(32'hba958a29),
	.w7(32'hbb041079),
	.w8(32'h3a8ced36),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f354e),
	.w1(32'hba3538f1),
	.w2(32'hbb000fdb),
	.w3(32'hba1f8878),
	.w4(32'hba9a7adc),
	.w5(32'hbaf4d8fc),
	.w6(32'hb9fe4c1b),
	.w7(32'hb9f7d9df),
	.w8(32'hb964e42d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd57ac),
	.w1(32'hba8270e8),
	.w2(32'h39aab69f),
	.w3(32'hbaa1557a),
	.w4(32'hbb72a92e),
	.w5(32'h3b54ddbe),
	.w6(32'hba1e6320),
	.w7(32'hba729f29),
	.w8(32'hbb9faddd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce6afe),
	.w1(32'h3ae0adf3),
	.w2(32'h3b9274cf),
	.w3(32'hbb1c66a3),
	.w4(32'h392588ce),
	.w5(32'h3b192d68),
	.w6(32'h3aaa7694),
	.w7(32'h3b70f9a6),
	.w8(32'h3b70f403),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67ceb1),
	.w1(32'hb9a1be33),
	.w2(32'h3b01706b),
	.w3(32'h3afcd8dd),
	.w4(32'h3a15b409),
	.w5(32'h3a53db54),
	.w6(32'h3a672068),
	.w7(32'h3a693911),
	.w8(32'h3b0c31fc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f000),
	.w1(32'hbaa39c86),
	.w2(32'hb890d577),
	.w3(32'h39ff0f46),
	.w4(32'hbb4fb92a),
	.w5(32'hb8d8208c),
	.w6(32'hbaf82b3c),
	.w7(32'hbaf1a136),
	.w8(32'hbb274672),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37e0ad),
	.w1(32'h3a473421),
	.w2(32'hbb2dece3),
	.w3(32'hba574727),
	.w4(32'hb8e7d62c),
	.w5(32'hbb5da8bc),
	.w6(32'h3a390f57),
	.w7(32'hbaff2930),
	.w8(32'h3a0be987),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3356d1),
	.w1(32'h3b299533),
	.w2(32'hbb65f091),
	.w3(32'h39f2b074),
	.w4(32'hbb85b69d),
	.w5(32'hbb129ffe),
	.w6(32'hba1dc874),
	.w7(32'hbb51a75a),
	.w8(32'hbac41e78),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c800b0),
	.w1(32'h39e636a7),
	.w2(32'h3a5890d6),
	.w3(32'h3a458b37),
	.w4(32'h3b087a0c),
	.w5(32'h3960b682),
	.w6(32'h3a470218),
	.w7(32'h39a9e33b),
	.w8(32'hb8cdec98),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946e5ce),
	.w1(32'h3b3e1c08),
	.w2(32'hbac474ad),
	.w3(32'hba4daf74),
	.w4(32'hbb4a914b),
	.w5(32'hbb8b9d3b),
	.w6(32'h3873efbb),
	.w7(32'hbb0b4be3),
	.w8(32'h3b351c2d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8a2d1),
	.w1(32'h3bbe688d),
	.w2(32'hbba95070),
	.w3(32'h3af9d6c2),
	.w4(32'h3b74d3be),
	.w5(32'hba9d3f3c),
	.w6(32'h3931a2f0),
	.w7(32'hbb743db1),
	.w8(32'hbaa68520),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7690),
	.w1(32'hbb8f3a35),
	.w2(32'h3bbc1f00),
	.w3(32'h3a9ab631),
	.w4(32'h3b86ec6e),
	.w5(32'hb90d0dfc),
	.w6(32'hbb6444b8),
	.w7(32'h3a536886),
	.w8(32'h3b6f8b85),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a71986),
	.w1(32'hbb09d084),
	.w2(32'hbb9108fd),
	.w3(32'h3b14d9c6),
	.w4(32'hbc010e5d),
	.w5(32'hba67ca37),
	.w6(32'h3aab6909),
	.w7(32'hbb9ea57c),
	.w8(32'hbb3db3a1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d1ae0),
	.w1(32'hba8d88e6),
	.w2(32'hba4b6a9a),
	.w3(32'h3b0144cd),
	.w4(32'hb96a6332),
	.w5(32'hb9c990e4),
	.w6(32'hbabcd7df),
	.w7(32'h3ac37f2b),
	.w8(32'h3ae00109),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3788db9b),
	.w1(32'hba3274d7),
	.w2(32'hba3f74c4),
	.w3(32'h3a29bdd8),
	.w4(32'h3a64580e),
	.w5(32'hba5f8acf),
	.w6(32'h3a1ff562),
	.w7(32'hb9e23a21),
	.w8(32'hba51ac2e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efddca),
	.w1(32'hbb0e7b25),
	.w2(32'hbb29737c),
	.w3(32'hb99012e5),
	.w4(32'hba953e2d),
	.w5(32'hbb1cafa5),
	.w6(32'hbaa29429),
	.w7(32'hbb22d2ad),
	.w8(32'h39abc3cb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b268c),
	.w1(32'hb9167f76),
	.w2(32'hba59ef54),
	.w3(32'hba42e403),
	.w4(32'hb918bfd6),
	.w5(32'hbac4ebae),
	.w6(32'h3b2d0141),
	.w7(32'hb8d4aed2),
	.w8(32'h3b522f5b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a280d),
	.w1(32'h3bdccd46),
	.w2(32'h3b22a5df),
	.w3(32'h3b6abfb0),
	.w4(32'hbabe9fb1),
	.w5(32'hb95e4ec7),
	.w6(32'h39b50b6e),
	.w7(32'h36c64ed3),
	.w8(32'h3b95b446),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0f2af),
	.w1(32'hb9f7674a),
	.w2(32'hbbe5550d),
	.w3(32'h3b09fe53),
	.w4(32'h3a870b13),
	.w5(32'hbb6a6ad6),
	.w6(32'h3b03ba31),
	.w7(32'hbb5824cf),
	.w8(32'hbaaa897c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266595),
	.w1(32'hbae5a359),
	.w2(32'h3cacc9f4),
	.w3(32'h37dd105f),
	.w4(32'h3bc1f26d),
	.w5(32'h3c1d9ece),
	.w6(32'h3b8ed43d),
	.w7(32'h3c2b0b3c),
	.w8(32'hbb11caec),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e570b),
	.w1(32'hb9cc3af7),
	.w2(32'h3b0f1a82),
	.w3(32'hbb28dbf9),
	.w4(32'hbafb326d),
	.w5(32'h3ab81554),
	.w6(32'hba0eca60),
	.w7(32'h3ae1a550),
	.w8(32'h3a64f535),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48a039),
	.w1(32'h3ad79660),
	.w2(32'hbb2e23ee),
	.w3(32'h3ac40125),
	.w4(32'h3a462234),
	.w5(32'hbb634834),
	.w6(32'h3aa3ebe3),
	.w7(32'hbb0505d6),
	.w8(32'hb988ce0b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc3c59),
	.w1(32'h3be3d4f8),
	.w2(32'h3b1002f0),
	.w3(32'h39f0a572),
	.w4(32'h3be67fa4),
	.w5(32'h3af6090b),
	.w6(32'h3c0bed9d),
	.w7(32'h3ba2ae70),
	.w8(32'h3b76436e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4aed9),
	.w1(32'hbc1bd0a9),
	.w2(32'h3ca9ba6a),
	.w3(32'h3b99cf33),
	.w4(32'h3ace67ee),
	.w5(32'h3bffbce7),
	.w6(32'h3b5dcfdc),
	.w7(32'h3bdcc734),
	.w8(32'h3c06f957),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94340),
	.w1(32'h3ae4ff57),
	.w2(32'hbb8196fb),
	.w3(32'h3be27efd),
	.w4(32'hbb4cb7c2),
	.w5(32'hbb49915b),
	.w6(32'hb9910de0),
	.w7(32'hbafc400e),
	.w8(32'h3acdaf21),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2c19d),
	.w1(32'hba56f2cd),
	.w2(32'h3a89b983),
	.w3(32'h3adc9cfc),
	.w4(32'h38579b8f),
	.w5(32'h38717061),
	.w6(32'h39fa61e4),
	.w7(32'hb98d636e),
	.w8(32'h3a8fd870),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1df8f),
	.w1(32'hb9226d95),
	.w2(32'hbaffcc4c),
	.w3(32'h38f8a592),
	.w4(32'hbb3a0840),
	.w5(32'hba87c58d),
	.w6(32'hbb12c8ee),
	.w7(32'hbaf83dc3),
	.w8(32'hba616460),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d7f64),
	.w1(32'hb8d666a8),
	.w2(32'hba960243),
	.w3(32'h39e850dd),
	.w4(32'h37ae53e0),
	.w5(32'hbaa27a81),
	.w6(32'hba92cb5d),
	.w7(32'hbb1bc8ca),
	.w8(32'hb92dca6f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba149259),
	.w1(32'h3b9788e9),
	.w2(32'h39439d7d),
	.w3(32'hbb2cb6e0),
	.w4(32'h3a4d6916),
	.w5(32'h3a69b0ea),
	.w6(32'h3a85cadb),
	.w7(32'h3adc30e3),
	.w8(32'hba944253),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a312784),
	.w1(32'h3af916aa),
	.w2(32'hbac6b353),
	.w3(32'hba3c81cf),
	.w4(32'hbb196917),
	.w5(32'hbb40e0f7),
	.w6(32'h38d60b78),
	.w7(32'hbac6b50d),
	.w8(32'h3aa1a510),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76d567),
	.w1(32'h3a57aa9d),
	.w2(32'hba5146f5),
	.w3(32'h3a6f20a4),
	.w4(32'hb9bec9b5),
	.w5(32'hb9b0eb1a),
	.w6(32'h3ab7af7e),
	.w7(32'hbb2328f0),
	.w8(32'hba0301d3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e9b2a),
	.w1(32'hbbce4124),
	.w2(32'h3c9217b5),
	.w3(32'hb9b8d805),
	.w4(32'h3bb33f96),
	.w5(32'h3b0da8a8),
	.w6(32'h3a8a4e98),
	.w7(32'h3b9494eb),
	.w8(32'h3bf4ff90),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1a56e),
	.w1(32'h3af4203f),
	.w2(32'h3b99931b),
	.w3(32'h3b680123),
	.w4(32'h3a9786e3),
	.w5(32'h3b22bfd0),
	.w6(32'h3b4274a3),
	.w7(32'h3b2ed4f9),
	.w8(32'h3b38fd28),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac566e1),
	.w1(32'h3a90fd5f),
	.w2(32'hb8662b0c),
	.w3(32'h3b0779e3),
	.w4(32'h3986b238),
	.w5(32'hbac91cb9),
	.w6(32'h38a5d518),
	.w7(32'h39c8865b),
	.w8(32'hb9e497cf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1939c),
	.w1(32'h39960862),
	.w2(32'hba846b1a),
	.w3(32'hb9ab47f1),
	.w4(32'h3aebde3c),
	.w5(32'hb9200a4a),
	.w6(32'h3a8f2418),
	.w7(32'hb9a877b3),
	.w8(32'h398b145c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04eeda),
	.w1(32'hbc384d71),
	.w2(32'h3c1da8b7),
	.w3(32'h3abbd3cb),
	.w4(32'hba10858c),
	.w5(32'h3b909003),
	.w6(32'hbb4d917f),
	.w7(32'h3b5aa6ed),
	.w8(32'h3bedb0b2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55a7a9),
	.w1(32'h3b1cf42a),
	.w2(32'hb92d1864),
	.w3(32'h3be83ebb),
	.w4(32'hba84fcc6),
	.w5(32'hba40e56f),
	.w6(32'h39a3c049),
	.w7(32'hb8d42771),
	.w8(32'h3b00313a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0197),
	.w1(32'hba4faaee),
	.w2(32'h3a8c237e),
	.w3(32'h3a89ab4c),
	.w4(32'hb9c3784a),
	.w5(32'hb7c27b16),
	.w6(32'h3aa51ed8),
	.w7(32'h398d7449),
	.w8(32'h3af45c5c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf44ac),
	.w1(32'h38b9afdc),
	.w2(32'h3ac0cd22),
	.w3(32'h3aa12c55),
	.w4(32'h3a62fbeb),
	.w5(32'h3a5a38ae),
	.w6(32'h3a84c4c5),
	.w7(32'h3a7ad9dd),
	.w8(32'h3ae9f876),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fbbc5),
	.w1(32'hba3e09b7),
	.w2(32'hbaa949d8),
	.w3(32'h39cf1ba8),
	.w4(32'hba282e6e),
	.w5(32'hbaf4c147),
	.w6(32'h39b6b558),
	.w7(32'hba2b0772),
	.w8(32'hb875a97c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba359946),
	.w1(32'hbb315205),
	.w2(32'hbbf19fc9),
	.w3(32'hba8290b5),
	.w4(32'hbbb4d753),
	.w5(32'hbbc28d94),
	.w6(32'hbb975cc4),
	.w7(32'hbbcd445f),
	.w8(32'hbb251665),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ba4a2),
	.w1(32'h3c360e72),
	.w2(32'hbbaf26ba),
	.w3(32'hbadfc93e),
	.w4(32'hbb8943d4),
	.w5(32'h3b717ff4),
	.w6(32'h3c10556d),
	.w7(32'h3b6c34d6),
	.w8(32'h3aafe1bd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc658b1),
	.w1(32'hbadcb2a0),
	.w2(32'h3abbcb17),
	.w3(32'hbad53183),
	.w4(32'h3957d343),
	.w5(32'hbad02cdc),
	.w6(32'hb9eb65f7),
	.w7(32'hba95b84b),
	.w8(32'h3b0df1cd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9dac3),
	.w1(32'h3bb28c63),
	.w2(32'hbae7f42f),
	.w3(32'h39a791b1),
	.w4(32'h3a2ccf83),
	.w5(32'h3a8afa98),
	.w6(32'h3a099d1f),
	.w7(32'h39a56708),
	.w8(32'h3bbd279e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36478f),
	.w1(32'hba0166b9),
	.w2(32'h3bfa1b40),
	.w3(32'h3b986604),
	.w4(32'hbabaf3e3),
	.w5(32'h3b28772a),
	.w6(32'hba148ce3),
	.w7(32'h3b8147c6),
	.w8(32'h3a905004),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c219),
	.w1(32'hb985d42f),
	.w2(32'h3b0922c8),
	.w3(32'h3b24e799),
	.w4(32'h3a7482d3),
	.w5(32'h3ad5b784),
	.w6(32'h398b5ade),
	.w7(32'h3a91b2c4),
	.w8(32'h39fcb4ba),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c678a7),
	.w1(32'h3991bdc4),
	.w2(32'hbae9b24b),
	.w3(32'h3a12ad66),
	.w4(32'h3995e482),
	.w5(32'hbb308a75),
	.w6(32'hb995973f),
	.w7(32'hba7780f2),
	.w8(32'hba83afcb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52e074),
	.w1(32'hbb0be6ce),
	.w2(32'hbb8c0acd),
	.w3(32'hba6d85ae),
	.w4(32'hbb0cf442),
	.w5(32'hbaee9e46),
	.w6(32'hbae4c7d4),
	.w7(32'hbb785fa4),
	.w8(32'h3a8eefc1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0834d1),
	.w1(32'hbadbf10e),
	.w2(32'hbb621373),
	.w3(32'h3ac83e5b),
	.w4(32'hba921738),
	.w5(32'hbb4f663c),
	.w6(32'hbb203411),
	.w7(32'hbaffb2bd),
	.w8(32'h3a9310bc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad46dcf),
	.w1(32'hbad0bc38),
	.w2(32'hbb9307fc),
	.w3(32'h3a32056b),
	.w4(32'hbb02492d),
	.w5(32'hbb334276),
	.w6(32'hbae46e7f),
	.w7(32'hbb0a8b61),
	.w8(32'h3aaaf217),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6d58),
	.w1(32'hbb0e4d22),
	.w2(32'h3b1bd724),
	.w3(32'hba89dba1),
	.w4(32'hbab95809),
	.w5(32'h3b2dcfc7),
	.w6(32'h38800805),
	.w7(32'h3baa7be2),
	.w8(32'h3a235161),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bce8fb),
	.w1(32'h3b491123),
	.w2(32'h3b15c7d2),
	.w3(32'h3a6ae98f),
	.w4(32'h3b9467a5),
	.w5(32'h3b961b15),
	.w6(32'h3b106534),
	.w7(32'h3b33cd98),
	.w8(32'h3bddac5d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb524a),
	.w1(32'h3c3de335),
	.w2(32'hbb0cbc1d),
	.w3(32'h3bcee983),
	.w4(32'h3bd62cf5),
	.w5(32'h3a2e0b8c),
	.w6(32'h3bed8993),
	.w7(32'h3b30409b),
	.w8(32'h3b37705c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82f64f),
	.w1(32'hb9972e35),
	.w2(32'hb9ad9201),
	.w3(32'h3abe8134),
	.w4(32'hb7e537a0),
	.w5(32'hb8fe2231),
	.w6(32'h39a2577a),
	.w7(32'hb98d1f74),
	.w8(32'h3996fce6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971d3bf),
	.w1(32'hbaf3c21a),
	.w2(32'hba8c85ea),
	.w3(32'hb9946845),
	.w4(32'hbb166a55),
	.w5(32'hb63efe97),
	.w6(32'hbabc87c6),
	.w7(32'h38e5095b),
	.w8(32'hb9b2018c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b8a1d),
	.w1(32'hba3e514b),
	.w2(32'h3a0a4e9f),
	.w3(32'h3a8c52c3),
	.w4(32'h3a28cb2c),
	.w5(32'h38889685),
	.w6(32'h38eca088),
	.w7(32'hb98aaf88),
	.w8(32'h39c44d6e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dee1b),
	.w1(32'hbb11ee09),
	.w2(32'hbae08d19),
	.w3(32'h3a355ca8),
	.w4(32'hba49dcd9),
	.w5(32'hbb114391),
	.w6(32'h398a06fa),
	.w7(32'hb95b516b),
	.w8(32'h3acdab69),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45c88f),
	.w1(32'h3ac09a02),
	.w2(32'h3b4a1644),
	.w3(32'h3a06cb56),
	.w4(32'h3a04dace),
	.w5(32'h3b485431),
	.w6(32'h3b4bb12a),
	.w7(32'h3b46a636),
	.w8(32'h3b5fd897),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516c4f),
	.w1(32'hbb2f4bae),
	.w2(32'hbbe66467),
	.w3(32'h3b8f6ffc),
	.w4(32'hbb821697),
	.w5(32'hbbad8f23),
	.w6(32'hbb18378b),
	.w7(32'hbb38570a),
	.w8(32'h3a103d2f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f7339),
	.w1(32'h3a926c88),
	.w2(32'hbb0989c1),
	.w3(32'hbb3b4a93),
	.w4(32'h39ce11d4),
	.w5(32'hbb36bc89),
	.w6(32'h39c98ca3),
	.w7(32'hbb05b395),
	.w8(32'hba508b43),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b77037),
	.w1(32'h3abfbe1d),
	.w2(32'h3a2e1d9e),
	.w3(32'hb9812737),
	.w4(32'h3a91bd05),
	.w5(32'hba3db9b1),
	.w6(32'hb910931a),
	.w7(32'hbac4f154),
	.w8(32'h393ad50f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5903),
	.w1(32'h3abcb847),
	.w2(32'h3c1a486e),
	.w3(32'hbac338c0),
	.w4(32'h3be0c7f0),
	.w5(32'hbbe2482b),
	.w6(32'h3b379b77),
	.w7(32'h3c02882c),
	.w8(32'h3bb5f10a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1640),
	.w1(32'h3b29c857),
	.w2(32'h3b399ae8),
	.w3(32'hbb9d6391),
	.w4(32'h3a929763),
	.w5(32'h3b403b06),
	.w6(32'h3afa4c81),
	.w7(32'h3b71c364),
	.w8(32'hb7f0fcad),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57ce33),
	.w1(32'h3b58de9e),
	.w2(32'h3a08204a),
	.w3(32'h38a9d3c6),
	.w4(32'h3a93704e),
	.w5(32'hbaa75b07),
	.w6(32'h3b3ba9bb),
	.w7(32'hbad61cd6),
	.w8(32'hb94fcb92),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10565d),
	.w1(32'hbb8ee77b),
	.w2(32'hbb892c68),
	.w3(32'hbb56bed3),
	.w4(32'hbb8b0cd4),
	.w5(32'hbb3b1213),
	.w6(32'hbb6caa79),
	.w7(32'hbb535e7a),
	.w8(32'hbb5ae2f2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc5d3),
	.w1(32'hba88db13),
	.w2(32'hbbbf4992),
	.w3(32'hba994bf1),
	.w4(32'hbb01371d),
	.w5(32'hbb32afeb),
	.w6(32'hba7ef6e7),
	.w7(32'hbbb5b42e),
	.w8(32'hbb265ab8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a184a94),
	.w1(32'hbc627ebf),
	.w2(32'h3c89f396),
	.w3(32'hba8ed511),
	.w4(32'hbbcb3d26),
	.w5(32'hbb929480),
	.w6(32'h3b59f219),
	.w7(32'hbb6adc99),
	.w8(32'h3b391764),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454e76),
	.w1(32'hbbe073b3),
	.w2(32'h3d17668d),
	.w3(32'h3b559953),
	.w4(32'h3c4ceb99),
	.w5(32'h3c3f39ad),
	.w6(32'h3af34aaa),
	.w7(32'h3c8d5959),
	.w8(32'h3bfb18f7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f89598),
	.w1(32'hbb899489),
	.w2(32'h3ac8e542),
	.w3(32'h3b25fbf0),
	.w4(32'h3a822aff),
	.w5(32'hbb226e16),
	.w6(32'h38e9f584),
	.w7(32'hbae20371),
	.w8(32'h3b6aacb8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe14dc),
	.w1(32'h398b2752),
	.w2(32'h3ab060cf),
	.w3(32'h3a32b125),
	.w4(32'h3a2f1f65),
	.w5(32'h3a07d5fa),
	.w6(32'h3b2d4483),
	.w7(32'h3aa52b5c),
	.w8(32'h3afefed8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae681ca),
	.w1(32'hbab42cba),
	.w2(32'h3a40d620),
	.w3(32'h3aa09c79),
	.w4(32'hb875a315),
	.w5(32'hbaa87605),
	.w6(32'hb80ffb57),
	.w7(32'hba727e0b),
	.w8(32'h3adcb5ef),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c89a),
	.w1(32'h38c3b95e),
	.w2(32'hba8f546a),
	.w3(32'h39b3b786),
	.w4(32'h392c895a),
	.w5(32'hba66bbb0),
	.w6(32'h3984b438),
	.w7(32'hba56eb4e),
	.w8(32'hb93d8c95),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0015e),
	.w1(32'h3ad89d0b),
	.w2(32'hbb7751fa),
	.w3(32'hba5caa9d),
	.w4(32'h3ae3c030),
	.w5(32'hbac7ad72),
	.w6(32'h3a3fae47),
	.w7(32'hb99f46c1),
	.w8(32'hbac8f25e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f8c95),
	.w1(32'hba5e7726),
	.w2(32'hbb03adbf),
	.w3(32'hba9bcf8b),
	.w4(32'hba1f515a),
	.w5(32'hbaf80106),
	.w6(32'h39eb2032),
	.w7(32'hb9990a25),
	.w8(32'h3aac32cd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f0899),
	.w1(32'hbaf4ed49),
	.w2(32'h3aa7dd4c),
	.w3(32'h3924eedd),
	.w4(32'h39a07995),
	.w5(32'hba9e7c3a),
	.w6(32'hb95ab6a9),
	.w7(32'hba3dea74),
	.w8(32'h3b06feb8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a628636),
	.w1(32'h3bb7742c),
	.w2(32'hbb3e6e78),
	.w3(32'h39aa78ac),
	.w4(32'h3b18b2df),
	.w5(32'h3910b6d2),
	.w6(32'h3b3d3940),
	.w7(32'hbaee64cf),
	.w8(32'h3920a603),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36acef),
	.w1(32'hbb01e6dc),
	.w2(32'hbaeca6d6),
	.w3(32'h39a3e7eb),
	.w4(32'hba8a6ba6),
	.w5(32'h38a2610c),
	.w6(32'hba9f3dd5),
	.w7(32'hba36aec1),
	.w8(32'h3ab9a0f1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab12e7),
	.w1(32'h3c307f15),
	.w2(32'h3b7e421b),
	.w3(32'h3a1e4dcf),
	.w4(32'h3b4da9f7),
	.w5(32'h3b6005a0),
	.w6(32'h3a6e1e02),
	.w7(32'h3a86a8b5),
	.w8(32'h3b3e18d0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b7f0d),
	.w1(32'hb9d4cc38),
	.w2(32'hbb2f637b),
	.w3(32'h3b894a2e),
	.w4(32'h39f091d0),
	.w5(32'h39a85426),
	.w6(32'h399e1df1),
	.w7(32'hbacf90a6),
	.w8(32'h39794628),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33c119),
	.w1(32'h3b44d351),
	.w2(32'hbaad17e3),
	.w3(32'h3b04f049),
	.w4(32'hbb3e5ad9),
	.w5(32'hb92d289c),
	.w6(32'h3aa70b52),
	.w7(32'hbb05b5d2),
	.w8(32'hb8f847f3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa70eb),
	.w1(32'h3b5aea3a),
	.w2(32'hbb7b0312),
	.w3(32'h3af71f11),
	.w4(32'h3b727e89),
	.w5(32'h3a1a3879),
	.w6(32'h3b49bef6),
	.w7(32'hbae26694),
	.w8(32'hb9b4913f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb361),
	.w1(32'hbb175435),
	.w2(32'h3aca0a24),
	.w3(32'h3a8bb0b7),
	.w4(32'h3964f7ff),
	.w5(32'hbae243a5),
	.w6(32'hb91b4c73),
	.w7(32'hba931a68),
	.w8(32'h3b351d0d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac780da),
	.w1(32'hba584ace),
	.w2(32'h3a9cd7ae),
	.w3(32'h39b703b1),
	.w4(32'h3858e93a),
	.w5(32'h39e3e124),
	.w6(32'h39d0def4),
	.w7(32'h396aaece),
	.w8(32'h3ab1dc41),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b82bf),
	.w1(32'hba17fc60),
	.w2(32'h3a0409eb),
	.w3(32'h3a44481e),
	.w4(32'h39685f80),
	.w5(32'hb9d501dd),
	.w6(32'h39f28896),
	.w7(32'hb9a3ec91),
	.w8(32'h3a99c61a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5148d9),
	.w1(32'hbae2a79b),
	.w2(32'h3bb04516),
	.w3(32'h394f6bf9),
	.w4(32'h3bb79556),
	.w5(32'hbb5029bc),
	.w6(32'hbaab04fb),
	.w7(32'hbb7a2d59),
	.w8(32'h393e1996),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b418e78),
	.w1(32'hbad779a8),
	.w2(32'h3c4ba852),
	.w3(32'hba637329),
	.w4(32'h3b503daa),
	.w5(32'h3b2eaf7b),
	.w6(32'h3ad1ae71),
	.w7(32'h3b332de8),
	.w8(32'h3bbe13ce),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ce874),
	.w1(32'h3a9fa6e6),
	.w2(32'hbb4095aa),
	.w3(32'h3a3e3f3f),
	.w4(32'h39675860),
	.w5(32'hb9fe5a54),
	.w6(32'h3b28adfc),
	.w7(32'hbb0c177a),
	.w8(32'hba881110),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada5d59),
	.w1(32'hbb05a3f4),
	.w2(32'hbb3c593b),
	.w3(32'h3a858b83),
	.w4(32'h38f51108),
	.w5(32'hba898f13),
	.w6(32'h3a1a70f3),
	.w7(32'hbaa9f640),
	.w8(32'h3b32b7a1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09fc8c),
	.w1(32'hba66772c),
	.w2(32'h3a8d8683),
	.w3(32'h3ab87cbc),
	.w4(32'h3987717d),
	.w5(32'h38964658),
	.w6(32'hb7deafdc),
	.w7(32'hb9332ef6),
	.w8(32'h3ae90d3f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae023bb),
	.w1(32'hbb9201f6),
	.w2(32'h3be9843a),
	.w3(32'h3a33a148),
	.w4(32'h3bae08c3),
	.w5(32'hbbc8370f),
	.w6(32'hbbceb57a),
	.w7(32'h3b5d584d),
	.w8(32'hba858107),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8fa52),
	.w1(32'h3b78e8ef),
	.w2(32'hbb896a2d),
	.w3(32'hbb40e5e1),
	.w4(32'h3b78603f),
	.w5(32'hbb1c3db6),
	.w6(32'h3bd336d1),
	.w7(32'h3af3fdb3),
	.w8(32'hbaad891e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25d63),
	.w1(32'hba8f6111),
	.w2(32'hbac73f32),
	.w3(32'hbba474d2),
	.w4(32'hb9cfb9e4),
	.w5(32'hba86f96f),
	.w6(32'hb8e6b6b1),
	.w7(32'hbaa0e5f0),
	.w8(32'hb9e98ad5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d5042),
	.w1(32'hbac54e65),
	.w2(32'hbb88e28d),
	.w3(32'hba791f9d),
	.w4(32'hb98719fc),
	.w5(32'hbb4bc14c),
	.w6(32'hb9481565),
	.w7(32'hbb174f97),
	.w8(32'hbb2979b8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb063d69),
	.w1(32'h3ac5a732),
	.w2(32'h39a51608),
	.w3(32'hbb16911d),
	.w4(32'h3b3a70f0),
	.w5(32'h3a96fcd7),
	.w6(32'h3a5711eb),
	.w7(32'h39aae3f5),
	.w8(32'hba41986e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule