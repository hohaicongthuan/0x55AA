module layer_10_featuremap_66(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a2565),
	.w1(32'h3c2a4ddf),
	.w2(32'hbc4a746c),
	.w3(32'hbb172715),
	.w4(32'hbc51023d),
	.w5(32'hbb153ad8),
	.w6(32'h3cbcabee),
	.w7(32'hbc38cec5),
	.w8(32'h3bd1ceaa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8f75),
	.w1(32'h3c488010),
	.w2(32'h39db80bb),
	.w3(32'hbbd35610),
	.w4(32'h3c919ae3),
	.w5(32'h3ba2bfd6),
	.w6(32'hbb12438f),
	.w7(32'h3abfeedd),
	.w8(32'h3c318d5f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760c4e),
	.w1(32'h3c97fc0b),
	.w2(32'h3c03126b),
	.w3(32'hbc7060dc),
	.w4(32'h3c509e9a),
	.w5(32'h3be9f73d),
	.w6(32'h3c55e8ea),
	.w7(32'hbc0bd910),
	.w8(32'h3ab05a2b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6a52c),
	.w1(32'h3ae2d5db),
	.w2(32'hbb473f56),
	.w3(32'h3bd0a5c8),
	.w4(32'hbb810e87),
	.w5(32'hbc1a8cbd),
	.w6(32'h3b5e2200),
	.w7(32'h3bc2d944),
	.w8(32'h3a6a7fc7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09fa85),
	.w1(32'hbb85b73a),
	.w2(32'hbb82103e),
	.w3(32'hbc89d04e),
	.w4(32'hbc103669),
	.w5(32'hbc78197a),
	.w6(32'h3b4114ef),
	.w7(32'hbc7c83a2),
	.w8(32'hbc4a7fdf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d2403),
	.w1(32'h3c4781ac),
	.w2(32'hbb3c2ddb),
	.w3(32'hbc268afd),
	.w4(32'h3b9e3f4b),
	.w5(32'hbae8c165),
	.w6(32'hbb182ed6),
	.w7(32'hbbc767ec),
	.w8(32'hbb93f355),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a5aa5),
	.w1(32'h3bc10910),
	.w2(32'hbb5c3d41),
	.w3(32'hbad1aa82),
	.w4(32'h3ae188e3),
	.w5(32'hbb722ec4),
	.w6(32'hbae4ce66),
	.w7(32'hbb54e082),
	.w8(32'h3b4edc0a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab83c6),
	.w1(32'hbb08eb37),
	.w2(32'hbbc2a9d9),
	.w3(32'hbb95c927),
	.w4(32'hbbd8f4e9),
	.w5(32'hbc6ad40e),
	.w6(32'h3bb9544f),
	.w7(32'hbba79d6f),
	.w8(32'hbc49f043),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1f39),
	.w1(32'hbc379c06),
	.w2(32'h3c36cf7d),
	.w3(32'hbbbf8831),
	.w4(32'hbcbe8d9c),
	.w5(32'h3bec0aad),
	.w6(32'h3add166f),
	.w7(32'hbc23301a),
	.w8(32'h3c054ac1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c01cf),
	.w1(32'h3c911bc0),
	.w2(32'h3b8b1174),
	.w3(32'h3b1a5f16),
	.w4(32'h3c89eca8),
	.w5(32'h3b4987d6),
	.w6(32'hb88fe266),
	.w7(32'h3c892e50),
	.w8(32'h3bd6be2c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d66be),
	.w1(32'h3aeec49c),
	.w2(32'h3a5205c2),
	.w3(32'hba86c197),
	.w4(32'h3b5721f7),
	.w5(32'h39b21a8f),
	.w6(32'hba9965ae),
	.w7(32'h3b90105d),
	.w8(32'h3b400db9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936816),
	.w1(32'hbba0f54e),
	.w2(32'h3ac451ca),
	.w3(32'hbc08bf8f),
	.w4(32'hbc2a44ca),
	.w5(32'h3a9ebb82),
	.w6(32'h3bdfc29c),
	.w7(32'h3b0a0f3f),
	.w8(32'h3acd695a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b361f55),
	.w1(32'h3b0dd2d1),
	.w2(32'h3c057937),
	.w3(32'h3bb4a9ea),
	.w4(32'h3b8d8aef),
	.w5(32'h3c0b0c3c),
	.w6(32'h3ac90424),
	.w7(32'h3bbc2d64),
	.w8(32'hb9508fc3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f7c1),
	.w1(32'h3bc1b933),
	.w2(32'h3c391ee2),
	.w3(32'h3c7064cb),
	.w4(32'h3bb6c54a),
	.w5(32'h3c18167e),
	.w6(32'h3ba48aa7),
	.w7(32'h3b42ca50),
	.w8(32'hbc159dcc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cc7abb),
	.w1(32'hba9a6136),
	.w2(32'hbb5b5154),
	.w3(32'h3c9bbc6f),
	.w4(32'h3b740b67),
	.w5(32'hbb09d340),
	.w6(32'h3c1766c9),
	.w7(32'h3c09e49a),
	.w8(32'h3c12ea34),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eeb3a),
	.w1(32'h3c1079d0),
	.w2(32'h3b284bc2),
	.w3(32'hbca3241d),
	.w4(32'h398a7866),
	.w5(32'h3a69e231),
	.w6(32'hbc9a67d4),
	.w7(32'hbc3ed695),
	.w8(32'h3baa51f6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5de6fd),
	.w1(32'h3afa0650),
	.w2(32'h3ae4e36e),
	.w3(32'h387415b9),
	.w4(32'h3b31e3af),
	.w5(32'h3b6d310d),
	.w6(32'hbb02a24e),
	.w7(32'h3afd15a6),
	.w8(32'h393161f0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1550),
	.w1(32'h3b8413f4),
	.w2(32'hbbabc5f5),
	.w3(32'hbc2ac65c),
	.w4(32'hba40633e),
	.w5(32'hbbe3f90e),
	.w6(32'hbc12c876),
	.w7(32'hbc607e7b),
	.w8(32'hbbd94837),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf86cc7),
	.w1(32'hbb729a93),
	.w2(32'h3c84fd47),
	.w3(32'h3b33534b),
	.w4(32'hbc03722b),
	.w5(32'h3b852402),
	.w6(32'h3c0f6e9f),
	.w7(32'hbb0e12ee),
	.w8(32'h3c622f9a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88031f),
	.w1(32'hbb91492e),
	.w2(32'hbb56c8e0),
	.w3(32'h3d3eca1e),
	.w4(32'h3c5a72bf),
	.w5(32'h3b6bfb9d),
	.w6(32'h3b5e0ca1),
	.w7(32'h3cc2436b),
	.w8(32'h3be0cdd2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4503),
	.w1(32'hba108719),
	.w2(32'h3c21025f),
	.w3(32'hbbcf60e1),
	.w4(32'hb904f2dd),
	.w5(32'hbb238276),
	.w6(32'hbc0f14aa),
	.w7(32'hbb337fe4),
	.w8(32'h3b32d117),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c8759),
	.w1(32'hbbd132ce),
	.w2(32'hbc179f60),
	.w3(32'h3cc99c96),
	.w4(32'h3bf458ae),
	.w5(32'hbbadb759),
	.w6(32'hbc2c19b4),
	.w7(32'h3c898f48),
	.w8(32'h3c26600d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b22dd),
	.w1(32'h3bbafb59),
	.w2(32'hbb3bdac7),
	.w3(32'hbc4ded87),
	.w4(32'hbbbeaa34),
	.w5(32'hbb00c63d),
	.w6(32'hbc3258b2),
	.w7(32'hbaf8102f),
	.w8(32'hba0ac47e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e561b),
	.w1(32'hb9db5a00),
	.w2(32'h3b60af36),
	.w3(32'h3b5cd480),
	.w4(32'h3b4838f4),
	.w5(32'h3ba84f33),
	.w6(32'h3a89f750),
	.w7(32'h3bcbd823),
	.w8(32'h3b99219e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4965),
	.w1(32'h3bb9749a),
	.w2(32'hbc46314c),
	.w3(32'h3ba0d895),
	.w4(32'h3bc54a47),
	.w5(32'hbbf009c5),
	.w6(32'h3c4bb423),
	.w7(32'h3889ddc1),
	.w8(32'hb9c487c8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc215f0c),
	.w1(32'hbb10167b),
	.w2(32'h3b1f5a02),
	.w3(32'hbc5ab935),
	.w4(32'hbc67a84f),
	.w5(32'h3bf5fd7f),
	.w6(32'hbc1dd194),
	.w7(32'hbc7ad011),
	.w8(32'h3b1cf3cb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada07f0),
	.w1(32'h3b690cb8),
	.w2(32'h3a6adf5e),
	.w3(32'h3b68550c),
	.w4(32'h3c00a8c3),
	.w5(32'h3b194ec5),
	.w6(32'h3b929c87),
	.w7(32'h3b101818),
	.w8(32'h39500c7c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c8f56),
	.w1(32'h3a86d7d5),
	.w2(32'h381b1130),
	.w3(32'h3a83e06a),
	.w4(32'h3b54b8e6),
	.w5(32'hbb69705e),
	.w6(32'hba231ae4),
	.w7(32'h3a1e1fdc),
	.w8(32'hba3d1f29),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71a629),
	.w1(32'h3b590c87),
	.w2(32'hbbd6f7b2),
	.w3(32'hba8f0b5b),
	.w4(32'h3c2678b1),
	.w5(32'h3c4446c1),
	.w6(32'h3a6c30a1),
	.w7(32'h3c4eeef9),
	.w8(32'h3c16893a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17da90),
	.w1(32'h3c8acdcb),
	.w2(32'h3922451c),
	.w3(32'h3ba9149c),
	.w4(32'h3ca5dec7),
	.w5(32'h3b466738),
	.w6(32'h3a90f03b),
	.w7(32'h3bb0a671),
	.w8(32'h3ab2e6c6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafec15f),
	.w1(32'hbb7b9346),
	.w2(32'hb9de8747),
	.w3(32'hbb374587),
	.w4(32'hbb98357d),
	.w5(32'h3cb49d7a),
	.w6(32'hbba40852),
	.w7(32'hbbfd18ab),
	.w8(32'h3cae9545),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb658119),
	.w1(32'h3b0e8a04),
	.w2(32'hbbc80b7c),
	.w3(32'hba21cf74),
	.w4(32'hbc2b31e2),
	.w5(32'h3b90cba4),
	.w6(32'hbaf0bb1f),
	.w7(32'hbcdbea24),
	.w8(32'h3c3d4512),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284dd0),
	.w1(32'h3bebf055),
	.w2(32'h39b09ed4),
	.w3(32'h3b91de40),
	.w4(32'hbbfd7a16),
	.w5(32'h3b0f07f1),
	.w6(32'h3ba0188c),
	.w7(32'hbc8d629b),
	.w8(32'h3b416471),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a57fa6),
	.w1(32'h3a87fa9d),
	.w2(32'hba9a4b92),
	.w3(32'h3afb228f),
	.w4(32'h38a5689d),
	.w5(32'h3c0da3eb),
	.w6(32'h3b2ce839),
	.w7(32'h3b2ce489),
	.w8(32'hbbeddd0c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26270a),
	.w1(32'h3bfc1e7a),
	.w2(32'hbb271d2a),
	.w3(32'h393ddba6),
	.w4(32'h3b2bd36c),
	.w5(32'hbb69dd22),
	.w6(32'hbbe05e1f),
	.w7(32'h39ba0cec),
	.w8(32'hba9b12c1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60915a),
	.w1(32'hbb599609),
	.w2(32'hbc80c6b6),
	.w3(32'hbb67fb22),
	.w4(32'hbac03a6f),
	.w5(32'hbc5a7cde),
	.w6(32'hbaf126d8),
	.w7(32'hba8b45a5),
	.w8(32'h3c88f465),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb455156),
	.w1(32'h3bee7444),
	.w2(32'hbab6d663),
	.w3(32'hbca4ebbf),
	.w4(32'hbab0dd73),
	.w5(32'hb9d79158),
	.w6(32'hbb19603d),
	.w7(32'hbcbd6025),
	.w8(32'h394f6e62),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32149),
	.w1(32'hbbd6fca7),
	.w2(32'h3c3bceda),
	.w3(32'hbb7da1ab),
	.w4(32'h39bd06ee),
	.w5(32'h3c92e8f7),
	.w6(32'hba019990),
	.w7(32'h3aa44647),
	.w8(32'h3a7b1762),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2825),
	.w1(32'hbaad1ba6),
	.w2(32'hbc810c53),
	.w3(32'h3bfac869),
	.w4(32'hbbc7b38f),
	.w5(32'h3aedaeab),
	.w6(32'h3ba97bd3),
	.w7(32'h3bbb8d05),
	.w8(32'h3a96fdfe),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c652b),
	.w1(32'h3bfce7bf),
	.w2(32'hba9eadc3),
	.w3(32'h3b76434d),
	.w4(32'h3c2163db),
	.w5(32'hba995727),
	.w6(32'h3be027eb),
	.w7(32'h3b85fced),
	.w8(32'hbb1491f0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba92b4),
	.w1(32'hbab141f9),
	.w2(32'h3bbc4482),
	.w3(32'hbbc9ca46),
	.w4(32'hbbe6866c),
	.w5(32'hbbb24b6b),
	.w6(32'hbc112849),
	.w7(32'hbbc03dea),
	.w8(32'hba7989fb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b3526),
	.w1(32'hba5aa235),
	.w2(32'h3b443d45),
	.w3(32'h3ad3c750),
	.w4(32'h3b1589ac),
	.w5(32'h3c2075d7),
	.w6(32'hbb89faeb),
	.w7(32'h3b9203d4),
	.w8(32'h3be2c384),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ab229),
	.w1(32'h3c3f97e2),
	.w2(32'hbb0979c4),
	.w3(32'h3c85805d),
	.w4(32'h3b312c54),
	.w5(32'hbb40c263),
	.w6(32'h3b3e90ac),
	.w7(32'hbb9a2196),
	.w8(32'hba155350),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449b1f),
	.w1(32'hbacc26bb),
	.w2(32'h3c01fe9b),
	.w3(32'hbb341b68),
	.w4(32'hb948d6d9),
	.w5(32'h3c11a97e),
	.w6(32'hb9f41d31),
	.w7(32'h3881d936),
	.w8(32'h3ada0e0c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd6887),
	.w1(32'h3adcca06),
	.w2(32'hbc6efacb),
	.w3(32'h3cdf0bea),
	.w4(32'h3cc5d75c),
	.w5(32'hbbb62a88),
	.w6(32'h3c627851),
	.w7(32'h3cd5444b),
	.w8(32'hbc0a476e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16a0fb),
	.w1(32'h3c86235b),
	.w2(32'h3c0dc6c3),
	.w3(32'hbab2b817),
	.w4(32'h3c95a630),
	.w5(32'hbc3587be),
	.w6(32'hba8b2baa),
	.w7(32'h3d056b5e),
	.w8(32'hbb51410f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305611),
	.w1(32'hbb504fa8),
	.w2(32'hbb0e7566),
	.w3(32'hbba8426f),
	.w4(32'hba961625),
	.w5(32'h3b39a8b1),
	.w6(32'hbb0ed632),
	.w7(32'hbb575c85),
	.w8(32'h3b401def),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab68e6),
	.w1(32'hbb9bc1a8),
	.w2(32'hbbe5d85b),
	.w3(32'hbc4d72fe),
	.w4(32'hbb0d0e35),
	.w5(32'hbbb46a1d),
	.w6(32'hbc2a71e1),
	.w7(32'h3b72659f),
	.w8(32'hbba0a481),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc12148),
	.w1(32'hbb15fc00),
	.w2(32'h3b2b7ea4),
	.w3(32'hbb6f17ee),
	.w4(32'h388a7077),
	.w5(32'h3c5372bf),
	.w6(32'hbb28e3a0),
	.w7(32'hbaa6eda7),
	.w8(32'h3aa08d99),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed7b69),
	.w1(32'hba4e0ae5),
	.w2(32'hbbd97e26),
	.w3(32'h3b94fa4e),
	.w4(32'hbc4eacf4),
	.w5(32'hbc42d198),
	.w6(32'h3ad1a9ec),
	.w7(32'hbb16a8b0),
	.w8(32'hbcaf5fbd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7f53),
	.w1(32'h3b99de06),
	.w2(32'hbbba5bbf),
	.w3(32'h3b38e2ff),
	.w4(32'h3c72dde3),
	.w5(32'hbba424b5),
	.w6(32'hbc12484a),
	.w7(32'h3bf2a3d9),
	.w8(32'hbc3447de),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce7da),
	.w1(32'h3aefaf6c),
	.w2(32'hbb0b0fe0),
	.w3(32'h3923ec26),
	.w4(32'h393a8a98),
	.w5(32'hbc91a84f),
	.w6(32'h3bb0559b),
	.w7(32'h3c0b01ae),
	.w8(32'hbcacc358),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e40c6),
	.w1(32'h3c0fa5bc),
	.w2(32'hba80cc2d),
	.w3(32'h3b82a051),
	.w4(32'h3c88f265),
	.w5(32'h3b245c42),
	.w6(32'hbb2d04ca),
	.w7(32'h3c5432e9),
	.w8(32'h3a1e8f5f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95594),
	.w1(32'hbb2e40d6),
	.w2(32'hbb97171a),
	.w3(32'h3bb67342),
	.w4(32'hbaca9503),
	.w5(32'hba295a6a),
	.w6(32'h3982d8e6),
	.w7(32'hbb80955b),
	.w8(32'h3c39226c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35da81),
	.w1(32'h3c758b78),
	.w2(32'hbc16920e),
	.w3(32'h3b10c736),
	.w4(32'h3c75ee64),
	.w5(32'h3c0d9a09),
	.w6(32'hbbb2fc17),
	.w7(32'hbbb6473e),
	.w8(32'h3ce680b4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f32e),
	.w1(32'h3b916b4c),
	.w2(32'hbba431ce),
	.w3(32'h3b53b905),
	.w4(32'h3ba552bb),
	.w5(32'hbb0b7f65),
	.w6(32'h3c66ea9d),
	.w7(32'hbc6ade0e),
	.w8(32'hbb3203b7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10b053),
	.w1(32'h395d2ca2),
	.w2(32'hbb79f5fc),
	.w3(32'h3c036764),
	.w4(32'h3c6d0207),
	.w5(32'h3a75259c),
	.w6(32'h3bdc2b3c),
	.w7(32'h3c0e6677),
	.w8(32'h3bbdc21e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa254),
	.w1(32'hbb104d7f),
	.w2(32'h3a2dd46d),
	.w3(32'hbb2cb652),
	.w4(32'hb9e36591),
	.w5(32'hbac49efe),
	.w6(32'h3a0d830c),
	.w7(32'h3b4423b0),
	.w8(32'h3b9b69db),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7cad1),
	.w1(32'h3c361789),
	.w2(32'hbb6f41c0),
	.w3(32'hbb38fc4d),
	.w4(32'h3c263640),
	.w5(32'h3b087604),
	.w6(32'h38318524),
	.w7(32'h3c873f25),
	.w8(32'hba947e18),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042381),
	.w1(32'h3bcffb19),
	.w2(32'hb92c49f7),
	.w3(32'h3bba89d1),
	.w4(32'h3b9cea3b),
	.w5(32'h3b8279f6),
	.w6(32'hba5ef4b2),
	.w7(32'hbb3488c2),
	.w8(32'hbb570711),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96000b),
	.w1(32'h3a1771dd),
	.w2(32'hbbb43024),
	.w3(32'hbbf1efc7),
	.w4(32'hbae4441f),
	.w5(32'hba6016ab),
	.w6(32'hbad65e69),
	.w7(32'h3bdae7e8),
	.w8(32'hbbfff324),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4188a2),
	.w1(32'hbaec5a22),
	.w2(32'hbc112828),
	.w3(32'h3b8f0b69),
	.w4(32'h3a96d811),
	.w5(32'hbcc160f8),
	.w6(32'h3c1d020f),
	.w7(32'h3c07150d),
	.w8(32'hbcbdebfa),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c763),
	.w1(32'hbb28d97f),
	.w2(32'hbb685263),
	.w3(32'h3b92a7d6),
	.w4(32'h3c9d221e),
	.w5(32'hbbcaeafd),
	.w6(32'h3bdec4bb),
	.w7(32'h3d025d7e),
	.w8(32'hbc084fdc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bffda),
	.w1(32'hbb0eb9e9),
	.w2(32'h3bd8c4c2),
	.w3(32'hbb72aa82),
	.w4(32'h3be7505e),
	.w5(32'h3c71a4cc),
	.w6(32'hbc1cf0da),
	.w7(32'hbbc059e0),
	.w8(32'h3cd8c438),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf74b69),
	.w1(32'hbb48d23a),
	.w2(32'hba5ccda8),
	.w3(32'hbb077bbb),
	.w4(32'hbca23b10),
	.w5(32'hb9c51cde),
	.w6(32'h3c0f565b),
	.w7(32'hbcc66d8d),
	.w8(32'h3b2aa17f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8ec29),
	.w1(32'hba503520),
	.w2(32'h3b1267b6),
	.w3(32'hbaece738),
	.w4(32'hbaaf5406),
	.w5(32'hb9bf6b4e),
	.w6(32'hbaaf6a91),
	.w7(32'h3aa5fea1),
	.w8(32'hba7bba4b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3fc2),
	.w1(32'hb81bfc9e),
	.w2(32'h3b9ff293),
	.w3(32'h3ad461e9),
	.w4(32'h3b702e1c),
	.w5(32'hbb546c02),
	.w6(32'h3b5062de),
	.w7(32'h3b5b84e0),
	.w8(32'hba35ea9a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64fe41),
	.w1(32'hbb2109e5),
	.w2(32'h39c51897),
	.w3(32'hbab7bce4),
	.w4(32'hbb807b94),
	.w5(32'hbbdf4a39),
	.w6(32'hbc1e30f8),
	.w7(32'hbab4e0d7),
	.w8(32'hbbc46814),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa9ce7),
	.w1(32'h3bcc70a8),
	.w2(32'hbae2fdd5),
	.w3(32'h3901e7b0),
	.w4(32'h3bcd8346),
	.w5(32'hbaada42b),
	.w6(32'hbb1b584c),
	.w7(32'h3c1601de),
	.w8(32'hba853a7a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace9c33),
	.w1(32'h3b8b8cbf),
	.w2(32'h3b692158),
	.w3(32'hbb0c60d4),
	.w4(32'h399f6901),
	.w5(32'h3bfa5585),
	.w6(32'hbb3f0b43),
	.w7(32'hba50c484),
	.w8(32'h3b9abb57),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd2008),
	.w1(32'h3b57ea26),
	.w2(32'h3a85947f),
	.w3(32'h3ba5ac16),
	.w4(32'h3b1d5228),
	.w5(32'hbb2de106),
	.w6(32'h3bc37c41),
	.w7(32'h3a2c61d2),
	.w8(32'hbb74d9af),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ff16),
	.w1(32'hba47537a),
	.w2(32'h3c01f615),
	.w3(32'h38ff17ba),
	.w4(32'h3a0861f0),
	.w5(32'h3b3761f3),
	.w6(32'hbb7e04d1),
	.w7(32'hbb06b62b),
	.w8(32'h3c423e65),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01065f),
	.w1(32'hbb333c16),
	.w2(32'hbb057e87),
	.w3(32'hbb85c25f),
	.w4(32'h3978e1d9),
	.w5(32'h3c8964f1),
	.w6(32'hbaf7b1a8),
	.w7(32'hba7cc07b),
	.w8(32'h3c90d792),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d250d),
	.w1(32'hb9f154b4),
	.w2(32'hbb1a3734),
	.w3(32'hbba4e09c),
	.w4(32'hbcd653bf),
	.w5(32'h39c12a2b),
	.w6(32'h3aff6f95),
	.w7(32'hbcd6e5b8),
	.w8(32'hba3f5f32),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18c961),
	.w1(32'h3b590b7b),
	.w2(32'h3bb12bb8),
	.w3(32'h3ab9c197),
	.w4(32'h3b8e3dd2),
	.w5(32'h3b8d224f),
	.w6(32'hbb4059a2),
	.w7(32'h397c1202),
	.w8(32'h3b2df7d6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33d9cb),
	.w1(32'hbbb3ee9b),
	.w2(32'hbb98d17d),
	.w3(32'h3b8691db),
	.w4(32'hbb89de94),
	.w5(32'hba5cb6c8),
	.w6(32'h3ba32f2f),
	.w7(32'hbb81821d),
	.w8(32'h3c23138e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1605e7),
	.w1(32'h3c199663),
	.w2(32'hbbdd09e1),
	.w3(32'h3c2435a6),
	.w4(32'h3c342e62),
	.w5(32'hba922ca4),
	.w6(32'h3cc0b91f),
	.w7(32'h3c9240e7),
	.w8(32'h3c159a1b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdf6b5),
	.w1(32'h3c1425fd),
	.w2(32'hbbc71b81),
	.w3(32'h3c1abd5b),
	.w4(32'h3c019b92),
	.w5(32'hbb8e0af2),
	.w6(32'h3cb406ae),
	.w7(32'h3c4ffbbe),
	.w8(32'hbb64a564),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3415a3),
	.w1(32'h3ae4a460),
	.w2(32'h3b6fdab7),
	.w3(32'h3b307d50),
	.w4(32'h3c256fe7),
	.w5(32'h3afa69fa),
	.w6(32'hbb3aa858),
	.w7(32'h3bdb7a04),
	.w8(32'h3a959439),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f1a49),
	.w1(32'h3abcf1cf),
	.w2(32'hbb0ae31a),
	.w3(32'hbb323fef),
	.w4(32'hbad1da30),
	.w5(32'hba42e1b3),
	.w6(32'hbab7aad4),
	.w7(32'hba0498a3),
	.w8(32'hbb13cd1c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3896b0e7),
	.w1(32'h3aff29a8),
	.w2(32'h3ae7a4c6),
	.w3(32'h3a4ada81),
	.w4(32'h3b709888),
	.w5(32'h3a83d59f),
	.w6(32'hba5b987d),
	.w7(32'h3a8ceb2f),
	.w8(32'hbb10b71a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b91f0),
	.w1(32'hbbd03cc4),
	.w2(32'h3be91476),
	.w3(32'hbaef1561),
	.w4(32'hbbbe137b),
	.w5(32'h3afb280b),
	.w6(32'hbba82068),
	.w7(32'hbbfecb54),
	.w8(32'h3bd83e0f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a8d27),
	.w1(32'h3b8974d6),
	.w2(32'hbc051a83),
	.w3(32'hbc6bc4be),
	.w4(32'hbc536ea2),
	.w5(32'hbb5b8bc4),
	.w6(32'hbbd4e608),
	.w7(32'h3b6072f7),
	.w8(32'hbb1bd249),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26ec7b),
	.w1(32'hbb4ad593),
	.w2(32'h3acbefa9),
	.w3(32'hbafafc5b),
	.w4(32'h3c1990ba),
	.w5(32'hbc796e0e),
	.w6(32'h3b315548),
	.w7(32'h3c6b036f),
	.w8(32'hbbbf6ff1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc840c07),
	.w1(32'hb9bbd99f),
	.w2(32'h3c845459),
	.w3(32'hbb8aa378),
	.w4(32'h3a387cf0),
	.w5(32'h3b310a84),
	.w6(32'h3c0332d7),
	.w7(32'h3c0b04e0),
	.w8(32'hbbb1ace3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d73d2),
	.w1(32'h3b79689d),
	.w2(32'hb9c602da),
	.w3(32'h3c03d1b8),
	.w4(32'h3b5fd125),
	.w5(32'h3ab94b18),
	.w6(32'h3c1c8cfb),
	.w7(32'h3be0c859),
	.w8(32'h3aad3662),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaa57d),
	.w1(32'h3bbfe7e0),
	.w2(32'h3b972bd1),
	.w3(32'hbb680181),
	.w4(32'h3be49175),
	.w5(32'h3b2b6252),
	.w6(32'hbbaead6c),
	.w7(32'h3c0c4d80),
	.w8(32'h3b8115ca),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa54ac),
	.w1(32'hbb2d3f26),
	.w2(32'hbc1b6862),
	.w3(32'h3aa60104),
	.w4(32'hbb3b7ea7),
	.w5(32'hbc9b950c),
	.w6(32'h39e50675),
	.w7(32'hbbaa383a),
	.w8(32'hbc8e3bfe),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0d184),
	.w1(32'h3c283e88),
	.w2(32'h3ba580ba),
	.w3(32'h3b8c1342),
	.w4(32'h3c600a68),
	.w5(32'hbbd41900),
	.w6(32'hbb8ce522),
	.w7(32'h3b45e903),
	.w8(32'h3b397746),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943d706),
	.w1(32'h38829c2d),
	.w2(32'hbb3414fc),
	.w3(32'hbb6af647),
	.w4(32'hbbd71226),
	.w5(32'hbb8e51d3),
	.w6(32'hbad39af9),
	.w7(32'hbbfa9387),
	.w8(32'hbb22ca39),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4490a7),
	.w1(32'h3b72db13),
	.w2(32'h398349e2),
	.w3(32'h3c02e15a),
	.w4(32'h3c58e05d),
	.w5(32'h3b08090f),
	.w6(32'h3a885372),
	.w7(32'h3bd4a577),
	.w8(32'h3b841da1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16a134),
	.w1(32'h3c0aaaed),
	.w2(32'h3b886d0b),
	.w3(32'h397479a0),
	.w4(32'h3c7de00c),
	.w5(32'h391f02b8),
	.w6(32'h3b1de75a),
	.w7(32'h3ca47410),
	.w8(32'hba0f859b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bb7ab),
	.w1(32'hbb1e5450),
	.w2(32'h39679a20),
	.w3(32'hbb68d01d),
	.w4(32'hbbd5cc24),
	.w5(32'h3a27f1a8),
	.w6(32'hbb1a6ca0),
	.w7(32'hbc0be0bf),
	.w8(32'h39c6efbd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ba726),
	.w1(32'h39c5a670),
	.w2(32'hbb543e3f),
	.w3(32'hbab61edb),
	.w4(32'hbac11cf2),
	.w5(32'hbc51ccb6),
	.w6(32'hba4eb3b5),
	.w7(32'h3991cfd7),
	.w8(32'hbc908f9a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5a3a),
	.w1(32'h3cbcd73c),
	.w2(32'h3ca87c75),
	.w3(32'h3beb2c9f),
	.w4(32'h3cda3a34),
	.w5(32'h3ccb3bae),
	.w6(32'h3bbe9cb5),
	.w7(32'h3c6aa0a2),
	.w8(32'h3b9d8358),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bab07),
	.w1(32'hbb2744cb),
	.w2(32'h3acba622),
	.w3(32'h3bbdcaf4),
	.w4(32'hbbef9b59),
	.w5(32'hbb1cb708),
	.w6(32'h3c2be9ce),
	.w7(32'h3c911757),
	.w8(32'h3a6e23d9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f55c1),
	.w1(32'h3b80c62e),
	.w2(32'hbc9ae9a9),
	.w3(32'hba8e2bea),
	.w4(32'h3b242cb5),
	.w5(32'hbcdc22c9),
	.w6(32'hbb896556),
	.w7(32'hbb2b47fc),
	.w8(32'hbc1598fe),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cc983),
	.w1(32'h3c28bf79),
	.w2(32'h3b02c687),
	.w3(32'h3c3a44fc),
	.w4(32'h3cbffe3f),
	.w5(32'h3bbe7d88),
	.w6(32'h3c6f1877),
	.w7(32'h3cc9152d),
	.w8(32'h3bbc2c6c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39022679),
	.w1(32'h3b7b37ba),
	.w2(32'h3a6fbe73),
	.w3(32'hbad34cf3),
	.w4(32'hbb8b3feb),
	.w5(32'hbad797f7),
	.w6(32'h3b2e0e35),
	.w7(32'h3adef91f),
	.w8(32'hb9cbe4ea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ff273),
	.w1(32'h3b81e31a),
	.w2(32'h3c0e7fe8),
	.w3(32'h3c05b5d4),
	.w4(32'h3c0b36c3),
	.w5(32'h3d195c83),
	.w6(32'h3c2ccaf4),
	.w7(32'h3c1cfd62),
	.w8(32'h3cf91a2f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948c1c),
	.w1(32'hbc1a7d9e),
	.w2(32'h3be5c789),
	.w3(32'h3b082755),
	.w4(32'hbd27b04d),
	.w5(32'h3ce07898),
	.w6(32'h3b073d73),
	.w7(32'hbd180535),
	.w8(32'h3d233d7d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7f3a9),
	.w1(32'hbbe48d34),
	.w2(32'h3a7166b2),
	.w3(32'hbb09a7c3),
	.w4(32'hbd147056),
	.w5(32'h3ad5196f),
	.w6(32'h3bc61c83),
	.w7(32'hbcd919de),
	.w8(32'h3bab73cf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad27ca3),
	.w1(32'hbb41d1c8),
	.w2(32'hbc00f8a5),
	.w3(32'hbad351a9),
	.w4(32'hbbea88ee),
	.w5(32'hbb99a923),
	.w6(32'h395f5dac),
	.w7(32'hbb9e49dc),
	.w8(32'hbb24b2bf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010501),
	.w1(32'h3acfab25),
	.w2(32'h3ab71bc9),
	.w3(32'h3a8f94ae),
	.w4(32'hba96aa1b),
	.w5(32'hbc167e37),
	.w6(32'h3a63c403),
	.w7(32'hbb639a42),
	.w8(32'hbc1e4192),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa55e61),
	.w1(32'hbb9b322d),
	.w2(32'hbbcad5ec),
	.w3(32'hbb7fd10b),
	.w4(32'hbbad102a),
	.w5(32'hbc062813),
	.w6(32'hbaa92d73),
	.w7(32'hbbcd19a3),
	.w8(32'hbb5d6d69),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e8f9a),
	.w1(32'h3a8fbf53),
	.w2(32'hbbc0f2fe),
	.w3(32'hbb3d4864),
	.w4(32'h3aba8ab9),
	.w5(32'hbbe186a8),
	.w6(32'hba85c5f2),
	.w7(32'h3a38118f),
	.w8(32'hbb81e641),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1fd3a),
	.w1(32'hb9cc21fe),
	.w2(32'h3a6ca98f),
	.w3(32'hbb1e63bf),
	.w4(32'h3bc95070),
	.w5(32'h3ad59503),
	.w6(32'hbbdf854f),
	.w7(32'h3b4f0e2c),
	.w8(32'hbb2d5f79),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05890a),
	.w1(32'h3a8b72d7),
	.w2(32'h391062b9),
	.w3(32'h3b08eb4c),
	.w4(32'h3b8d7337),
	.w5(32'hbc40eddb),
	.w6(32'h3b856894),
	.w7(32'hba9d6c08),
	.w8(32'hbc080a01),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f3e38),
	.w1(32'h3b470770),
	.w2(32'h3beb5c3f),
	.w3(32'hb82d8d65),
	.w4(32'h3c8f9d07),
	.w5(32'h3cb0ab1d),
	.w6(32'h3c78d5c3),
	.w7(32'h3c643d20),
	.w8(32'h3cd1ba16),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbccda0),
	.w1(32'h3b2f1579),
	.w2(32'hbbe289eb),
	.w3(32'h3ba9f381),
	.w4(32'hbc079f8f),
	.w5(32'hbc14ed7f),
	.w6(32'h3a29f9e7),
	.w7(32'hbca0873f),
	.w8(32'hbc3895e5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1062cd),
	.w1(32'h3bc79372),
	.w2(32'h3b81f821),
	.w3(32'h3c803df1),
	.w4(32'h3ca48def),
	.w5(32'h3ada82ad),
	.w6(32'h3c547d3e),
	.w7(32'h3c987f2a),
	.w8(32'hbbfd1fce),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d40f),
	.w1(32'hbb4922a8),
	.w2(32'h3b107e22),
	.w3(32'hbbc8d7b0),
	.w4(32'hbc280fa9),
	.w5(32'hbae8df51),
	.w6(32'hbbf947c8),
	.w7(32'hbbc2ef40),
	.w8(32'h3ad60e2c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bd8a0),
	.w1(32'hbbdfcf3f),
	.w2(32'hbbcb0de7),
	.w3(32'hbbd62dcd),
	.w4(32'hbb90ddb3),
	.w5(32'h3c443682),
	.w6(32'hbc8be2da),
	.w7(32'hbba9f79d),
	.w8(32'h3c3c4407),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b992400),
	.w1(32'h3c15b6fa),
	.w2(32'hbbd9886a),
	.w3(32'h3b8111a1),
	.w4(32'h3aa1bb91),
	.w5(32'h3af4f4cd),
	.w6(32'hbb85eb16),
	.w7(32'hbc4e8b82),
	.w8(32'h3aaa1ff3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42ba5c),
	.w1(32'hb62fa4e3),
	.w2(32'hb9fb75e7),
	.w3(32'h3be11c60),
	.w4(32'h3c07c0c7),
	.w5(32'hbb8f174e),
	.w6(32'h3b52e1a5),
	.w7(32'h3b5fc652),
	.w8(32'hbb9ef379),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15799d),
	.w1(32'h3a68b896),
	.w2(32'hbb2822dc),
	.w3(32'hbb55d6e0),
	.w4(32'h3b0cf246),
	.w5(32'h3af1a33f),
	.w6(32'hba0737b0),
	.w7(32'h3bf98a34),
	.w8(32'h39bdd901),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63548d),
	.w1(32'h3b8e09f5),
	.w2(32'hba7fe814),
	.w3(32'h3ad81f25),
	.w4(32'h3b96e136),
	.w5(32'hb8f455e7),
	.w6(32'hbb868493),
	.w7(32'hbb943598),
	.w8(32'hba546773),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd7839),
	.w1(32'h3a28e828),
	.w2(32'hbb1f4929),
	.w3(32'h3ac1f903),
	.w4(32'hbb3a6d6d),
	.w5(32'h3c8830b7),
	.w6(32'h3ab124dd),
	.w7(32'hbb2cbe4c),
	.w8(32'h3ca535c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b249),
	.w1(32'h3b7a6de6),
	.w2(32'h3c3788fc),
	.w3(32'hb9e9265d),
	.w4(32'hbc70bd37),
	.w5(32'h3d10aa67),
	.w6(32'h3abc45de),
	.w7(32'hbc82b1c1),
	.w8(32'h3d25a5e9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1167d1),
	.w1(32'hbbce2850),
	.w2(32'h3ba75882),
	.w3(32'hbb6f7492),
	.w4(32'hbd1eb2e1),
	.w5(32'hbc16571d),
	.w6(32'hbb8b146d),
	.w7(32'hbd1ef919),
	.w8(32'hbbe352b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7c293),
	.w1(32'hba656ae9),
	.w2(32'hbb5a5777),
	.w3(32'h39da0ab1),
	.w4(32'h3c57aaed),
	.w5(32'hbb145550),
	.w6(32'h3a2468da),
	.w7(32'h3c3721d4),
	.w8(32'hbb8c8c78),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0acc8d),
	.w1(32'hbb38f59f),
	.w2(32'hba9a761e),
	.w3(32'hbb788f46),
	.w4(32'hbb955fd2),
	.w5(32'hba1a3e4f),
	.w6(32'hbbaf558c),
	.w7(32'hbbc28905),
	.w8(32'h3a3cb6e1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9843e7),
	.w1(32'hb9f67635),
	.w2(32'hbbb8aa8b),
	.w3(32'h3a8c5ff5),
	.w4(32'h397d2535),
	.w5(32'h3b178ba3),
	.w6(32'hb89f7ee5),
	.w7(32'h3acd63d7),
	.w8(32'h3b27a178),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ab2d),
	.w1(32'hbbc9c24b),
	.w2(32'hba852a01),
	.w3(32'hbc7ed119),
	.w4(32'h3b366fdd),
	.w5(32'hb9c14d50),
	.w6(32'hbc4cfb78),
	.w7(32'h3a55c725),
	.w8(32'hba41c3c0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab14b1e),
	.w1(32'h3ae69e47),
	.w2(32'hbb54d061),
	.w3(32'hb964ed16),
	.w4(32'hbab1cdb4),
	.w5(32'hbc485eb1),
	.w6(32'hba9c21f9),
	.w7(32'hba56b7a7),
	.w8(32'hbc0c94c5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934b529),
	.w1(32'h3a9ad43d),
	.w2(32'h3c257afd),
	.w3(32'hbc23317b),
	.w4(32'h373e2752),
	.w5(32'hbbfc4dba),
	.w6(32'hbc3ad311),
	.w7(32'h3c1ecc32),
	.w8(32'hbb7291f6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2f311),
	.w1(32'hbc341dd9),
	.w2(32'h3c0989cc),
	.w3(32'hbaec54e3),
	.w4(32'hbb463d8f),
	.w5(32'hbc025f7a),
	.w6(32'hbb38c17b),
	.w7(32'hba6b48cc),
	.w8(32'hbba1bd69),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd08ad),
	.w1(32'hbc26041c),
	.w2(32'hbaa4564e),
	.w3(32'h370bf2ed),
	.w4(32'hbc022192),
	.w5(32'h3af032d1),
	.w6(32'hbafe1222),
	.w7(32'hba07141c),
	.w8(32'h3abcca9d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac428fc),
	.w1(32'h3b8c00c0),
	.w2(32'h3b5858eb),
	.w3(32'h3b1c2134),
	.w4(32'hb93e5592),
	.w5(32'hba83dd6b),
	.w6(32'h3bcbd04c),
	.w7(32'h3af19b31),
	.w8(32'hbbd76a22),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f2f9a),
	.w1(32'h3b8b89da),
	.w2(32'h3c47ab3d),
	.w3(32'h3a5294ad),
	.w4(32'hb8b87bf5),
	.w5(32'h3cc714d2),
	.w6(32'h3bdf449e),
	.w7(32'h3bc14362),
	.w8(32'h3cde45ba),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99aa14),
	.w1(32'hbc7a8c38),
	.w2(32'h3bf2e38b),
	.w3(32'hbba46b3d),
	.w4(32'hbc9b2c7b),
	.w5(32'h3c152b3a),
	.w6(32'h3ab19ac4),
	.w7(32'hbc731c57),
	.w8(32'h3b990b89),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf27769),
	.w1(32'h3c170076),
	.w2(32'hbc01cc0d),
	.w3(32'h3cc56ec2),
	.w4(32'h3c247761),
	.w5(32'h3bd21486),
	.w6(32'h3c61398c),
	.w7(32'hbb523f71),
	.w8(32'hbb7bf54c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6f740),
	.w1(32'h3a782c58),
	.w2(32'h3c62058d),
	.w3(32'hbc0f621a),
	.w4(32'hbb8722e5),
	.w5(32'h3cf891c5),
	.w6(32'hba990995),
	.w7(32'h3bf4e8ac),
	.w8(32'h3c873147),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe165f),
	.w1(32'hbbebc099),
	.w2(32'hbad03de4),
	.w3(32'h3c535243),
	.w4(32'hba41a8f2),
	.w5(32'h3b4ab2c2),
	.w6(32'h3c5498d4),
	.w7(32'hbc072809),
	.w8(32'hbb28bcd2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81d7a2),
	.w1(32'hbb242a63),
	.w2(32'h3af2f35b),
	.w3(32'hbabd372f),
	.w4(32'hbb49873a),
	.w5(32'h3adf9e23),
	.w6(32'hbb861904),
	.w7(32'hbb853d69),
	.w8(32'h3a96546c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846b54),
	.w1(32'h3bb342e7),
	.w2(32'h397c7354),
	.w3(32'h3b400bb8),
	.w4(32'h39b714de),
	.w5(32'h3ad19cb5),
	.w6(32'h3b511053),
	.w7(32'hbb945d11),
	.w8(32'hba6ab4b0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d889b),
	.w1(32'h3a2554f1),
	.w2(32'h3a8ebeb5),
	.w3(32'hbb6f4287),
	.w4(32'h3bc7e380),
	.w5(32'hbbf41cb2),
	.w6(32'hbc239aa5),
	.w7(32'hbb729b0a),
	.w8(32'h38d1435c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952ef23),
	.w1(32'hbbd809ff),
	.w2(32'h3b0d1823),
	.w3(32'hbac4739c),
	.w4(32'hbb5fd70f),
	.w5(32'h3a053e11),
	.w6(32'hbb4a882a),
	.w7(32'hbb70927a),
	.w8(32'hba6d23b7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0a6e9),
	.w1(32'h396ddade),
	.w2(32'h3aa09433),
	.w3(32'h3a3d1678),
	.w4(32'hba9b9ef4),
	.w5(32'h3ca38e11),
	.w6(32'h3a2fbc45),
	.w7(32'h3a96a133),
	.w8(32'h3c5429a2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baa3d1),
	.w1(32'h3bfd9225),
	.w2(32'h388399aa),
	.w3(32'h3bfcbd3f),
	.w4(32'h3c26587b),
	.w5(32'h3b171442),
	.w6(32'h3b9c061a),
	.w7(32'hbc2d3cdd),
	.w8(32'h3b1cd3cb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8596e),
	.w1(32'h3afaaeae),
	.w2(32'hbb19c597),
	.w3(32'hb9bd4854),
	.w4(32'h3b296b3d),
	.w5(32'hbb37e2fd),
	.w6(32'h3ac38830),
	.w7(32'h3b2c541e),
	.w8(32'hba636cbc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605b8a),
	.w1(32'hb879c450),
	.w2(32'h3c121b73),
	.w3(32'hba9d12a2),
	.w4(32'h3c3cc85d),
	.w5(32'h3cd8d973),
	.w6(32'h3b595abc),
	.w7(32'h3c348f2d),
	.w8(32'h3aa8ca59),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32b01),
	.w1(32'hbcb3b1ce),
	.w2(32'h39ccda43),
	.w3(32'h379f4908),
	.w4(32'hbcefab94),
	.w5(32'h3b6a2c90),
	.w6(32'h3b63967b),
	.w7(32'h3b825aad),
	.w8(32'h3b1e8c8e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4bb9),
	.w1(32'h3b700bde),
	.w2(32'h3b2b0f40),
	.w3(32'h3b2a593b),
	.w4(32'h397a1e32),
	.w5(32'h3b27c1b6),
	.w6(32'h3b2c6cfa),
	.w7(32'h3b24a7a7),
	.w8(32'h3a5b437d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39226d),
	.w1(32'h397ccb47),
	.w2(32'h398db799),
	.w3(32'h3ae744df),
	.w4(32'hb895a13d),
	.w5(32'h3b593bac),
	.w6(32'h3a869c9a),
	.w7(32'h3aa21e24),
	.w8(32'hbb98d31c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701087),
	.w1(32'h3b1eafe9),
	.w2(32'h3b4bfa8e),
	.w3(32'h3abfc454),
	.w4(32'h3b3d27d1),
	.w5(32'hb8b9414f),
	.w6(32'hbb1a544a),
	.w7(32'h3a26165f),
	.w8(32'h3b84ddef),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb307a49),
	.w1(32'hba888be4),
	.w2(32'hbb735231),
	.w3(32'hba6dce5e),
	.w4(32'h3b4caae9),
	.w5(32'h39d303c5),
	.w6(32'h3b8fe103),
	.w7(32'h3bc02ec2),
	.w8(32'h3a573f52),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f92b9),
	.w1(32'h3c09f77c),
	.w2(32'hbb1d1b6e),
	.w3(32'h3c6087e2),
	.w4(32'h3bc680cf),
	.w5(32'hbab069bf),
	.w6(32'h3c18d49b),
	.w7(32'h3c3663ed),
	.w8(32'h3b3bc118),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834f89),
	.w1(32'hbb65cdd1),
	.w2(32'hbc9d52ae),
	.w3(32'h3aa04853),
	.w4(32'hbb00c162),
	.w5(32'hbc92895a),
	.w6(32'h3b3dbce6),
	.w7(32'hbb301454),
	.w8(32'hbc9af888),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31869f),
	.w1(32'h3c13a4a6),
	.w2(32'h3a682a45),
	.w3(32'hbc1b9d8f),
	.w4(32'h3cb9f85c),
	.w5(32'h3814f970),
	.w6(32'h3b8a56eb),
	.w7(32'h3ce18c70),
	.w8(32'h3bffcae2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb470b2b),
	.w1(32'h3bbe9d42),
	.w2(32'h3b293c38),
	.w3(32'h3b3670f9),
	.w4(32'hbb56f33a),
	.w5(32'h38a9bd73),
	.w6(32'h3a6ae318),
	.w7(32'hbb0bfcbf),
	.w8(32'h3a5e22e0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c7de7),
	.w1(32'hbb225298),
	.w2(32'hbb143d40),
	.w3(32'hbb5b9cb0),
	.w4(32'hbbdd9519),
	.w5(32'hbbbaee90),
	.w6(32'hbb8197f1),
	.w7(32'hbbbadc1f),
	.w8(32'hbb6190e7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9461812),
	.w1(32'h3a277498),
	.w2(32'h3c12b868),
	.w3(32'hbb41173b),
	.w4(32'h3bf27389),
	.w5(32'h3c8dd3df),
	.w6(32'hbb431d53),
	.w7(32'h3b70d730),
	.w8(32'hbb7085fa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66f3c5),
	.w1(32'hba2acefc),
	.w2(32'hbc27425d),
	.w3(32'h3c511ed4),
	.w4(32'hba0135a4),
	.w5(32'hbbbaef46),
	.w6(32'hbbc46827),
	.w7(32'h3c666770),
	.w8(32'hbbb626a9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ba65),
	.w1(32'h3c72aa64),
	.w2(32'h3a1f66f8),
	.w3(32'h3c429edd),
	.w4(32'h3cae89f5),
	.w5(32'h3b7a09d9),
	.w6(32'h3c39af07),
	.w7(32'h3c99ef10),
	.w8(32'h38d4610c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b82af),
	.w1(32'h3a7f582e),
	.w2(32'hbb0f2d62),
	.w3(32'h3c1662ae),
	.w4(32'h3ac4460f),
	.w5(32'h3bb02d6d),
	.w6(32'h3a26b955),
	.w7(32'hba88dcaf),
	.w8(32'h3bb27553),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2033ae),
	.w1(32'hbc008459),
	.w2(32'hbca5a58b),
	.w3(32'h3b191cf5),
	.w4(32'hbaaa8d71),
	.w5(32'hbc6d7a5e),
	.w6(32'h3a8b7fd7),
	.w7(32'h3b8afa9f),
	.w8(32'h3b79c6cb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9af6ed),
	.w1(32'hb94e8822),
	.w2(32'hbb02d622),
	.w3(32'hbc270aae),
	.w4(32'h390f6268),
	.w5(32'h39f24894),
	.w6(32'hbb81f46f),
	.w7(32'hbb895df9),
	.w8(32'h3ad5a6d2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae58843),
	.w1(32'hbb249e9a),
	.w2(32'hbc4c2033),
	.w3(32'h3b4d8bca),
	.w4(32'hba7535f5),
	.w5(32'hbcb28118),
	.w6(32'h3b8f7b6e),
	.w7(32'hba1f92ad),
	.w8(32'hbc881ae6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc1a0b),
	.w1(32'h3c3a3c2f),
	.w2(32'h3c169b9a),
	.w3(32'hbc14b747),
	.w4(32'h3c6a2fa8),
	.w5(32'hbc61ac40),
	.w6(32'hbbf90cd3),
	.w7(32'h3c7a9bf5),
	.w8(32'hbc9eaa23),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84282),
	.w1(32'h3c32189b),
	.w2(32'hb9e21bd9),
	.w3(32'h3acc127d),
	.w4(32'h3c4f23f3),
	.w5(32'hbabdcd2c),
	.w6(32'h3ac5f320),
	.w7(32'h3ba22b70),
	.w8(32'h3b0facab),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dad988),
	.w1(32'hbab49607),
	.w2(32'h3b040662),
	.w3(32'hbb5d0a78),
	.w4(32'hbbb9c65b),
	.w5(32'h3b57f156),
	.w6(32'hbada1ae4),
	.w7(32'hbb72b9f7),
	.w8(32'h3bf3e503),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5f777),
	.w1(32'h3c2b0dd3),
	.w2(32'h39160bf3),
	.w3(32'h3c392ad6),
	.w4(32'h3c3888fd),
	.w5(32'hba399534),
	.w6(32'hbad9602d),
	.w7(32'h3aa7d3fe),
	.w8(32'hb96bb77a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26a6bc),
	.w1(32'h3a08cd27),
	.w2(32'h3cca84a5),
	.w3(32'hbb2cdd39),
	.w4(32'hbac359a7),
	.w5(32'h3cb7c28a),
	.w6(32'hbb17550b),
	.w7(32'h3748f3fd),
	.w8(32'h3cb84eea),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bd3a5),
	.w1(32'h3cc6276c),
	.w2(32'hbbb143c0),
	.w3(32'h3d0d6074),
	.w4(32'h3ccac16b),
	.w5(32'h3c005b50),
	.w6(32'h3cb9c2bb),
	.w7(32'h3c923587),
	.w8(32'h3c06ca70),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9c24),
	.w1(32'hbc39a4ba),
	.w2(32'hbc31ba0a),
	.w3(32'h3c1089cb),
	.w4(32'h3b10c731),
	.w5(32'hbb66b73a),
	.w6(32'h3c4223fe),
	.w7(32'h3b277b77),
	.w8(32'hbac91193),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49fe2),
	.w1(32'hbb95f830),
	.w2(32'h39cd5831),
	.w3(32'hbbf758e9),
	.w4(32'h3c2b2c16),
	.w5(32'h3bcde7dd),
	.w6(32'hb9576200),
	.w7(32'h3b3ff963),
	.w8(32'h3b862171),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fd80a),
	.w1(32'hbaa70aac),
	.w2(32'h3aa93fc5),
	.w3(32'h3c16ceb5),
	.w4(32'hb8d06a21),
	.w5(32'hbb27bf6c),
	.w6(32'h3b690003),
	.w7(32'hbbb8a7c3),
	.w8(32'hbb23b519),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d8358),
	.w1(32'hba0b4afd),
	.w2(32'h3c11bd9e),
	.w3(32'hba3a189a),
	.w4(32'hbad2cf87),
	.w5(32'h3c52b02b),
	.w6(32'h3b03f427),
	.w7(32'h39b86b42),
	.w8(32'h3bfbc5cb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd1fd),
	.w1(32'hbac9d2f8),
	.w2(32'hbcbc0e37),
	.w3(32'h3b883ee5),
	.w4(32'h3bd02c10),
	.w5(32'hbce84730),
	.w6(32'h3bd39346),
	.w7(32'h3c365cb0),
	.w8(32'hbc0b11fe),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91d246),
	.w1(32'hbbb4d7fc),
	.w2(32'h3990e5fc),
	.w3(32'hbccee794),
	.w4(32'hba997b6b),
	.w5(32'h3b3de5e8),
	.w6(32'hbc14811f),
	.w7(32'hb9cb12a0),
	.w8(32'h3b76e231),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43c44f),
	.w1(32'hbac661c0),
	.w2(32'hbc53211e),
	.w3(32'h3ac57100),
	.w4(32'h3bc4eae3),
	.w5(32'hbb8bd2ea),
	.w6(32'h3b27ad12),
	.w7(32'h3b7f4c48),
	.w8(32'hbbb91d6a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb12a8e),
	.w1(32'hbcc49b1c),
	.w2(32'h3b00cbad),
	.w3(32'hbd295794),
	.w4(32'hbcbc03da),
	.w5(32'h3b4f3ce1),
	.w6(32'hbd099de3),
	.w7(32'hbcdfd85f),
	.w8(32'hbb8ee26a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1053e0),
	.w1(32'h3c15cfed),
	.w2(32'h3b9e1cea),
	.w3(32'h3c8df8ce),
	.w4(32'h3c284e3d),
	.w5(32'h3b9bb03e),
	.w6(32'h3b5601d3),
	.w7(32'h3b7eac70),
	.w8(32'h3ba9b459),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1acf2d),
	.w1(32'h3be8dc46),
	.w2(32'h3c4d2ef5),
	.w3(32'h3bf1340c),
	.w4(32'h3bde6adb),
	.w5(32'h3c83df87),
	.w6(32'h3c1f68fb),
	.w7(32'h3b24f8dc),
	.w8(32'h3c814c2f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72e8fc),
	.w1(32'hbb94c069),
	.w2(32'hbaa3fb9b),
	.w3(32'hbaeb8d5a),
	.w4(32'h3bbffd54),
	.w5(32'h3b01ca1e),
	.w6(32'h3b801241),
	.w7(32'hbc1bfc78),
	.w8(32'h3b0000a1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19bb3),
	.w1(32'hbb14aa5e),
	.w2(32'h3b75e2bd),
	.w3(32'h3b82e0fc),
	.w4(32'h3b87c403),
	.w5(32'hbc1531a3),
	.w6(32'h3ba804d0),
	.w7(32'h3bb24b21),
	.w8(32'hbc596304),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7150),
	.w1(32'hbb92fdb6),
	.w2(32'h3b9bc460),
	.w3(32'h3b4cc425),
	.w4(32'h3b41b286),
	.w5(32'h3c7e4c24),
	.w6(32'hbb3d3e3f),
	.w7(32'hbacd3477),
	.w8(32'h3c149f06),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb57b7d),
	.w1(32'h3c00d7e2),
	.w2(32'h3c018d1b),
	.w3(32'h3ccd2455),
	.w4(32'h3caf3272),
	.w5(32'hbc2a1f0d),
	.w6(32'h3c85a7a2),
	.w7(32'h3c58d934),
	.w8(32'hbc19fc3c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e92e),
	.w1(32'hbbdbca04),
	.w2(32'h3bf17bbe),
	.w3(32'h39a48dbc),
	.w4(32'hbb992337),
	.w5(32'h3c84c340),
	.w6(32'hbac7f788),
	.w7(32'hbaaff97e),
	.w8(32'h3c2d972b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e8830),
	.w1(32'hba8883e5),
	.w2(32'hbab44ff5),
	.w3(32'h3ce6605b),
	.w4(32'h3cb32839),
	.w5(32'hbbe93231),
	.w6(32'h3ccd4e6c),
	.w7(32'h3c8ce39f),
	.w8(32'hbbb94af1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8184),
	.w1(32'h3c2c3bd4),
	.w2(32'hbc2a92fb),
	.w3(32'hbb6763f8),
	.w4(32'h3b5936e3),
	.w5(32'hbc1d4e2a),
	.w6(32'h3b96817c),
	.w7(32'h3c33dbba),
	.w8(32'h3a1db9cc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a62404),
	.w1(32'h3bf9e4a9),
	.w2(32'h3c142d21),
	.w3(32'h3a091a01),
	.w4(32'h3c5f9c87),
	.w5(32'hbc3a7ee4),
	.w6(32'h3a30adb9),
	.w7(32'hbb6ec391),
	.w8(32'hbcc120e3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152d14),
	.w1(32'h3bbcbbeb),
	.w2(32'hba82df87),
	.w3(32'hbc440175),
	.w4(32'h3ba0e441),
	.w5(32'h3b2f1b6b),
	.w6(32'hbccd29c6),
	.w7(32'h3b11475c),
	.w8(32'h3c0302cd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5279bf),
	.w1(32'hbb3e02c6),
	.w2(32'hbc4cf0d6),
	.w3(32'h3c4cedde),
	.w4(32'hbb8e169f),
	.w5(32'hbbdae9b0),
	.w6(32'h3c434ea9),
	.w7(32'hbae3651b),
	.w8(32'hbbb2df3a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63928c),
	.w1(32'hbbfd7dfa),
	.w2(32'hbb6853c3),
	.w3(32'h39ccd086),
	.w4(32'hba55aeee),
	.w5(32'hbbe5efb7),
	.w6(32'h3b1f0905),
	.w7(32'h3a7b05b3),
	.w8(32'h3c53fd03),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c299c5),
	.w1(32'hbc7afa66),
	.w2(32'hbaf13d24),
	.w3(32'h3b6857ae),
	.w4(32'hbca7c94b),
	.w5(32'hbc7f36a8),
	.w6(32'h3c8e259e),
	.w7(32'hbb5567d5),
	.w8(32'hbc102628),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b59b9),
	.w1(32'h3c00ec8a),
	.w2(32'hbb727ea6),
	.w3(32'h3b1ceae5),
	.w4(32'h3c04ad8e),
	.w5(32'hbbfb3160),
	.w6(32'h3be21c0c),
	.w7(32'h3c312226),
	.w8(32'hbb7b5d9b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f412b),
	.w1(32'hbb0b1b8b),
	.w2(32'hbad8a414),
	.w3(32'hbb0f6b44),
	.w4(32'h3b30a492),
	.w5(32'hbbb70289),
	.w6(32'hbbb450b9),
	.w7(32'h3bdb1d2a),
	.w8(32'h3b741d9c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4bc4),
	.w1(32'h3c3a072f),
	.w2(32'hbbbb4134),
	.w3(32'h3ba21258),
	.w4(32'h3c34ace7),
	.w5(32'hbb402bab),
	.w6(32'h3acf0877),
	.w7(32'h3c0c7397),
	.w8(32'hbbf04407),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932538),
	.w1(32'h3bbe2524),
	.w2(32'h3a4a536a),
	.w3(32'h3b81ee39),
	.w4(32'h3b9ea0ba),
	.w5(32'h3c47f44e),
	.w6(32'h3b69f2bb),
	.w7(32'h3c555f0b),
	.w8(32'h3b204c69),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5f30),
	.w1(32'h3b405552),
	.w2(32'hbc16d7eb),
	.w3(32'h3c029fe5),
	.w4(32'h3bae9235),
	.w5(32'hbcbef3da),
	.w6(32'h3a6b21ce),
	.w7(32'h3b3f5a7f),
	.w8(32'hbd0d98f2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba400240),
	.w1(32'h3c054727),
	.w2(32'h3ba83f25),
	.w3(32'hbcd0fcc7),
	.w4(32'hba839e9c),
	.w5(32'h3b7a140a),
	.w6(32'hbd13ff09),
	.w7(32'hbc4605f7),
	.w8(32'h3a2ae4db),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd26389),
	.w1(32'h3b3f84db),
	.w2(32'hbb844692),
	.w3(32'h3bc163f7),
	.w4(32'h39519878),
	.w5(32'h3a8849df),
	.w6(32'h3add8f18),
	.w7(32'hba9ff54f),
	.w8(32'h3b21f842),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc82715),
	.w1(32'hbbdd5afb),
	.w2(32'hba9d2f24),
	.w3(32'h39eca8d8),
	.w4(32'h3b1581fc),
	.w5(32'h3c06db99),
	.w6(32'h3aa281d6),
	.w7(32'hbaa27de3),
	.w8(32'h3ac74a46),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72623),
	.w1(32'hbcaff6e5),
	.w2(32'h3b23c32c),
	.w3(32'hbc023425),
	.w4(32'hbc30dbd2),
	.w5(32'hbb9fe2a5),
	.w6(32'h3b51d9ec),
	.w7(32'hbb18469b),
	.w8(32'hbba386c3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b2dc),
	.w1(32'h3c4e41b5),
	.w2(32'h3c054216),
	.w3(32'h3c8c34d9),
	.w4(32'h3c94318e),
	.w5(32'h3c0ffe00),
	.w6(32'h3bd4c584),
	.w7(32'h3aee2f59),
	.w8(32'h3c289b52),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf8bdf),
	.w1(32'h3bb19387),
	.w2(32'h3b17d9ca),
	.w3(32'h3c06f19a),
	.w4(32'h3b62e27b),
	.w5(32'h3c0aa0ad),
	.w6(32'h3c23d83d),
	.w7(32'h3bb5bc4e),
	.w8(32'h3baef63d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc380e6c),
	.w1(32'hbb672a73),
	.w2(32'h396542a6),
	.w3(32'h3a571206),
	.w4(32'h3afe4ef5),
	.w5(32'h3b54ba4b),
	.w6(32'hba706a3c),
	.w7(32'h3b327fc3),
	.w8(32'h3ba467be),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1b90),
	.w1(32'h3adc2177),
	.w2(32'hbbf1cce8),
	.w3(32'hb9e7d9f8),
	.w4(32'h3b045228),
	.w5(32'hbbaf20c3),
	.w6(32'h3b4b0762),
	.w7(32'h3ae3e93b),
	.w8(32'hb9a4b464),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cd121),
	.w1(32'hbc57ac78),
	.w2(32'hbca14fe4),
	.w3(32'hbc54a5b4),
	.w4(32'hbce02b52),
	.w5(32'hbd1a56b2),
	.w6(32'hbb434447),
	.w7(32'hbc79578a),
	.w8(32'hbd013766),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf14b96),
	.w1(32'h3c847865),
	.w2(32'hb9f12cd9),
	.w3(32'h3b8c3de3),
	.w4(32'h3c85d797),
	.w5(32'h3a61e135),
	.w6(32'hb97140de),
	.w7(32'h3beec381),
	.w8(32'h3a452b54),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92962f2),
	.w1(32'h3aaaa63d),
	.w2(32'hbb8227c4),
	.w3(32'h3be231cf),
	.w4(32'h3bd5bad8),
	.w5(32'hbbc561fd),
	.w6(32'h3bb5879b),
	.w7(32'h3b2365eb),
	.w8(32'hbba658f5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0106b8),
	.w1(32'h3b74c480),
	.w2(32'hbc256bcc),
	.w3(32'hbc121115),
	.w4(32'h3b231e00),
	.w5(32'hbd0b1edf),
	.w6(32'hbc230aca),
	.w7(32'h3b0b6976),
	.w8(32'hbcf2e47e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab052ea),
	.w1(32'h3c67ad02),
	.w2(32'hbbba1b87),
	.w3(32'hbcc9fed2),
	.w4(32'h3c0e3e1b),
	.w5(32'hbd03230f),
	.w6(32'hbc986416),
	.w7(32'h3bd9367b),
	.w8(32'hbce3aeab),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03a302),
	.w1(32'h3ca4cdc5),
	.w2(32'h3b7f7607),
	.w3(32'hbc6961a5),
	.w4(32'h3c5064f0),
	.w5(32'h3c81eb8f),
	.w6(32'hbc74b791),
	.w7(32'hba1c304d),
	.w8(32'h3c737734),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97f88a),
	.w1(32'h3c1f503a),
	.w2(32'h3ae3a166),
	.w3(32'h3bbca739),
	.w4(32'h3b51194c),
	.w5(32'h3b9c1582),
	.w6(32'h3c80395c),
	.w7(32'h3c1eaabc),
	.w8(32'h3ae53000),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bbbab),
	.w1(32'h3b2e1c04),
	.w2(32'h3b1c7e3a),
	.w3(32'h3c14fbc9),
	.w4(32'h3b9cbe3c),
	.w5(32'h3bbacad5),
	.w6(32'hbb6370dc),
	.w7(32'h3ab79549),
	.w8(32'h399c3760),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5689d),
	.w1(32'hb9a2b0db),
	.w2(32'hba5354c6),
	.w3(32'hbb09555d),
	.w4(32'hbad0afcd),
	.w5(32'h3b5e85ac),
	.w6(32'hbbed0df8),
	.w7(32'hbb934717),
	.w8(32'h3b2a34d3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9ee8f),
	.w1(32'hba9b171c),
	.w2(32'h3c92620e),
	.w3(32'h3ba0a859),
	.w4(32'h3b915157),
	.w5(32'h3c6e2b8e),
	.w6(32'h3b058e8a),
	.w7(32'hba2d78e9),
	.w8(32'h3c92ce47),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fde5d),
	.w1(32'hbc549a3d),
	.w2(32'h3be317da),
	.w3(32'h3cf75474),
	.w4(32'hbae72b94),
	.w5(32'h3c7f6f2a),
	.w6(32'h3ced9b6f),
	.w7(32'hbb6f5fb7),
	.w8(32'h3bfb7fe6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf157db),
	.w1(32'h3bf8c957),
	.w2(32'hbbae9b65),
	.w3(32'h3b069455),
	.w4(32'h3bfec8f4),
	.w5(32'h3c42b07e),
	.w6(32'h3ad0f1b8),
	.w7(32'hb94a9be8),
	.w8(32'h3c0752bf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f538c),
	.w1(32'h3c08d2bc),
	.w2(32'h3b965762),
	.w3(32'h3c0ec73c),
	.w4(32'h3b4c804b),
	.w5(32'h3a8c2efc),
	.w6(32'h3c82fa91),
	.w7(32'h3c4399ce),
	.w8(32'hbaeabd7c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f07d5),
	.w1(32'hbc3d1df0),
	.w2(32'hbb156063),
	.w3(32'h3b49cc65),
	.w4(32'hbcba6805),
	.w5(32'hbbb068e8),
	.w6(32'h39b1c406),
	.w7(32'hbc807c6a),
	.w8(32'h3a007180),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344d82),
	.w1(32'hbbf11fd1),
	.w2(32'hbb1fc6b5),
	.w3(32'h3b916060),
	.w4(32'hbbf1adfa),
	.w5(32'hbb8e7b17),
	.w6(32'h3c155206),
	.w7(32'hbba85adb),
	.w8(32'hbb99e539),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165112),
	.w1(32'h3a615df4),
	.w2(32'h3c1df1dc),
	.w3(32'hbb65bf81),
	.w4(32'hbaec6e2a),
	.w5(32'h3c0d20e2),
	.w6(32'hbb872279),
	.w7(32'hbb2a531f),
	.w8(32'h3b19b37c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c675056),
	.w1(32'h3699c481),
	.w2(32'h3c5aaac6),
	.w3(32'h3cc26c9d),
	.w4(32'h3c540ebc),
	.w5(32'h3b9d88b5),
	.w6(32'h3c8416b4),
	.w7(32'h3c1e5623),
	.w8(32'h3b699826),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8525bb),
	.w1(32'h3c143659),
	.w2(32'h3b522c01),
	.w3(32'h3c4d5454),
	.w4(32'h3be1737e),
	.w5(32'hbb0c6f60),
	.w6(32'hbb18fa08),
	.w7(32'hba926af4),
	.w8(32'hba5e17f8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1e153),
	.w1(32'hbb9b2070),
	.w2(32'hbc080e15),
	.w3(32'hb92b107d),
	.w4(32'hbb05044e),
	.w5(32'h3b63dea1),
	.w6(32'h3bc1e8f0),
	.w7(32'hb9ab2332),
	.w8(32'h3ad93ed2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc434f19),
	.w1(32'hbc0b9527),
	.w2(32'h3b2e0a6f),
	.w3(32'h3bf98f23),
	.w4(32'h3b179dde),
	.w5(32'h3b10e793),
	.w6(32'h3c1af59e),
	.w7(32'h3c147bc9),
	.w8(32'h3a356bf5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8b6c),
	.w1(32'hbb71bf69),
	.w2(32'hbb87faf3),
	.w3(32'hbb3f0468),
	.w4(32'hbb90832f),
	.w5(32'hbb4596f0),
	.w6(32'hbb620ac9),
	.w7(32'hbb821dce),
	.w8(32'h3958801a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc157f41),
	.w1(32'hbb9c316e),
	.w2(32'h3a8a105b),
	.w3(32'hbac0cf61),
	.w4(32'hba206e84),
	.w5(32'h3abe5695),
	.w6(32'h399e4109),
	.w7(32'h3b1ee419),
	.w8(32'hba36d267),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59a9f8),
	.w1(32'h3c1cd809),
	.w2(32'h3b73f9f3),
	.w3(32'h3c8f8200),
	.w4(32'h3c899c3c),
	.w5(32'hbbe69ff2),
	.w6(32'h3bb43f67),
	.w7(32'h3b335546),
	.w8(32'hbc70f79d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf400ef),
	.w1(32'hbc3485ac),
	.w2(32'h3c0f24de),
	.w3(32'hbbf6529b),
	.w4(32'hbc25a50a),
	.w5(32'h3bc7f9c6),
	.w6(32'hbbc6f038),
	.w7(32'hbbe7c8f1),
	.w8(32'h3b8d98ba),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08063a),
	.w1(32'hbbcb6c73),
	.w2(32'hbc1a601c),
	.w3(32'h3b49dc53),
	.w4(32'hba911b71),
	.w5(32'hbc719f5f),
	.w6(32'hbb28361b),
	.w7(32'hbbfce7cb),
	.w8(32'h3af94cee),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe41084),
	.w1(32'hbb5578a7),
	.w2(32'h3b5f329c),
	.w3(32'h3c1484d0),
	.w4(32'h3c71e5e9),
	.w5(32'hbbb576df),
	.w6(32'h3c3e9fa3),
	.w7(32'h3c9ff939),
	.w8(32'hbc50b579),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d7f8b),
	.w1(32'h3c533c51),
	.w2(32'hbbe45822),
	.w3(32'h3aae85ad),
	.w4(32'h3cc3a987),
	.w5(32'h3b894d09),
	.w6(32'hbbabd31d),
	.w7(32'h3c696718),
	.w8(32'hbac5a6be),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1ec52),
	.w1(32'hbbaffbb4),
	.w2(32'hbce6bb10),
	.w3(32'hb9f09d56),
	.w4(32'h3c089b2b),
	.w5(32'hbd1d1a13),
	.w6(32'hbb2ca763),
	.w7(32'h3aad3f92),
	.w8(32'hbcabce8b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceafeed),
	.w1(32'hbc196560),
	.w2(32'hbc92f271),
	.w3(32'hbd6a74e8),
	.w4(32'hbcbef300),
	.w5(32'hbd245b98),
	.w6(32'hbd091228),
	.w7(32'hbbfb5bff),
	.w8(32'hbd327ee9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc931e39),
	.w1(32'hbab5380c),
	.w2(32'hbbac5c29),
	.w3(32'hbd662d0a),
	.w4(32'hbc810ef9),
	.w5(32'hbae506fa),
	.w6(32'hbd30bfa7),
	.w7(32'hbc952a4b),
	.w8(32'h3a695041),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba865320),
	.w1(32'h3a0072a2),
	.w2(32'h3b179120),
	.w3(32'h3b285d02),
	.w4(32'hba66fa30),
	.w5(32'hbbbdc594),
	.w6(32'h3b754c01),
	.w7(32'hbb6d427a),
	.w8(32'hbc4228a0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0291e3),
	.w1(32'h3bcc5bf1),
	.w2(32'h3c004096),
	.w3(32'hbc0d4d03),
	.w4(32'hbb7392ba),
	.w5(32'h3b85babb),
	.w6(32'hbb95b83b),
	.w7(32'hba964d34),
	.w8(32'h3b0feba1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4148d9),
	.w1(32'h3b02fbcb),
	.w2(32'h3bbedf0f),
	.w3(32'h3b6e49ce),
	.w4(32'h3c03731b),
	.w5(32'h3b4be4a4),
	.w6(32'hbac6c172),
	.w7(32'h3af63017),
	.w8(32'h3b173a97),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c056874),
	.w1(32'h3c2130f3),
	.w2(32'h3b506aec),
	.w3(32'h3bce98fd),
	.w4(32'h3b7b2b89),
	.w5(32'h3c0686eb),
	.w6(32'h3ad9ce65),
	.w7(32'h39f74791),
	.w8(32'h3b273fa4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae85ef8),
	.w1(32'hbbc344de),
	.w2(32'hbc3fcb6f),
	.w3(32'h3b6a2355),
	.w4(32'hbc2d2e32),
	.w5(32'hbaf49ed4),
	.w6(32'h3a235247),
	.w7(32'hbc33707f),
	.w8(32'hbaede255),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad907f),
	.w1(32'hba509cac),
	.w2(32'hbbe5871d),
	.w3(32'h3b232eac),
	.w4(32'h3be0e8e1),
	.w5(32'h3b0b68b0),
	.w6(32'hbaa2192a),
	.w7(32'h3a8a5d71),
	.w8(32'h3c594366),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7175),
	.w1(32'h3c47fde7),
	.w2(32'hba9f2fff),
	.w3(32'h3c64efbb),
	.w4(32'h3c163f28),
	.w5(32'hbc814d4f),
	.w6(32'h3c385217),
	.w7(32'hba761271),
	.w8(32'hbc733120),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227ad1),
	.w1(32'h3bf8c291),
	.w2(32'hbcc73c31),
	.w3(32'hbc40b0eb),
	.w4(32'h3aafbd45),
	.w5(32'hbca8e014),
	.w6(32'hbc0dbfde),
	.w7(32'h3b95fad5),
	.w8(32'hbc530263),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3ec57),
	.w1(32'hbbab2d5c),
	.w2(32'h3c1abde0),
	.w3(32'hbc4d8624),
	.w4(32'hbc0ab4e3),
	.w5(32'h3b04c4c7),
	.w6(32'hbc2cb0c0),
	.w7(32'h3c15eb9f),
	.w8(32'h3909dc7e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab230f2),
	.w1(32'hbb999ce1),
	.w2(32'h3ca69adf),
	.w3(32'h3b8923fd),
	.w4(32'h3bb40acd),
	.w5(32'h3cc7c145),
	.w6(32'hbbb2b033),
	.w7(32'h3addd86c),
	.w8(32'h3c509787),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35a810),
	.w1(32'hbbf8d269),
	.w2(32'hbc2ac737),
	.w3(32'h3c4388f8),
	.w4(32'hbb1d62d4),
	.w5(32'hbc1b7a13),
	.w6(32'h3ad9b0bc),
	.w7(32'h3acbd1fd),
	.w8(32'hbbed7fda),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83661c),
	.w1(32'h3bb1b8d9),
	.w2(32'h3b8e185a),
	.w3(32'h3b870f79),
	.w4(32'h3c55f919),
	.w5(32'hbc64fe54),
	.w6(32'h3b27fd3a),
	.w7(32'h3c32bf46),
	.w8(32'hbc490847),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1580df),
	.w1(32'hbbe385bc),
	.w2(32'hbad1e525),
	.w3(32'hbc40443d),
	.w4(32'hbb6b57f7),
	.w5(32'h3b00eb98),
	.w6(32'hbcaaec88),
	.w7(32'hbbc1b9a2),
	.w8(32'h3ba424ca),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae96af),
	.w1(32'hbbef87fd),
	.w2(32'hb8dcf1f8),
	.w3(32'hbafc96a4),
	.w4(32'hbb97c34d),
	.w5(32'hba535006),
	.w6(32'h39d6d222),
	.w7(32'hbbafa5d5),
	.w8(32'hbb7a29c6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc36a),
	.w1(32'hbb08b7f1),
	.w2(32'hbb1e3eee),
	.w3(32'h3bd246e7),
	.w4(32'h39952aaf),
	.w5(32'hbba78fa3),
	.w6(32'h3945b373),
	.w7(32'h3b11ecf8),
	.w8(32'hbafe7dca),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50640c),
	.w1(32'h3a32bb19),
	.w2(32'hbbc6fa35),
	.w3(32'hba1a83cd),
	.w4(32'h3b282c87),
	.w5(32'hbd0a5dba),
	.w6(32'h3512d78a),
	.w7(32'h3b9c0495),
	.w8(32'hbc9f085f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605ddb),
	.w1(32'h3c651d19),
	.w2(32'hbcaaf8d2),
	.w3(32'hbb90e49f),
	.w4(32'h3c757852),
	.w5(32'hbd387c7f),
	.w6(32'hbc124f4b),
	.w7(32'h3c0be6dc),
	.w8(32'hbd29bf6e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6a2f6),
	.w1(32'hbbc055d2),
	.w2(32'hbc12ccd2),
	.w3(32'hbd56aa58),
	.w4(32'hbcd1a309),
	.w5(32'hbc8ef05c),
	.w6(32'hbd3117a0),
	.w7(32'hbcc0bfb9),
	.w8(32'hbc712087),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23cba5),
	.w1(32'hbc0ab1fb),
	.w2(32'h3b7b4824),
	.w3(32'hbc35b777),
	.w4(32'hbbc378fd),
	.w5(32'h3b4d90dd),
	.w6(32'hbad0fa4a),
	.w7(32'h3ba99365),
	.w8(32'h3b3c148b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cae7f),
	.w1(32'h3b0c2400),
	.w2(32'hbaa42281),
	.w3(32'h3b60f765),
	.w4(32'h3a921819),
	.w5(32'hbb06d6d2),
	.w6(32'h3afedc13),
	.w7(32'h3b7ebd01),
	.w8(32'hba71ecd1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09ac4c),
	.w1(32'hbb39040f),
	.w2(32'h3b6716c1),
	.w3(32'hbae30f6b),
	.w4(32'hbb5d45ce),
	.w5(32'h3b552825),
	.w6(32'hbb0ca309),
	.w7(32'hbb0f8054),
	.w8(32'h3bc41828),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67161c),
	.w1(32'h3bde486c),
	.w2(32'hbb71e225),
	.w3(32'hbc3d7244),
	.w4(32'hbad13a52),
	.w5(32'hbb6bf66f),
	.w6(32'hbc1f97a5),
	.w7(32'hbb8364a3),
	.w8(32'hbaa48509),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cded0f),
	.w1(32'h3ac9b35f),
	.w2(32'h3c12fb9f),
	.w3(32'hba4ef03c),
	.w4(32'h3a8e4996),
	.w5(32'h38f2f5ce),
	.w6(32'h3b1a5e10),
	.w7(32'h3ae66f3b),
	.w8(32'h3ba3578d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be19dfe),
	.w1(32'hb9a418a9),
	.w2(32'hbc05d51d),
	.w3(32'h3c49aaa9),
	.w4(32'h3c060c4a),
	.w5(32'hbb7224ef),
	.w6(32'h3bbabbdd),
	.w7(32'h3c08f803),
	.w8(32'h3a2c05c4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cc837),
	.w1(32'hbca5420f),
	.w2(32'hbabed728),
	.w3(32'hbc95aa5d),
	.w4(32'hbc473942),
	.w5(32'hbb63de16),
	.w6(32'hbc4c9662),
	.w7(32'hbc463501),
	.w8(32'hbb4212ff),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc778560),
	.w1(32'hbc9de486),
	.w2(32'h3b61afd9),
	.w3(32'hbc98b0b1),
	.w4(32'hbcd0dc63),
	.w5(32'h384ced94),
	.w6(32'hbc81be21),
	.w7(32'hbc6a0e12),
	.w8(32'h3c049830),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule