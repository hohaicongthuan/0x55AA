module layer_11 (
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 16384;
	parameter IMG_SIZE = 13;

	wire	valid_out_0,
		valid_out_1,
		valid_out_2,
		valid_out_3,
		valid_out_4,
		valid_out_5,
		valid_out_6,
		valid_out_7,
		valid_out_8,
		valid_out_9,
		valid_out_10,
		valid_out_11,
		valid_out_12,
		valid_out_13,
		valid_out_14,
		valid_out_15,
		valid_out_16,
		valid_out_17,
		valid_out_18,
		valid_out_19,
		valid_out_20,
		valid_out_21,
		valid_out_22,
		valid_out_23,
		valid_out_24,
		valid_out_25,
		valid_out_26,
		valid_out_27,
		valid_out_28,
		valid_out_29,
		valid_out_30,
		valid_out_31,
		valid_out_32,
		valid_out_33,
		valid_out_34,
		valid_out_35,
		valid_out_36,
		valid_out_37,
		valid_out_38,
		valid_out_39,
		valid_out_40,
		valid_out_41,
		valid_out_42,
		valid_out_43,
		valid_out_44,
		valid_out_45,
		valid_out_46,
		valid_out_47,
		valid_out_48,
		valid_out_49,
		valid_out_50,
		valid_out_51,
		valid_out_52,
		valid_out_53,
		valid_out_54,
		valid_out_55,
		valid_out_56,
		valid_out_57,
		valid_out_58,
		valid_out_59,
		valid_out_60,
		valid_out_61,
		valid_out_62,
		valid_out_63,
		valid_out_64,
		valid_out_65,
		valid_out_66,
		valid_out_67,
		valid_out_68,
		valid_out_69,
		valid_out_70,
		valid_out_71,
		valid_out_72,
		valid_out_73,
		valid_out_74,
		valid_out_75,
		valid_out_76,
		valid_out_77,
		valid_out_78,
		valid_out_79,
		valid_out_80,
		valid_out_81,
		valid_out_82,
		valid_out_83,
		valid_out_84,
		valid_out_85,
		valid_out_86,
		valid_out_87,
		valid_out_88,
		valid_out_89,
		valid_out_90,
		valid_out_91,
		valid_out_92,
		valid_out_93,
		valid_out_94,
		valid_out_95,
		valid_out_96,
		valid_out_97,
		valid_out_98,
		valid_out_99,
		valid_out_100,
		valid_out_101,
		valid_out_102,
		valid_out_103,
		valid_out_104,
		valid_out_105,
		valid_out_106,
		valid_out_107,
		valid_out_108,
		valid_out_109,
		valid_out_110,
		valid_out_111,
		valid_out_112,
		valid_out_113,
		valid_out_114,
		valid_out_115,
		valid_out_116,
		valid_out_117,
		valid_out_118,
		valid_out_119,
		valid_out_120,
		valid_out_121,
		valid_out_122,
		valid_out_123,
		valid_out_124,
		valid_out_125,
		valid_out_126,
		valid_out_127,
		valid_out_128,
		valid_out_129,
		valid_out_130,
		valid_out_131,
		valid_out_132,
		valid_out_133,
		valid_out_134,
		valid_out_135,
		valid_out_136,
		valid_out_137,
		valid_out_138,
		valid_out_139,
		valid_out_140,
		valid_out_141,
		valid_out_142,
		valid_out_143,
		valid_out_144,
		valid_out_145,
		valid_out_146,
		valid_out_147,
		valid_out_148,
		valid_out_149,
		valid_out_150,
		valid_out_151,
		valid_out_152,
		valid_out_153,
		valid_out_154,
		valid_out_155,
		valid_out_156,
		valid_out_157,
		valid_out_158,
		valid_out_159,
		valid_out_160,
		valid_out_161,
		valid_out_162,
		valid_out_163,
		valid_out_164,
		valid_out_165,
		valid_out_166,
		valid_out_167,
		valid_out_168,
		valid_out_169,
		valid_out_170,
		valid_out_171,
		valid_out_172,
		valid_out_173,
		valid_out_174,
		valid_out_175,
		valid_out_176,
		valid_out_177,
		valid_out_178,
		valid_out_179,
		valid_out_180,
		valid_out_181,
		valid_out_182,
		valid_out_183,
		valid_out_184,
		valid_out_185,
		valid_out_186,
		valid_out_187,
		valid_out_188,
		valid_out_189,
		valid_out_190,
		valid_out_191,
		valid_out_192,
		valid_out_193,
		valid_out_194,
		valid_out_195,
		valid_out_196,
		valid_out_197,
		valid_out_198,
		valid_out_199,
		valid_out_200,
		valid_out_201,
		valid_out_202,
		valid_out_203,
		valid_out_204,
		valid_out_205,
		valid_out_206,
		valid_out_207,
		valid_out_208,
		valid_out_209,
		valid_out_210,
		valid_out_211,
		valid_out_212,
		valid_out_213,
		valid_out_214,
		valid_out_215,
		valid_out_216,
		valid_out_217,
		valid_out_218,
		valid_out_219,
		valid_out_220,
		valid_out_221,
		valid_out_222,
		valid_out_223,
		valid_out_224,
		valid_out_225,
		valid_out_226,
		valid_out_227,
		valid_out_228,
		valid_out_229,
		valid_out_230,
		valid_out_231,
		valid_out_232,
		valid_out_233,
		valid_out_234,
		valid_out_235,
		valid_out_236,
		valid_out_237,
		valid_out_238,
		valid_out_239,
		valid_out_240,
		valid_out_241,
		valid_out_242,
		valid_out_243,
		valid_out_244,
		valid_out_245,
		valid_out_246,
		valid_out_247,
		valid_out_248,
		valid_out_249,
		valid_out_250,
		valid_out_251,
		valid_out_252,
		valid_out_253,
		valid_out_254,
		valid_out_255,
		valid_out_256,
		valid_out_257,
		valid_out_258,
		valid_out_259,
		valid_out_260,
		valid_out_261,
		valid_out_262,
		valid_out_263,
		valid_out_264,
		valid_out_265,
		valid_out_266,
		valid_out_267,
		valid_out_268,
		valid_out_269,
		valid_out_270,
		valid_out_271,
		valid_out_272,
		valid_out_273,
		valid_out_274,
		valid_out_275,
		valid_out_276,
		valid_out_277,
		valid_out_278,
		valid_out_279,
		valid_out_280,
		valid_out_281,
		valid_out_282,
		valid_out_283,
		valid_out_284,
		valid_out_285,
		valid_out_286,
		valid_out_287,
		valid_out_288,
		valid_out_289,
		valid_out_290,
		valid_out_291,
		valid_out_292,
		valid_out_293,
		valid_out_294,
		valid_out_295,
		valid_out_296,
		valid_out_297,
		valid_out_298,
		valid_out_299,
		valid_out_300,
		valid_out_301,
		valid_out_302,
		valid_out_303,
		valid_out_304,
		valid_out_305,
		valid_out_306,
		valid_out_307,
		valid_out_308,
		valid_out_309,
		valid_out_310,
		valid_out_311,
		valid_out_312,
		valid_out_313,
		valid_out_314,
		valid_out_315,
		valid_out_316,
		valid_out_317,
		valid_out_318,
		valid_out_319,
		valid_out_320,
		valid_out_321,
		valid_out_322,
		valid_out_323,
		valid_out_324,
		valid_out_325,
		valid_out_326,
		valid_out_327,
		valid_out_328,
		valid_out_329,
		valid_out_330,
		valid_out_331,
		valid_out_332,
		valid_out_333,
		valid_out_334,
		valid_out_335,
		valid_out_336,
		valid_out_337,
		valid_out_338,
		valid_out_339,
		valid_out_340,
		valid_out_341,
		valid_out_342,
		valid_out_343,
		valid_out_344,
		valid_out_345,
		valid_out_346,
		valid_out_347,
		valid_out_348,
		valid_out_349,
		valid_out_350,
		valid_out_351,
		valid_out_352,
		valid_out_353,
		valid_out_354,
		valid_out_355,
		valid_out_356,
		valid_out_357,
		valid_out_358,
		valid_out_359,
		valid_out_360,
		valid_out_361,
		valid_out_362,
		valid_out_363,
		valid_out_364,
		valid_out_365,
		valid_out_366,
		valid_out_367,
		valid_out_368,
		valid_out_369,
		valid_out_370,
		valid_out_371,
		valid_out_372,
		valid_out_373,
		valid_out_374,
		valid_out_375,
		valid_out_376,
		valid_out_377,
		valid_out_378,
		valid_out_379,
		valid_out_380,
		valid_out_381,
		valid_out_382,
		valid_out_383,
		valid_out_384,
		valid_out_385,
		valid_out_386,
		valid_out_387,
		valid_out_388,
		valid_out_389,
		valid_out_390,
		valid_out_391,
		valid_out_392,
		valid_out_393,
		valid_out_394,
		valid_out_395,
		valid_out_396,
		valid_out_397,
		valid_out_398,
		valid_out_399,
		valid_out_400,
		valid_out_401,
		valid_out_402,
		valid_out_403,
		valid_out_404,
		valid_out_405,
		valid_out_406,
		valid_out_407,
		valid_out_408,
		valid_out_409,
		valid_out_410,
		valid_out_411,
		valid_out_412,
		valid_out_413,
		valid_out_414,
		valid_out_415,
		valid_out_416,
		valid_out_417,
		valid_out_418,
		valid_out_419,
		valid_out_420,
		valid_out_421,
		valid_out_422,
		valid_out_423,
		valid_out_424,
		valid_out_425,
		valid_out_426,
		valid_out_427,
		valid_out_428,
		valid_out_429,
		valid_out_430,
		valid_out_431,
		valid_out_432,
		valid_out_433,
		valid_out_434,
		valid_out_435,
		valid_out_436,
		valid_out_437,
		valid_out_438,
		valid_out_439,
		valid_out_440,
		valid_out_441,
		valid_out_442,
		valid_out_443,
		valid_out_444,
		valid_out_445,
		valid_out_446,
		valid_out_447,
		valid_out_448,
		valid_out_449,
		valid_out_450,
		valid_out_451,
		valid_out_452,
		valid_out_453,
		valid_out_454,
		valid_out_455,
		valid_out_456,
		valid_out_457,
		valid_out_458,
		valid_out_459,
		valid_out_460,
		valid_out_461,
		valid_out_462,
		valid_out_463,
		valid_out_464,
		valid_out_465,
		valid_out_466,
		valid_out_467,
		valid_out_468,
		valid_out_469,
		valid_out_470,
		valid_out_471,
		valid_out_472,
		valid_out_473,
		valid_out_474,
		valid_out_475,
		valid_out_476,
		valid_out_477,
		valid_out_478,
		valid_out_479,
		valid_out_480,
		valid_out_481,
		valid_out_482,
		valid_out_483,
		valid_out_484,
		valid_out_485,
		valid_out_486,
		valid_out_487,
		valid_out_488,
		valid_out_489,
		valid_out_490,
		valid_out_491,
		valid_out_492,
		valid_out_493,
		valid_out_494,
		valid_out_495,
		valid_out_496,
		valid_out_497,
		valid_out_498,
		valid_out_499,
		valid_out_500,
		valid_out_501,
		valid_out_502,
		valid_out_503,
		valid_out_504,
		valid_out_505,
		valid_out_506,
		valid_out_507,
		valid_out_508,
		valid_out_509,
		valid_out_510,
		valid_out_511;
Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(data_out[31:0]),
	.valid_out(valid_out_0)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(data_out[63:32]),
	.valid_out(valid_out_1)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(data_out[95:64]),
	.valid_out(valid_out_2)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(data_out[127:96]),
	.valid_out(valid_out_3)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(data_out[159:128]),
	.valid_out(valid_out_4)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(data_out[191:160]),
	.valid_out(valid_out_5)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(data_out[223:192]),
	.valid_out(valid_out_6)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(data_out[255:224]),
	.valid_out(valid_out_7)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(data_out[287:256]),
	.valid_out(valid_out_8)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(data_out[319:288]),
	.valid_out(valid_out_9)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(data_out[351:320]),
	.valid_out(valid_out_10)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(data_out[383:352]),
	.valid_out(valid_out_11)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(data_out[415:384]),
	.valid_out(valid_out_12)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(data_out[447:416]),
	.valid_out(valid_out_13)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(data_out[479:448]),
	.valid_out(valid_out_14)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(data_out[511:480]),
	.valid_out(valid_out_15)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(data_out[543:512]),
	.valid_out(valid_out_16)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(data_out[575:544]),
	.valid_out(valid_out_17)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(data_out[607:576]),
	.valid_out(valid_out_18)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(data_out[639:608]),
	.valid_out(valid_out_19)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(data_out[671:640]),
	.valid_out(valid_out_20)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(data_out[703:672]),
	.valid_out(valid_out_21)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(data_out[735:704]),
	.valid_out(valid_out_22)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(data_out[767:736]),
	.valid_out(valid_out_23)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(data_out[799:768]),
	.valid_out(valid_out_24)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(data_out[831:800]),
	.valid_out(valid_out_25)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(data_out[863:832]),
	.valid_out(valid_out_26)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(data_out[895:864]),
	.valid_out(valid_out_27)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(data_out[927:896]),
	.valid_out(valid_out_28)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(data_out[959:928]),
	.valid_out(valid_out_29)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(data_out[991:960]),
	.valid_out(valid_out_30)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(data_out[1023:992]),
	.valid_out(valid_out_31)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(data_out[1055:1024]),
	.valid_out(valid_out_32)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(data_out[1087:1056]),
	.valid_out(valid_out_33)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(data_out[1119:1088]),
	.valid_out(valid_out_34)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(data_out[1151:1120]),
	.valid_out(valid_out_35)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(data_out[1183:1152]),
	.valid_out(valid_out_36)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(data_out[1215:1184]),
	.valid_out(valid_out_37)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(data_out[1247:1216]),
	.valid_out(valid_out_38)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(data_out[1279:1248]),
	.valid_out(valid_out_39)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(data_out[1311:1280]),
	.valid_out(valid_out_40)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(data_out[1343:1312]),
	.valid_out(valid_out_41)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(data_out[1375:1344]),
	.valid_out(valid_out_42)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(data_out[1407:1376]),
	.valid_out(valid_out_43)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(data_out[1439:1408]),
	.valid_out(valid_out_44)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(data_out[1471:1440]),
	.valid_out(valid_out_45)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(data_out[1503:1472]),
	.valid_out(valid_out_46)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(data_out[1535:1504]),
	.valid_out(valid_out_47)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(data_out[1567:1536]),
	.valid_out(valid_out_48)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(data_out[1599:1568]),
	.valid_out(valid_out_49)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(data_out[1631:1600]),
	.valid_out(valid_out_50)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(data_out[1663:1632]),
	.valid_out(valid_out_51)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(data_out[1695:1664]),
	.valid_out(valid_out_52)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(data_out[1727:1696]),
	.valid_out(valid_out_53)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(data_out[1759:1728]),
	.valid_out(valid_out_54)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(data_out[1791:1760]),
	.valid_out(valid_out_55)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(data_out[1823:1792]),
	.valid_out(valid_out_56)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(data_out[1855:1824]),
	.valid_out(valid_out_57)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(data_out[1887:1856]),
	.valid_out(valid_out_58)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(data_out[1919:1888]),
	.valid_out(valid_out_59)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(data_out[1951:1920]),
	.valid_out(valid_out_60)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(data_out[1983:1952]),
	.valid_out(valid_out_61)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(data_out[2015:1984]),
	.valid_out(valid_out_62)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(data_out[2047:2016]),
	.valid_out(valid_out_63)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(data_out[2079:2048]),
	.valid_out(valid_out_64)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(data_out[2111:2080]),
	.valid_out(valid_out_65)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(data_out[2143:2112]),
	.valid_out(valid_out_66)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(data_out[2175:2144]),
	.valid_out(valid_out_67)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(data_out[2207:2176]),
	.valid_out(valid_out_68)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(data_out[2239:2208]),
	.valid_out(valid_out_69)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(data_out[2271:2240]),
	.valid_out(valid_out_70)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(data_out[2303:2272]),
	.valid_out(valid_out_71)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(data_out[2335:2304]),
	.valid_out(valid_out_72)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(data_out[2367:2336]),
	.valid_out(valid_out_73)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(data_out[2399:2368]),
	.valid_out(valid_out_74)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(data_out[2431:2400]),
	.valid_out(valid_out_75)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(data_out[2463:2432]),
	.valid_out(valid_out_76)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(data_out[2495:2464]),
	.valid_out(valid_out_77)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(data_out[2527:2496]),
	.valid_out(valid_out_78)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(data_out[2559:2528]),
	.valid_out(valid_out_79)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(data_out[2591:2560]),
	.valid_out(valid_out_80)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(data_out[2623:2592]),
	.valid_out(valid_out_81)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(data_out[2655:2624]),
	.valid_out(valid_out_82)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(data_out[2687:2656]),
	.valid_out(valid_out_83)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(data_out[2719:2688]),
	.valid_out(valid_out_84)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(data_out[2751:2720]),
	.valid_out(valid_out_85)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(data_out[2783:2752]),
	.valid_out(valid_out_86)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(data_out[2815:2784]),
	.valid_out(valid_out_87)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(data_out[2847:2816]),
	.valid_out(valid_out_88)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(data_out[2879:2848]),
	.valid_out(valid_out_89)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(data_out[2911:2880]),
	.valid_out(valid_out_90)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(data_out[2943:2912]),
	.valid_out(valid_out_91)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(data_out[2975:2944]),
	.valid_out(valid_out_92)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(data_out[3007:2976]),
	.valid_out(valid_out_93)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(data_out[3039:3008]),
	.valid_out(valid_out_94)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(data_out[3071:3040]),
	.valid_out(valid_out_95)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(data_out[3103:3072]),
	.valid_out(valid_out_96)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(data_out[3135:3104]),
	.valid_out(valid_out_97)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(data_out[3167:3136]),
	.valid_out(valid_out_98)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(data_out[3199:3168]),
	.valid_out(valid_out_99)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(data_out[3231:3200]),
	.valid_out(valid_out_100)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(data_out[3263:3232]),
	.valid_out(valid_out_101)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(data_out[3295:3264]),
	.valid_out(valid_out_102)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(data_out[3327:3296]),
	.valid_out(valid_out_103)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(data_out[3359:3328]),
	.valid_out(valid_out_104)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(data_out[3391:3360]),
	.valid_out(valid_out_105)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(data_out[3423:3392]),
	.valid_out(valid_out_106)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(data_out[3455:3424]),
	.valid_out(valid_out_107)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(data_out[3487:3456]),
	.valid_out(valid_out_108)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(data_out[3519:3488]),
	.valid_out(valid_out_109)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(data_out[3551:3520]),
	.valid_out(valid_out_110)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(data_out[3583:3552]),
	.valid_out(valid_out_111)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(data_out[3615:3584]),
	.valid_out(valid_out_112)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(data_out[3647:3616]),
	.valid_out(valid_out_113)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(data_out[3679:3648]),
	.valid_out(valid_out_114)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(data_out[3711:3680]),
	.valid_out(valid_out_115)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(data_out[3743:3712]),
	.valid_out(valid_out_116)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(data_out[3775:3744]),
	.valid_out(valid_out_117)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(data_out[3807:3776]),
	.valid_out(valid_out_118)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(data_out[3839:3808]),
	.valid_out(valid_out_119)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(data_out[3871:3840]),
	.valid_out(valid_out_120)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(data_out[3903:3872]),
	.valid_out(valid_out_121)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(data_out[3935:3904]),
	.valid_out(valid_out_122)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(data_out[3967:3936]),
	.valid_out(valid_out_123)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(data_out[3999:3968]),
	.valid_out(valid_out_124)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(data_out[4031:4000]),
	.valid_out(valid_out_125)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(data_out[4063:4032]),
	.valid_out(valid_out_126)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(data_out[4095:4064]),
	.valid_out(valid_out_127)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(data_out[4127:4096]),
	.valid_out(valid_out_128)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(data_out[4159:4128]),
	.valid_out(valid_out_129)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(data_out[4191:4160]),
	.valid_out(valid_out_130)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(data_out[4223:4192]),
	.valid_out(valid_out_131)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(data_out[4255:4224]),
	.valid_out(valid_out_132)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(data_out[4287:4256]),
	.valid_out(valid_out_133)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(data_out[4319:4288]),
	.valid_out(valid_out_134)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(data_out[4351:4320]),
	.valid_out(valid_out_135)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(data_out[4383:4352]),
	.valid_out(valid_out_136)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(data_out[4415:4384]),
	.valid_out(valid_out_137)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(data_out[4447:4416]),
	.valid_out(valid_out_138)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(data_out[4479:4448]),
	.valid_out(valid_out_139)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(data_out[4511:4480]),
	.valid_out(valid_out_140)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(data_out[4543:4512]),
	.valid_out(valid_out_141)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(data_out[4575:4544]),
	.valid_out(valid_out_142)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(data_out[4607:4576]),
	.valid_out(valid_out_143)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(data_out[4639:4608]),
	.valid_out(valid_out_144)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(data_out[4671:4640]),
	.valid_out(valid_out_145)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(data_out[4703:4672]),
	.valid_out(valid_out_146)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(data_out[4735:4704]),
	.valid_out(valid_out_147)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(data_out[4767:4736]),
	.valid_out(valid_out_148)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(data_out[4799:4768]),
	.valid_out(valid_out_149)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(data_out[4831:4800]),
	.valid_out(valid_out_150)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(data_out[4863:4832]),
	.valid_out(valid_out_151)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(data_out[4895:4864]),
	.valid_out(valid_out_152)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(data_out[4927:4896]),
	.valid_out(valid_out_153)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(data_out[4959:4928]),
	.valid_out(valid_out_154)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(data_out[4991:4960]),
	.valid_out(valid_out_155)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(data_out[5023:4992]),
	.valid_out(valid_out_156)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(data_out[5055:5024]),
	.valid_out(valid_out_157)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(data_out[5087:5056]),
	.valid_out(valid_out_158)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(data_out[5119:5088]),
	.valid_out(valid_out_159)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(data_out[5151:5120]),
	.valid_out(valid_out_160)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(data_out[5183:5152]),
	.valid_out(valid_out_161)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(data_out[5215:5184]),
	.valid_out(valid_out_162)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(data_out[5247:5216]),
	.valid_out(valid_out_163)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(data_out[5279:5248]),
	.valid_out(valid_out_164)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(data_out[5311:5280]),
	.valid_out(valid_out_165)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(data_out[5343:5312]),
	.valid_out(valid_out_166)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(data_out[5375:5344]),
	.valid_out(valid_out_167)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(data_out[5407:5376]),
	.valid_out(valid_out_168)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(data_out[5439:5408]),
	.valid_out(valid_out_169)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(data_out[5471:5440]),
	.valid_out(valid_out_170)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(data_out[5503:5472]),
	.valid_out(valid_out_171)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(data_out[5535:5504]),
	.valid_out(valid_out_172)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(data_out[5567:5536]),
	.valid_out(valid_out_173)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(data_out[5599:5568]),
	.valid_out(valid_out_174)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(data_out[5631:5600]),
	.valid_out(valid_out_175)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(data_out[5663:5632]),
	.valid_out(valid_out_176)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(data_out[5695:5664]),
	.valid_out(valid_out_177)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(data_out[5727:5696]),
	.valid_out(valid_out_178)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(data_out[5759:5728]),
	.valid_out(valid_out_179)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(data_out[5791:5760]),
	.valid_out(valid_out_180)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(data_out[5823:5792]),
	.valid_out(valid_out_181)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(data_out[5855:5824]),
	.valid_out(valid_out_182)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(data_out[5887:5856]),
	.valid_out(valid_out_183)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(data_out[5919:5888]),
	.valid_out(valid_out_184)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(data_out[5951:5920]),
	.valid_out(valid_out_185)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(data_out[5983:5952]),
	.valid_out(valid_out_186)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(data_out[6015:5984]),
	.valid_out(valid_out_187)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(data_out[6047:6016]),
	.valid_out(valid_out_188)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(data_out[6079:6048]),
	.valid_out(valid_out_189)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(data_out[6111:6080]),
	.valid_out(valid_out_190)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(data_out[6143:6112]),
	.valid_out(valid_out_191)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(data_out[6175:6144]),
	.valid_out(valid_out_192)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(data_out[6207:6176]),
	.valid_out(valid_out_193)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(data_out[6239:6208]),
	.valid_out(valid_out_194)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(data_out[6271:6240]),
	.valid_out(valid_out_195)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(data_out[6303:6272]),
	.valid_out(valid_out_196)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(data_out[6335:6304]),
	.valid_out(valid_out_197)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(data_out[6367:6336]),
	.valid_out(valid_out_198)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(data_out[6399:6368]),
	.valid_out(valid_out_199)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(data_out[6431:6400]),
	.valid_out(valid_out_200)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(data_out[6463:6432]),
	.valid_out(valid_out_201)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(data_out[6495:6464]),
	.valid_out(valid_out_202)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(data_out[6527:6496]),
	.valid_out(valid_out_203)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(data_out[6559:6528]),
	.valid_out(valid_out_204)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(data_out[6591:6560]),
	.valid_out(valid_out_205)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(data_out[6623:6592]),
	.valid_out(valid_out_206)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(data_out[6655:6624]),
	.valid_out(valid_out_207)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(data_out[6687:6656]),
	.valid_out(valid_out_208)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(data_out[6719:6688]),
	.valid_out(valid_out_209)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(data_out[6751:6720]),
	.valid_out(valid_out_210)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(data_out[6783:6752]),
	.valid_out(valid_out_211)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(data_out[6815:6784]),
	.valid_out(valid_out_212)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(data_out[6847:6816]),
	.valid_out(valid_out_213)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(data_out[6879:6848]),
	.valid_out(valid_out_214)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(data_out[6911:6880]),
	.valid_out(valid_out_215)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(data_out[6943:6912]),
	.valid_out(valid_out_216)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(data_out[6975:6944]),
	.valid_out(valid_out_217)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(data_out[7007:6976]),
	.valid_out(valid_out_218)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(data_out[7039:7008]),
	.valid_out(valid_out_219)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(data_out[7071:7040]),
	.valid_out(valid_out_220)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(data_out[7103:7072]),
	.valid_out(valid_out_221)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(data_out[7135:7104]),
	.valid_out(valid_out_222)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(data_out[7167:7136]),
	.valid_out(valid_out_223)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(data_out[7199:7168]),
	.valid_out(valid_out_224)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(data_out[7231:7200]),
	.valid_out(valid_out_225)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(data_out[7263:7232]),
	.valid_out(valid_out_226)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(data_out[7295:7264]),
	.valid_out(valid_out_227)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(data_out[7327:7296]),
	.valid_out(valid_out_228)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(data_out[7359:7328]),
	.valid_out(valid_out_229)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(data_out[7391:7360]),
	.valid_out(valid_out_230)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(data_out[7423:7392]),
	.valid_out(valid_out_231)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(data_out[7455:7424]),
	.valid_out(valid_out_232)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(data_out[7487:7456]),
	.valid_out(valid_out_233)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(data_out[7519:7488]),
	.valid_out(valid_out_234)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(data_out[7551:7520]),
	.valid_out(valid_out_235)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(data_out[7583:7552]),
	.valid_out(valid_out_236)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(data_out[7615:7584]),
	.valid_out(valid_out_237)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(data_out[7647:7616]),
	.valid_out(valid_out_238)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(data_out[7679:7648]),
	.valid_out(valid_out_239)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(data_out[7711:7680]),
	.valid_out(valid_out_240)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(data_out[7743:7712]),
	.valid_out(valid_out_241)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(data_out[7775:7744]),
	.valid_out(valid_out_242)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(data_out[7807:7776]),
	.valid_out(valid_out_243)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(data_out[7839:7808]),
	.valid_out(valid_out_244)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(data_out[7871:7840]),
	.valid_out(valid_out_245)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(data_out[7903:7872]),
	.valid_out(valid_out_246)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(data_out[7935:7904]),
	.valid_out(valid_out_247)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(data_out[7967:7936]),
	.valid_out(valid_out_248)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(data_out[7999:7968]),
	.valid_out(valid_out_249)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(data_out[8031:8000]),
	.valid_out(valid_out_250)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(data_out[8063:8032]),
	.valid_out(valid_out_251)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(data_out[8095:8064]),
	.valid_out(valid_out_252)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(data_out[8127:8096]),
	.valid_out(valid_out_253)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(data_out[8159:8128]),
	.valid_out(valid_out_254)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(data_out[8191:8160]),
	.valid_out(valid_out_255)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst256(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8223:8192]),
	.valid_in(valid_in),
	.data_out(data_out[8223:8192]),
	.valid_out(valid_out_256)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst257(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8255:8224]),
	.valid_in(valid_in),
	.data_out(data_out[8255:8224]),
	.valid_out(valid_out_257)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst258(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8287:8256]),
	.valid_in(valid_in),
	.data_out(data_out[8287:8256]),
	.valid_out(valid_out_258)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst259(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8319:8288]),
	.valid_in(valid_in),
	.data_out(data_out[8319:8288]),
	.valid_out(valid_out_259)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst260(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8351:8320]),
	.valid_in(valid_in),
	.data_out(data_out[8351:8320]),
	.valid_out(valid_out_260)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst261(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8383:8352]),
	.valid_in(valid_in),
	.data_out(data_out[8383:8352]),
	.valid_out(valid_out_261)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst262(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8415:8384]),
	.valid_in(valid_in),
	.data_out(data_out[8415:8384]),
	.valid_out(valid_out_262)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst263(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8447:8416]),
	.valid_in(valid_in),
	.data_out(data_out[8447:8416]),
	.valid_out(valid_out_263)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst264(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8479:8448]),
	.valid_in(valid_in),
	.data_out(data_out[8479:8448]),
	.valid_out(valid_out_264)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst265(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8511:8480]),
	.valid_in(valid_in),
	.data_out(data_out[8511:8480]),
	.valid_out(valid_out_265)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst266(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8543:8512]),
	.valid_in(valid_in),
	.data_out(data_out[8543:8512]),
	.valid_out(valid_out_266)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst267(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8575:8544]),
	.valid_in(valid_in),
	.data_out(data_out[8575:8544]),
	.valid_out(valid_out_267)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst268(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8607:8576]),
	.valid_in(valid_in),
	.data_out(data_out[8607:8576]),
	.valid_out(valid_out_268)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst269(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8639:8608]),
	.valid_in(valid_in),
	.data_out(data_out[8639:8608]),
	.valid_out(valid_out_269)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst270(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8671:8640]),
	.valid_in(valid_in),
	.data_out(data_out[8671:8640]),
	.valid_out(valid_out_270)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst271(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8703:8672]),
	.valid_in(valid_in),
	.data_out(data_out[8703:8672]),
	.valid_out(valid_out_271)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst272(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8735:8704]),
	.valid_in(valid_in),
	.data_out(data_out[8735:8704]),
	.valid_out(valid_out_272)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst273(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8767:8736]),
	.valid_in(valid_in),
	.data_out(data_out[8767:8736]),
	.valid_out(valid_out_273)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst274(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8799:8768]),
	.valid_in(valid_in),
	.data_out(data_out[8799:8768]),
	.valid_out(valid_out_274)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst275(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8831:8800]),
	.valid_in(valid_in),
	.data_out(data_out[8831:8800]),
	.valid_out(valid_out_275)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst276(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8863:8832]),
	.valid_in(valid_in),
	.data_out(data_out[8863:8832]),
	.valid_out(valid_out_276)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst277(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8895:8864]),
	.valid_in(valid_in),
	.data_out(data_out[8895:8864]),
	.valid_out(valid_out_277)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst278(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8927:8896]),
	.valid_in(valid_in),
	.data_out(data_out[8927:8896]),
	.valid_out(valid_out_278)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst279(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8959:8928]),
	.valid_in(valid_in),
	.data_out(data_out[8959:8928]),
	.valid_out(valid_out_279)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst280(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8991:8960]),
	.valid_in(valid_in),
	.data_out(data_out[8991:8960]),
	.valid_out(valid_out_280)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst281(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9023:8992]),
	.valid_in(valid_in),
	.data_out(data_out[9023:8992]),
	.valid_out(valid_out_281)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst282(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9055:9024]),
	.valid_in(valid_in),
	.data_out(data_out[9055:9024]),
	.valid_out(valid_out_282)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst283(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9087:9056]),
	.valid_in(valid_in),
	.data_out(data_out[9087:9056]),
	.valid_out(valid_out_283)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst284(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9119:9088]),
	.valid_in(valid_in),
	.data_out(data_out[9119:9088]),
	.valid_out(valid_out_284)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst285(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9151:9120]),
	.valid_in(valid_in),
	.data_out(data_out[9151:9120]),
	.valid_out(valid_out_285)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst286(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9183:9152]),
	.valid_in(valid_in),
	.data_out(data_out[9183:9152]),
	.valid_out(valid_out_286)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst287(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9215:9184]),
	.valid_in(valid_in),
	.data_out(data_out[9215:9184]),
	.valid_out(valid_out_287)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst288(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9247:9216]),
	.valid_in(valid_in),
	.data_out(data_out[9247:9216]),
	.valid_out(valid_out_288)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst289(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9279:9248]),
	.valid_in(valid_in),
	.data_out(data_out[9279:9248]),
	.valid_out(valid_out_289)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst290(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9311:9280]),
	.valid_in(valid_in),
	.data_out(data_out[9311:9280]),
	.valid_out(valid_out_290)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst291(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9343:9312]),
	.valid_in(valid_in),
	.data_out(data_out[9343:9312]),
	.valid_out(valid_out_291)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst292(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9375:9344]),
	.valid_in(valid_in),
	.data_out(data_out[9375:9344]),
	.valid_out(valid_out_292)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst293(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9407:9376]),
	.valid_in(valid_in),
	.data_out(data_out[9407:9376]),
	.valid_out(valid_out_293)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst294(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9439:9408]),
	.valid_in(valid_in),
	.data_out(data_out[9439:9408]),
	.valid_out(valid_out_294)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst295(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9471:9440]),
	.valid_in(valid_in),
	.data_out(data_out[9471:9440]),
	.valid_out(valid_out_295)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst296(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9503:9472]),
	.valid_in(valid_in),
	.data_out(data_out[9503:9472]),
	.valid_out(valid_out_296)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst297(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9535:9504]),
	.valid_in(valid_in),
	.data_out(data_out[9535:9504]),
	.valid_out(valid_out_297)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst298(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9567:9536]),
	.valid_in(valid_in),
	.data_out(data_out[9567:9536]),
	.valid_out(valid_out_298)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst299(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9599:9568]),
	.valid_in(valid_in),
	.data_out(data_out[9599:9568]),
	.valid_out(valid_out_299)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst300(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9631:9600]),
	.valid_in(valid_in),
	.data_out(data_out[9631:9600]),
	.valid_out(valid_out_300)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst301(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9663:9632]),
	.valid_in(valid_in),
	.data_out(data_out[9663:9632]),
	.valid_out(valid_out_301)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst302(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9695:9664]),
	.valid_in(valid_in),
	.data_out(data_out[9695:9664]),
	.valid_out(valid_out_302)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst303(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9727:9696]),
	.valid_in(valid_in),
	.data_out(data_out[9727:9696]),
	.valid_out(valid_out_303)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst304(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9759:9728]),
	.valid_in(valid_in),
	.data_out(data_out[9759:9728]),
	.valid_out(valid_out_304)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst305(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9791:9760]),
	.valid_in(valid_in),
	.data_out(data_out[9791:9760]),
	.valid_out(valid_out_305)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst306(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9823:9792]),
	.valid_in(valid_in),
	.data_out(data_out[9823:9792]),
	.valid_out(valid_out_306)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst307(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9855:9824]),
	.valid_in(valid_in),
	.data_out(data_out[9855:9824]),
	.valid_out(valid_out_307)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst308(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9887:9856]),
	.valid_in(valid_in),
	.data_out(data_out[9887:9856]),
	.valid_out(valid_out_308)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst309(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9919:9888]),
	.valid_in(valid_in),
	.data_out(data_out[9919:9888]),
	.valid_out(valid_out_309)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst310(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9951:9920]),
	.valid_in(valid_in),
	.data_out(data_out[9951:9920]),
	.valid_out(valid_out_310)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst311(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[9983:9952]),
	.valid_in(valid_in),
	.data_out(data_out[9983:9952]),
	.valid_out(valid_out_311)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst312(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10015:9984]),
	.valid_in(valid_in),
	.data_out(data_out[10015:9984]),
	.valid_out(valid_out_312)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst313(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10047:10016]),
	.valid_in(valid_in),
	.data_out(data_out[10047:10016]),
	.valid_out(valid_out_313)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst314(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10079:10048]),
	.valid_in(valid_in),
	.data_out(data_out[10079:10048]),
	.valid_out(valid_out_314)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst315(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10111:10080]),
	.valid_in(valid_in),
	.data_out(data_out[10111:10080]),
	.valid_out(valid_out_315)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst316(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10143:10112]),
	.valid_in(valid_in),
	.data_out(data_out[10143:10112]),
	.valid_out(valid_out_316)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst317(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10175:10144]),
	.valid_in(valid_in),
	.data_out(data_out[10175:10144]),
	.valid_out(valid_out_317)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst318(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10207:10176]),
	.valid_in(valid_in),
	.data_out(data_out[10207:10176]),
	.valid_out(valid_out_318)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst319(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10239:10208]),
	.valid_in(valid_in),
	.data_out(data_out[10239:10208]),
	.valid_out(valid_out_319)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst320(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10271:10240]),
	.valid_in(valid_in),
	.data_out(data_out[10271:10240]),
	.valid_out(valid_out_320)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst321(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10303:10272]),
	.valid_in(valid_in),
	.data_out(data_out[10303:10272]),
	.valid_out(valid_out_321)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst322(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10335:10304]),
	.valid_in(valid_in),
	.data_out(data_out[10335:10304]),
	.valid_out(valid_out_322)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst323(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10367:10336]),
	.valid_in(valid_in),
	.data_out(data_out[10367:10336]),
	.valid_out(valid_out_323)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst324(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10399:10368]),
	.valid_in(valid_in),
	.data_out(data_out[10399:10368]),
	.valid_out(valid_out_324)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst325(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10431:10400]),
	.valid_in(valid_in),
	.data_out(data_out[10431:10400]),
	.valid_out(valid_out_325)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst326(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10463:10432]),
	.valid_in(valid_in),
	.data_out(data_out[10463:10432]),
	.valid_out(valid_out_326)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst327(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10495:10464]),
	.valid_in(valid_in),
	.data_out(data_out[10495:10464]),
	.valid_out(valid_out_327)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst328(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10527:10496]),
	.valid_in(valid_in),
	.data_out(data_out[10527:10496]),
	.valid_out(valid_out_328)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst329(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10559:10528]),
	.valid_in(valid_in),
	.data_out(data_out[10559:10528]),
	.valid_out(valid_out_329)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst330(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10591:10560]),
	.valid_in(valid_in),
	.data_out(data_out[10591:10560]),
	.valid_out(valid_out_330)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst331(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10623:10592]),
	.valid_in(valid_in),
	.data_out(data_out[10623:10592]),
	.valid_out(valid_out_331)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst332(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10655:10624]),
	.valid_in(valid_in),
	.data_out(data_out[10655:10624]),
	.valid_out(valid_out_332)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst333(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10687:10656]),
	.valid_in(valid_in),
	.data_out(data_out[10687:10656]),
	.valid_out(valid_out_333)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst334(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10719:10688]),
	.valid_in(valid_in),
	.data_out(data_out[10719:10688]),
	.valid_out(valid_out_334)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst335(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10751:10720]),
	.valid_in(valid_in),
	.data_out(data_out[10751:10720]),
	.valid_out(valid_out_335)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst336(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10783:10752]),
	.valid_in(valid_in),
	.data_out(data_out[10783:10752]),
	.valid_out(valid_out_336)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst337(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10815:10784]),
	.valid_in(valid_in),
	.data_out(data_out[10815:10784]),
	.valid_out(valid_out_337)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst338(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10847:10816]),
	.valid_in(valid_in),
	.data_out(data_out[10847:10816]),
	.valid_out(valid_out_338)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst339(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10879:10848]),
	.valid_in(valid_in),
	.data_out(data_out[10879:10848]),
	.valid_out(valid_out_339)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst340(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10911:10880]),
	.valid_in(valid_in),
	.data_out(data_out[10911:10880]),
	.valid_out(valid_out_340)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst341(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10943:10912]),
	.valid_in(valid_in),
	.data_out(data_out[10943:10912]),
	.valid_out(valid_out_341)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst342(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[10975:10944]),
	.valid_in(valid_in),
	.data_out(data_out[10975:10944]),
	.valid_out(valid_out_342)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst343(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11007:10976]),
	.valid_in(valid_in),
	.data_out(data_out[11007:10976]),
	.valid_out(valid_out_343)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst344(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11039:11008]),
	.valid_in(valid_in),
	.data_out(data_out[11039:11008]),
	.valid_out(valid_out_344)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst345(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11071:11040]),
	.valid_in(valid_in),
	.data_out(data_out[11071:11040]),
	.valid_out(valid_out_345)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst346(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11103:11072]),
	.valid_in(valid_in),
	.data_out(data_out[11103:11072]),
	.valid_out(valid_out_346)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst347(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11135:11104]),
	.valid_in(valid_in),
	.data_out(data_out[11135:11104]),
	.valid_out(valid_out_347)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst348(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11167:11136]),
	.valid_in(valid_in),
	.data_out(data_out[11167:11136]),
	.valid_out(valid_out_348)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst349(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11199:11168]),
	.valid_in(valid_in),
	.data_out(data_out[11199:11168]),
	.valid_out(valid_out_349)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst350(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11231:11200]),
	.valid_in(valid_in),
	.data_out(data_out[11231:11200]),
	.valid_out(valid_out_350)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst351(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11263:11232]),
	.valid_in(valid_in),
	.data_out(data_out[11263:11232]),
	.valid_out(valid_out_351)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst352(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11295:11264]),
	.valid_in(valid_in),
	.data_out(data_out[11295:11264]),
	.valid_out(valid_out_352)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst353(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11327:11296]),
	.valid_in(valid_in),
	.data_out(data_out[11327:11296]),
	.valid_out(valid_out_353)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst354(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11359:11328]),
	.valid_in(valid_in),
	.data_out(data_out[11359:11328]),
	.valid_out(valid_out_354)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst355(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11391:11360]),
	.valid_in(valid_in),
	.data_out(data_out[11391:11360]),
	.valid_out(valid_out_355)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst356(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11423:11392]),
	.valid_in(valid_in),
	.data_out(data_out[11423:11392]),
	.valid_out(valid_out_356)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst357(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11455:11424]),
	.valid_in(valid_in),
	.data_out(data_out[11455:11424]),
	.valid_out(valid_out_357)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst358(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11487:11456]),
	.valid_in(valid_in),
	.data_out(data_out[11487:11456]),
	.valid_out(valid_out_358)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst359(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11519:11488]),
	.valid_in(valid_in),
	.data_out(data_out[11519:11488]),
	.valid_out(valid_out_359)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst360(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11551:11520]),
	.valid_in(valid_in),
	.data_out(data_out[11551:11520]),
	.valid_out(valid_out_360)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst361(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11583:11552]),
	.valid_in(valid_in),
	.data_out(data_out[11583:11552]),
	.valid_out(valid_out_361)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst362(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11615:11584]),
	.valid_in(valid_in),
	.data_out(data_out[11615:11584]),
	.valid_out(valid_out_362)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst363(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11647:11616]),
	.valid_in(valid_in),
	.data_out(data_out[11647:11616]),
	.valid_out(valid_out_363)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst364(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11679:11648]),
	.valid_in(valid_in),
	.data_out(data_out[11679:11648]),
	.valid_out(valid_out_364)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst365(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11711:11680]),
	.valid_in(valid_in),
	.data_out(data_out[11711:11680]),
	.valid_out(valid_out_365)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst366(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11743:11712]),
	.valid_in(valid_in),
	.data_out(data_out[11743:11712]),
	.valid_out(valid_out_366)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst367(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11775:11744]),
	.valid_in(valid_in),
	.data_out(data_out[11775:11744]),
	.valid_out(valid_out_367)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst368(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11807:11776]),
	.valid_in(valid_in),
	.data_out(data_out[11807:11776]),
	.valid_out(valid_out_368)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst369(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11839:11808]),
	.valid_in(valid_in),
	.data_out(data_out[11839:11808]),
	.valid_out(valid_out_369)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst370(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11871:11840]),
	.valid_in(valid_in),
	.data_out(data_out[11871:11840]),
	.valid_out(valid_out_370)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst371(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11903:11872]),
	.valid_in(valid_in),
	.data_out(data_out[11903:11872]),
	.valid_out(valid_out_371)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst372(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11935:11904]),
	.valid_in(valid_in),
	.data_out(data_out[11935:11904]),
	.valid_out(valid_out_372)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst373(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11967:11936]),
	.valid_in(valid_in),
	.data_out(data_out[11967:11936]),
	.valid_out(valid_out_373)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst374(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[11999:11968]),
	.valid_in(valid_in),
	.data_out(data_out[11999:11968]),
	.valid_out(valid_out_374)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst375(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12031:12000]),
	.valid_in(valid_in),
	.data_out(data_out[12031:12000]),
	.valid_out(valid_out_375)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst376(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12063:12032]),
	.valid_in(valid_in),
	.data_out(data_out[12063:12032]),
	.valid_out(valid_out_376)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst377(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12095:12064]),
	.valid_in(valid_in),
	.data_out(data_out[12095:12064]),
	.valid_out(valid_out_377)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst378(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12127:12096]),
	.valid_in(valid_in),
	.data_out(data_out[12127:12096]),
	.valid_out(valid_out_378)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst379(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12159:12128]),
	.valid_in(valid_in),
	.data_out(data_out[12159:12128]),
	.valid_out(valid_out_379)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst380(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12191:12160]),
	.valid_in(valid_in),
	.data_out(data_out[12191:12160]),
	.valid_out(valid_out_380)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst381(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12223:12192]),
	.valid_in(valid_in),
	.data_out(data_out[12223:12192]),
	.valid_out(valid_out_381)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst382(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12255:12224]),
	.valid_in(valid_in),
	.data_out(data_out[12255:12224]),
	.valid_out(valid_out_382)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst383(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12287:12256]),
	.valid_in(valid_in),
	.data_out(data_out[12287:12256]),
	.valid_out(valid_out_383)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst384(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12319:12288]),
	.valid_in(valid_in),
	.data_out(data_out[12319:12288]),
	.valid_out(valid_out_384)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst385(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12351:12320]),
	.valid_in(valid_in),
	.data_out(data_out[12351:12320]),
	.valid_out(valid_out_385)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst386(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12383:12352]),
	.valid_in(valid_in),
	.data_out(data_out[12383:12352]),
	.valid_out(valid_out_386)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst387(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12415:12384]),
	.valid_in(valid_in),
	.data_out(data_out[12415:12384]),
	.valid_out(valid_out_387)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst388(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12447:12416]),
	.valid_in(valid_in),
	.data_out(data_out[12447:12416]),
	.valid_out(valid_out_388)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst389(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12479:12448]),
	.valid_in(valid_in),
	.data_out(data_out[12479:12448]),
	.valid_out(valid_out_389)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst390(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12511:12480]),
	.valid_in(valid_in),
	.data_out(data_out[12511:12480]),
	.valid_out(valid_out_390)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst391(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12543:12512]),
	.valid_in(valid_in),
	.data_out(data_out[12543:12512]),
	.valid_out(valid_out_391)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst392(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12575:12544]),
	.valid_in(valid_in),
	.data_out(data_out[12575:12544]),
	.valid_out(valid_out_392)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst393(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12607:12576]),
	.valid_in(valid_in),
	.data_out(data_out[12607:12576]),
	.valid_out(valid_out_393)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst394(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12639:12608]),
	.valid_in(valid_in),
	.data_out(data_out[12639:12608]),
	.valid_out(valid_out_394)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst395(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12671:12640]),
	.valid_in(valid_in),
	.data_out(data_out[12671:12640]),
	.valid_out(valid_out_395)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst396(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12703:12672]),
	.valid_in(valid_in),
	.data_out(data_out[12703:12672]),
	.valid_out(valid_out_396)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst397(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12735:12704]),
	.valid_in(valid_in),
	.data_out(data_out[12735:12704]),
	.valid_out(valid_out_397)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst398(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12767:12736]),
	.valid_in(valid_in),
	.data_out(data_out[12767:12736]),
	.valid_out(valid_out_398)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst399(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12799:12768]),
	.valid_in(valid_in),
	.data_out(data_out[12799:12768]),
	.valid_out(valid_out_399)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst400(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12831:12800]),
	.valid_in(valid_in),
	.data_out(data_out[12831:12800]),
	.valid_out(valid_out_400)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst401(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12863:12832]),
	.valid_in(valid_in),
	.data_out(data_out[12863:12832]),
	.valid_out(valid_out_401)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst402(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12895:12864]),
	.valid_in(valid_in),
	.data_out(data_out[12895:12864]),
	.valid_out(valid_out_402)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst403(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12927:12896]),
	.valid_in(valid_in),
	.data_out(data_out[12927:12896]),
	.valid_out(valid_out_403)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst404(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12959:12928]),
	.valid_in(valid_in),
	.data_out(data_out[12959:12928]),
	.valid_out(valid_out_404)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst405(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[12991:12960]),
	.valid_in(valid_in),
	.data_out(data_out[12991:12960]),
	.valid_out(valid_out_405)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst406(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13023:12992]),
	.valid_in(valid_in),
	.data_out(data_out[13023:12992]),
	.valid_out(valid_out_406)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst407(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13055:13024]),
	.valid_in(valid_in),
	.data_out(data_out[13055:13024]),
	.valid_out(valid_out_407)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst408(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13087:13056]),
	.valid_in(valid_in),
	.data_out(data_out[13087:13056]),
	.valid_out(valid_out_408)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst409(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13119:13088]),
	.valid_in(valid_in),
	.data_out(data_out[13119:13088]),
	.valid_out(valid_out_409)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst410(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13151:13120]),
	.valid_in(valid_in),
	.data_out(data_out[13151:13120]),
	.valid_out(valid_out_410)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst411(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13183:13152]),
	.valid_in(valid_in),
	.data_out(data_out[13183:13152]),
	.valid_out(valid_out_411)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst412(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13215:13184]),
	.valid_in(valid_in),
	.data_out(data_out[13215:13184]),
	.valid_out(valid_out_412)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst413(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13247:13216]),
	.valid_in(valid_in),
	.data_out(data_out[13247:13216]),
	.valid_out(valid_out_413)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst414(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13279:13248]),
	.valid_in(valid_in),
	.data_out(data_out[13279:13248]),
	.valid_out(valid_out_414)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst415(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13311:13280]),
	.valid_in(valid_in),
	.data_out(data_out[13311:13280]),
	.valid_out(valid_out_415)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst416(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13343:13312]),
	.valid_in(valid_in),
	.data_out(data_out[13343:13312]),
	.valid_out(valid_out_416)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst417(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13375:13344]),
	.valid_in(valid_in),
	.data_out(data_out[13375:13344]),
	.valid_out(valid_out_417)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst418(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13407:13376]),
	.valid_in(valid_in),
	.data_out(data_out[13407:13376]),
	.valid_out(valid_out_418)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst419(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13439:13408]),
	.valid_in(valid_in),
	.data_out(data_out[13439:13408]),
	.valid_out(valid_out_419)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst420(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13471:13440]),
	.valid_in(valid_in),
	.data_out(data_out[13471:13440]),
	.valid_out(valid_out_420)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst421(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13503:13472]),
	.valid_in(valid_in),
	.data_out(data_out[13503:13472]),
	.valid_out(valid_out_421)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst422(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13535:13504]),
	.valid_in(valid_in),
	.data_out(data_out[13535:13504]),
	.valid_out(valid_out_422)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst423(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13567:13536]),
	.valid_in(valid_in),
	.data_out(data_out[13567:13536]),
	.valid_out(valid_out_423)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst424(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13599:13568]),
	.valid_in(valid_in),
	.data_out(data_out[13599:13568]),
	.valid_out(valid_out_424)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst425(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13631:13600]),
	.valid_in(valid_in),
	.data_out(data_out[13631:13600]),
	.valid_out(valid_out_425)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst426(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13663:13632]),
	.valid_in(valid_in),
	.data_out(data_out[13663:13632]),
	.valid_out(valid_out_426)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst427(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13695:13664]),
	.valid_in(valid_in),
	.data_out(data_out[13695:13664]),
	.valid_out(valid_out_427)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst428(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13727:13696]),
	.valid_in(valid_in),
	.data_out(data_out[13727:13696]),
	.valid_out(valid_out_428)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst429(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13759:13728]),
	.valid_in(valid_in),
	.data_out(data_out[13759:13728]),
	.valid_out(valid_out_429)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst430(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13791:13760]),
	.valid_in(valid_in),
	.data_out(data_out[13791:13760]),
	.valid_out(valid_out_430)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst431(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13823:13792]),
	.valid_in(valid_in),
	.data_out(data_out[13823:13792]),
	.valid_out(valid_out_431)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst432(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13855:13824]),
	.valid_in(valid_in),
	.data_out(data_out[13855:13824]),
	.valid_out(valid_out_432)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst433(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13887:13856]),
	.valid_in(valid_in),
	.data_out(data_out[13887:13856]),
	.valid_out(valid_out_433)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst434(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13919:13888]),
	.valid_in(valid_in),
	.data_out(data_out[13919:13888]),
	.valid_out(valid_out_434)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst435(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13951:13920]),
	.valid_in(valid_in),
	.data_out(data_out[13951:13920]),
	.valid_out(valid_out_435)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst436(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[13983:13952]),
	.valid_in(valid_in),
	.data_out(data_out[13983:13952]),
	.valid_out(valid_out_436)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst437(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14015:13984]),
	.valid_in(valid_in),
	.data_out(data_out[14015:13984]),
	.valid_out(valid_out_437)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst438(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14047:14016]),
	.valid_in(valid_in),
	.data_out(data_out[14047:14016]),
	.valid_out(valid_out_438)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst439(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14079:14048]),
	.valid_in(valid_in),
	.data_out(data_out[14079:14048]),
	.valid_out(valid_out_439)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst440(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14111:14080]),
	.valid_in(valid_in),
	.data_out(data_out[14111:14080]),
	.valid_out(valid_out_440)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst441(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14143:14112]),
	.valid_in(valid_in),
	.data_out(data_out[14143:14112]),
	.valid_out(valid_out_441)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst442(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14175:14144]),
	.valid_in(valid_in),
	.data_out(data_out[14175:14144]),
	.valid_out(valid_out_442)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst443(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14207:14176]),
	.valid_in(valid_in),
	.data_out(data_out[14207:14176]),
	.valid_out(valid_out_443)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst444(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14239:14208]),
	.valid_in(valid_in),
	.data_out(data_out[14239:14208]),
	.valid_out(valid_out_444)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst445(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14271:14240]),
	.valid_in(valid_in),
	.data_out(data_out[14271:14240]),
	.valid_out(valid_out_445)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst446(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14303:14272]),
	.valid_in(valid_in),
	.data_out(data_out[14303:14272]),
	.valid_out(valid_out_446)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst447(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14335:14304]),
	.valid_in(valid_in),
	.data_out(data_out[14335:14304]),
	.valid_out(valid_out_447)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst448(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14367:14336]),
	.valid_in(valid_in),
	.data_out(data_out[14367:14336]),
	.valid_out(valid_out_448)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst449(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14399:14368]),
	.valid_in(valid_in),
	.data_out(data_out[14399:14368]),
	.valid_out(valid_out_449)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst450(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14431:14400]),
	.valid_in(valid_in),
	.data_out(data_out[14431:14400]),
	.valid_out(valid_out_450)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst451(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14463:14432]),
	.valid_in(valid_in),
	.data_out(data_out[14463:14432]),
	.valid_out(valid_out_451)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst452(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14495:14464]),
	.valid_in(valid_in),
	.data_out(data_out[14495:14464]),
	.valid_out(valid_out_452)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst453(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14527:14496]),
	.valid_in(valid_in),
	.data_out(data_out[14527:14496]),
	.valid_out(valid_out_453)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst454(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14559:14528]),
	.valid_in(valid_in),
	.data_out(data_out[14559:14528]),
	.valid_out(valid_out_454)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst455(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14591:14560]),
	.valid_in(valid_in),
	.data_out(data_out[14591:14560]),
	.valid_out(valid_out_455)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst456(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14623:14592]),
	.valid_in(valid_in),
	.data_out(data_out[14623:14592]),
	.valid_out(valid_out_456)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst457(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14655:14624]),
	.valid_in(valid_in),
	.data_out(data_out[14655:14624]),
	.valid_out(valid_out_457)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst458(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14687:14656]),
	.valid_in(valid_in),
	.data_out(data_out[14687:14656]),
	.valid_out(valid_out_458)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst459(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14719:14688]),
	.valid_in(valid_in),
	.data_out(data_out[14719:14688]),
	.valid_out(valid_out_459)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst460(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14751:14720]),
	.valid_in(valid_in),
	.data_out(data_out[14751:14720]),
	.valid_out(valid_out_460)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst461(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14783:14752]),
	.valid_in(valid_in),
	.data_out(data_out[14783:14752]),
	.valid_out(valid_out_461)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst462(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14815:14784]),
	.valid_in(valid_in),
	.data_out(data_out[14815:14784]),
	.valid_out(valid_out_462)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst463(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14847:14816]),
	.valid_in(valid_in),
	.data_out(data_out[14847:14816]),
	.valid_out(valid_out_463)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst464(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14879:14848]),
	.valid_in(valid_in),
	.data_out(data_out[14879:14848]),
	.valid_out(valid_out_464)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst465(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14911:14880]),
	.valid_in(valid_in),
	.data_out(data_out[14911:14880]),
	.valid_out(valid_out_465)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst466(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14943:14912]),
	.valid_in(valid_in),
	.data_out(data_out[14943:14912]),
	.valid_out(valid_out_466)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst467(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[14975:14944]),
	.valid_in(valid_in),
	.data_out(data_out[14975:14944]),
	.valid_out(valid_out_467)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst468(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15007:14976]),
	.valid_in(valid_in),
	.data_out(data_out[15007:14976]),
	.valid_out(valid_out_468)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst469(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15039:15008]),
	.valid_in(valid_in),
	.data_out(data_out[15039:15008]),
	.valid_out(valid_out_469)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst470(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15071:15040]),
	.valid_in(valid_in),
	.data_out(data_out[15071:15040]),
	.valid_out(valid_out_470)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst471(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15103:15072]),
	.valid_in(valid_in),
	.data_out(data_out[15103:15072]),
	.valid_out(valid_out_471)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst472(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15135:15104]),
	.valid_in(valid_in),
	.data_out(data_out[15135:15104]),
	.valid_out(valid_out_472)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst473(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15167:15136]),
	.valid_in(valid_in),
	.data_out(data_out[15167:15136]),
	.valid_out(valid_out_473)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst474(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15199:15168]),
	.valid_in(valid_in),
	.data_out(data_out[15199:15168]),
	.valid_out(valid_out_474)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst475(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15231:15200]),
	.valid_in(valid_in),
	.data_out(data_out[15231:15200]),
	.valid_out(valid_out_475)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst476(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15263:15232]),
	.valid_in(valid_in),
	.data_out(data_out[15263:15232]),
	.valid_out(valid_out_476)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst477(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15295:15264]),
	.valid_in(valid_in),
	.data_out(data_out[15295:15264]),
	.valid_out(valid_out_477)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst478(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15327:15296]),
	.valid_in(valid_in),
	.data_out(data_out[15327:15296]),
	.valid_out(valid_out_478)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst479(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15359:15328]),
	.valid_in(valid_in),
	.data_out(data_out[15359:15328]),
	.valid_out(valid_out_479)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst480(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15391:15360]),
	.valid_in(valid_in),
	.data_out(data_out[15391:15360]),
	.valid_out(valid_out_480)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst481(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15423:15392]),
	.valid_in(valid_in),
	.data_out(data_out[15423:15392]),
	.valid_out(valid_out_481)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst482(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15455:15424]),
	.valid_in(valid_in),
	.data_out(data_out[15455:15424]),
	.valid_out(valid_out_482)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst483(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15487:15456]),
	.valid_in(valid_in),
	.data_out(data_out[15487:15456]),
	.valid_out(valid_out_483)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst484(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15519:15488]),
	.valid_in(valid_in),
	.data_out(data_out[15519:15488]),
	.valid_out(valid_out_484)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst485(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15551:15520]),
	.valid_in(valid_in),
	.data_out(data_out[15551:15520]),
	.valid_out(valid_out_485)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst486(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15583:15552]),
	.valid_in(valid_in),
	.data_out(data_out[15583:15552]),
	.valid_out(valid_out_486)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst487(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15615:15584]),
	.valid_in(valid_in),
	.data_out(data_out[15615:15584]),
	.valid_out(valid_out_487)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst488(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15647:15616]),
	.valid_in(valid_in),
	.data_out(data_out[15647:15616]),
	.valid_out(valid_out_488)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst489(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15679:15648]),
	.valid_in(valid_in),
	.data_out(data_out[15679:15648]),
	.valid_out(valid_out_489)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst490(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15711:15680]),
	.valid_in(valid_in),
	.data_out(data_out[15711:15680]),
	.valid_out(valid_out_490)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst491(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15743:15712]),
	.valid_in(valid_in),
	.data_out(data_out[15743:15712]),
	.valid_out(valid_out_491)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst492(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15775:15744]),
	.valid_in(valid_in),
	.data_out(data_out[15775:15744]),
	.valid_out(valid_out_492)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst493(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15807:15776]),
	.valid_in(valid_in),
	.data_out(data_out[15807:15776]),
	.valid_out(valid_out_493)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst494(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15839:15808]),
	.valid_in(valid_in),
	.data_out(data_out[15839:15808]),
	.valid_out(valid_out_494)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst495(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15871:15840]),
	.valid_in(valid_in),
	.data_out(data_out[15871:15840]),
	.valid_out(valid_out_495)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst496(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15903:15872]),
	.valid_in(valid_in),
	.data_out(data_out[15903:15872]),
	.valid_out(valid_out_496)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst497(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15935:15904]),
	.valid_in(valid_in),
	.data_out(data_out[15935:15904]),
	.valid_out(valid_out_497)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst498(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15967:15936]),
	.valid_in(valid_in),
	.data_out(data_out[15967:15936]),
	.valid_out(valid_out_498)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst499(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15999:15968]),
	.valid_in(valid_in),
	.data_out(data_out[15999:15968]),
	.valid_out(valid_out_499)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst500(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16031:16000]),
	.valid_in(valid_in),
	.data_out(data_out[16031:16000]),
	.valid_out(valid_out_500)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst501(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16063:16032]),
	.valid_in(valid_in),
	.data_out(data_out[16063:16032]),
	.valid_out(valid_out_501)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst502(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16095:16064]),
	.valid_in(valid_in),
	.data_out(data_out[16095:16064]),
	.valid_out(valid_out_502)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst503(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16127:16096]),
	.valid_in(valid_in),
	.data_out(data_out[16127:16096]),
	.valid_out(valid_out_503)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst504(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16159:16128]),
	.valid_in(valid_in),
	.data_out(data_out[16159:16128]),
	.valid_out(valid_out_504)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst505(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16191:16160]),
	.valid_in(valid_in),
	.data_out(data_out[16191:16160]),
	.valid_out(valid_out_505)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst506(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16223:16192]),
	.valid_in(valid_in),
	.data_out(data_out[16223:16192]),
	.valid_out(valid_out_506)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst507(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16255:16224]),
	.valid_in(valid_in),
	.data_out(data_out[16255:16224]),
	.valid_out(valid_out_507)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst508(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16287:16256]),
	.valid_in(valid_in),
	.data_out(data_out[16287:16256]),
	.valid_out(valid_out_508)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst509(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16319:16288]),
	.valid_in(valid_in),
	.data_out(data_out[16319:16288]),
	.valid_out(valid_out_509)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst510(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16351:16320]),
	.valid_in(valid_in),
	.data_out(data_out[16351:16320]),
	.valid_out(valid_out_510)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst511(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[16383:16352]),
	.valid_in(valid_in),
	.data_out(data_out[16383:16352]),
	.valid_out(valid_out_511)
);

	assign valid_out = valid_out_0 & valid_out_1 & valid_out_2 & valid_out_3 & valid_out_4 & valid_out_5 & valid_out_6 & valid_out_7 & valid_out_8 & valid_out_9 & valid_out_10 & valid_out_11 & valid_out_12 & valid_out_13 & valid_out_14 & valid_out_15 & valid_out_16 & valid_out_17 & valid_out_18 & valid_out_19 & valid_out_20 & valid_out_21 & valid_out_22 & valid_out_23 & valid_out_24 & valid_out_25 & valid_out_26 & valid_out_27 & valid_out_28 & valid_out_29 & valid_out_30 & valid_out_31 & valid_out_32 & valid_out_33 & valid_out_34 & valid_out_35 & valid_out_36 & valid_out_37 & valid_out_38 & valid_out_39 & valid_out_40 & valid_out_41 & valid_out_42 & valid_out_43 & valid_out_44 & valid_out_45 & valid_out_46 & valid_out_47 & valid_out_48 & valid_out_49 & valid_out_50 & valid_out_51 & valid_out_52 & valid_out_53 & valid_out_54 & valid_out_55 & valid_out_56 & valid_out_57 & valid_out_58 & valid_out_59 & valid_out_60 & valid_out_61 & valid_out_62 & valid_out_63 & valid_out_64 & valid_out_65 & valid_out_66 & valid_out_67 & valid_out_68 & valid_out_69 & valid_out_70 & valid_out_71 & valid_out_72 & valid_out_73 & valid_out_74 & valid_out_75 & valid_out_76 & valid_out_77 & valid_out_78 & valid_out_79 & valid_out_80 & valid_out_81 & valid_out_82 & valid_out_83 & valid_out_84 & valid_out_85 & valid_out_86 & valid_out_87 & valid_out_88 & valid_out_89 & valid_out_90 & valid_out_91 & valid_out_92 & valid_out_93 & valid_out_94 & valid_out_95 & valid_out_96 & valid_out_97 & valid_out_98 & valid_out_99 & valid_out_100 & valid_out_101 & valid_out_102 & valid_out_103 & valid_out_104 & valid_out_105 & valid_out_106 & valid_out_107 & valid_out_108 & valid_out_109 & valid_out_110 & valid_out_111 & valid_out_112 & valid_out_113 & valid_out_114 & valid_out_115 & valid_out_116 & valid_out_117 & valid_out_118 & valid_out_119 & valid_out_120 & valid_out_121 & valid_out_122 & valid_out_123 & valid_out_124 & valid_out_125 & valid_out_126 & valid_out_127 & valid_out_128 & valid_out_129 & valid_out_130 & valid_out_131 & valid_out_132 & valid_out_133 & valid_out_134 & valid_out_135 & valid_out_136 & valid_out_137 & valid_out_138 & valid_out_139 & valid_out_140 & valid_out_141 & valid_out_142 & valid_out_143 & valid_out_144 & valid_out_145 & valid_out_146 & valid_out_147 & valid_out_148 & valid_out_149 & valid_out_150 & valid_out_151 & valid_out_152 & valid_out_153 & valid_out_154 & valid_out_155 & valid_out_156 & valid_out_157 & valid_out_158 & valid_out_159 & valid_out_160 & valid_out_161 & valid_out_162 & valid_out_163 & valid_out_164 & valid_out_165 & valid_out_166 & valid_out_167 & valid_out_168 & valid_out_169 & valid_out_170 & valid_out_171 & valid_out_172 & valid_out_173 & valid_out_174 & valid_out_175 & valid_out_176 & valid_out_177 & valid_out_178 & valid_out_179 & valid_out_180 & valid_out_181 & valid_out_182 & valid_out_183 & valid_out_184 & valid_out_185 & valid_out_186 & valid_out_187 & valid_out_188 & valid_out_189 & valid_out_190 & valid_out_191 & valid_out_192 & valid_out_193 & valid_out_194 & valid_out_195 & valid_out_196 & valid_out_197 & valid_out_198 & valid_out_199 & valid_out_200 & valid_out_201 & valid_out_202 & valid_out_203 & valid_out_204 & valid_out_205 & valid_out_206 & valid_out_207 & valid_out_208 & valid_out_209 & valid_out_210 & valid_out_211 & valid_out_212 & valid_out_213 & valid_out_214 & valid_out_215 & valid_out_216 & valid_out_217 & valid_out_218 & valid_out_219 & valid_out_220 & valid_out_221 & valid_out_222 & valid_out_223 & valid_out_224 & valid_out_225 & valid_out_226 & valid_out_227 & valid_out_228 & valid_out_229 & valid_out_230 & valid_out_231 & valid_out_232 & valid_out_233 & valid_out_234 & valid_out_235 & valid_out_236 & valid_out_237 & valid_out_238 & valid_out_239 & valid_out_240 & valid_out_241 & valid_out_242 & valid_out_243 & valid_out_244 & valid_out_245 & valid_out_246 & valid_out_247 & valid_out_248 & valid_out_249 & valid_out_250 & valid_out_251 & valid_out_252 & valid_out_253 & valid_out_254 & valid_out_255 & valid_out_256 & valid_out_257 & valid_out_258 & valid_out_259 & valid_out_260 & valid_out_261 & valid_out_262 & valid_out_263 & valid_out_264 & valid_out_265 & valid_out_266 & valid_out_267 & valid_out_268 & valid_out_269 & valid_out_270 & valid_out_271 & valid_out_272 & valid_out_273 & valid_out_274 & valid_out_275 & valid_out_276 & valid_out_277 & valid_out_278 & valid_out_279 & valid_out_280 & valid_out_281 & valid_out_282 & valid_out_283 & valid_out_284 & valid_out_285 & valid_out_286 & valid_out_287 & valid_out_288 & valid_out_289 & valid_out_290 & valid_out_291 & valid_out_292 & valid_out_293 & valid_out_294 & valid_out_295 & valid_out_296 & valid_out_297 & valid_out_298 & valid_out_299 & valid_out_300 & valid_out_301 & valid_out_302 & valid_out_303 & valid_out_304 & valid_out_305 & valid_out_306 & valid_out_307 & valid_out_308 & valid_out_309 & valid_out_310 & valid_out_311 & valid_out_312 & valid_out_313 & valid_out_314 & valid_out_315 & valid_out_316 & valid_out_317 & valid_out_318 & valid_out_319 & valid_out_320 & valid_out_321 & valid_out_322 & valid_out_323 & valid_out_324 & valid_out_325 & valid_out_326 & valid_out_327 & valid_out_328 & valid_out_329 & valid_out_330 & valid_out_331 & valid_out_332 & valid_out_333 & valid_out_334 & valid_out_335 & valid_out_336 & valid_out_337 & valid_out_338 & valid_out_339 & valid_out_340 & valid_out_341 & valid_out_342 & valid_out_343 & valid_out_344 & valid_out_345 & valid_out_346 & valid_out_347 & valid_out_348 & valid_out_349 & valid_out_350 & valid_out_351 & valid_out_352 & valid_out_353 & valid_out_354 & valid_out_355 & valid_out_356 & valid_out_357 & valid_out_358 & valid_out_359 & valid_out_360 & valid_out_361 & valid_out_362 & valid_out_363 & valid_out_364 & valid_out_365 & valid_out_366 & valid_out_367 & valid_out_368 & valid_out_369 & valid_out_370 & valid_out_371 & valid_out_372 & valid_out_373 & valid_out_374 & valid_out_375 & valid_out_376 & valid_out_377 & valid_out_378 & valid_out_379 & valid_out_380 & valid_out_381 & valid_out_382 & valid_out_383 & valid_out_384 & valid_out_385 & valid_out_386 & valid_out_387 & valid_out_388 & valid_out_389 & valid_out_390 & valid_out_391 & valid_out_392 & valid_out_393 & valid_out_394 & valid_out_395 & valid_out_396 & valid_out_397 & valid_out_398 & valid_out_399 & valid_out_400 & valid_out_401 & valid_out_402 & valid_out_403 & valid_out_404 & valid_out_405 & valid_out_406 & valid_out_407 & valid_out_408 & valid_out_409 & valid_out_410 & valid_out_411 & valid_out_412 & valid_out_413 & valid_out_414 & valid_out_415 & valid_out_416 & valid_out_417 & valid_out_418 & valid_out_419 & valid_out_420 & valid_out_421 & valid_out_422 & valid_out_423 & valid_out_424 & valid_out_425 & valid_out_426 & valid_out_427 & valid_out_428 & valid_out_429 & valid_out_430 & valid_out_431 & valid_out_432 & valid_out_433 & valid_out_434 & valid_out_435 & valid_out_436 & valid_out_437 & valid_out_438 & valid_out_439 & valid_out_440 & valid_out_441 & valid_out_442 & valid_out_443 & valid_out_444 & valid_out_445 & valid_out_446 & valid_out_447 & valid_out_448 & valid_out_449 & valid_out_450 & valid_out_451 & valid_out_452 & valid_out_453 & valid_out_454 & valid_out_455 & valid_out_456 & valid_out_457 & valid_out_458 & valid_out_459 & valid_out_460 & valid_out_461 & valid_out_462 & valid_out_463 & valid_out_464 & valid_out_465 & valid_out_466 & valid_out_467 & valid_out_468 & valid_out_469 & valid_out_470 & valid_out_471 & valid_out_472 & valid_out_473 & valid_out_474 & valid_out_475 & valid_out_476 & valid_out_477 & valid_out_478 & valid_out_479 & valid_out_480 & valid_out_481 & valid_out_482 & valid_out_483 & valid_out_484 & valid_out_485 & valid_out_486 & valid_out_487 & valid_out_488 & valid_out_489 & valid_out_490 & valid_out_491 & valid_out_492 & valid_out_493 & valid_out_494 & valid_out_495 & valid_out_496 & valid_out_497 & valid_out_498 & valid_out_499 & valid_out_500 & valid_out_501 & valid_out_502 & valid_out_503 & valid_out_504 & valid_out_505 & valid_out_506 & valid_out_507 & valid_out_508 & valid_out_509 & valid_out_510 & valid_out_511;
endmodule