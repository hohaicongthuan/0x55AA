module layer_10_featuremap_130(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdcbb5),
	.w1(32'h3c590182),
	.w2(32'hbc9e1f2e),
	.w3(32'hba080417),
	.w4(32'h3a768b73),
	.w5(32'hb9989f54),
	.w6(32'h3afd3ea5),
	.w7(32'hbc106dcd),
	.w8(32'hba4c1d1e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac99a39),
	.w1(32'h3c2a320f),
	.w2(32'hbb40ef0b),
	.w3(32'hbb8084aa),
	.w4(32'h3ba4f015),
	.w5(32'h39f6189c),
	.w6(32'h3b9d8101),
	.w7(32'hba04dee0),
	.w8(32'hbbbb776f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc586cdc),
	.w1(32'hba7c4b66),
	.w2(32'hbb62a556),
	.w3(32'hbb76aada),
	.w4(32'hb8e28c39),
	.w5(32'hbb563270),
	.w6(32'hb6b1a048),
	.w7(32'hbbd16ea0),
	.w8(32'hbba05475),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba233470),
	.w1(32'h3b97aa03),
	.w2(32'hbc4f24b8),
	.w3(32'hbb302014),
	.w4(32'h3be00c53),
	.w5(32'hbbdbc319),
	.w6(32'hb71fe0dc),
	.w7(32'h38364b56),
	.w8(32'hba87dc1e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1921),
	.w1(32'hbb3f8817),
	.w2(32'h3cbe7d8d),
	.w3(32'hbb8b08dd),
	.w4(32'hbb503aa0),
	.w5(32'hbbcefd19),
	.w6(32'hb9b072b1),
	.w7(32'hbafbf8b1),
	.w8(32'hbc005950),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0202cd),
	.w1(32'h3bc1db91),
	.w2(32'h3a94035e),
	.w3(32'hbb1f117e),
	.w4(32'h3bc810c8),
	.w5(32'hba8265af),
	.w6(32'h3bd15bd4),
	.w7(32'h3a303041),
	.w8(32'hbb9fa8a0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d1ceb),
	.w1(32'hbacf81d2),
	.w2(32'h3ba5633e),
	.w3(32'hbbdd1773),
	.w4(32'hbb220eae),
	.w5(32'hbad16370),
	.w6(32'hbb0bcafc),
	.w7(32'hbb4bf0e4),
	.w8(32'hbad192f1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff24cf),
	.w1(32'hbbc6f37b),
	.w2(32'h3ac07594),
	.w3(32'hbab23537),
	.w4(32'hba8f6d0f),
	.w5(32'hbb6189a9),
	.w6(32'hbb306827),
	.w7(32'hba85b5d3),
	.w8(32'h3aedb1d9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5cf16),
	.w1(32'hbb73d60c),
	.w2(32'hbb26dfe5),
	.w3(32'h39ee88de),
	.w4(32'hba6fc6a2),
	.w5(32'h3ac90858),
	.w6(32'hbb9a1839),
	.w7(32'h3a1560ab),
	.w8(32'h3954ed97),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81ef69),
	.w1(32'h3c08846c),
	.w2(32'h39eb2567),
	.w3(32'h3a39bbac),
	.w4(32'h3b89ffdc),
	.w5(32'hbb0a956e),
	.w6(32'h3af3d3c1),
	.w7(32'hbb3d4020),
	.w8(32'h3a7f8540),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19574),
	.w1(32'h3b46fba7),
	.w2(32'h3a909591),
	.w3(32'h3984eb66),
	.w4(32'h3bb4597b),
	.w5(32'hba9d76c9),
	.w6(32'h3b895414),
	.w7(32'hbb472909),
	.w8(32'hbc2815f2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3394),
	.w1(32'hbc93181d),
	.w2(32'hbbc93b2a),
	.w3(32'hbbb9973e),
	.w4(32'hbc0101da),
	.w5(32'hbbd8116b),
	.w6(32'hbc6f8657),
	.w7(32'hbbcd49c1),
	.w8(32'hbc1e1fc1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcfe3),
	.w1(32'hbaa94828),
	.w2(32'hbaa80e39),
	.w3(32'hbb429896),
	.w4(32'hbb2ec3f5),
	.w5(32'hbb379f0d),
	.w6(32'hbacec564),
	.w7(32'hbb64a798),
	.w8(32'hba944761),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab945d3),
	.w1(32'hbcdc1955),
	.w2(32'hbb9a9f58),
	.w3(32'hba726cfe),
	.w4(32'hbc905711),
	.w5(32'hbc3c2598),
	.w6(32'hbc95bf5e),
	.w7(32'hbc2e89c8),
	.w8(32'h3b8c649e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d179ea0),
	.w1(32'hbc84ced9),
	.w2(32'h3b818bc9),
	.w3(32'h3ad164a2),
	.w4(32'hba60a987),
	.w5(32'hbc0569f8),
	.w6(32'hbc1da39b),
	.w7(32'h3bc4ad59),
	.w8(32'hbc2cc5ea),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e1730),
	.w1(32'hbb3b069c),
	.w2(32'hbb3358c0),
	.w3(32'hbafefc10),
	.w4(32'hbb04ea0f),
	.w5(32'h3aa83f4f),
	.w6(32'hbb7c5558),
	.w7(32'h3b330d62),
	.w8(32'hbb157e91),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b7b7),
	.w1(32'h3bbbe884),
	.w2(32'hbc181d2b),
	.w3(32'h38efa7f2),
	.w4(32'hbbc9e9fc),
	.w5(32'hbb828de2),
	.w6(32'h3b81b122),
	.w7(32'hbb8e3811),
	.w8(32'h3a8b2c28),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5c2cd),
	.w1(32'h3c164312),
	.w2(32'hbb1006ed),
	.w3(32'h3929dd1f),
	.w4(32'h3b728468),
	.w5(32'hbaca18e3),
	.w6(32'h3b343f5e),
	.w7(32'h3af7d012),
	.w8(32'h3981206d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1e06),
	.w1(32'hbb761d5e),
	.w2(32'hbb995d1d),
	.w3(32'h3add2a19),
	.w4(32'hbade57ec),
	.w5(32'hbb9be014),
	.w6(32'hbb7277f8),
	.w7(32'hbb360794),
	.w8(32'hbac952b4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390e1f),
	.w1(32'hbba15ffe),
	.w2(32'hbb299181),
	.w3(32'hbae0a3da),
	.w4(32'hba598e3c),
	.w5(32'h39d1e89e),
	.w6(32'hbb856afd),
	.w7(32'h38e964a7),
	.w8(32'h3865d9a9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a3b2),
	.w1(32'hbb6a44c0),
	.w2(32'hbb9bc5bc),
	.w3(32'h3a241fca),
	.w4(32'hbb2b036b),
	.w5(32'hbb1ff099),
	.w6(32'hbb930cf1),
	.w7(32'hbb524ae0),
	.w8(32'hbb0db0ce),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad38756),
	.w1(32'hbc90f806),
	.w2(32'h3b8696b8),
	.w3(32'h39c9f6b1),
	.w4(32'hbc37707a),
	.w5(32'h3aacaffd),
	.w6(32'h3b1f7933),
	.w7(32'hbc391c63),
	.w8(32'h3b02777e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf48335),
	.w1(32'hba545198),
	.w2(32'hb98634f1),
	.w3(32'hbb957e12),
	.w4(32'h3b0619cd),
	.w5(32'hba219530),
	.w6(32'h3b45489a),
	.w7(32'h3b619671),
	.w8(32'h3aa7c7a1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba78b99),
	.w1(32'hbb8d9a73),
	.w2(32'hbaea229d),
	.w3(32'hbb9e7da5),
	.w4(32'hba8ccc32),
	.w5(32'hbaaec1fd),
	.w6(32'hbb2cd552),
	.w7(32'hbaa0ac65),
	.w8(32'hb9ef4ea3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72b04),
	.w1(32'h3b6e9f3e),
	.w2(32'hbb3f7507),
	.w3(32'h39ecfea7),
	.w4(32'hbb3e56c4),
	.w5(32'h3a85ca09),
	.w6(32'hba830bfe),
	.w7(32'h3b975743),
	.w8(32'hbb81cec0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b706),
	.w1(32'h3bedf8fb),
	.w2(32'h3bc4a964),
	.w3(32'hba14a44f),
	.w4(32'h3ba87863),
	.w5(32'h3ac5b069),
	.w6(32'h3c070c71),
	.w7(32'h3add53fe),
	.w8(32'h3ba75acc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2073a),
	.w1(32'hbad33a44),
	.w2(32'hbaad49ce),
	.w3(32'h3a76ce1d),
	.w4(32'h39fd69ff),
	.w5(32'h3b030b55),
	.w6(32'hbb1ed49f),
	.w7(32'hb916ae44),
	.w8(32'h3a3769d4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eb8df),
	.w1(32'h3b3ad92e),
	.w2(32'h39231706),
	.w3(32'h395604cd),
	.w4(32'h3b961c58),
	.w5(32'h3bb6de6d),
	.w6(32'hbb9bbc30),
	.w7(32'hbaf06584),
	.w8(32'hba4b4dda),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57ca8f),
	.w1(32'hbaf55665),
	.w2(32'hbbfc8204),
	.w3(32'h3aa73ca3),
	.w4(32'hbb68a653),
	.w5(32'hbc0b28ba),
	.w6(32'hbb5b069e),
	.w7(32'hbbf383ab),
	.w8(32'hbb177b80),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab12b81),
	.w1(32'hba3a56d8),
	.w2(32'hbbc7c070),
	.w3(32'hbb919c9b),
	.w4(32'hbb4534ca),
	.w5(32'hbb899eab),
	.w6(32'hb9c83cc4),
	.w7(32'hbbacdda5),
	.w8(32'h39b14cc6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62794d),
	.w1(32'hb835cd7e),
	.w2(32'h394b10e9),
	.w3(32'hbb1651ad),
	.w4(32'h3a5f62b4),
	.w5(32'h3ac68721),
	.w6(32'hba47ecb1),
	.w7(32'h3758ee56),
	.w8(32'h3aa55ba9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affbed9),
	.w1(32'h3a03d88f),
	.w2(32'h397bfacf),
	.w3(32'h3a8b5e3f),
	.w4(32'h3aa3b03d),
	.w5(32'h3b2b60a8),
	.w6(32'hb9c98274),
	.w7(32'h3acd637a),
	.w8(32'h3b622639),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b235af3),
	.w1(32'h39e033e5),
	.w2(32'h3c2a946c),
	.w3(32'h3b1392f2),
	.w4(32'h3b477a54),
	.w5(32'h3c7e98dd),
	.w6(32'hbb66df8d),
	.w7(32'h3c1f38e1),
	.w8(32'h3ba26495),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d9926),
	.w1(32'hbc18cd7c),
	.w2(32'hbbdf4b7a),
	.w3(32'h3b6abf2d),
	.w4(32'hbbc67ed3),
	.w5(32'hbc441922),
	.w6(32'hba90cb0f),
	.w7(32'hbb7639f0),
	.w8(32'h3bf6aa68),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8392),
	.w1(32'h3c356546),
	.w2(32'hbbb14b52),
	.w3(32'h3bf02369),
	.w4(32'h3babd8bd),
	.w5(32'hbb9e1736),
	.w6(32'h3b635f9f),
	.w7(32'hbb501d63),
	.w8(32'hbb8ef06d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ffef3),
	.w1(32'hbb2e59d4),
	.w2(32'hbb19b078),
	.w3(32'hbb5be779),
	.w4(32'hb9523b46),
	.w5(32'h3b08e8a6),
	.w6(32'hbb8d6832),
	.w7(32'hbb7c4d05),
	.w8(32'hbb1f2c54),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c9af),
	.w1(32'h3c6c1b28),
	.w2(32'h3bcedeb7),
	.w3(32'hb9903879),
	.w4(32'h3bf03bb8),
	.w5(32'h3b01bd59),
	.w6(32'h3be82943),
	.w7(32'h3bdd98d5),
	.w8(32'hbb3fe990),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e963e),
	.w1(32'hbae34193),
	.w2(32'hbb818819),
	.w3(32'hbaa42471),
	.w4(32'hbb0499db),
	.w5(32'hbb839d93),
	.w6(32'hbb2506e4),
	.w7(32'hbb8ce612),
	.w8(32'hbb8031b1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12607b),
	.w1(32'h3a35370c),
	.w2(32'hba71287e),
	.w3(32'hbba7d1e2),
	.w4(32'h3ad0793d),
	.w5(32'h39cff926),
	.w6(32'h39ec5b4c),
	.w7(32'h3b149e8b),
	.w8(32'hb91dcfe3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b5998),
	.w1(32'hbaa606bd),
	.w2(32'h3b83968c),
	.w3(32'h3a3398de),
	.w4(32'hbb1a30a5),
	.w5(32'hb88a1f87),
	.w6(32'hbaa1e311),
	.w7(32'h39fb55be),
	.w8(32'hbab0f7d6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d82c),
	.w1(32'h3b0e0263),
	.w2(32'hba407286),
	.w3(32'hb9f6572b),
	.w4(32'hbb1cc694),
	.w5(32'h3974856b),
	.w6(32'h3ad256bd),
	.w7(32'h390d9f31),
	.w8(32'hba34fbe0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4fad9),
	.w1(32'hba72993d),
	.w2(32'hbaf66880),
	.w3(32'hbb24e394),
	.w4(32'hb9fd1b26),
	.w5(32'hbb1c42d4),
	.w6(32'hbbe29efc),
	.w7(32'hbb68cd7a),
	.w8(32'hbc1a41fc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc696),
	.w1(32'hbb32b5d0),
	.w2(32'hb8ed0fc0),
	.w3(32'hbb411dfc),
	.w4(32'hba9330a9),
	.w5(32'h3aa97963),
	.w6(32'hbae15402),
	.w7(32'h398ed562),
	.w8(32'h3b8aae84),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf86b),
	.w1(32'h3c7b3cd9),
	.w2(32'hbb6f3eca),
	.w3(32'h3b8500dc),
	.w4(32'h3bf3d01b),
	.w5(32'hbbd08fc4),
	.w6(32'h3ba0ce54),
	.w7(32'hbc102cbc),
	.w8(32'h3bb5fe72),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec5ea),
	.w1(32'hbc4eca41),
	.w2(32'hbc12be62),
	.w3(32'h3be9b17a),
	.w4(32'hbb8329a9),
	.w5(32'h3aabf4d8),
	.w6(32'hbbeb199c),
	.w7(32'hbbae339e),
	.w8(32'h3c12aeeb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05f9d3),
	.w1(32'hbc0d28c1),
	.w2(32'h3c1875d4),
	.w3(32'h36bdc2dd),
	.w4(32'hbbc6771b),
	.w5(32'hbbae20fb),
	.w6(32'hbab3daab),
	.w7(32'hbc15c92f),
	.w8(32'h3b62b257),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c465849),
	.w1(32'hbba6df3c),
	.w2(32'h3b9ec54b),
	.w3(32'h3a9affb2),
	.w4(32'h3bb3e5a8),
	.w5(32'hb9ddd44a),
	.w6(32'hbbd7af2b),
	.w7(32'h3bcfb731),
	.w8(32'hbbade777),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e70a),
	.w1(32'h3ab575fa),
	.w2(32'hbb482cb6),
	.w3(32'hbb130d2c),
	.w4(32'h3ac07650),
	.w5(32'h3a11399a),
	.w6(32'hba4b642e),
	.w7(32'hba18de4f),
	.w8(32'h3b5e9a0f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3ba0e),
	.w1(32'hbb0d18c4),
	.w2(32'hba8e8c69),
	.w3(32'h3b0c5ab5),
	.w4(32'hba9616af),
	.w5(32'h3a4bced5),
	.w6(32'hbabcb1c8),
	.w7(32'h395c1782),
	.w8(32'h3b4137a7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41d366),
	.w1(32'hbbe674f1),
	.w2(32'h3b7c66f8),
	.w3(32'h3aa49438),
	.w4(32'hbb120e78),
	.w5(32'hba6c5c4f),
	.w6(32'hbb883f3b),
	.w7(32'h39fef575),
	.w8(32'h3b142a53),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3746c4),
	.w1(32'hbc691377),
	.w2(32'h3c055395),
	.w3(32'h3b00e19c),
	.w4(32'hbc3acc06),
	.w5(32'hbc068525),
	.w6(32'hbc38db60),
	.w7(32'hbc15db4b),
	.w8(32'hbb8fe43c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d4777),
	.w1(32'hbb962c41),
	.w2(32'hbd1392ca),
	.w3(32'hbb0b9ba3),
	.w4(32'hbb360c9e),
	.w5(32'hbb842243),
	.w6(32'hbb9eda29),
	.w7(32'hbc1ca730),
	.w8(32'hbc705897),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06dd23),
	.w1(32'h3bdeef9a),
	.w2(32'hbc0d1a70),
	.w3(32'h3a3241ab),
	.w4(32'h3b0d413b),
	.w5(32'hbaa1fdd8),
	.w6(32'h3bb3a590),
	.w7(32'h3b542151),
	.w8(32'hbb4a7be1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc616fa6),
	.w1(32'h3a96281f),
	.w2(32'h3c362c50),
	.w3(32'hbba4e615),
	.w4(32'hbb8dc1ca),
	.w5(32'hba9a1f46),
	.w6(32'hbb97ec6d),
	.w7(32'hbae8a11c),
	.w8(32'hbb6f40f1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936531),
	.w1(32'h3b9456e9),
	.w2(32'hbc2e4049),
	.w3(32'h391bdcf2),
	.w4(32'hba309f91),
	.w5(32'hbb277bab),
	.w6(32'h3a43a81d),
	.w7(32'hbaeaee3a),
	.w8(32'h383f34ce),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c6a06),
	.w1(32'h3be7766c),
	.w2(32'hbb5e7a16),
	.w3(32'hba4c2fd6),
	.w4(32'h3b11102d),
	.w5(32'hbb6740d5),
	.w6(32'hbafc60d7),
	.w7(32'hba00c2f6),
	.w8(32'hbb24da16),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf930fb),
	.w1(32'hbbd5071c),
	.w2(32'hb9ec0149),
	.w3(32'hbba4d398),
	.w4(32'hba97cb22),
	.w5(32'hbb15025b),
	.w6(32'hbb400ab5),
	.w7(32'hbbbdae87),
	.w8(32'hba3db65c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bacba),
	.w1(32'hbbcc0346),
	.w2(32'h3a8b729f),
	.w3(32'h3aaebf7b),
	.w4(32'hbc2ad1c4),
	.w5(32'hbcdbec92),
	.w6(32'hbc112a44),
	.w7(32'hbcce6981),
	.w8(32'hbc101393),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af2690),
	.w1(32'h3b438c10),
	.w2(32'hbb8ecba6),
	.w3(32'hbc241add),
	.w4(32'h3a318f97),
	.w5(32'hbaf65d27),
	.w6(32'hbaa41843),
	.w7(32'h388e377a),
	.w8(32'hbaff43f1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5f54),
	.w1(32'hbace3fbc),
	.w2(32'hbb856558),
	.w3(32'hba3a92b6),
	.w4(32'h39cf70b7),
	.w5(32'hba2be439),
	.w6(32'hbaf8c24b),
	.w7(32'hb7dd34de),
	.w8(32'h3a89ff10),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5230),
	.w1(32'hbabf82ed),
	.w2(32'hb8279779),
	.w3(32'h39f94aa5),
	.w4(32'hbaf0f180),
	.w5(32'hba627ba5),
	.w6(32'hbbb66fc5),
	.w7(32'hbb15b635),
	.w8(32'hbaefc1e5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d39b5),
	.w1(32'hbb6a80a1),
	.w2(32'hbb8b734a),
	.w3(32'hbaa26ed3),
	.w4(32'hbb1d6d6a),
	.w5(32'hba1b5dc7),
	.w6(32'hb9c2d563),
	.w7(32'hb91c8897),
	.w8(32'h3b494532),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d3a1),
	.w1(32'hbb77b098),
	.w2(32'h3c62a3f0),
	.w3(32'h39fc8a74),
	.w4(32'hbbddc828),
	.w5(32'h3c70746d),
	.w6(32'hbb0b76a1),
	.w7(32'h3ba253f7),
	.w8(32'hbbb8827f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd84fe),
	.w1(32'h3c33a124),
	.w2(32'hbaf9730e),
	.w3(32'hbac141ad),
	.w4(32'h3b9ecdec),
	.w5(32'hbb541622),
	.w6(32'h3b683177),
	.w7(32'hbbb26a19),
	.w8(32'h3b0ed3cc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038e9b),
	.w1(32'h3b8bf11a),
	.w2(32'h3bf54a2b),
	.w3(32'h3b94d2fa),
	.w4(32'h3a58a233),
	.w5(32'h3b851733),
	.w6(32'h3b1ad4a9),
	.w7(32'h3bfd6cc8),
	.w8(32'hbb38088b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64bb4),
	.w1(32'hbbd65d98),
	.w2(32'hbbfa02e0),
	.w3(32'hbba6332c),
	.w4(32'hbc608c94),
	.w5(32'hbcd5e372),
	.w6(32'hbbd60d3b),
	.w7(32'hbcff40d4),
	.w8(32'hbc2d17f5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ab2c1),
	.w1(32'h3ba80003),
	.w2(32'hbbf888ac),
	.w3(32'hbb5e44f8),
	.w4(32'h3b19a555),
	.w5(32'hbb65779b),
	.w6(32'h3b8fae4b),
	.w7(32'hbb10ed0b),
	.w8(32'hbadf9bfc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb76f80),
	.w1(32'hbaf2b850),
	.w2(32'hbb234ce9),
	.w3(32'hbbf03b21),
	.w4(32'hbb962777),
	.w5(32'hbb97fe2e),
	.w6(32'hbb298686),
	.w7(32'hbb4b4c7c),
	.w8(32'hbb2ee8a5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0648),
	.w1(32'h3b28fd9b),
	.w2(32'hba01dd52),
	.w3(32'hbb7dc484),
	.w4(32'h39e5b9d5),
	.w5(32'h3bad9118),
	.w6(32'h3b4be908),
	.w7(32'h3bc92a66),
	.w8(32'h3aaf5e1c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18f03e),
	.w1(32'hbca44046),
	.w2(32'h3cd7c363),
	.w3(32'h3b94f967),
	.w4(32'hbc8c5648),
	.w5(32'hbc8103fb),
	.w6(32'hbc7192a2),
	.w7(32'hbc7d5c7c),
	.w8(32'h3a069969),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c977a67),
	.w1(32'h3c071ab4),
	.w2(32'hbc1a42ab),
	.w3(32'hba9dc4ad),
	.w4(32'h3ba7fc25),
	.w5(32'hbb47c170),
	.w6(32'h3b860072),
	.w7(32'hbb2e36ae),
	.w8(32'hbb2749c8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46b46),
	.w1(32'h3b079b38),
	.w2(32'hbada5082),
	.w3(32'h3ab4e184),
	.w4(32'h3ac34dce),
	.w5(32'hbb018a8c),
	.w6(32'h38c80a3c),
	.w7(32'hbb0d4467),
	.w8(32'hbb4387ec),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dbc62),
	.w1(32'h3a814e5e),
	.w2(32'hbb480ef7),
	.w3(32'hba1022ea),
	.w4(32'h3ae2373f),
	.w5(32'h3a2cda5d),
	.w6(32'h3a04b7a1),
	.w7(32'h3a88ba34),
	.w8(32'h39ad2f5c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994f4d3),
	.w1(32'hba2e9cba),
	.w2(32'hbaa9ed74),
	.w3(32'h3abe1d79),
	.w4(32'hba02e3e5),
	.w5(32'h3adc7e24),
	.w6(32'hbb1c0016),
	.w7(32'hba070b08),
	.w8(32'h3b072198),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16943d),
	.w1(32'h3bcfaa70),
	.w2(32'hbbc1c826),
	.w3(32'h3b0c64d8),
	.w4(32'h3b26d593),
	.w5(32'h3b4f4571),
	.w6(32'h3a200f9c),
	.w7(32'h3b55692f),
	.w8(32'hbb603fd0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb313d00),
	.w1(32'hbc5749e6),
	.w2(32'h3aebdbf5),
	.w3(32'h3bc36fbb),
	.w4(32'h3a092e9b),
	.w5(32'hbb5a604e),
	.w6(32'hbca09fba),
	.w7(32'hbb4763a7),
	.w8(32'hbc3b2b58),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc095ef),
	.w1(32'hbbc59138),
	.w2(32'h3a86e64e),
	.w3(32'hbba7e804),
	.w4(32'hbad5e758),
	.w5(32'hbbafd43f),
	.w6(32'hbb345325),
	.w7(32'hbb4b0e00),
	.w8(32'h3bb7254f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e7685),
	.w1(32'hbbb74bab),
	.w2(32'hba7c881d),
	.w3(32'h3a487aa1),
	.w4(32'hbb18b8a2),
	.w5(32'h3b0a7dc6),
	.w6(32'hbbab507b),
	.w7(32'h3ae30627),
	.w8(32'hbbb8b302),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38836),
	.w1(32'hb9cbe36b),
	.w2(32'hbc970df0),
	.w3(32'hbb62cd24),
	.w4(32'h3a3fa9ac),
	.w5(32'h3aff2dbf),
	.w6(32'h3b9a644f),
	.w7(32'hbb9f0a7e),
	.w8(32'h3b11dd2e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac86f62),
	.w1(32'hba21364c),
	.w2(32'hbb61259e),
	.w3(32'h3b6e8e7d),
	.w4(32'hb8d645ef),
	.w5(32'hba0256b7),
	.w6(32'hbaa8e490),
	.w7(32'hbb1a59da),
	.w8(32'h39604dca),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8618),
	.w1(32'h3b7e1329),
	.w2(32'hbb343c95),
	.w3(32'h3ac1f2ca),
	.w4(32'h3a759192),
	.w5(32'hbae04571),
	.w6(32'h3b1ae749),
	.w7(32'h3910e351),
	.w8(32'hba0ce622),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5cb7),
	.w1(32'h3bf0b27b),
	.w2(32'h3b66a463),
	.w3(32'hba269006),
	.w4(32'h3b64143f),
	.w5(32'h3ba5193d),
	.w6(32'h3b704289),
	.w7(32'h3b8f8cd3),
	.w8(32'hbb1b5b4d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc52eb),
	.w1(32'h3bbaca16),
	.w2(32'hbb40f9aa),
	.w3(32'hbaef8983),
	.w4(32'hba33a2ff),
	.w5(32'h3a15f8c5),
	.w6(32'h3b20f7d0),
	.w7(32'h3ade575e),
	.w8(32'hbaeb17f8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ab658),
	.w1(32'h3b85fe01),
	.w2(32'hbb6811bc),
	.w3(32'hbaba99fe),
	.w4(32'hb9c0a12e),
	.w5(32'h3a6c176a),
	.w6(32'hbaa4c095),
	.w7(32'hbb04c65e),
	.w8(32'hbaccad6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5497),
	.w1(32'hbb7b87db),
	.w2(32'h3b8f02c7),
	.w3(32'hbb64e821),
	.w4(32'h3b570d17),
	.w5(32'h3b2ff227),
	.w6(32'hbb1f317d),
	.w7(32'hba87e160),
	.w8(32'hbba6a8d1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb958b65),
	.w1(32'h3b29b3d3),
	.w2(32'hbbb76950),
	.w3(32'hbb3e5fb9),
	.w4(32'h3a96878b),
	.w5(32'hbb56cc5d),
	.w6(32'h3b5ffe5c),
	.w7(32'hbb08d348),
	.w8(32'hbb5d7409),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef1a18),
	.w1(32'hbb9cd28e),
	.w2(32'hbad02ea4),
	.w3(32'hbbc93d85),
	.w4(32'hbb7ccb58),
	.w5(32'hbb58debc),
	.w6(32'hbc0586cd),
	.w7(32'hbaa9660f),
	.w8(32'hbb89f839),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caaf81a),
	.w1(32'h380e0fe2),
	.w2(32'hbaa3a913),
	.w3(32'hba31445f),
	.w4(32'hb9ab2825),
	.w5(32'h3a259ce7),
	.w6(32'hba8dd294),
	.w7(32'hb9d3b21d),
	.w8(32'h398d7a1f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a7ecf),
	.w1(32'h3b7e5f5e),
	.w2(32'hbbfadec4),
	.w3(32'h3a910e85),
	.w4(32'hba82be5e),
	.w5(32'hbb03c1fa),
	.w6(32'h39c1aa60),
	.w7(32'hbad5861f),
	.w8(32'hbb22b2c7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcae02e),
	.w1(32'hba55c179),
	.w2(32'hba6bc1d5),
	.w3(32'hba9b8f33),
	.w4(32'h39e1474b),
	.w5(32'h3a8ff9d2),
	.w6(32'hbb098601),
	.w7(32'hb9d8d93b),
	.w8(32'h3acb4cf5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2447f9),
	.w1(32'hbabc1d7c),
	.w2(32'hbac2d6d7),
	.w3(32'h3b1a82c2),
	.w4(32'hb864b7ae),
	.w5(32'h3aadae7b),
	.w6(32'hbac41ad4),
	.w7(32'hb9bf945e),
	.w8(32'h39a125ce),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1ab4d),
	.w1(32'hbaa75c17),
	.w2(32'hbb088ef0),
	.w3(32'h3a28345c),
	.w4(32'hba454845),
	.w5(32'hbb20c4e2),
	.w6(32'hbb3fff12),
	.w7(32'hbb99cddb),
	.w8(32'h39fb4706),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5212ad),
	.w1(32'h3c8f0b84),
	.w2(32'hbc494308),
	.w3(32'h3a4ca247),
	.w4(32'h3c566166),
	.w5(32'hba9b7a7e),
	.w6(32'h3bfbb60a),
	.w7(32'hbafe0a81),
	.w8(32'hbc23df06),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe4c2a),
	.w1(32'h3b290518),
	.w2(32'hba513556),
	.w3(32'hbc146d52),
	.w4(32'hba45333e),
	.w5(32'hbac90542),
	.w6(32'h37dd4b05),
	.w7(32'h3a74e703),
	.w8(32'h3a1a9aa6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ce445),
	.w1(32'h3a9f5c1e),
	.w2(32'h39fb1474),
	.w3(32'hbacac6a5),
	.w4(32'h3a194e14),
	.w5(32'hbb6b4f43),
	.w6(32'h3b2c5f87),
	.w7(32'hbb13c6ab),
	.w8(32'hbb64cdb8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28277b),
	.w1(32'hb91d77f9),
	.w2(32'h3c0c093b),
	.w3(32'hbb92c3ec),
	.w4(32'h3b70cbf5),
	.w5(32'h3bfd2acf),
	.w6(32'hbb8806e4),
	.w7(32'h3b030ada),
	.w8(32'h39c38b73),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0081c6),
	.w1(32'hb9dc5f2f),
	.w2(32'hbb9ead35),
	.w3(32'hbbbbcc45),
	.w4(32'h3b4535b7),
	.w5(32'hbb8f3d56),
	.w6(32'h3b98b70b),
	.w7(32'h393e242e),
	.w8(32'hbab2d521),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1be4b),
	.w1(32'hbb3050ba),
	.w2(32'hbb3d68ee),
	.w3(32'hbac2b361),
	.w4(32'hb9cd2da7),
	.w5(32'h3b7d10ca),
	.w6(32'hbb0ac3f1),
	.w7(32'hbb55b1a8),
	.w8(32'hbb09a797),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27eea8),
	.w1(32'h3b0b50e4),
	.w2(32'hbb4ec0fd),
	.w3(32'hbab6702d),
	.w4(32'hb98a78d7),
	.w5(32'hbb0bab33),
	.w6(32'h3b1cfcda),
	.w7(32'hbac1c2dd),
	.w8(32'hbb9a1857),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a9ae9),
	.w1(32'h3c3ce193),
	.w2(32'hbc43e47d),
	.w3(32'hbb858d30),
	.w4(32'h3b387b9a),
	.w5(32'hbba5ffb6),
	.w6(32'h3b81d302),
	.w7(32'h3a87d1fe),
	.w8(32'hbc10a172),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca95b5f),
	.w1(32'hbc34ffd3),
	.w2(32'h3b91f640),
	.w3(32'hbb97d14f),
	.w4(32'hbc16dc59),
	.w5(32'hbccb48b8),
	.w6(32'hbc1e0675),
	.w7(32'hbcae1e9e),
	.w8(32'hbb9c0eb0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8732db),
	.w1(32'hbba779ad),
	.w2(32'hbb290834),
	.w3(32'hbb45447d),
	.w4(32'hbc195a47),
	.w5(32'hbb9e9168),
	.w6(32'hbc06d227),
	.w7(32'hbc992841),
	.w8(32'hbc867d52),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d3480),
	.w1(32'hbc1a8f1c),
	.w2(32'h3afe3d62),
	.w3(32'hbb972028),
	.w4(32'hbb1ad0aa),
	.w5(32'hbc0be2e3),
	.w6(32'hbb874abf),
	.w7(32'hbb9a2e37),
	.w8(32'h3c16138b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2c9b8),
	.w1(32'h3bb3473e),
	.w2(32'h3b983a9f),
	.w3(32'h3ab903a9),
	.w4(32'h3bdd0efb),
	.w5(32'h3b420847),
	.w6(32'h3b490124),
	.w7(32'h3a7f8899),
	.w8(32'h398fc2e4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb711c30),
	.w1(32'hbb7213fe),
	.w2(32'h39b94eea),
	.w3(32'h3a8b3854),
	.w4(32'hba42f5f8),
	.w5(32'hbb671fc5),
	.w6(32'hbabef989),
	.w7(32'hbb01de52),
	.w8(32'h3b804106),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d9a77),
	.w1(32'hbb962c1a),
	.w2(32'hb9b4e9a1),
	.w3(32'h3a74a6a8),
	.w4(32'h3961c6fe),
	.w5(32'h3b5bed60),
	.w6(32'hbb87e13d),
	.w7(32'h3a8aca3a),
	.w8(32'h3b0a699f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc883e4),
	.w1(32'h38aa4eec),
	.w2(32'hb9fcdaea),
	.w3(32'h3a9b3d8d),
	.w4(32'h3a313018),
	.w5(32'hbb3667db),
	.w6(32'h3b1aa7cd),
	.w7(32'hbb23caa6),
	.w8(32'hbb80a248),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e36cf),
	.w1(32'hbb061b83),
	.w2(32'hbb2b587a),
	.w3(32'hbb7b34ba),
	.w4(32'hbae5ed78),
	.w5(32'hba3a4bce),
	.w6(32'hbb53b9f2),
	.w7(32'hba9d17c6),
	.w8(32'hba788365),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b41c2f),
	.w1(32'hbbaf2f0b),
	.w2(32'h3ac8c09c),
	.w3(32'hbab84dd8),
	.w4(32'hbabf7f6f),
	.w5(32'hbb98d41a),
	.w6(32'hbb1e1f77),
	.w7(32'hbb35465a),
	.w8(32'h3b978336),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2996dd),
	.w1(32'hbc0537e5),
	.w2(32'hbbb5da5f),
	.w3(32'h39370826),
	.w4(32'hbb8b4335),
	.w5(32'hbaad49c5),
	.w6(32'hbbf86237),
	.w7(32'hbb3b3043),
	.w8(32'h39a3872f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c857c18),
	.w1(32'hbb491d38),
	.w2(32'hbbbe9697),
	.w3(32'hbbbce8c6),
	.w4(32'hbb102e57),
	.w5(32'h39c11df4),
	.w6(32'h39865755),
	.w7(32'h3b03142d),
	.w8(32'hbb090fe1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87796f),
	.w1(32'hbc76bfd2),
	.w2(32'hbc662b14),
	.w3(32'h3b07f30e),
	.w4(32'hbc4b41db),
	.w5(32'h3be8ddd3),
	.w6(32'hbc1949f4),
	.w7(32'hbbdf33ef),
	.w8(32'hbc90bb60),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dc122),
	.w1(32'h3b229e28),
	.w2(32'hbb7b09f4),
	.w3(32'hbc1a83ff),
	.w4(32'h3a7bd096),
	.w5(32'h3b69f517),
	.w6(32'h3b5401d9),
	.w7(32'h3b80fa67),
	.w8(32'hbad8c5fd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ee88e),
	.w1(32'hbabe460d),
	.w2(32'hb9d9d952),
	.w3(32'h3b84747e),
	.w4(32'h3abfcd19),
	.w5(32'hbb279726),
	.w6(32'hbb2b9981),
	.w7(32'hbb711e3b),
	.w8(32'hbbf23b3e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8fb8c),
	.w1(32'hbbfb7697),
	.w2(32'h3b73929a),
	.w3(32'hbac6ba68),
	.w4(32'hbb7b93fa),
	.w5(32'h3b599963),
	.w6(32'hbb9df1c2),
	.w7(32'hbb22e4f2),
	.w8(32'hb949901f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c933ce0),
	.w1(32'hbbe2c874),
	.w2(32'h3aaad6e9),
	.w3(32'hbadded38),
	.w4(32'hbae7d561),
	.w5(32'hbbc51ed6),
	.w6(32'hbb415718),
	.w7(32'hbb5b13ec),
	.w8(32'h3bd77325),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ab69b),
	.w1(32'hb908605b),
	.w2(32'h39af4fde),
	.w3(32'h3a6f5196),
	.w4(32'h3a9d29d4),
	.w5(32'hba126c87),
	.w6(32'h3b087022),
	.w7(32'hba50e472),
	.w8(32'hba1ee164),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72d13),
	.w1(32'h3a72447e),
	.w2(32'hb98c4a98),
	.w3(32'hb96786e5),
	.w4(32'h3b2dcf4d),
	.w5(32'hba11e42d),
	.w6(32'h3b271176),
	.w7(32'h38b9da29),
	.w8(32'h3a27e25b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08bcca),
	.w1(32'hbc750327),
	.w2(32'hbc0f7660),
	.w3(32'h3983261e),
	.w4(32'hbc3d4a69),
	.w5(32'hbb0d059a),
	.w6(32'hbbbf9722),
	.w7(32'hbc3b6fd8),
	.w8(32'h3b68e49b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ca088),
	.w1(32'hbbc5317b),
	.w2(32'hbb213643),
	.w3(32'hbbb3f883),
	.w4(32'hbbbaa8fb),
	.w5(32'hbc2c0dd2),
	.w6(32'hbb6b0014),
	.w7(32'hbc438598),
	.w8(32'hbb356e04),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0294bb),
	.w1(32'h3ad18c72),
	.w2(32'h3ba726bf),
	.w3(32'h3b2b1d6c),
	.w4(32'h3c1300dc),
	.w5(32'h3bb9e1b6),
	.w6(32'hb9f48ed5),
	.w7(32'h392c8f43),
	.w8(32'hba2faee0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcdcf),
	.w1(32'hba9c6b01),
	.w2(32'hbb510fa6),
	.w3(32'hba7cbcce),
	.w4(32'hbb344b54),
	.w5(32'h3a8364bd),
	.w6(32'hbadfd0c8),
	.w7(32'h3b7431eb),
	.w8(32'hbae10178),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31e46b),
	.w1(32'hbb3bb663),
	.w2(32'hba1f419c),
	.w3(32'hba9d537f),
	.w4(32'h39af332a),
	.w5(32'hba0eb8bf),
	.w6(32'hbadaa86c),
	.w7(32'hb91c6a6f),
	.w8(32'h3a53693f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d385b),
	.w1(32'hbbc8c1e6),
	.w2(32'hbb6c1c2f),
	.w3(32'h38bf5645),
	.w4(32'hbc478e5a),
	.w5(32'h3b00ace2),
	.w6(32'h3b0c7fde),
	.w7(32'hbc14842d),
	.w8(32'h3b3b736a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfcfd9),
	.w1(32'h3c82c2de),
	.w2(32'hba5b86f7),
	.w3(32'hbb5829e3),
	.w4(32'h3c27b9e6),
	.w5(32'h3ad63672),
	.w6(32'h3c1fe207),
	.w7(32'h3c04b176),
	.w8(32'hbaa99538),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd14c65),
	.w1(32'h39c76536),
	.w2(32'hbb01e73c),
	.w3(32'hbb6e985c),
	.w4(32'hb986e59b),
	.w5(32'h3ad077d4),
	.w6(32'hbabf2bd2),
	.w7(32'hb72ae1fb),
	.w8(32'h3a8cabab),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbda49),
	.w1(32'h3788fea7),
	.w2(32'h37ee38e6),
	.w3(32'h3b12b140),
	.w4(32'h36b9b5ea),
	.w5(32'h3724fdde),
	.w6(32'h37ae0115),
	.w7(32'h37ee94ed),
	.w8(32'h3752cd37),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c2739c),
	.w1(32'h37d57a4a),
	.w2(32'hb6871a80),
	.w3(32'h37553983),
	.w4(32'h3826e286),
	.w5(32'h37e2cad2),
	.w6(32'hb859d35b),
	.w7(32'hb790a762),
	.w8(32'hb6bb1f29),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38950433),
	.w1(32'h3827ea75),
	.w2(32'hb85b721f),
	.w3(32'h38420aba),
	.w4(32'h3885414f),
	.w5(32'hb7b82a88),
	.w6(32'hb8c183e3),
	.w7(32'hb89d7c1a),
	.w8(32'h37c6a429),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70677c1),
	.w1(32'h368fbaa1),
	.w2(32'h368dbeb1),
	.w3(32'hb3ba832f),
	.w4(32'hb705f3b7),
	.w5(32'hb735dc54),
	.w6(32'h36404d28),
	.w7(32'hb6289125),
	.w8(32'hb5d3a810),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82918ed),
	.w1(32'hb7fb371f),
	.w2(32'hb40805ff),
	.w3(32'hb88bd575),
	.w4(32'hb89f5ffd),
	.w5(32'hb806888d),
	.w6(32'hb7c958f3),
	.w7(32'hb83ed553),
	.w8(32'hb76e005a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379daed0),
	.w1(32'h378d4a8c),
	.w2(32'h35f8e61a),
	.w3(32'h35dcee2f),
	.w4(32'h36e13f82),
	.w5(32'h3705b614),
	.w6(32'hb7c5451c),
	.w7(32'hb7c9118b),
	.w8(32'hb839b4b7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d34f50),
	.w1(32'h37e8ab11),
	.w2(32'h377fa972),
	.w3(32'hb7d4b84e),
	.w4(32'h3800f2b8),
	.w5(32'h38086806),
	.w6(32'hb8842843),
	.w7(32'hb82cb3f3),
	.w8(32'hb857b2a8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76b6c8c),
	.w1(32'hb728ef0f),
	.w2(32'h371baba0),
	.w3(32'h3710fc3b),
	.w4(32'hb7ded461),
	.w5(32'hb70cc468),
	.w6(32'hb80c0e94),
	.w7(32'hb751e548),
	.w8(32'hb6416cc4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387483ce),
	.w1(32'h38a92031),
	.w2(32'h382a56b0),
	.w3(32'h3895e99b),
	.w4(32'h38aa546f),
	.w5(32'h38455cf3),
	.w6(32'hb7855286),
	.w7(32'h381342c6),
	.w8(32'h383b51a7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378fb418),
	.w1(32'h38673dc5),
	.w2(32'h38c6d561),
	.w3(32'hb8145572),
	.w4(32'h38426f6f),
	.w5(32'h38120459),
	.w6(32'hb87e11f3),
	.w7(32'hb5ee2347),
	.w8(32'hb820eef8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b3fac1),
	.w1(32'h381470d2),
	.w2(32'h3830fa3d),
	.w3(32'h382177c8),
	.w4(32'h37d6d61d),
	.w5(32'h383dab99),
	.w6(32'h37d94e22),
	.w7(32'h38796d49),
	.w8(32'h382d5a83),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb67bb),
	.w1(32'h392fed67),
	.w2(32'h38e85b5a),
	.w3(32'h381f1307),
	.w4(32'h390e2fff),
	.w5(32'h38ecb356),
	.w6(32'h379dfa71),
	.w7(32'h382ad821),
	.w8(32'h3895ede2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a98b09),
	.w1(32'hb6e66a36),
	.w2(32'h36f6606e),
	.w3(32'h384fccd6),
	.w4(32'h3806fb28),
	.w5(32'hb8b9e0e6),
	.w6(32'hb829bbb2),
	.w7(32'hb841779b),
	.w8(32'hb7140f88),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386204ce),
	.w1(32'h38d08c0d),
	.w2(32'h37fe7641),
	.w3(32'h37140c6b),
	.w4(32'h39011ac6),
	.w5(32'h380cfd2b),
	.w6(32'hb847b5e9),
	.w7(32'h380f0cf9),
	.w8(32'h370962d1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d40939),
	.w1(32'h36d6cae3),
	.w2(32'h371db695),
	.w3(32'h370fb67d),
	.w4(32'h37c54faf),
	.w5(32'h379ca48f),
	.w6(32'hb7e31394),
	.w7(32'hb749e7a5),
	.w8(32'h36100db8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843e5ce),
	.w1(32'h38d0caf2),
	.w2(32'h384bb9ee),
	.w3(32'hb80d5adb),
	.w4(32'h38ae5aba),
	.w5(32'h37b6339d),
	.w6(32'hb850b0ab),
	.w7(32'h38088fe8),
	.w8(32'h3792f334),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954a580),
	.w1(32'h394de996),
	.w2(32'h38bbbe6e),
	.w3(32'h392bb9ca),
	.w4(32'h3944b832),
	.w5(32'hb70e19ba),
	.w6(32'h390d0196),
	.w7(32'h38fe2937),
	.w8(32'hb880dd30),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78b73da),
	.w1(32'hb765a0f2),
	.w2(32'hb6637185),
	.w3(32'hb49d8c8b),
	.w4(32'hb783a79a),
	.w5(32'hb6c18e39),
	.w6(32'hb7ac07f4),
	.w7(32'hb72df015),
	.w8(32'hb6da313f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70e520e),
	.w1(32'h36bae3a4),
	.w2(32'hb67a36fe),
	.w3(32'hb6a36066),
	.w4(32'h353946d2),
	.w5(32'hb740dcf0),
	.w6(32'hb6011adf),
	.w7(32'hb7577f8a),
	.w8(32'hb7920314),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71cdc80),
	.w1(32'h366ffe65),
	.w2(32'h375c24a7),
	.w3(32'hb7653789),
	.w4(32'hb72be87f),
	.w5(32'hb6e98bc7),
	.w6(32'h342c9dcd),
	.w7(32'hb789064a),
	.w8(32'hb743a836),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930a952),
	.w1(32'h39790b79),
	.w2(32'h3959515a),
	.w3(32'h38dee468),
	.w4(32'h394384bb),
	.w5(32'h38a3c7cf),
	.w6(32'h38ef28da),
	.w7(32'h390a5b84),
	.w8(32'h38a086ff),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d0ca88),
	.w1(32'hb91f9875),
	.w2(32'hb8ef4e6d),
	.w3(32'hb9335352),
	.w4(32'hb88b7853),
	.w5(32'h379fec40),
	.w6(32'hb9ac68dd),
	.w7(32'hb98305f3),
	.w8(32'hb9080eb8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36daaf2e),
	.w1(32'h3720eed6),
	.w2(32'h378077d0),
	.w3(32'h3682d2ad),
	.w4(32'hb6b11690),
	.w5(32'h362d3019),
	.w6(32'h3699c35c),
	.w7(32'h37a91cfa),
	.w8(32'h3688a055),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c153ff),
	.w1(32'h38390ced),
	.w2(32'h36d65979),
	.w3(32'h387d4ba2),
	.w4(32'h38f4074e),
	.w5(32'h3707cbc3),
	.w6(32'hb8db3e8b),
	.w7(32'hb804b0c9),
	.w8(32'h372017a1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38580be4),
	.w1(32'h378c7704),
	.w2(32'hb5cdb1f2),
	.w3(32'h378f6d16),
	.w4(32'h38333c3e),
	.w5(32'h374c06d0),
	.w6(32'hb8792a21),
	.w7(32'hb5d0f0f5),
	.w8(32'h373d9795),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37964c4f),
	.w1(32'h38830ae3),
	.w2(32'h38249747),
	.w3(32'h36b46f01),
	.w4(32'h38b2e513),
	.w5(32'h38bf3f7e),
	.w6(32'hb7b46fb9),
	.w7(32'h382ae310),
	.w8(32'h38868298),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed7290),
	.w1(32'h385b30ed),
	.w2(32'h37d38398),
	.w3(32'hb6c98515),
	.w4(32'h37f0f688),
	.w5(32'h379abcd8),
	.w6(32'hb8350560),
	.w7(32'hb813559c),
	.w8(32'hb7f03c36),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384fd459),
	.w1(32'h38c57011),
	.w2(32'h389bf4bc),
	.w3(32'h38d4f727),
	.w4(32'h38aa9534),
	.w5(32'h38a02b59),
	.w6(32'h38aa7672),
	.w7(32'h38988069),
	.w8(32'h383548d6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374288f1),
	.w1(32'h36bee7cf),
	.w2(32'h37f506e9),
	.w3(32'h38032821),
	.w4(32'hb75b39a7),
	.w5(32'h37e43e76),
	.w6(32'h368ee661),
	.w7(32'h374aebb2),
	.w8(32'h3822eb70),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5922012),
	.w1(32'h37f40659),
	.w2(32'hb724537e),
	.w3(32'hb6dc1f46),
	.w4(32'h3851e361),
	.w5(32'h36bc6834),
	.w6(32'hb89e3bd2),
	.w7(32'hb7e07609),
	.w8(32'hb7fe3ee4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817720a),
	.w1(32'h38310049),
	.w2(32'hb80a3d76),
	.w3(32'h36fc35f7),
	.w4(32'h3704e2d3),
	.w5(32'hb8848de6),
	.w6(32'h382c4161),
	.w7(32'h38b74c90),
	.w8(32'hb8c9218a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83de5c9),
	.w1(32'hb8675c40),
	.w2(32'hb87dbbe2),
	.w3(32'hb8a370d9),
	.w4(32'hb8bdd84c),
	.w5(32'hb8314072),
	.w6(32'hb7bd5f9f),
	.w7(32'hb83fc011),
	.w8(32'hb7972f0d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72a3a4a),
	.w1(32'h372537f8),
	.w2(32'h3784dfef),
	.w3(32'hb7718c5b),
	.w4(32'hb5e22afd),
	.w5(32'h37141601),
	.w6(32'h369c031a),
	.w7(32'h3764e3b5),
	.w8(32'h37484f80),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fe909a),
	.w1(32'h36515b98),
	.w2(32'h36c6467f),
	.w3(32'h36c5e9ed),
	.w4(32'hb6a33092),
	.w5(32'h3530b913),
	.w6(32'hb5e41e30),
	.w7(32'hb502173f),
	.w8(32'h362de213),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828af16),
	.w1(32'h380fcc11),
	.w2(32'h370c3843),
	.w3(32'h37f13fad),
	.w4(32'h368c9b55),
	.w5(32'h375bcc70),
	.w6(32'h373adb4f),
	.w7(32'h36bc80e5),
	.w8(32'h37f6d945),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3558f93f),
	.w1(32'hb7bacb91),
	.w2(32'h38071066),
	.w3(32'h370790e3),
	.w4(32'hb7ec4957),
	.w5(32'h3776488f),
	.w6(32'hb7a079fd),
	.w7(32'hb6a04756),
	.w8(32'h3630080f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68c71c1),
	.w1(32'h387f33ae),
	.w2(32'h374f5c52),
	.w3(32'hb79e73a6),
	.w4(32'h3866b212),
	.w5(32'h37f1dc1f),
	.w6(32'hb84a9a37),
	.w7(32'hb88126d7),
	.w8(32'h377df499),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368928a7),
	.w1(32'hb6488d9d),
	.w2(32'h376af3b0),
	.w3(32'hb7acdd9f),
	.w4(32'hb7a18ff9),
	.w5(32'h37091987),
	.w6(32'hb706638e),
	.w7(32'hb7363415),
	.w8(32'h36e954e6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3844c020),
	.w1(32'hb8ad5670),
	.w2(32'hb81994cf),
	.w3(32'h380b6619),
	.w4(32'hb911b517),
	.w5(32'hb87f02db),
	.w6(32'h36c1a8a4),
	.w7(32'h372b7539),
	.w8(32'h3780aa39),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3640d891),
	.w1(32'h3796ffe0),
	.w2(32'h37ab5565),
	.w3(32'hb717147f),
	.w4(32'h36c545a4),
	.w5(32'h364a1376),
	.w6(32'h3786cb92),
	.w7(32'h37698015),
	.w8(32'h36a6a4ea),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372a3823),
	.w1(32'h361bccb9),
	.w2(32'h377a2d82),
	.w3(32'hb6a2e05b),
	.w4(32'hb6f45c00),
	.w5(32'h3693005c),
	.w6(32'h36bb39a6),
	.w7(32'h3759371d),
	.w8(32'h37653323),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881bcca),
	.w1(32'h3899b0e8),
	.w2(32'h3881f190),
	.w3(32'hb63359f9),
	.w4(32'h37e07d46),
	.w5(32'h36a1b483),
	.w6(32'hb7f6204c),
	.w7(32'hb86d79f6),
	.w8(32'hb78fe76e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39239acc),
	.w1(32'h390d2945),
	.w2(32'h375671dd),
	.w3(32'h392829a2),
	.w4(32'h38d78dc3),
	.w5(32'hb88be2e6),
	.w6(32'hb79bed37),
	.w7(32'h383d7017),
	.w8(32'hb8798475),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d04e56),
	.w1(32'hb8a857eb),
	.w2(32'hb7ed0800),
	.w3(32'hb8502d06),
	.w4(32'hb8be4d21),
	.w5(32'hb653c00a),
	.w6(32'hb818eb27),
	.w7(32'hb820ab64),
	.w8(32'hb732eb44),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38033566),
	.w1(32'h384e62e2),
	.w2(32'h380d0a27),
	.w3(32'h3783dae9),
	.w4(32'h38e5e008),
	.w5(32'h387ca6c2),
	.w6(32'hb854b0e7),
	.w7(32'hb7dfb3af),
	.w8(32'hb7914154),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3629e2d3),
	.w1(32'h370acca7),
	.w2(32'h365cfad3),
	.w3(32'hb659b708),
	.w4(32'hb7b4c7ec),
	.w5(32'hb784f409),
	.w6(32'hb77fec1d),
	.w7(32'hb7f831a4),
	.w8(32'hb770a551),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81876e4),
	.w1(32'hb91eef8f),
	.w2(32'hb91bd39d),
	.w3(32'hb895ed9f),
	.w4(32'hb90443a2),
	.w5(32'hb9390907),
	.w6(32'hb8e02709),
	.w7(32'hb91315b1),
	.w8(32'hb8fb505e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ded3f2),
	.w1(32'h382450c5),
	.w2(32'h389f8110),
	.w3(32'hb5d021fe),
	.w4(32'hb74d4c74),
	.w5(32'h3840dcf0),
	.w6(32'h371df66e),
	.w7(32'hb6e3ef5d),
	.w8(32'h37b20802),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e0e1e),
	.w1(32'h38453e39),
	.w2(32'h37578b6f),
	.w3(32'h3827882d),
	.w4(32'h3901f99a),
	.w5(32'h3868dcbd),
	.w6(32'hb9050dcb),
	.w7(32'hb7ebd90e),
	.w8(32'hb839c1b0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73eaed7),
	.w1(32'h374cb447),
	.w2(32'hb4dbe805),
	.w3(32'h364915ba),
	.w4(32'hb7086b70),
	.w5(32'hb79d2098),
	.w6(32'hb67d51d8),
	.w7(32'hb695215f),
	.w8(32'h3715aedd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900b9ef),
	.w1(32'h38c4218b),
	.w2(32'h3882c626),
	.w3(32'h38d048db),
	.w4(32'h38911aa3),
	.w5(32'hb7ce65e0),
	.w6(32'h383ef020),
	.w7(32'h3883b5cf),
	.w8(32'h375ee3bf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364222ba),
	.w1(32'hb5c5ffeb),
	.w2(32'h361b005b),
	.w3(32'h36948fb3),
	.w4(32'hb6e58afb),
	.w5(32'hb67a995f),
	.w6(32'hb7019184),
	.w7(32'h3621c6e4),
	.w8(32'hb5d09a3d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da8758),
	.w1(32'h36b58f79),
	.w2(32'hb7b1a5d0),
	.w3(32'hb6998192),
	.w4(32'h36c3c123),
	.w5(32'hb71b825b),
	.w6(32'hb7c731e1),
	.w7(32'hb7d39928),
	.w8(32'hb8906d40),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb771331a),
	.w1(32'h37f721ff),
	.w2(32'h3761d10b),
	.w3(32'hb72a62ec),
	.w4(32'h35b23b8d),
	.w5(32'h375a7edb),
	.w6(32'hb647c342),
	.w7(32'hb7be9506),
	.w8(32'h361d86d5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6833561),
	.w1(32'hb86a8794),
	.w2(32'hb89ba0de),
	.w3(32'hb732718d),
	.w4(32'hb842d514),
	.w5(32'hb8829da1),
	.w6(32'hb8220d43),
	.w7(32'h36cca2ce),
	.w8(32'hb6e04bc1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7407f4a),
	.w1(32'hb708d099),
	.w2(32'h37184ad7),
	.w3(32'hb7960b63),
	.w4(32'hb6d05800),
	.w5(32'hb745c34f),
	.w6(32'hb74c71a9),
	.w7(32'h36e4e1fd),
	.w8(32'hb745def3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375a4fbc),
	.w1(32'h368acf82),
	.w2(32'h368cdec1),
	.w3(32'hb6143bb3),
	.w4(32'h359be9f7),
	.w5(32'h37256e79),
	.w6(32'h361e4452),
	.w7(32'hb61f821c),
	.w8(32'hb4c70f6c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb618ac56),
	.w1(32'hb71760c4),
	.w2(32'hb669322d),
	.w3(32'h369d7c14),
	.w4(32'h3559622d),
	.w5(32'hb7744f61),
	.w6(32'hb7474cba),
	.w7(32'hb6c2928c),
	.w8(32'h3699afc7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f9bd1b),
	.w1(32'h35b64f28),
	.w2(32'h3784a6ee),
	.w3(32'hb8a9257b),
	.w4(32'hb7d8e108),
	.w5(32'h38004f92),
	.w6(32'hb7e262f5),
	.w7(32'h3673e726),
	.w8(32'h38416357),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d1caa5),
	.w1(32'hb75e8d23),
	.w2(32'h37d827a0),
	.w3(32'hb6875df4),
	.w4(32'hb63179dc),
	.w5(32'h37bcd736),
	.w6(32'hb6978f7c),
	.w7(32'hb7175cd4),
	.w8(32'hb8325504),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3538fdd3),
	.w1(32'hb7ab47a4),
	.w2(32'hb685367c),
	.w3(32'h37a06421),
	.w4(32'hb828c5b0),
	.w5(32'hb7941f3d),
	.w6(32'h36ce7aca),
	.w7(32'hb608b5f7),
	.w8(32'hb7639228),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954110b),
	.w1(32'hb8d30fa4),
	.w2(32'hb93bc816),
	.w3(32'hb8bde682),
	.w4(32'h38e4de11),
	.w5(32'h38a0a3b2),
	.w6(32'hb9ed4f33),
	.w7(32'hb94d53b0),
	.w8(32'hb8eb3c39),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b28802),
	.w1(32'h37e068ba),
	.w2(32'hb6214355),
	.w3(32'h3890c259),
	.w4(32'h3745afbd),
	.w5(32'hb6ea136b),
	.w6(32'h388a5c97),
	.w7(32'h38f84908),
	.w8(32'hb6f56c8b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377757e5),
	.w1(32'hb75c4d29),
	.w2(32'h36e10a00),
	.w3(32'h373526a8),
	.w4(32'hb719d359),
	.w5(32'h3731f39b),
	.w6(32'hb73a889b),
	.w7(32'hb6fb8d8a),
	.w8(32'h375f4013),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34174552),
	.w1(32'h36f2b49f),
	.w2(32'h37ca96c1),
	.w3(32'h364ea8ad),
	.w4(32'hb789165b),
	.w5(32'h3748822d),
	.w6(32'h3787ebfc),
	.w7(32'hb7aece90),
	.w8(32'h38211e0d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a0dc0d),
	.w1(32'hb63da29e),
	.w2(32'hb5841738),
	.w3(32'h37e64d6a),
	.w4(32'hb7a53f78),
	.w5(32'hb75df72b),
	.w6(32'hb6d80d48),
	.w7(32'hb7ae362e),
	.w8(32'hb71ccf59),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b0f7ea),
	.w1(32'h36aaacba),
	.w2(32'h3517c890),
	.w3(32'hb797e91f),
	.w4(32'h3703ec63),
	.w5(32'h36a92dbd),
	.w6(32'h36ef3431),
	.w7(32'hb689400b),
	.w8(32'h3460df40),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c55a6e),
	.w1(32'h371a73d7),
	.w2(32'h38258e94),
	.w3(32'h367be737),
	.w4(32'h373cc2bb),
	.w5(32'h382d4885),
	.w6(32'hb6f66733),
	.w7(32'h36f80f67),
	.w8(32'h377bdc71),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a63f3),
	.w1(32'h3941d43c),
	.w2(32'h377da063),
	.w3(32'h3994efcd),
	.w4(32'h3987f63a),
	.w5(32'h389c1e46),
	.w6(32'h38a60ad0),
	.w7(32'h39226cc3),
	.w8(32'h38f54352),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387282a4),
	.w1(32'h38ad18a3),
	.w2(32'h3875caa1),
	.w3(32'h3841b5e3),
	.w4(32'h38987b76),
	.w5(32'h377c88a1),
	.w6(32'hb8823ac2),
	.w7(32'hb878d279),
	.w8(32'hb89c003e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6888e07),
	.w1(32'hb791e0c9),
	.w2(32'h379ec617),
	.w3(32'hb87883b3),
	.w4(32'hb6c46390),
	.w5(32'h37d729c9),
	.w6(32'hb78a4792),
	.w7(32'hb7bedac4),
	.w8(32'hb54c1b89),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80db8d8),
	.w1(32'h386f1037),
	.w2(32'h3714c55a),
	.w3(32'hb8b5d585),
	.w4(32'h38b39b50),
	.w5(32'h38b7f6a1),
	.w6(32'hb9346daf),
	.w7(32'hb8ef3b96),
	.w8(32'hb75bef24),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d293f5),
	.w1(32'h35fec958),
	.w2(32'h379ca250),
	.w3(32'hb7a89cca),
	.w4(32'hb7f89f53),
	.w5(32'hb6a4a85b),
	.w6(32'hb7444ad8),
	.w7(32'hb8010d73),
	.w8(32'hb7019c58),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37367482),
	.w1(32'hb6899ea2),
	.w2(32'h3700e362),
	.w3(32'hb6bf2350),
	.w4(32'hb6046f39),
	.w5(32'hb392b882),
	.w6(32'hb70e5aea),
	.w7(32'h36021f47),
	.w8(32'hb6122228),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c8e768),
	.w1(32'hb73aaaf5),
	.w2(32'hb66b0184),
	.w3(32'h364fb1cb),
	.w4(32'hb7519d20),
	.w5(32'hb723290f),
	.w6(32'hb75ab2cc),
	.w7(32'hb72c2d5c),
	.w8(32'h3618ed14),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370976cd),
	.w1(32'h368609bd),
	.w2(32'h3705cd8a),
	.w3(32'h3688aae0),
	.w4(32'hb6cb059f),
	.w5(32'hb673720c),
	.w6(32'hb5e57236),
	.w7(32'h3667afc3),
	.w8(32'h362815e2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cc2d6),
	.w1(32'h38511d6c),
	.w2(32'h36dd3c4f),
	.w3(32'hb6fde6d9),
	.w4(32'h38212ead),
	.w5(32'hb6c4157b),
	.w6(32'hb8b72299),
	.w7(32'hb8da6f1c),
	.w8(32'hb8996db0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395262cd),
	.w1(32'h396e3ab2),
	.w2(32'h38a945e4),
	.w3(32'h3966002f),
	.w4(32'h38d65971),
	.w5(32'h381798cd),
	.w6(32'h399db829),
	.w7(32'h396ac778),
	.w8(32'h38031353),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d85480),
	.w1(32'h388c1ecd),
	.w2(32'h385fbb1b),
	.w3(32'h381e2b00),
	.w4(32'h38a07ed7),
	.w5(32'h3851e67c),
	.w6(32'hb7d90e83),
	.w7(32'h37768cf8),
	.w8(32'hb7124209),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7baaa44),
	.w1(32'hb7fef3ff),
	.w2(32'hb6bf93fa),
	.w3(32'hb81073df),
	.w4(32'hb8847a57),
	.w5(32'hb72782a1),
	.w6(32'hb7d146aa),
	.w7(32'hb7f5077c),
	.w8(32'hb6face41),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843ec07),
	.w1(32'h388a01d5),
	.w2(32'h37924174),
	.w3(32'h37348491),
	.w4(32'h37e48736),
	.w5(32'h37c0ed5e),
	.w6(32'hb86335fc),
	.w7(32'hb8a013a1),
	.w8(32'hb8aa396c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7487375),
	.w1(32'h3776f69b),
	.w2(32'hb6cf006e),
	.w3(32'h37f42958),
	.w4(32'h383926e1),
	.w5(32'h37a8363e),
	.w6(32'hb8b76458),
	.w7(32'hb8025279),
	.w8(32'hb75b9259),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9111fcc),
	.w1(32'hb933825c),
	.w2(32'hb8d42724),
	.w3(32'hb8c47515),
	.w4(32'hb86e5f09),
	.w5(32'h3788048c),
	.w6(32'hb9345cb1),
	.w7(32'hb84db291),
	.w8(32'hb7869b7c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb762940f),
	.w1(32'h361cbc6d),
	.w2(32'h36691988),
	.w3(32'hb7f357ab),
	.w4(32'hb2d62ff9),
	.w5(32'h36f5eaf6),
	.w6(32'hb5868948),
	.w7(32'hb65c8562),
	.w8(32'h370147ee),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fa9eb9),
	.w1(32'hb699a62e),
	.w2(32'h358aca5e),
	.w3(32'h36b315b3),
	.w4(32'hb6f5e539),
	.w5(32'hb6484193),
	.w6(32'hb5c681c2),
	.w7(32'hb6c2da96),
	.w8(32'hb6a54442),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38956b1f),
	.w1(32'h38c4da4a),
	.w2(32'h38a27db1),
	.w3(32'h36822161),
	.w4(32'hb7dc3bca),
	.w5(32'h37d3245c),
	.w6(32'h3892dd43),
	.w7(32'h3748b6c8),
	.w8(32'h37f023fb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904125f),
	.w1(32'h38e1b397),
	.w2(32'h3878fc1b),
	.w3(32'h389bf97d),
	.w4(32'h38d0de32),
	.w5(32'h3764bf69),
	.w6(32'hb820ecde),
	.w7(32'h3749f2c4),
	.w8(32'h36f82312),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3253e),
	.w1(32'h386d5260),
	.w2(32'h3810d25f),
	.w3(32'h38191f70),
	.w4(32'h38a8a468),
	.w5(32'h34612642),
	.w6(32'hb82c0763),
	.w7(32'hb832b24a),
	.w8(32'hb87b253c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b52366),
	.w1(32'h380d5c03),
	.w2(32'h36a57103),
	.w3(32'h37b25172),
	.w4(32'h377e09f9),
	.w5(32'h36d39851),
	.w6(32'h377b4731),
	.w7(32'h366079f4),
	.w8(32'hb6c0777c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36152ad1),
	.w1(32'h37050327),
	.w2(32'h36dac959),
	.w3(32'h36ab76f3),
	.w4(32'h35e57b65),
	.w5(32'hb5de9782),
	.w6(32'h368afd05),
	.w7(32'h36d65b20),
	.w8(32'hb64cf53d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3625abfd),
	.w1(32'h35cb1a1d),
	.w2(32'hb6805a8b),
	.w3(32'h3638f505),
	.w4(32'h369247b8),
	.w5(32'hb6c144eb),
	.w6(32'h36aaa805),
	.w7(32'hb666c0ca),
	.w8(32'hb6581122),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa2d2e),
	.w1(32'h366565db),
	.w2(32'h3889743e),
	.w3(32'hb81215e8),
	.w4(32'hb8020855),
	.w5(32'h383c72ef),
	.w6(32'hb714bd1f),
	.w7(32'hb77f9764),
	.w8(32'h37cb86db),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b0a3a),
	.w1(32'h377a7fa6),
	.w2(32'hb98f950b),
	.w3(32'h3916950e),
	.w4(32'h38e56cb8),
	.w5(32'hb8a646bb),
	.w6(32'hb93e84f1),
	.w7(32'hb90d8e8f),
	.w8(32'hb7aab8e6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387808e2),
	.w1(32'h3893885e),
	.w2(32'h384d5e04),
	.w3(32'h37e8f078),
	.w4(32'h388ce3b7),
	.w5(32'h37f5fba4),
	.w6(32'h3882f315),
	.w7(32'h388f8ed0),
	.w8(32'h380c0cb4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b953d9),
	.w1(32'h37311359),
	.w2(32'h3865800b),
	.w3(32'hb8481174),
	.w4(32'hb8a09c1d),
	.w5(32'hb83665fb),
	.w6(32'h383320da),
	.w7(32'hb8214e55),
	.w8(32'hb6fe4f43),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78356a4),
	.w1(32'hb7bb1695),
	.w2(32'hb60c6efb),
	.w3(32'hb860f26c),
	.w4(32'hb8a0a821),
	.w5(32'hb7f7f5e6),
	.w6(32'hb84f1e68),
	.w7(32'hb893b3fd),
	.w8(32'hb832ae19),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76390ed),
	.w1(32'h356d2ca4),
	.w2(32'h36d9e075),
	.w3(32'hb7edb276),
	.w4(32'hb716a9fd),
	.w5(32'hb71e1f71),
	.w6(32'h360a40fc),
	.w7(32'h35b149af),
	.w8(32'h363f5f64),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365312a1),
	.w1(32'hb7f11dcc),
	.w2(32'hb720b026),
	.w3(32'hb6851d3c),
	.w4(32'hb78d34f2),
	.w5(32'hb70d37a6),
	.w6(32'hb7b72924),
	.w7(32'hb6ea9c1b),
	.w8(32'hb72ea153),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c4fa8),
	.w1(32'hb4c6be9f),
	.w2(32'hb7170c5d),
	.w3(32'hb7a189e7),
	.w4(32'hb7e872fd),
	.w5(32'hb616c305),
	.w6(32'hb69abee0),
	.w7(32'hb68eacac),
	.w8(32'h36d5f96c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bb97ac),
	.w1(32'h370bd907),
	.w2(32'h3780e06c),
	.w3(32'hb721a51a),
	.w4(32'hb729e393),
	.w5(32'h36cc2664),
	.w6(32'hb6dd5009),
	.w7(32'hb78caa82),
	.w8(32'hb62115d3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797df88),
	.w1(32'hb6f22445),
	.w2(32'hb68d97e8),
	.w3(32'hb706f609),
	.w4(32'hb77130f3),
	.w5(32'h36c11c13),
	.w6(32'hb5b19bec),
	.w7(32'hb6a6babb),
	.w8(32'h3769db0d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881c02e),
	.w1(32'h38972625),
	.w2(32'hb6dd38d8),
	.w3(32'hb6e3f81d),
	.w4(32'h38e71f3b),
	.w5(32'h35e15385),
	.w6(32'hb867587a),
	.w7(32'hb837878e),
	.w8(32'hb6f46778),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3d06978),
	.w1(32'hb79aaca9),
	.w2(32'h38046b2b),
	.w3(32'hb69dcf95),
	.w4(32'h37939c8c),
	.w5(32'h38254cec),
	.w6(32'hb8695d1f),
	.w7(32'h3653305f),
	.w8(32'hb8a3bff8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7518b98),
	.w1(32'hb77448f7),
	.w2(32'hb5784524),
	.w3(32'h35ca3afa),
	.w4(32'h358731fb),
	.w5(32'h37c12f9f),
	.w6(32'hb5982a22),
	.w7(32'hb7caf809),
	.w8(32'hb6c076f4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38630eee),
	.w1(32'h38045166),
	.w2(32'h34b08d13),
	.w3(32'hb3897f62),
	.w4(32'h38025663),
	.w5(32'h382ccfb4),
	.w6(32'hb88cba79),
	.w7(32'hb7c4053a),
	.w8(32'h38318533),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38832fcf),
	.w1(32'h3837c63e),
	.w2(32'h381b8f5e),
	.w3(32'h3851ee09),
	.w4(32'h3844e14e),
	.w5(32'h37372b53),
	.w6(32'hb5f55f1e),
	.w7(32'h37ae5458),
	.w8(32'hb71c5631),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3694fef5),
	.w1(32'hb6eefd24),
	.w2(32'hb65e468e),
	.w3(32'hb655c201),
	.w4(32'hb73ec184),
	.w5(32'hb6e4a096),
	.w6(32'hb76f1a33),
	.w7(32'hb5dce76d),
	.w8(32'hb65c29f4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8523de0),
	.w1(32'hb82903c3),
	.w2(32'hb6bc4ea9),
	.w3(32'hb88dd747),
	.w4(32'hb753c6f7),
	.w5(32'h386b66a0),
	.w6(32'hb8c84185),
	.w7(32'hb855d28f),
	.w8(32'h386798f7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3665ea2b),
	.w1(32'h36d40e9f),
	.w2(32'h3777ffaf),
	.w3(32'h35de826d),
	.w4(32'hb6527439),
	.w5(32'h35a48925),
	.w6(32'hb5187b9b),
	.w7(32'hb6430b85),
	.w8(32'h371a3160),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37176d41),
	.w1(32'h36ed7c1f),
	.w2(32'h377a4207),
	.w3(32'hb68b4afe),
	.w4(32'hb6d86e82),
	.w5(32'h3528638a),
	.w6(32'h359d478f),
	.w7(32'h373d07ee),
	.w8(32'h3706e90b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3762e631),
	.w1(32'hb719eeb6),
	.w2(32'hb65deb55),
	.w3(32'h36953eab),
	.w4(32'hb73d4df4),
	.w5(32'hb6d1a7f4),
	.w6(32'hb744c8d1),
	.w7(32'h35177658),
	.w8(32'hb684e622),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362021fc),
	.w1(32'h37ab710d),
	.w2(32'h3690a5a8),
	.w3(32'h35ed9a92),
	.w4(32'h3737b181),
	.w5(32'hb583094a),
	.w6(32'h3781e8ca),
	.w7(32'hb71f263c),
	.w8(32'h369ea01b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb871469f),
	.w1(32'hb8329413),
	.w2(32'hb6745184),
	.w3(32'hb8888f25),
	.w4(32'hb80dbebf),
	.w5(32'h37905752),
	.w6(32'hb8296883),
	.w7(32'hb80750f1),
	.w8(32'hb3089833),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcb3e7),
	.w1(32'h38fb0e97),
	.w2(32'h37959010),
	.w3(32'h38bb78f9),
	.w4(32'h393059d3),
	.w5(32'h38341600),
	.w6(32'hb818f3b0),
	.w7(32'h3789552d),
	.w8(32'h37e4dd8b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f1279),
	.w1(32'h378b9f25),
	.w2(32'hb68fb6c2),
	.w3(32'h3780f7d0),
	.w4(32'h380dd8dd),
	.w5(32'h36f36773),
	.w6(32'hb8c3c400),
	.w7(32'hb85f0337),
	.w8(32'h36065e40),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37993394),
	.w1(32'h3796de16),
	.w2(32'hb58a1e23),
	.w3(32'h3805c9b0),
	.w4(32'h38719329),
	.w5(32'h379b45d2),
	.w6(32'hb84aeb06),
	.w7(32'h364af730),
	.w8(32'hb7653624),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eadf98),
	.w1(32'hb629eaaa),
	.w2(32'h3784c959),
	.w3(32'hb61bffea),
	.w4(32'hb7c5cb1f),
	.w5(32'hb60352a0),
	.w6(32'h371afdda),
	.w7(32'h3726375b),
	.w8(32'h375ec808),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b0209),
	.w1(32'hb746ef24),
	.w2(32'hb696f095),
	.w3(32'h360e07bb),
	.w4(32'hb78d13bf),
	.w5(32'hb7229c69),
	.w6(32'hb78c94f9),
	.w7(32'h345cdcb5),
	.w8(32'hb6b4f96b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ad3135),
	.w1(32'hb72772bf),
	.w2(32'hb4adea10),
	.w3(32'h36430e24),
	.w4(32'hb6c12c7b),
	.w5(32'hb5dfda0a),
	.w6(32'hb719e6b5),
	.w7(32'h36b6697f),
	.w8(32'h3617ac5f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36785016),
	.w1(32'hb74ddb24),
	.w2(32'hb638b695),
	.w3(32'h3595f0d0),
	.w4(32'hb71c7343),
	.w5(32'hb690a21e),
	.w6(32'hb76a6fc8),
	.w7(32'h36267d93),
	.w8(32'h35830a4a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39321f9d),
	.w1(32'h38663096),
	.w2(32'hb7e2f169),
	.w3(32'h390cf006),
	.w4(32'h3910638a),
	.w5(32'hb86d4f2f),
	.w6(32'h361c732b),
	.w7(32'h3730e588),
	.w8(32'hb7990cb1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dcaf08),
	.w1(32'h3621e1dc),
	.w2(32'h37aa545c),
	.w3(32'hb74d91cc),
	.w4(32'hb6cf5e07),
	.w5(32'h379a25cb),
	.w6(32'hb6b8877d),
	.w7(32'h35c1a425),
	.w8(32'hb729bb9c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb639c2c2),
	.w1(32'hb871b404),
	.w2(32'hb801dcd8),
	.w3(32'hb73c54a3),
	.w4(32'hb8ae9f71),
	.w5(32'hb7345b28),
	.w6(32'hb7bbc659),
	.w7(32'hb7144dc9),
	.w8(32'hb712e185),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73a92c7),
	.w1(32'hb82ab75b),
	.w2(32'hb7aa3f3b),
	.w3(32'hb7a39dbf),
	.w4(32'hb82fc4c0),
	.w5(32'hb7a7c8cc),
	.w6(32'hb7a939d9),
	.w7(32'hb7cf31e3),
	.w8(32'hb7e35c83),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74ac4d5),
	.w1(32'hb677d4af),
	.w2(32'h36c385a5),
	.w3(32'hb7b09baa),
	.w4(32'hb68945bf),
	.w5(32'h36058281),
	.w6(32'hb73ffa55),
	.w7(32'h3665da47),
	.w8(32'h36c3a0e1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378525e7),
	.w1(32'hb7c3512c),
	.w2(32'hb78b327d),
	.w3(32'h3727f066),
	.w4(32'h3610354d),
	.w5(32'h37513de3),
	.w6(32'hb777c7ed),
	.w7(32'hb82fbf45),
	.w8(32'h36366561),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c639e3),
	.w1(32'hb74b3f20),
	.w2(32'h34d7608e),
	.w3(32'hb6316c36),
	.w4(32'hb68ab5a5),
	.w5(32'h343cf283),
	.w6(32'hb6e3d685),
	.w7(32'h36b59d80),
	.w8(32'h36e91630),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842d6fa),
	.w1(32'h382a73ac),
	.w2(32'h36d35f4b),
	.w3(32'h38311836),
	.w4(32'h37e5b9cd),
	.w5(32'hb48b18f9),
	.w6(32'h3824032a),
	.w7(32'h3806e6d7),
	.w8(32'h37d1db63),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363ada2b),
	.w1(32'h3a3db288),
	.w2(32'h3b21bd8d),
	.w3(32'h35e740c9),
	.w4(32'h39965345),
	.w5(32'h3b06e4d6),
	.w6(32'hb6b11efa),
	.w7(32'h3a9318eb),
	.w8(32'h3a419f94),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bcc06),
	.w1(32'hb94e7aa4),
	.w2(32'hba28bb5d),
	.w3(32'h3a1339ac),
	.w4(32'hba3cf12d),
	.w5(32'hba8b7892),
	.w6(32'hb954946b),
	.w7(32'hba3dd0be),
	.w8(32'hb9c7ae2e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule