module layer_10_featuremap_508(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eb552),
	.w1(32'h3bc38a3e),
	.w2(32'h3c91079e),
	.w3(32'hbaf42b26),
	.w4(32'h3bac02b3),
	.w5(32'h3b25e6c7),
	.w6(32'hbba3068b),
	.w7(32'hbc49bd91),
	.w8(32'h3bfc6cb0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939bf06),
	.w1(32'hb98db1cd),
	.w2(32'h3c7cb775),
	.w3(32'hbc12eed2),
	.w4(32'hbc7eff9b),
	.w5(32'h3b9b2149),
	.w6(32'h3bc773de),
	.w7(32'hbd3173bc),
	.w8(32'hbc4aa2bc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a69e6),
	.w1(32'h3c045200),
	.w2(32'hbcb0f300),
	.w3(32'h3bf6efac),
	.w4(32'h3c51d924),
	.w5(32'h3abc8aa4),
	.w6(32'hbb26664f),
	.w7(32'hbc42cec0),
	.w8(32'h3c2da885),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c927527),
	.w1(32'hbb1785d3),
	.w2(32'hbb1b80aa),
	.w3(32'h3be10606),
	.w4(32'hbb853c65),
	.w5(32'h3987ab95),
	.w6(32'hbb4601fa),
	.w7(32'hbc9cdb18),
	.w8(32'h3c27cb17),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe07dba),
	.w1(32'hbcb38aed),
	.w2(32'h3c2eb058),
	.w3(32'hbb4b47fa),
	.w4(32'h3d005dc6),
	.w5(32'hbae14dcf),
	.w6(32'h3bf290b4),
	.w7(32'hbba657b3),
	.w8(32'hbbd71876),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2120bc),
	.w1(32'h3b39e9a7),
	.w2(32'hbc2dbfdc),
	.w3(32'h3c637788),
	.w4(32'h38ba3483),
	.w5(32'h3a41dbc3),
	.w6(32'h3b358415),
	.w7(32'h3c90dad1),
	.w8(32'hbcd87cdc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c27d7),
	.w1(32'h3b8c666e),
	.w2(32'hbc0a819d),
	.w3(32'hbc6bcd97),
	.w4(32'h3b46e557),
	.w5(32'hbb764761),
	.w6(32'hbb738bc4),
	.w7(32'hbbd2c87d),
	.w8(32'h3bf3120c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3f2d),
	.w1(32'h3b879500),
	.w2(32'h3b90a69a),
	.w3(32'hbc1a6940),
	.w4(32'hbc65105f),
	.w5(32'h3ae4d753),
	.w6(32'hbc2874e4),
	.w7(32'hbc151a6e),
	.w8(32'h3c56c2b0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade0640),
	.w1(32'h3aa8e4ae),
	.w2(32'hbc02c3f6),
	.w3(32'hbbe1fd1c),
	.w4(32'hbcc3bbcd),
	.w5(32'h3b2696db),
	.w6(32'h3bba1a1f),
	.w7(32'h3c0935b2),
	.w8(32'hba34000a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2aa6b),
	.w1(32'h3bca10ab),
	.w2(32'h3c3aded8),
	.w3(32'h3aa72fa2),
	.w4(32'h3bcd75b0),
	.w5(32'hbb0254dc),
	.w6(32'hbc06d32d),
	.w7(32'h3ae628be),
	.w8(32'h3ce22299),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef52d),
	.w1(32'hbb99423e),
	.w2(32'h3d11d3d8),
	.w3(32'hbc69db4e),
	.w4(32'hbb54432b),
	.w5(32'hba9ea3f7),
	.w6(32'hba0fd683),
	.w7(32'hbca22d5b),
	.w8(32'h3a997872),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28a610),
	.w1(32'hbbcd5421),
	.w2(32'h3b941d12),
	.w3(32'hbc2986ed),
	.w4(32'hba4e72e6),
	.w5(32'h3bb2ce38),
	.w6(32'hba463f23),
	.w7(32'h3a327cb8),
	.w8(32'hbcf75d49),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bab28),
	.w1(32'h3bf2404e),
	.w2(32'h3d08675b),
	.w3(32'h3ced765f),
	.w4(32'h3d045af2),
	.w5(32'hbc8c01d2),
	.w6(32'h3b32c090),
	.w7(32'h3c47e34b),
	.w8(32'hbb671a10),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb2001),
	.w1(32'h3a9edeeb),
	.w2(32'hbb041148),
	.w3(32'h3bc1cb28),
	.w4(32'h3ba443a9),
	.w5(32'h3b3248f4),
	.w6(32'hbbbae67b),
	.w7(32'hbc149ce7),
	.w8(32'hbba38187),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c940695),
	.w1(32'h3c8622e0),
	.w2(32'h3b8310ce),
	.w3(32'h3c0278ac),
	.w4(32'hbb2195fe),
	.w5(32'h3c1e2d4d),
	.w6(32'hbc83ed70),
	.w7(32'hbcb98e16),
	.w8(32'h3c4ed9b8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49a9a1),
	.w1(32'h3ba32710),
	.w2(32'hbbdb9916),
	.w3(32'h3aac6809),
	.w4(32'h3a02bcad),
	.w5(32'hbaf48126),
	.w6(32'hbb885af7),
	.w7(32'h3b8b6960),
	.w8(32'hbaddcacf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094ae5),
	.w1(32'h396c3f78),
	.w2(32'h3c7352fd),
	.w3(32'h3b9ff7eb),
	.w4(32'h3a11a555),
	.w5(32'hbbe5ddcc),
	.w6(32'hbabfc2c2),
	.w7(32'hbbdafab1),
	.w8(32'h3bf29398),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2af5c),
	.w1(32'hbc41e4b1),
	.w2(32'hbc522019),
	.w3(32'hbc3bd216),
	.w4(32'h3a98bf61),
	.w5(32'hbc0e97fa),
	.w6(32'hbcbd7fc7),
	.w7(32'hbc6e94a6),
	.w8(32'hbc803e7d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10b4d4),
	.w1(32'hbb6ed34c),
	.w2(32'hbc1dd31e),
	.w3(32'hbc0496df),
	.w4(32'hbc2520c1),
	.w5(32'hbb43b50f),
	.w6(32'hbc1fc9e9),
	.w7(32'hbc68f79c),
	.w8(32'h3c1e0479),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeab1a),
	.w1(32'hbb0fad96),
	.w2(32'h3acc1450),
	.w3(32'hbaa21d8e),
	.w4(32'hbbb70583),
	.w5(32'hb90a4b52),
	.w6(32'h3b0a9def),
	.w7(32'h3a03dc42),
	.w8(32'h3b382f04),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60346b),
	.w1(32'hbb6d63ad),
	.w2(32'hbb7b813f),
	.w3(32'h3a94cf14),
	.w4(32'hbb7e0a1e),
	.w5(32'h3c0ae8e2),
	.w6(32'hbc107d73),
	.w7(32'h3c20832c),
	.w8(32'h3bf4dee9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ea9bd),
	.w1(32'h3c359c6f),
	.w2(32'h3cba2382),
	.w3(32'h3b4115cc),
	.w4(32'hb9a5d3fb),
	.w5(32'hbb843d4a),
	.w6(32'hbb55a7a5),
	.w7(32'hba924646),
	.w8(32'h3c11010e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbeea4),
	.w1(32'hbc881c06),
	.w2(32'hbb65ff68),
	.w3(32'h3b57a751),
	.w4(32'h3c39822f),
	.w5(32'h3bee03f6),
	.w6(32'hbc517c51),
	.w7(32'hbc720798),
	.w8(32'h3c099527),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aadc7),
	.w1(32'h3add9919),
	.w2(32'h3a1d861f),
	.w3(32'hbc4147f4),
	.w4(32'h3daf62bb),
	.w5(32'h3cd1a8e8),
	.w6(32'hbcb7ad73),
	.w7(32'h3bba5102),
	.w8(32'hbc7213ca),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab131),
	.w1(32'hbbc93506),
	.w2(32'hbc611816),
	.w3(32'hbc65a52a),
	.w4(32'h3ba3ab65),
	.w5(32'hbc039a08),
	.w6(32'h3bb99379),
	.w7(32'hbb70c7e2),
	.w8(32'hbc9f2fee),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bcefd),
	.w1(32'hbaef0180),
	.w2(32'hbc9aea4e),
	.w3(32'hbad1bf05),
	.w4(32'hbcd9f441),
	.w5(32'h3c5482a8),
	.w6(32'h3a0d2992),
	.w7(32'h3c342122),
	.w8(32'hbb192991),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccdb24),
	.w1(32'h3bb8964e),
	.w2(32'hbc5c2f94),
	.w3(32'hbc0999bb),
	.w4(32'hbb8a008c),
	.w5(32'hbb33c6bb),
	.w6(32'h3bb18572),
	.w7(32'hbbbbb81d),
	.w8(32'h3b061bd8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7da6c0),
	.w1(32'h3bf5c0bb),
	.w2(32'h3b6487fe),
	.w3(32'h3c9a306b),
	.w4(32'hbb8970a6),
	.w5(32'hbb7dd0ef),
	.w6(32'hbb08c9e8),
	.w7(32'hbc076611),
	.w8(32'hbae17bea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d0829),
	.w1(32'hbbc76449),
	.w2(32'hbb4ebddd),
	.w3(32'h3d525304),
	.w4(32'hbb59e445),
	.w5(32'hbb95bd59),
	.w6(32'hbac49ce5),
	.w7(32'hbb2a18e5),
	.w8(32'hb7ed22ad),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6c609),
	.w1(32'h3be3d621),
	.w2(32'hbbfd08b1),
	.w3(32'h3cd1e828),
	.w4(32'h3c39809d),
	.w5(32'hba4d0b9c),
	.w6(32'h3c5c4f71),
	.w7(32'h3c601c8b),
	.w8(32'hbb481508),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4c1d),
	.w1(32'hbb21f026),
	.w2(32'hbc2b3720),
	.w3(32'h3c44a5e7),
	.w4(32'h3c0c7090),
	.w5(32'h3bc5223d),
	.w6(32'hbc8b893b),
	.w7(32'h3c531c67),
	.w8(32'h391cd37c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d31c0),
	.w1(32'hbc324c40),
	.w2(32'hbcbc5628),
	.w3(32'h3cccafb5),
	.w4(32'hbb94715d),
	.w5(32'hbb9ce36a),
	.w6(32'hb9c84fe2),
	.w7(32'h3cb1c04f),
	.w8(32'h3c369626),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b589e22),
	.w1(32'hbc0b6f97),
	.w2(32'h3c4751cb),
	.w3(32'hbb17e1fb),
	.w4(32'hbc906688),
	.w5(32'hbb075883),
	.w6(32'hbbf3468a),
	.w7(32'h3b6ab407),
	.w8(32'hbc86a56a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6fdd),
	.w1(32'h3bba22c9),
	.w2(32'h3be6e4a0),
	.w3(32'hbc39022d),
	.w4(32'h3bf92115),
	.w5(32'hb920ad42),
	.w6(32'h3b944b2b),
	.w7(32'hbb5605ca),
	.w8(32'h3ab3a104),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1625f0),
	.w1(32'hbb09ba71),
	.w2(32'hbb426e51),
	.w3(32'h3aa83e83),
	.w4(32'hbcc83659),
	.w5(32'h3bffab57),
	.w6(32'h3b57029d),
	.w7(32'hbc2e664e),
	.w8(32'h3b9fadb4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ff83a),
	.w1(32'h3b464ecf),
	.w2(32'h397da8d5),
	.w3(32'h3b327f9f),
	.w4(32'hbbff9ab5),
	.w5(32'hbac3d792),
	.w6(32'h3c6a8472),
	.w7(32'hbc875464),
	.w8(32'h3b669055),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d2a16),
	.w1(32'hbb4fdf8f),
	.w2(32'h3bf4f0f1),
	.w3(32'hbc0a7a7d),
	.w4(32'hbc01588e),
	.w5(32'h3b897735),
	.w6(32'hbc3b6be5),
	.w7(32'h39e374b5),
	.w8(32'h3c25b932),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9755bba),
	.w1(32'hbbd7436e),
	.w2(32'h3b8a3366),
	.w3(32'h3b21fbda),
	.w4(32'hbc1b68f7),
	.w5(32'h3c56c45b),
	.w6(32'h3b2ad608),
	.w7(32'hbc02b333),
	.w8(32'hbb08dc93),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f7ac9),
	.w1(32'hbb3da37b),
	.w2(32'h3abe08be),
	.w3(32'hbbf2b9fb),
	.w4(32'h3c08ce15),
	.w5(32'hbbb8b60b),
	.w6(32'hbb186ead),
	.w7(32'hbc7e5f9f),
	.w8(32'hbbb77afc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d4eae),
	.w1(32'hbb6b07de),
	.w2(32'hbc17954a),
	.w3(32'hba821175),
	.w4(32'hbc1e3b94),
	.w5(32'h3bc0a8c3),
	.w6(32'hbc09ab64),
	.w7(32'h3c523862),
	.w8(32'h3b299589),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba4188),
	.w1(32'hbbd2fdbf),
	.w2(32'hba1e92f5),
	.w3(32'h3bf6c883),
	.w4(32'hbca57e07),
	.w5(32'h3c5c18ce),
	.w6(32'h3b6dca19),
	.w7(32'h3b7bb0cb),
	.w8(32'h3af217f8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf68d99),
	.w1(32'hbbc77069),
	.w2(32'h3d031cbc),
	.w3(32'hbb246983),
	.w4(32'hbc8aaf18),
	.w5(32'hbb9c0c61),
	.w6(32'hbcf75680),
	.w7(32'hba805b10),
	.w8(32'hbc2535dd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8edb96),
	.w1(32'h398bce67),
	.w2(32'h3c26b17a),
	.w3(32'hbc0b249f),
	.w4(32'h3c2f3f10),
	.w5(32'hbbc4c140),
	.w6(32'h3c501626),
	.w7(32'h3c193d20),
	.w8(32'hbc391934),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8403),
	.w1(32'h3c0f1499),
	.w2(32'hbba16c8e),
	.w3(32'hbb38980e),
	.w4(32'h3b71eabd),
	.w5(32'h3aa660cb),
	.w6(32'hbb85a6e0),
	.w7(32'h3b3fb97e),
	.w8(32'h3b65933f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf55b8),
	.w1(32'hbba8423b),
	.w2(32'h3b6be0a9),
	.w3(32'hb9c6008a),
	.w4(32'h3b323858),
	.w5(32'hba38fb1c),
	.w6(32'hbb661550),
	.w7(32'h3b95f6c6),
	.w8(32'h3b411c21),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89aed7),
	.w1(32'h3bc85b2c),
	.w2(32'hbb9f36ba),
	.w3(32'hbb800748),
	.w4(32'h3cc2f730),
	.w5(32'h3ae65be8),
	.w6(32'hbc3ad0ad),
	.w7(32'hb7c87384),
	.w8(32'hbc64da0e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c4d1),
	.w1(32'hbad3f9a1),
	.w2(32'hbb4c050a),
	.w3(32'hbc88bc03),
	.w4(32'h3bf2bba0),
	.w5(32'hbb82c30b),
	.w6(32'hbbd19b2e),
	.w7(32'hbc88218d),
	.w8(32'hbb222b2f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7fab),
	.w1(32'hbc86cbf0),
	.w2(32'hbc975caa),
	.w3(32'hbbd88056),
	.w4(32'h3b9de560),
	.w5(32'hbc1d02c9),
	.w6(32'hbd93ca10),
	.w7(32'hbc25ef23),
	.w8(32'hbc1e5ba1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc24df9),
	.w1(32'hbb019f28),
	.w2(32'hbc87b92f),
	.w3(32'h3b9abb3d),
	.w4(32'hbbc8fa7e),
	.w5(32'hbc14059e),
	.w6(32'hbb7f315a),
	.w7(32'h3a9002a5),
	.w8(32'h39759723),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddf7e2),
	.w1(32'hbb822092),
	.w2(32'hbc275aca),
	.w3(32'hbb70ac2a),
	.w4(32'hbbb4faa5),
	.w5(32'h3ccb06b3),
	.w6(32'h3c9ec3ef),
	.w7(32'h3b0360fb),
	.w8(32'h38c51db7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a854a),
	.w1(32'h3c3406b8),
	.w2(32'h3bc81f30),
	.w3(32'hbbcf428f),
	.w4(32'hbc4a800b),
	.w5(32'hbad3c84d),
	.w6(32'hbc18e9c1),
	.w7(32'hbc0b8b03),
	.w8(32'h3b978cdf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb97161),
	.w1(32'hbc280d50),
	.w2(32'hbc1f0169),
	.w3(32'h3b8cde31),
	.w4(32'hbb22f3b6),
	.w5(32'hbc215b5f),
	.w6(32'hbbd96cd5),
	.w7(32'h3b8511cf),
	.w8(32'h39f73573),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4af30),
	.w1(32'h38fa2837),
	.w2(32'hba9a1b17),
	.w3(32'hbbfd3ffa),
	.w4(32'h3ba19f5b),
	.w5(32'hbb9059f3),
	.w6(32'hbc26d241),
	.w7(32'hbc29f73b),
	.w8(32'hbd244c02),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861789),
	.w1(32'hbb4e9e70),
	.w2(32'hbc4daf24),
	.w3(32'hbc88a6bd),
	.w4(32'hbc21caa5),
	.w5(32'hbc4d8bef),
	.w6(32'hba1d73e1),
	.w7(32'hbc84898e),
	.w8(32'hbb03e96b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b591e0d),
	.w1(32'h3ab66240),
	.w2(32'hbb59858b),
	.w3(32'h3c0c6160),
	.w4(32'h3c18cd4f),
	.w5(32'h3ca3f28a),
	.w6(32'hbc413d17),
	.w7(32'hbc42ba0f),
	.w8(32'hbbfcc048),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e8c67),
	.w1(32'hbb0094b9),
	.w2(32'h3bf4307a),
	.w3(32'hbba97fb1),
	.w4(32'hbd1b49e2),
	.w5(32'h3c299c5c),
	.w6(32'hba7e39eb),
	.w7(32'hbc853585),
	.w8(32'h3c7e2588),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35fb8d),
	.w1(32'hbbb198eb),
	.w2(32'h3b05286a),
	.w3(32'hbceaf27d),
	.w4(32'hbceaa11a),
	.w5(32'h3acd8074),
	.w6(32'hba077c0a),
	.w7(32'h3b0a76bf),
	.w8(32'hbc759de4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64660d),
	.w1(32'hbc4bb428),
	.w2(32'hbc717d1b),
	.w3(32'h397f5e5b),
	.w4(32'h3b805c30),
	.w5(32'hbc22152b),
	.w6(32'h3ba28b08),
	.w7(32'hbb0e7f6c),
	.w8(32'hbc3eeccf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf3815e),
	.w1(32'h3c3fdc41),
	.w2(32'h3c2afa06),
	.w3(32'h3b8232da),
	.w4(32'hbcf1881d),
	.w5(32'h3a6b52b9),
	.w6(32'h3c3080c7),
	.w7(32'h3b7fb5dd),
	.w8(32'h3cfd47db),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2dd9),
	.w1(32'hba30cd2f),
	.w2(32'hbcad5f74),
	.w3(32'hbb99e7db),
	.w4(32'hbba4d7cd),
	.w5(32'h3c8507d0),
	.w6(32'hbad1384f),
	.w7(32'hba11ce50),
	.w8(32'h3bc49045),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507b32),
	.w1(32'hbae25fee),
	.w2(32'hbc254716),
	.w3(32'hbca3e8b3),
	.w4(32'hbc82d008),
	.w5(32'hbd07d6b7),
	.w6(32'hba1e8dd0),
	.w7(32'hbbc2d2bc),
	.w8(32'h3cbdec2e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38be82),
	.w1(32'h3bea03b0),
	.w2(32'hbb7344c1),
	.w3(32'hbbcd9569),
	.w4(32'hbad057f3),
	.w5(32'hbb8e940b),
	.w6(32'hbc25acbf),
	.w7(32'h3a5d79c4),
	.w8(32'h3c208068),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca185a0),
	.w1(32'h3b331f6f),
	.w2(32'hbafd5ceb),
	.w3(32'h3af1896c),
	.w4(32'h3b281a70),
	.w5(32'hbc9ecebe),
	.w6(32'h3bdd1f05),
	.w7(32'h3c30dd40),
	.w8(32'h3c37edcf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102bc4),
	.w1(32'hbc00ef50),
	.w2(32'h3b8d8b66),
	.w3(32'h3b2c5f20),
	.w4(32'h3d0a8e1b),
	.w5(32'hbc07b6ca),
	.w6(32'hbc817f13),
	.w7(32'hbb616647),
	.w8(32'h3d6da28c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e0d4),
	.w1(32'h3b8169ef),
	.w2(32'hbb2965c7),
	.w3(32'hbc714e96),
	.w4(32'hbc917db4),
	.w5(32'hbc189505),
	.w6(32'h3b636c3d),
	.w7(32'h3c993c7e),
	.w8(32'hbb177f50),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc02dc2),
	.w1(32'hbc5acc95),
	.w2(32'hb9ad0244),
	.w3(32'h3b4c3f02),
	.w4(32'hbc8b17a3),
	.w5(32'hbc50e74f),
	.w6(32'h39489cd1),
	.w7(32'h3c065ec0),
	.w8(32'hbbc5829f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8007e3),
	.w1(32'h3b8f37f0),
	.w2(32'h3c73e6bc),
	.w3(32'hbb1abd3f),
	.w4(32'hbad217ae),
	.w5(32'hbd4ec5b3),
	.w6(32'h3c2f39da),
	.w7(32'hbb97501e),
	.w8(32'h3c35b75d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9ff38),
	.w1(32'h3bdf1c4d),
	.w2(32'hb92c2848),
	.w3(32'h3b3db704),
	.w4(32'hbad7fa9b),
	.w5(32'h3933f806),
	.w6(32'h380ea63d),
	.w7(32'h3b89e613),
	.w8(32'h3a8689eb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc612d31),
	.w1(32'hbc13df37),
	.w2(32'hbb76a225),
	.w3(32'h3c695aae),
	.w4(32'hbbbc5b2b),
	.w5(32'hbcac4856),
	.w6(32'h398f98fa),
	.w7(32'hbc9d6c54),
	.w8(32'hbc67a57c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8671dd),
	.w1(32'h3b85c115),
	.w2(32'hbc47c9cc),
	.w3(32'hbc06b027),
	.w4(32'h3ca14e1c),
	.w5(32'h3c36ff33),
	.w6(32'hbc8d62c8),
	.w7(32'hbc00ea4d),
	.w8(32'hb8d70889),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb000fb),
	.w1(32'hbb7fb0f2),
	.w2(32'hbc24e133),
	.w3(32'h3b8dc3d3),
	.w4(32'h3b541b00),
	.w5(32'hbb37302c),
	.w6(32'h3c0c496b),
	.w7(32'h3ad710ae),
	.w8(32'h3ccdae4b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae8a0),
	.w1(32'hbc02db31),
	.w2(32'hbc4e2fdf),
	.w3(32'h3b8e3a74),
	.w4(32'hbcd78006),
	.w5(32'hbbe031fc),
	.w6(32'hbc429599),
	.w7(32'h3c1b2300),
	.w8(32'hbbd009a2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb96739),
	.w1(32'hb8ede80f),
	.w2(32'h3bb02285),
	.w3(32'h3bbd37f8),
	.w4(32'h3b7eef56),
	.w5(32'hbb27ac8b),
	.w6(32'hbbf15331),
	.w7(32'hbc426b3e),
	.w8(32'h3c62cfcf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d6ae),
	.w1(32'hb8c746da),
	.w2(32'h3abd8f72),
	.w3(32'h3bace4f1),
	.w4(32'hbbf87c27),
	.w5(32'hbc4d4b34),
	.w6(32'hbade03c2),
	.w7(32'hbb92ea3a),
	.w8(32'hbb4f28f2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc357a71),
	.w1(32'hbbd8d1a9),
	.w2(32'hbb1e13a7),
	.w3(32'hbc0226f5),
	.w4(32'hbbe8455d),
	.w5(32'h3a84c36d),
	.w6(32'h3a932ae9),
	.w7(32'hba87d3ab),
	.w8(32'hbb727343),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0485),
	.w1(32'h3b8197ab),
	.w2(32'hbc0f4c0c),
	.w3(32'h393e8754),
	.w4(32'hbbdb20b8),
	.w5(32'h3b567207),
	.w6(32'hbb8e1595),
	.w7(32'hbaccdd47),
	.w8(32'hbc0d1ef5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce5b4),
	.w1(32'hbc911ca1),
	.w2(32'hbb47a204),
	.w3(32'h3c7ff632),
	.w4(32'hbb8cc2b2),
	.w5(32'hb991322c),
	.w6(32'hbc9bf87a),
	.w7(32'hbb90321f),
	.w8(32'hbd016eea),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2871c1),
	.w1(32'hbb9a6bc8),
	.w2(32'hbc6f75c5),
	.w3(32'hba99d83e),
	.w4(32'h3c97970b),
	.w5(32'h3c5aa310),
	.w6(32'h3ad828a6),
	.w7(32'h3b6d4e86),
	.w8(32'h3b84d2c2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb397473),
	.w1(32'h3b98559c),
	.w2(32'hbbe6acc8),
	.w3(32'hbad00583),
	.w4(32'hbb620ec1),
	.w5(32'hbc821cb7),
	.w6(32'h38022d90),
	.w7(32'h3c3fe42f),
	.w8(32'h3a88532c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7cb92),
	.w1(32'hb9cfd776),
	.w2(32'hbc915aca),
	.w3(32'hbb827baa),
	.w4(32'h3bfa7bd5),
	.w5(32'h3c7e7a08),
	.w6(32'hbc1eb5dc),
	.w7(32'h3be096d0),
	.w8(32'h3c5da8c6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc091b7d),
	.w1(32'h3ce8d0f5),
	.w2(32'hb915bc0b),
	.w3(32'h3c007c62),
	.w4(32'h3bf23d57),
	.w5(32'hbb48665f),
	.w6(32'h3c127f5d),
	.w7(32'h3cb21184),
	.w8(32'h3c0704a9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceb764e),
	.w1(32'hbb8c6770),
	.w2(32'h3a43fc2d),
	.w3(32'h3c5dbf24),
	.w4(32'hbbecfaeb),
	.w5(32'h3c01f08b),
	.w6(32'hbbcb7fea),
	.w7(32'hbbc60eeb),
	.w8(32'hbbb05e2a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39265f3d),
	.w1(32'h3c8277f6),
	.w2(32'h3c1202e7),
	.w3(32'hbc3ec77c),
	.w4(32'h3ac49e6e),
	.w5(32'h3b4ef74c),
	.w6(32'h3cf2a39b),
	.w7(32'hbc9d35bd),
	.w8(32'h3c5ca0c2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccba19a),
	.w1(32'h3b155bb6),
	.w2(32'h3aeb8e56),
	.w3(32'hbc130f99),
	.w4(32'hbc7e78ab),
	.w5(32'hb945b12d),
	.w6(32'h3bcdba0f),
	.w7(32'hbc01a36e),
	.w8(32'hbb048170),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fe329),
	.w1(32'hbb212627),
	.w2(32'h3b984c31),
	.w3(32'h3aa4b0f4),
	.w4(32'h3b7b57eb),
	.w5(32'hbaedea04),
	.w6(32'hb9aed75e),
	.w7(32'h3a5abac7),
	.w8(32'h3b7edfe1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6a9285),
	.w1(32'h3cc9b8c7),
	.w2(32'hba7396c8),
	.w3(32'h3b57e3b9),
	.w4(32'hbb2ddaeb),
	.w5(32'h3b230ccb),
	.w6(32'hbbf7fe48),
	.w7(32'hbbe53a0d),
	.w8(32'hba3030eb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4476),
	.w1(32'h3c83e298),
	.w2(32'h3bf9413e),
	.w3(32'h3d00056a),
	.w4(32'hbb351dca),
	.w5(32'h3b3f74d1),
	.w6(32'h3c67138f),
	.w7(32'hbb9ef63d),
	.w8(32'h3b72a8a3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09200d),
	.w1(32'hbb6301b0),
	.w2(32'h3c6fa49c),
	.w3(32'hbb8eb540),
	.w4(32'h3d008b09),
	.w5(32'hbc2dd79a),
	.w6(32'hbc3b8e02),
	.w7(32'h3c7754b2),
	.w8(32'hb995380d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97ecef),
	.w1(32'h3cd30e5e),
	.w2(32'hbb8087ef),
	.w3(32'h3a37dd12),
	.w4(32'h3c901bf8),
	.w5(32'hbb2fe5bc),
	.w6(32'h3c138d91),
	.w7(32'h3b85f65c),
	.w8(32'hbb4e0ac6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40615b),
	.w1(32'hbab7572b),
	.w2(32'hbb526bc0),
	.w3(32'hbb24afdc),
	.w4(32'hbc45de93),
	.w5(32'h3d574fa6),
	.w6(32'hbc7b6a74),
	.w7(32'h3c1316c7),
	.w8(32'hbb90dfae),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e9913),
	.w1(32'h3b81e23b),
	.w2(32'h3bb7a8b9),
	.w3(32'h3ab07e6d),
	.w4(32'h3ab7f5de),
	.w5(32'hb98b1ccb),
	.w6(32'hbbc0c409),
	.w7(32'h3b9b9091),
	.w8(32'h3bc76d26),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc469ce),
	.w1(32'hbc42cf63),
	.w2(32'hbb8bd2cb),
	.w3(32'hbc6ede88),
	.w4(32'hbc52f5c9),
	.w5(32'hbc46fccd),
	.w6(32'hbbd961aa),
	.w7(32'hbbe710ab),
	.w8(32'hbb853fec),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb26e6),
	.w1(32'h3c261f58),
	.w2(32'h3b737961),
	.w3(32'hbb8af79b),
	.w4(32'h3b5a8c5a),
	.w5(32'h3b2be86a),
	.w6(32'hb978cd6f),
	.w7(32'hbbc620c6),
	.w8(32'hbb089e11),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e9a0),
	.w1(32'hbc094367),
	.w2(32'hbc5d3c08),
	.w3(32'hbb49313a),
	.w4(32'h3c10ee30),
	.w5(32'h3bcaa59c),
	.w6(32'hbc72082f),
	.w7(32'hbbd1e368),
	.w8(32'h3b41a996),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9f754),
	.w1(32'h3c30d9b7),
	.w2(32'hbb9e81bd),
	.w3(32'hbba34ddb),
	.w4(32'h3c2b567d),
	.w5(32'hbb8d5679),
	.w6(32'h3bbb1848),
	.w7(32'hbba63a39),
	.w8(32'h3b86e3e5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90ea9f),
	.w1(32'hbb68795c),
	.w2(32'hba57b523),
	.w3(32'hbb1858ac),
	.w4(32'h3c1b7f1a),
	.w5(32'hbbf3af7c),
	.w6(32'h3a07cde3),
	.w7(32'h3c11e779),
	.w8(32'hbb902872),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cee28),
	.w1(32'hbbaaf1ac),
	.w2(32'h391b937f),
	.w3(32'h3c10fc23),
	.w4(32'h3afc063c),
	.w5(32'hbb9c2e1b),
	.w6(32'h3c6bca1c),
	.w7(32'h3b08f157),
	.w8(32'hb9621961),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62e0d6),
	.w1(32'h3c19ce7a),
	.w2(32'h3b89be01),
	.w3(32'h3bc3e5d4),
	.w4(32'h3bd84ffa),
	.w5(32'h3ba8cefa),
	.w6(32'hbcb85837),
	.w7(32'h3cb37215),
	.w8(32'hbacfe618),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f26e),
	.w1(32'h3ad5f410),
	.w2(32'h3b0578f5),
	.w3(32'hbc9ab064),
	.w4(32'hbc06031e),
	.w5(32'hbb879755),
	.w6(32'hbcaaac0a),
	.w7(32'hbb61e16c),
	.w8(32'hbc81b74c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f768),
	.w1(32'h3d2de5b9),
	.w2(32'hbb143905),
	.w3(32'hbbf7c6f8),
	.w4(32'hbc2489d2),
	.w5(32'hbc05fa6a),
	.w6(32'hbc1727b8),
	.w7(32'hbb8dda9c),
	.w8(32'h3b83aade),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0ce0),
	.w1(32'hbbe4ae3f),
	.w2(32'h3c8ada4a),
	.w3(32'hbc2e3c63),
	.w4(32'hbc1136fb),
	.w5(32'h3c48f73f),
	.w6(32'h38a803a2),
	.w7(32'hbab93bae),
	.w8(32'h3b5b84f3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5ec5),
	.w1(32'h3b034f9b),
	.w2(32'h3bdc5011),
	.w3(32'hbba013b4),
	.w4(32'h3c295df4),
	.w5(32'h3bd215d1),
	.w6(32'h3b0e5ce6),
	.w7(32'h3c3ebae3),
	.w8(32'hbba5641f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192c64),
	.w1(32'h3bc4fe53),
	.w2(32'hbbd3f732),
	.w3(32'hbc83a2b9),
	.w4(32'hbc401e5f),
	.w5(32'hbb44eefc),
	.w6(32'hbc2e17b6),
	.w7(32'h3ac87532),
	.w8(32'hbbb1a8dd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce8a46),
	.w1(32'h3c82ebc1),
	.w2(32'hbbda5413),
	.w3(32'h3b81363c),
	.w4(32'hbc0339ec),
	.w5(32'hbae0e66c),
	.w6(32'hbb9200a9),
	.w7(32'h3bff0b57),
	.w8(32'hbba308dd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81463),
	.w1(32'hbc6854c1),
	.w2(32'hbca1ec80),
	.w3(32'h3c24b701),
	.w4(32'hbc9250d6),
	.w5(32'hbc0932d4),
	.w6(32'hbc2f9e2d),
	.w7(32'hbc77c5f1),
	.w8(32'hbaa7c507),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bc6cc),
	.w1(32'h3c645390),
	.w2(32'h3c2fdabb),
	.w3(32'h3c2736d3),
	.w4(32'hbc26d5cb),
	.w5(32'hba81f8cb),
	.w6(32'h3b13f453),
	.w7(32'hbbc1592f),
	.w8(32'h3bbe773d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe14512),
	.w1(32'h3c3b9c3c),
	.w2(32'hb9f67838),
	.w3(32'hbc9e1405),
	.w4(32'h3b8fe35a),
	.w5(32'h3bd312a1),
	.w6(32'h3b3efed5),
	.w7(32'hbb9e7a58),
	.w8(32'hb91bd6e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb80f9),
	.w1(32'h3c8f32df),
	.w2(32'h3b2354d5),
	.w3(32'h3a07d588),
	.w4(32'h3c027653),
	.w5(32'h3aefcfcc),
	.w6(32'h3b45ca8e),
	.w7(32'h3b3b7924),
	.w8(32'hba9e7e1a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8fac),
	.w1(32'h3b6b590d),
	.w2(32'h3c1690a8),
	.w3(32'hbc8869eb),
	.w4(32'h39c4de57),
	.w5(32'h3c253d06),
	.w6(32'hbb05ec43),
	.w7(32'h3cbdb71d),
	.w8(32'h3d120173),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0294c),
	.w1(32'h3b9042a0),
	.w2(32'hba3ae077),
	.w3(32'hbb88b16f),
	.w4(32'hbaa07d38),
	.w5(32'h3c08b0b8),
	.w6(32'h3baab7b8),
	.w7(32'h3a409132),
	.w8(32'hbaab1074),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d59d),
	.w1(32'hbb7bf900),
	.w2(32'hbb01ba81),
	.w3(32'h3bb73a5b),
	.w4(32'h3b061b00),
	.w5(32'hbbb2c450),
	.w6(32'hbbd85596),
	.w7(32'hbc412c0d),
	.w8(32'h3cdc40e1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71aeee),
	.w1(32'h3be7e657),
	.w2(32'h3c893ca4),
	.w3(32'hbb417108),
	.w4(32'h3ae719e5),
	.w5(32'hb90e9da9),
	.w6(32'hbba1fbba),
	.w7(32'h3b220a78),
	.w8(32'hbac09830),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e4b71),
	.w1(32'h3b8fe079),
	.w2(32'hbb3d3fcb),
	.w3(32'hb9dde53b),
	.w4(32'hb9f7099c),
	.w5(32'hbb85de25),
	.w6(32'hbbf83c21),
	.w7(32'hbc137713),
	.w8(32'hbb3a328f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe018b1),
	.w1(32'hbc11d97b),
	.w2(32'hbb6cfb67),
	.w3(32'hbac1fc32),
	.w4(32'hba7cd9ef),
	.w5(32'hbbaae3c1),
	.w6(32'h3cd16c7f),
	.w7(32'h3b367542),
	.w8(32'hbc67d894),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c26a2),
	.w1(32'hbca4caa1),
	.w2(32'hbc016e9e),
	.w3(32'hbb54fd9d),
	.w4(32'hbc4fe3c4),
	.w5(32'h3b5a119b),
	.w6(32'h3bb398fc),
	.w7(32'h3ae01256),
	.w8(32'h3c40d8f6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73902c),
	.w1(32'h3c0197e4),
	.w2(32'h3c63d5a5),
	.w3(32'hbb9020db),
	.w4(32'h3c0a65b4),
	.w5(32'hbc2a71b8),
	.w6(32'h39d9be6b),
	.w7(32'hbc3f9f97),
	.w8(32'hbc28884f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e59dc7),
	.w1(32'h3b6b128c),
	.w2(32'hbba86258),
	.w3(32'h3aa0eeb1),
	.w4(32'hbc4bd528),
	.w5(32'h3b5af60d),
	.w6(32'hb98c3389),
	.w7(32'h3b51ffa1),
	.w8(32'h3c96dfa3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068414),
	.w1(32'h3baa7e75),
	.w2(32'hb96d8021),
	.w3(32'hbc29e558),
	.w4(32'hbba1afa0),
	.w5(32'h3c512ad6),
	.w6(32'h3cd7e975),
	.w7(32'hbcaace9b),
	.w8(32'hbb8d251d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e2e64),
	.w1(32'hb956f698),
	.w2(32'h3b687a59),
	.w3(32'hbb4c7c55),
	.w4(32'hbc331772),
	.w5(32'hbce25f74),
	.w6(32'hbb358e0a),
	.w7(32'h3b4193ab),
	.w8(32'hbc56ecd6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc220bc6),
	.w1(32'h386f69f6),
	.w2(32'hbbbd244a),
	.w3(32'h3bcb8b6d),
	.w4(32'hbc39ef11),
	.w5(32'h3c8327b8),
	.w6(32'h3b1adaee),
	.w7(32'h3c680e78),
	.w8(32'h3cd15546),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d70d2),
	.w1(32'h3bb4fb56),
	.w2(32'hba62200d),
	.w3(32'hba20e319),
	.w4(32'hbbd4c121),
	.w5(32'hbc0f9aab),
	.w6(32'hbc3e13ca),
	.w7(32'h3b589457),
	.w8(32'hbbb052aa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f2c5),
	.w1(32'h3ae0b230),
	.w2(32'h3cbab410),
	.w3(32'hbbebac4a),
	.w4(32'hbbe72b75),
	.w5(32'hba8c6e50),
	.w6(32'hbb829af7),
	.w7(32'hb994fc22),
	.w8(32'hbb5c0f10),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa901b),
	.w1(32'h3bd1be0c),
	.w2(32'h3b6cbd32),
	.w3(32'h3c2d2569),
	.w4(32'hbc91f944),
	.w5(32'h3ba81277),
	.w6(32'h3cdb59af),
	.w7(32'h3a70c7ed),
	.w8(32'hbc49eda5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc520c6d),
	.w1(32'h3ab77c26),
	.w2(32'h3ba9f448),
	.w3(32'h39718ec5),
	.w4(32'hbb015cc9),
	.w5(32'h3aadaa6c),
	.w6(32'h3c363fda),
	.w7(32'h3cfbdeee),
	.w8(32'h3aef2176),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bede11f),
	.w1(32'hbc05715d),
	.w2(32'hbbb7961e),
	.w3(32'hbb588d8d),
	.w4(32'hbc32faee),
	.w5(32'hbbd25469),
	.w6(32'hbb4e87c4),
	.w7(32'hba7edd1a),
	.w8(32'h3ba62546),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba018fa4),
	.w1(32'h39c82759),
	.w2(32'hba0407fd),
	.w3(32'hbad62204),
	.w4(32'h3bb22cef),
	.w5(32'h398c9d80),
	.w6(32'h39f88243),
	.w7(32'hba1353f5),
	.w8(32'hbb9f4e2e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43288),
	.w1(32'hbc054653),
	.w2(32'h3c12b2be),
	.w3(32'hbaa5c6ac),
	.w4(32'h3d01b501),
	.w5(32'h3b8e101b),
	.w6(32'h39a97b53),
	.w7(32'h3c357ea1),
	.w8(32'h3b41acdf),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bfbcc),
	.w1(32'hba69b778),
	.w2(32'h3cf89ec1),
	.w3(32'h3b698036),
	.w4(32'h3bb4245e),
	.w5(32'hbb230deb),
	.w6(32'h3b5e7906),
	.w7(32'hbc4d6768),
	.w8(32'hbc8126a0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32b936),
	.w1(32'h3bac9818),
	.w2(32'hbc0aa37d),
	.w3(32'h3c8cc68b),
	.w4(32'hbb91fde6),
	.w5(32'hbb33597d),
	.w6(32'hbaa92816),
	.w7(32'h3956b8b8),
	.w8(32'hbb756aac),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbca57f),
	.w1(32'hbbfd0d57),
	.w2(32'h3af58cf9),
	.w3(32'hbb454ab5),
	.w4(32'hbb0e25f0),
	.w5(32'h3af6b0f6),
	.w6(32'h3ab155ed),
	.w7(32'h3bfc896f),
	.w8(32'hbc1a4b28),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4aca41),
	.w1(32'h3b08339c),
	.w2(32'hbb8e0817),
	.w3(32'h3beceffd),
	.w4(32'hbc385636),
	.w5(32'h3c259fca),
	.w6(32'hbae3d5a6),
	.w7(32'hbc6a3bba),
	.w8(32'hbc548891),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66bdd2),
	.w1(32'h3babfbb5),
	.w2(32'hbb67ee2b),
	.w3(32'hb8694364),
	.w4(32'hbb889dd2),
	.w5(32'h3b7b58e8),
	.w6(32'hbb84edb0),
	.w7(32'h3c10d2ea),
	.w8(32'hbb743aef),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2240e5),
	.w1(32'hbc57cbd5),
	.w2(32'h3986b20b),
	.w3(32'h3b2cde1e),
	.w4(32'hbb27f164),
	.w5(32'h3c0b567c),
	.w6(32'hb9fa1d81),
	.w7(32'hbccae0bf),
	.w8(32'h3c97419e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda7e1a),
	.w1(32'h3acd6414),
	.w2(32'hbb9551eb),
	.w3(32'h3c1c29ae),
	.w4(32'h3a46c69f),
	.w5(32'h3b41f92f),
	.w6(32'hbb281e86),
	.w7(32'hbb7392d0),
	.w8(32'hbbe1251f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4996a7),
	.w1(32'h3ae36c5e),
	.w2(32'h3c85f7f2),
	.w3(32'hbc423f57),
	.w4(32'h3a38f548),
	.w5(32'h3a58b0f8),
	.w6(32'hb94b29ee),
	.w7(32'hbc1d1eff),
	.w8(32'h3c2dc5dd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09c408),
	.w1(32'h3b7e91a3),
	.w2(32'hbc02fa80),
	.w3(32'h3c6ab125),
	.w4(32'h3c1fe202),
	.w5(32'h3c105be5),
	.w6(32'h3c006fad),
	.w7(32'h3c0d810a),
	.w8(32'h3bb3d839),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa3460),
	.w1(32'hbce3ff81),
	.w2(32'h3be68846),
	.w3(32'hbb198072),
	.w4(32'h3b9c8f38),
	.w5(32'h3b850090),
	.w6(32'hbc1a356a),
	.w7(32'hbb58e0b0),
	.w8(32'h3b77f4a5),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dfaad),
	.w1(32'hba2466bf),
	.w2(32'hbb47edec),
	.w3(32'h3b8e1518),
	.w4(32'hbbe4d4d1),
	.w5(32'hbbfaae51),
	.w6(32'hbc6a6a09),
	.w7(32'hbcd15152),
	.w8(32'hbc11276a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d9acc),
	.w1(32'h3a7663fe),
	.w2(32'hbc00d388),
	.w3(32'h3b97c98e),
	.w4(32'hbb0b76e6),
	.w5(32'hbaaf5c3b),
	.w6(32'hbd0af18c),
	.w7(32'hbb8d3f1a),
	.w8(32'h3cc75639),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e9bd),
	.w1(32'h3b05fa0b),
	.w2(32'hbc3100cb),
	.w3(32'hb805ccb2),
	.w4(32'h3b9cd3ea),
	.w5(32'h3b36d949),
	.w6(32'hbbcb5df6),
	.w7(32'h3c039771),
	.w8(32'hbb3a2a24),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb51f77),
	.w1(32'h39bf10fe),
	.w2(32'hba0d9895),
	.w3(32'hba7a9b5e),
	.w4(32'hbbe26a88),
	.w5(32'h3bd20276),
	.w6(32'h3ba7e183),
	.w7(32'h3b806397),
	.w8(32'hbc7da7b2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409f10),
	.w1(32'hbc349568),
	.w2(32'h3c063505),
	.w3(32'hbb061c65),
	.w4(32'hbb84de8f),
	.w5(32'hbc9eeaf0),
	.w6(32'h3c66193c),
	.w7(32'h3c1d2bb9),
	.w8(32'h3b9d175c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b14b1),
	.w1(32'hbc4fe969),
	.w2(32'hb99894a5),
	.w3(32'h3bde0b47),
	.w4(32'h3b75612e),
	.w5(32'h3bc21ab8),
	.w6(32'h3b818097),
	.w7(32'h3c59766d),
	.w8(32'h3b5ab265),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9792f),
	.w1(32'h3ba33d91),
	.w2(32'h3c98c85d),
	.w3(32'hbc32bea9),
	.w4(32'h3b3d6c23),
	.w5(32'h3c19bd94),
	.w6(32'h3c02e6a3),
	.w7(32'h3c4bb3f3),
	.w8(32'h3c0e2b95),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d388),
	.w1(32'h3d3a53a2),
	.w2(32'hbb40b4ee),
	.w3(32'h3b88460a),
	.w4(32'hbbd7afe2),
	.w5(32'h3adc599d),
	.w6(32'hbc930e60),
	.w7(32'hbc4fb066),
	.w8(32'h3c057be4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f1b7),
	.w1(32'h3c4d8076),
	.w2(32'hba0a3cad),
	.w3(32'h3c1d6ea6),
	.w4(32'h3c9ee372),
	.w5(32'hbc71cfbf),
	.w6(32'hbcec78dc),
	.w7(32'hbbf5a642),
	.w8(32'hbc3f9917),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f34b8),
	.w1(32'hbbc64139),
	.w2(32'hbbe34aa8),
	.w3(32'h3ce0a592),
	.w4(32'hbc721a1b),
	.w5(32'h3c694367),
	.w6(32'h3ba88b73),
	.w7(32'hba354f46),
	.w8(32'hbc20d6ad),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d1924),
	.w1(32'hbc529026),
	.w2(32'hbcb07f27),
	.w3(32'h3af57f13),
	.w4(32'h3beb9daa),
	.w5(32'hbc810473),
	.w6(32'hbc101128),
	.w7(32'h3cd40560),
	.w8(32'hbb638055),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc8a13),
	.w1(32'hbc0c040b),
	.w2(32'h3b5556c6),
	.w3(32'hbc2d6e13),
	.w4(32'h3c09f43c),
	.w5(32'h3c487312),
	.w6(32'h3c3c9c44),
	.w7(32'hbcd52f32),
	.w8(32'h3c57533a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1910ea),
	.w1(32'hbb8de57d),
	.w2(32'h3c708ca6),
	.w3(32'hbbc63f07),
	.w4(32'h3d05bfa8),
	.w5(32'hbb22388f),
	.w6(32'h3d5539f5),
	.w7(32'h3c0e93a5),
	.w8(32'h3c1da9cc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca9c5a),
	.w1(32'hb7deac1e),
	.w2(32'h3b82133d),
	.w3(32'hbd095f41),
	.w4(32'h3bce7ed4),
	.w5(32'h3a6e41e6),
	.w6(32'h3c1fbf03),
	.w7(32'h3c41ccc8),
	.w8(32'hbbdf458b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af91c48),
	.w1(32'hbc92f9aa),
	.w2(32'hba9e81b8),
	.w3(32'hbba75915),
	.w4(32'hbbd8546e),
	.w5(32'hbc2c1ce5),
	.w6(32'hb957d764),
	.w7(32'hbcac9b13),
	.w8(32'hbc76a179),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2ddb),
	.w1(32'h3c8130f2),
	.w2(32'hbb790bb0),
	.w3(32'hbc7806d3),
	.w4(32'hbc27cde7),
	.w5(32'h3b956cb8),
	.w6(32'hbc0ef221),
	.w7(32'hbb83e4f2),
	.w8(32'h3993ecab),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c8563),
	.w1(32'hbc65e0f4),
	.w2(32'hbb87f342),
	.w3(32'h3b12ac4a),
	.w4(32'hbc74167d),
	.w5(32'h3adb055c),
	.w6(32'h3bef2e21),
	.w7(32'hbbbe51bb),
	.w8(32'hbbbe1919),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28613d),
	.w1(32'hbc3a37aa),
	.w2(32'hbb8dab01),
	.w3(32'h3b7f1a4c),
	.w4(32'h3c9cfe14),
	.w5(32'h3b90227f),
	.w6(32'h3c1ecb59),
	.w7(32'hbbdc0ae2),
	.w8(32'h3bda25ca),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d98a),
	.w1(32'h3c3f4e46),
	.w2(32'h3ba0ee39),
	.w3(32'hbc702a7c),
	.w4(32'hbbc8bef1),
	.w5(32'hbb57ae65),
	.w6(32'h3c3ed9ae),
	.w7(32'h3c966a9c),
	.w8(32'h3c054c51),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce4ec2),
	.w1(32'h3b150428),
	.w2(32'hbbd1c0f9),
	.w3(32'hbc3ea504),
	.w4(32'h3c7a50be),
	.w5(32'hbbb7e762),
	.w6(32'h3c8b6ba7),
	.w7(32'h3c79e2a9),
	.w8(32'h3b113ca1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3073),
	.w1(32'h3b7ea1ab),
	.w2(32'h3b94a949),
	.w3(32'hbbc286ca),
	.w4(32'h3c420e67),
	.w5(32'h3b7d5381),
	.w6(32'hbc4e019d),
	.w7(32'h3b78532f),
	.w8(32'hbb4b4a39),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee912),
	.w1(32'h3be84eb2),
	.w2(32'h39b263f0),
	.w3(32'h3bd91c7b),
	.w4(32'hbc3070c9),
	.w5(32'hbc70ceff),
	.w6(32'hbc460261),
	.w7(32'hbbcb6799),
	.w8(32'hbbe37d98),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b06a),
	.w1(32'hbc1f10f7),
	.w2(32'hbbacc850),
	.w3(32'hbc14e33a),
	.w4(32'h3b5796b3),
	.w5(32'hbc2b4412),
	.w6(32'hbbccc3a1),
	.w7(32'h3b4662ae),
	.w8(32'hbcaed8cb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cf01e),
	.w1(32'h3b91ccda),
	.w2(32'h3aee0c80),
	.w3(32'hbc2d891c),
	.w4(32'h3cc31889),
	.w5(32'h3b23b83c),
	.w6(32'h3c8f2fe3),
	.w7(32'hbbdbcfb1),
	.w8(32'hbc021bc5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09409),
	.w1(32'hbc911d2f),
	.w2(32'h3a59ce3a),
	.w3(32'hbc468c31),
	.w4(32'hbc028147),
	.w5(32'h3c900b0c),
	.w6(32'h3ac138fa),
	.w7(32'hbc2c020b),
	.w8(32'hbc05b339),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cca6e),
	.w1(32'h3be8d6a6),
	.w2(32'hbbc4051f),
	.w3(32'h3c943707),
	.w4(32'hbae77a39),
	.w5(32'hbb9fd4b4),
	.w6(32'hbcef0912),
	.w7(32'hbb59e725),
	.w8(32'h3a4b040b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc23882),
	.w1(32'hbc739ad9),
	.w2(32'hbb337295),
	.w3(32'hbb6a8140),
	.w4(32'h3c82c968),
	.w5(32'hbacc4371),
	.w6(32'h39f76f7e),
	.w7(32'hbc9ab0b3),
	.w8(32'h3c845621),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2adfec),
	.w1(32'hbc742340),
	.w2(32'h3b384191),
	.w3(32'hbc1055f6),
	.w4(32'hba3abda1),
	.w5(32'h3c5e765c),
	.w6(32'hbc99e414),
	.w7(32'hbc92ab97),
	.w8(32'h3c3fc6fa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c148bb5),
	.w1(32'hbbbe5abd),
	.w2(32'h3d61498c),
	.w3(32'h3bfc17a9),
	.w4(32'h3cdfe359),
	.w5(32'h3cfb976d),
	.w6(32'hbbb97d0f),
	.w7(32'h3b9a6af7),
	.w8(32'hba581fd5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83be22),
	.w1(32'h3ccc8678),
	.w2(32'h3bb79ab4),
	.w3(32'hbbc84ecc),
	.w4(32'hbc1b931b),
	.w5(32'hbc542c00),
	.w6(32'h3c9086a1),
	.w7(32'hba5eedd1),
	.w8(32'h3bb8d117),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95657e),
	.w1(32'hbaea05ef),
	.w2(32'h3d65a72a),
	.w3(32'h3bc49bcd),
	.w4(32'hbbb3ea05),
	.w5(32'h3c818bf4),
	.w6(32'hbc37b686),
	.w7(32'h3cd72190),
	.w8(32'h3c7cc080),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc681055),
	.w1(32'hbc71ced8),
	.w2(32'hbc29e50b),
	.w3(32'hbc73498b),
	.w4(32'hb983ea0f),
	.w5(32'hbcc8f92a),
	.w6(32'h3cfa1b33),
	.w7(32'h3c3859c2),
	.w8(32'hbc8beb3b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf4f47),
	.w1(32'h3c71b5bd),
	.w2(32'h3c93a094),
	.w3(32'h3ba1cb3f),
	.w4(32'hbc8d70ed),
	.w5(32'hbb8572eb),
	.w6(32'hba9c0e33),
	.w7(32'hbb28e909),
	.w8(32'h3c0a8cab),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae91cfd),
	.w1(32'h3c84d5af),
	.w2(32'hbc2e3731),
	.w3(32'hb9587d19),
	.w4(32'h3b79fc2f),
	.w5(32'hbac801b4),
	.w6(32'hbc431d50),
	.w7(32'hbbb2452b),
	.w8(32'hb9d7e5ea),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1470e7),
	.w1(32'hbb90a550),
	.w2(32'hbb5b549d),
	.w3(32'h3a3c4361),
	.w4(32'h3a460b93),
	.w5(32'hba864ef3),
	.w6(32'h3c7b1d87),
	.w7(32'h3b2c22ed),
	.w8(32'hba97b95c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0f349),
	.w1(32'h3bdbd6a9),
	.w2(32'h3c9a2a7d),
	.w3(32'hbc64c2d8),
	.w4(32'hbb918725),
	.w5(32'hbbbf8a34),
	.w6(32'hbd07df23),
	.w7(32'h3b96d14e),
	.w8(32'hbb1d98ee),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde2767),
	.w1(32'hbb962701),
	.w2(32'h3beae060),
	.w3(32'hbb8fcb8f),
	.w4(32'hbb7b3575),
	.w5(32'hbc89cfa7),
	.w6(32'hbc4e7090),
	.w7(32'hbb4752c7),
	.w8(32'hbd04588c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a6ae4),
	.w1(32'h3aaea515),
	.w2(32'hbc67bfff),
	.w3(32'hbbe1ed6a),
	.w4(32'h3c38e005),
	.w5(32'hbb8034fa),
	.w6(32'hbc07e802),
	.w7(32'hbba54567),
	.w8(32'h3b2c952e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574960),
	.w1(32'hbbad9828),
	.w2(32'h3c165682),
	.w3(32'h3c003e1e),
	.w4(32'h386dcb35),
	.w5(32'hbaa13c4f),
	.w6(32'hbb807e43),
	.w7(32'hbbb5941c),
	.w8(32'h3c966c69),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd606ae),
	.w1(32'h38af50ac),
	.w2(32'hbc1dc035),
	.w3(32'h3a51efd1),
	.w4(32'h3b43b061),
	.w5(32'hbbb23247),
	.w6(32'hbb15bd86),
	.w7(32'hbc0577ec),
	.w8(32'hbc048f27),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866893),
	.w1(32'h3c2d797b),
	.w2(32'hbb414577),
	.w3(32'h3c16d4bb),
	.w4(32'h3bed7544),
	.w5(32'hbc4105dd),
	.w6(32'h3c28a4dc),
	.w7(32'h3aecdeb2),
	.w8(32'hbc14f5f7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb564b6d),
	.w1(32'h3ba1c05c),
	.w2(32'hba45b54e),
	.w3(32'hbbf5f3a8),
	.w4(32'h3b65a2c4),
	.w5(32'hbb70c4a2),
	.w6(32'hbb50338d),
	.w7(32'hbb8b58e6),
	.w8(32'hbbef06d8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a862fd5),
	.w1(32'h3cbbfeb6),
	.w2(32'hbb7eb5ae),
	.w3(32'h3ac2b956),
	.w4(32'hbaf27a47),
	.w5(32'hbb17796d),
	.w6(32'h3bb83c8e),
	.w7(32'hbc8f28bd),
	.w8(32'hbc8dfac0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc7b15),
	.w1(32'h3cafdd41),
	.w2(32'h3c264bb4),
	.w3(32'hbc419ff1),
	.w4(32'hbc24ab1d),
	.w5(32'hbc4e4054),
	.w6(32'hbc176813),
	.w7(32'hbb352410),
	.w8(32'h3cb07247),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99500c),
	.w1(32'hbbbcf444),
	.w2(32'h3acea559),
	.w3(32'h3bf0dbd0),
	.w4(32'hbb3cf36c),
	.w5(32'h3b1da306),
	.w6(32'hbc11bd6b),
	.w7(32'hba7887d1),
	.w8(32'hbbd8d2ed),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1710d),
	.w1(32'hbcc2c7fe),
	.w2(32'hbc980611),
	.w3(32'h3bc036a8),
	.w4(32'h3b4c004a),
	.w5(32'hbb1bc9c0),
	.w6(32'h38d15a3b),
	.w7(32'hbb1deabc),
	.w8(32'hbae0b0cd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990561c),
	.w1(32'h3b5fe3cf),
	.w2(32'hbbef19ee),
	.w3(32'hbc5f00b1),
	.w4(32'hbbe0fd34),
	.w5(32'h3be311e0),
	.w6(32'h3b0c513b),
	.w7(32'h3c6cbbad),
	.w8(32'hb99921e4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af63e4e),
	.w1(32'h3c7627ba),
	.w2(32'hbbd8f3ea),
	.w3(32'hbba54f77),
	.w4(32'hbb92c1e2),
	.w5(32'hbbc335e9),
	.w6(32'h3bf1f290),
	.w7(32'h3b45d8f3),
	.w8(32'h3cc84910),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de10b),
	.w1(32'h3a74bdeb),
	.w2(32'hbc96388b),
	.w3(32'hbc765e29),
	.w4(32'h398cf33e),
	.w5(32'hbc511b5b),
	.w6(32'h3b5bdaa9),
	.w7(32'h3c5c1f9f),
	.w8(32'hbb6c9935),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe42f61),
	.w1(32'h3c0c2fd1),
	.w2(32'hbac6f325),
	.w3(32'hbb8d8551),
	.w4(32'h3a6c9772),
	.w5(32'hbc77830c),
	.w6(32'hbc56c730),
	.w7(32'hbc38b66a),
	.w8(32'hbb59570c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25f2e3),
	.w1(32'h3a6754cf),
	.w2(32'h3b66f038),
	.w3(32'h3bb50b18),
	.w4(32'h3c0efc84),
	.w5(32'hbc0432d5),
	.w6(32'hba810efc),
	.w7(32'h3b3e1503),
	.w8(32'hbc5465a6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb426b03),
	.w1(32'hbb9bfb1d),
	.w2(32'h3bba8d41),
	.w3(32'hbcaef816),
	.w4(32'h39a819df),
	.w5(32'h3c079a17),
	.w6(32'h3c22937d),
	.w7(32'h3b99ea9a),
	.w8(32'hba83d2ae),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4df5a3),
	.w1(32'hbbee9058),
	.w2(32'hbad80ca2),
	.w3(32'hbb2915e7),
	.w4(32'h3c7fbc12),
	.w5(32'hbb3c2236),
	.w6(32'hbb9e739a),
	.w7(32'hbb8cca0a),
	.w8(32'hb8f26641),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96f031),
	.w1(32'h3b32e680),
	.w2(32'h3b1114bc),
	.w3(32'h3b98a060),
	.w4(32'hbb97816c),
	.w5(32'hba174a4a),
	.w6(32'h3c8874c6),
	.w7(32'hbb5b4541),
	.w8(32'hbbcd44d4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7abbf3),
	.w1(32'h3b8329cf),
	.w2(32'hbc111682),
	.w3(32'hbaa73120),
	.w4(32'h3c679685),
	.w5(32'hb9e23d32),
	.w6(32'h3c19a3ab),
	.w7(32'h3bdeb958),
	.w8(32'hbc2a7839),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26aa45),
	.w1(32'hbb8c90ae),
	.w2(32'hbc33df72),
	.w3(32'hb85a8b54),
	.w4(32'hbc4f790d),
	.w5(32'h3acb0d20),
	.w6(32'hba96c1fd),
	.w7(32'h399e7409),
	.w8(32'hbac316d4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfaf6),
	.w1(32'hbc2b2dd8),
	.w2(32'h3b4d71cd),
	.w3(32'hbb78983b),
	.w4(32'h3c2c0b40),
	.w5(32'hbb169631),
	.w6(32'h3afbc6cc),
	.w7(32'hbb87a4b7),
	.w8(32'hbc1d25c8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302e17),
	.w1(32'hbb090cf5),
	.w2(32'hbbd7b65e),
	.w3(32'h3bf9a96f),
	.w4(32'hbc498319),
	.w5(32'hbc460b9d),
	.w6(32'hbb3a8b25),
	.w7(32'h38f1d7ba),
	.w8(32'hbb6245d0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2444e1),
	.w1(32'hba53a529),
	.w2(32'h3aaeda48),
	.w3(32'h3c95b33c),
	.w4(32'h3bb30848),
	.w5(32'hbc7cbbd0),
	.w6(32'hbb7bd7d3),
	.w7(32'hbbee2133),
	.w8(32'h3c6f1c6b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99709d7),
	.w1(32'hbc55fae2),
	.w2(32'hbbbad3ab),
	.w3(32'h3b47f04c),
	.w4(32'hbc2b4963),
	.w5(32'hbc10ef0d),
	.w6(32'hbb3f604a),
	.w7(32'hbb69f081),
	.w8(32'hbb0beeb4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81b834),
	.w1(32'h3c8acb29),
	.w2(32'hbb01cf77),
	.w3(32'hbb0fc1c1),
	.w4(32'h3b36d98f),
	.w5(32'hbb879321),
	.w6(32'hbc825f83),
	.w7(32'hbbd0111e),
	.w8(32'hbbb36bff),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1eaf),
	.w1(32'h3b6c6a01),
	.w2(32'h3b9e333f),
	.w3(32'hbc27dc4f),
	.w4(32'hbb6be681),
	.w5(32'hbc33168c),
	.w6(32'h3bb7e779),
	.w7(32'h393df605),
	.w8(32'h3baaca06),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432c55),
	.w1(32'h39fb9ea6),
	.w2(32'hbc63bf34),
	.w3(32'hbb5ea561),
	.w4(32'h3bc2e8b5),
	.w5(32'hbbd98e7c),
	.w6(32'hbb2087d1),
	.w7(32'h3c2388d8),
	.w8(32'h3ccf6c65),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbdcc4),
	.w1(32'hbb03154f),
	.w2(32'hbbc55f05),
	.w3(32'h3c15a6c0),
	.w4(32'hbb883ef1),
	.w5(32'h3c466709),
	.w6(32'h3b38ea59),
	.w7(32'h3bcaf523),
	.w8(32'hbb1e76d0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d177b5),
	.w1(32'h39d36bb1),
	.w2(32'hbc6d95a5),
	.w3(32'h3b927321),
	.w4(32'h3bac173f),
	.w5(32'hbbe31413),
	.w6(32'hb9251100),
	.w7(32'hb9ae608f),
	.w8(32'hb99bbd7d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a35d),
	.w1(32'h3bfd8904),
	.w2(32'hbaff76eb),
	.w3(32'hbbeaa54b),
	.w4(32'h3b8680ee),
	.w5(32'hbba76c26),
	.w6(32'hbd35e973),
	.w7(32'hbc83d150),
	.w8(32'hbb161deb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd5656),
	.w1(32'h3c8f473f),
	.w2(32'h3c22761d),
	.w3(32'hbc5b81e9),
	.w4(32'h3b39e706),
	.w5(32'h3b33dab7),
	.w6(32'h3c0f7cf5),
	.w7(32'h3b1bc363),
	.w8(32'h3b81dc03),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7caa0),
	.w1(32'h3ab8c57c),
	.w2(32'hbbc7f885),
	.w3(32'hb9563232),
	.w4(32'h3b67a45f),
	.w5(32'h39db8d65),
	.w6(32'h3b83d086),
	.w7(32'h3b91c1d7),
	.w8(32'h3b4ed473),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52ae2),
	.w1(32'hbb9748aa),
	.w2(32'hbb9bca3a),
	.w3(32'h3bab2881),
	.w4(32'hba8d52f3),
	.w5(32'hbb532a98),
	.w6(32'hba993475),
	.w7(32'h39a944ff),
	.w8(32'hbaacb8af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4366d7),
	.w1(32'hbbdb18da),
	.w2(32'h3bdaa5d4),
	.w3(32'hbb039714),
	.w4(32'h3c95038f),
	.w5(32'h3b84fc06),
	.w6(32'h3c49c3d1),
	.w7(32'h3b3b431c),
	.w8(32'hb993fe4f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06d971),
	.w1(32'h3be5ed24),
	.w2(32'h3b89cad6),
	.w3(32'h3aecfc8e),
	.w4(32'hb9fa2f51),
	.w5(32'h3ab303fc),
	.w6(32'h3ba4090b),
	.w7(32'hbbaa94e8),
	.w8(32'hbc24abe0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c774658),
	.w1(32'h3c5d6579),
	.w2(32'h3adf2ad1),
	.w3(32'h3bfe4795),
	.w4(32'h3b7fdbfe),
	.w5(32'hbb70b26f),
	.w6(32'h3c18a5f1),
	.w7(32'hba8713c7),
	.w8(32'hbbe5619c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cd424),
	.w1(32'h3b51b00f),
	.w2(32'hbb5a26cd),
	.w3(32'h3be98337),
	.w4(32'hbbdf0068),
	.w5(32'hba6bb324),
	.w6(32'hba490061),
	.w7(32'hbbe5e153),
	.w8(32'hbb947497),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981fc4e),
	.w1(32'h3a5a552f),
	.w2(32'h389f54b8),
	.w3(32'h3b8c546a),
	.w4(32'hbbd6e7c3),
	.w5(32'h3bab91e5),
	.w6(32'h3c650a54),
	.w7(32'hbacf5ae1),
	.w8(32'h3b9dc373),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed929b),
	.w1(32'h3b65259e),
	.w2(32'h3b60ff0a),
	.w3(32'hbb1a75da),
	.w4(32'hb717e786),
	.w5(32'h3b5a5d5a),
	.w6(32'hbad17b6e),
	.w7(32'h3ae8c3f1),
	.w8(32'h3b91701f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d257e),
	.w1(32'hbb4413b6),
	.w2(32'hbad87cf5),
	.w3(32'hba028864),
	.w4(32'hbc02ccd9),
	.w5(32'hbc9338c1),
	.w6(32'hbbba68b6),
	.w7(32'hbbe45596),
	.w8(32'hb8813fca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c94926),
	.w1(32'hbbf81bcf),
	.w2(32'h3ae75e67),
	.w3(32'h3c85cee5),
	.w4(32'h3b51eb23),
	.w5(32'hbb15b20a),
	.w6(32'hbb1ae03a),
	.w7(32'h3a4264f5),
	.w8(32'hbb3941aa),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f58f),
	.w1(32'h3baf383b),
	.w2(32'h3c02ce12),
	.w3(32'h390c382c),
	.w4(32'hba291453),
	.w5(32'h3a675494),
	.w6(32'h3b8404e8),
	.w7(32'h3afc0990),
	.w8(32'hb94ed669),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc638),
	.w1(32'h3b8cf2c5),
	.w2(32'h3bf769e7),
	.w3(32'h3b5742d6),
	.w4(32'h3b7f0d94),
	.w5(32'h3c8402d7),
	.w6(32'hbbd7c2b6),
	.w7(32'h3a0cfddb),
	.w8(32'hbb7aaf6a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74a095),
	.w1(32'hbaef9555),
	.w2(32'hbbd1b5b0),
	.w3(32'h3c44db30),
	.w4(32'h3bb39478),
	.w5(32'hbbc1ab75),
	.w6(32'hbc462934),
	.w7(32'hbc01510d),
	.w8(32'hbb06bfb9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c49c3),
	.w1(32'hbb995ac6),
	.w2(32'h3b05d2ad),
	.w3(32'h3bb68150),
	.w4(32'hbbd64f96),
	.w5(32'h3b24c910),
	.w6(32'h3bf12b49),
	.w7(32'hbbc317df),
	.w8(32'h3cb67769),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9d5ed),
	.w1(32'hbc7c4a2c),
	.w2(32'hbbdc008b),
	.w3(32'hbc15ad02),
	.w4(32'hbce7fb01),
	.w5(32'hbc06c64d),
	.w6(32'hba129add),
	.w7(32'hbc0b2cae),
	.w8(32'hbc049358),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7398f),
	.w1(32'hbbb93d39),
	.w2(32'hbb95cbb5),
	.w3(32'hbc0098c2),
	.w4(32'h39b8ae33),
	.w5(32'hbb2716be),
	.w6(32'hbca70555),
	.w7(32'hbbc1e567),
	.w8(32'h3ba7530a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15aee5),
	.w1(32'h390150ae),
	.w2(32'h3b9a1502),
	.w3(32'hbc1b5963),
	.w4(32'hbc0681ae),
	.w5(32'h3a68a2d6),
	.w6(32'hba533abb),
	.w7(32'h3b649353),
	.w8(32'hbb96198d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff3d4),
	.w1(32'h3bf6612b),
	.w2(32'hbb4b5eb4),
	.w3(32'h3b851d29),
	.w4(32'hb9201629),
	.w5(32'h3c0dc5b5),
	.w6(32'h3ae5a72f),
	.w7(32'h3b4a17d6),
	.w8(32'hbc025514),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf89923),
	.w1(32'h3bfda9c2),
	.w2(32'h3c1374dd),
	.w3(32'h3b86e5a6),
	.w4(32'h3ba81ad9),
	.w5(32'hbb793df3),
	.w6(32'h3c4760cb),
	.w7(32'hbbf16fc1),
	.w8(32'hbbdb6a85),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103284),
	.w1(32'hbba2d3c2),
	.w2(32'hbbc7d628),
	.w3(32'hbb3aa194),
	.w4(32'h3aff16f6),
	.w5(32'h393e801b),
	.w6(32'h3b1bcb42),
	.w7(32'h3c9cc810),
	.w8(32'hbbf10f1c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b212f9c),
	.w1(32'hbbf14fc0),
	.w2(32'hba2ca353),
	.w3(32'hbbd7b33c),
	.w4(32'h3b532cc1),
	.w5(32'h3c566cd7),
	.w6(32'hbc3e2821),
	.w7(32'hbc46755d),
	.w8(32'h3bc584ad),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdfe00),
	.w1(32'h3b4745fc),
	.w2(32'h3b9a0ae5),
	.w3(32'h3a39f6e8),
	.w4(32'h362877a1),
	.w5(32'hbb297f05),
	.w6(32'h3be799f3),
	.w7(32'hbbcf7ed6),
	.w8(32'hbb226357),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadadb2),
	.w1(32'h3c02b909),
	.w2(32'h3c00edd2),
	.w3(32'hbbd38725),
	.w4(32'h3b084627),
	.w5(32'hbc4da963),
	.w6(32'hbaae7fd6),
	.w7(32'hbc16c1a7),
	.w8(32'h3aa1927c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28622f),
	.w1(32'hba321861),
	.w2(32'h3c0124d8),
	.w3(32'hbc65248c),
	.w4(32'hbc7ecc9d),
	.w5(32'h3abe0cd2),
	.w6(32'h3aef52a2),
	.w7(32'hbb7c2d91),
	.w8(32'h3c03b9f3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4149),
	.w1(32'h3d4395b8),
	.w2(32'h3adcf0a1),
	.w3(32'hbc77a970),
	.w4(32'hba8f566d),
	.w5(32'h3b896b35),
	.w6(32'h3a29d2ba),
	.w7(32'hbbe2009d),
	.w8(32'h3c114319),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3723b1),
	.w1(32'h3aea2aa5),
	.w2(32'hbc306178),
	.w3(32'hb9eda2bf),
	.w4(32'hb8c97840),
	.w5(32'h3bf39e6d),
	.w6(32'hbc22a4ec),
	.w7(32'h3bbdd934),
	.w8(32'hbb26584f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1a62),
	.w1(32'hbb1b46a1),
	.w2(32'hbb6cdfaa),
	.w3(32'hbb8ae2ce),
	.w4(32'hbab46a9b),
	.w5(32'h3c6ce9ee),
	.w6(32'hbcaec80c),
	.w7(32'hbbd092cc),
	.w8(32'hbc859bca),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f6fab),
	.w1(32'h3b7c7311),
	.w2(32'hba72e9cd),
	.w3(32'h3c1bbaeb),
	.w4(32'hbc1f140a),
	.w5(32'h3c2fd14d),
	.w6(32'hbbeb9a89),
	.w7(32'hbadab66b),
	.w8(32'hbb44516e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39134358),
	.w1(32'h3c10712f),
	.w2(32'hbae76540),
	.w3(32'h3b95160b),
	.w4(32'hbc0ba582),
	.w5(32'h3bcd61e9),
	.w6(32'h3be8d8c8),
	.w7(32'hbbde4bae),
	.w8(32'hbc2d80a2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dec98),
	.w1(32'h3c93ad36),
	.w2(32'hba409d0c),
	.w3(32'hbc37550a),
	.w4(32'h3a2bafcd),
	.w5(32'hbbb547b2),
	.w6(32'hbbebd40f),
	.w7(32'hba4683cd),
	.w8(32'h3cf3b42d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b2c8a),
	.w1(32'h3abb8980),
	.w2(32'hb9832b79),
	.w3(32'hbc247be3),
	.w4(32'h3b938678),
	.w5(32'hbc999de0),
	.w6(32'hbb882146),
	.w7(32'h3b39fbe0),
	.w8(32'hbb0f9485),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b27f),
	.w1(32'h3aea4d2e),
	.w2(32'h3cd5fd34),
	.w3(32'h3b973ac9),
	.w4(32'hbae955f2),
	.w5(32'hbad45e6b),
	.w6(32'h3cc6bacf),
	.w7(32'h3b6c4be7),
	.w8(32'h3c23eb3e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8ba4),
	.w1(32'h3a0845a1),
	.w2(32'h3c0c08d3),
	.w3(32'hbc1f3313),
	.w4(32'hbbf8717a),
	.w5(32'h3bdeddb9),
	.w6(32'hb95bc907),
	.w7(32'hb8ffacd9),
	.w8(32'h3aab816a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d182a),
	.w1(32'hbc8d52e2),
	.w2(32'hbbd107a6),
	.w3(32'hbad3d802),
	.w4(32'h3cc70d4e),
	.w5(32'hbc57f705),
	.w6(32'hbcb1d88b),
	.w7(32'h3b1d04ee),
	.w8(32'h3b99f6e6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f256f),
	.w1(32'h3a474718),
	.w2(32'h3c98b114),
	.w3(32'h3b8b78e4),
	.w4(32'hbbdf441b),
	.w5(32'h3a255b4c),
	.w6(32'h3b38cc15),
	.w7(32'hbc5fe408),
	.w8(32'hbb9fe026),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2921a),
	.w1(32'h3bb6a96a),
	.w2(32'h3c064344),
	.w3(32'hbacf70d3),
	.w4(32'hbbe62601),
	.w5(32'h3ba33b52),
	.w6(32'h3b75f5c7),
	.w7(32'h3c368ab5),
	.w8(32'h3c065403),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cf11),
	.w1(32'hbc8daa9c),
	.w2(32'h3b0d3072),
	.w3(32'hbb2439b3),
	.w4(32'hbc366644),
	.w5(32'hb74cca09),
	.w6(32'hbc2bdbd2),
	.w7(32'h39fe326a),
	.w8(32'hbb9b659f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2626eb),
	.w1(32'hbc235b91),
	.w2(32'hbc3752c5),
	.w3(32'h3b3779cc),
	.w4(32'hbb8e0707),
	.w5(32'hbc8aa2f8),
	.w6(32'hbc1b5aae),
	.w7(32'hbc46c286),
	.w8(32'hbb7a46ac),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb291d84),
	.w1(32'hbb208563),
	.w2(32'h3c1a8cd1),
	.w3(32'hbc2bdb2d),
	.w4(32'hbc52916c),
	.w5(32'h3b644635),
	.w6(32'hb830c0bf),
	.w7(32'hbb998b9a),
	.w8(32'h3c13262b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643aa3),
	.w1(32'hbc0aea05),
	.w2(32'h3c3dc5ec),
	.w3(32'hbb8a2831),
	.w4(32'hbb7b1f77),
	.w5(32'h3b9d8221),
	.w6(32'hbb22ea6c),
	.w7(32'h3b8323ab),
	.w8(32'h3b9a3425),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef59b),
	.w1(32'hbc461851),
	.w2(32'h3b486504),
	.w3(32'hbacf775c),
	.w4(32'hb987530c),
	.w5(32'hbbc154cf),
	.w6(32'h3a482b7c),
	.w7(32'h3c000f93),
	.w8(32'hbb39041b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80ab47),
	.w1(32'hbaa35a0a),
	.w2(32'hbbab5965),
	.w3(32'h3b26ac5a),
	.w4(32'hbac9e789),
	.w5(32'hbbf464f2),
	.w6(32'h3a4170b7),
	.w7(32'h3cb12128),
	.w8(32'hbc0f0620),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c605),
	.w1(32'h3b357d4c),
	.w2(32'h3bfe508a),
	.w3(32'hbb29c280),
	.w4(32'h3b862a53),
	.w5(32'hbb9dbfc6),
	.w6(32'hbacb5235),
	.w7(32'hb9962ff1),
	.w8(32'h3a3ca213),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a355658),
	.w1(32'h3ae5c231),
	.w2(32'hbc36ee5b),
	.w3(32'hbbe40c17),
	.w4(32'hbaae29ab),
	.w5(32'hba0e7211),
	.w6(32'h3ca302b8),
	.w7(32'h3b3f7baf),
	.w8(32'h3b06c869),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b0f03),
	.w1(32'hbb69ff68),
	.w2(32'hbb291ed3),
	.w3(32'hba262bd8),
	.w4(32'hb9dd1088),
	.w5(32'hbc254c00),
	.w6(32'h3bb7733d),
	.w7(32'hbb730780),
	.w8(32'h39d0f5e6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf29864),
	.w1(32'h3bef1d57),
	.w2(32'h3a94d914),
	.w3(32'h3b26bf67),
	.w4(32'hba84f7b7),
	.w5(32'h3bca230f),
	.w6(32'hbc0478b2),
	.w7(32'h3beea81b),
	.w8(32'hbbdbd16e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea0e7e),
	.w1(32'hbb2338be),
	.w2(32'h3cb76e32),
	.w3(32'hbc1a0ab9),
	.w4(32'h3b088b2e),
	.w5(32'hbbe467c8),
	.w6(32'h3b22202e),
	.w7(32'hbc6b4858),
	.w8(32'hbb2a1985),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87f6e5),
	.w1(32'h3b93ee9e),
	.w2(32'hbbcacf65),
	.w3(32'hbc8bd67b),
	.w4(32'hbc080e8e),
	.w5(32'hbaad163a),
	.w6(32'hbbdf5723),
	.w7(32'hbb59fdc0),
	.w8(32'hbbf97b6e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a337ed6),
	.w1(32'hbbe51283),
	.w2(32'hbc217fe4),
	.w3(32'hbba34747),
	.w4(32'hbbd9bd21),
	.w5(32'h39fda2ce),
	.w6(32'h3c834e90),
	.w7(32'hbb93c109),
	.w8(32'hbc5fa09a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc664950),
	.w1(32'h3baf0af4),
	.w2(32'hbc2bd48d),
	.w3(32'hbc0520b3),
	.w4(32'hbb954305),
	.w5(32'h3beb66eb),
	.w6(32'h3c980439),
	.w7(32'hbcb72121),
	.w8(32'hbc9cc513),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0260dc),
	.w1(32'hbb341e42),
	.w2(32'h3b0a2a69),
	.w3(32'h3bbe6049),
	.w4(32'h3d55221a),
	.w5(32'h3c8fbd73),
	.w6(32'h3a932d29),
	.w7(32'hbcdab066),
	.w8(32'h3c88877f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d2699),
	.w1(32'h3b06ea80),
	.w2(32'h3aade3b7),
	.w3(32'hbb8d9124),
	.w4(32'h3aaf9b2a),
	.w5(32'hbc0a342d),
	.w6(32'hbc0eeca0),
	.w7(32'hbbee51d6),
	.w8(32'h3d262360),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule