module layer_10_featuremap_81(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c00ac),
	.w1(32'hbbf0bf8e),
	.w2(32'hbb979869),
	.w3(32'hbb96cdd9),
	.w4(32'hbba8f339),
	.w5(32'hbb2244be),
	.w6(32'h3a25947e),
	.w7(32'hbbd89c65),
	.w8(32'hbc2407a7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ab348),
	.w1(32'hbada4d61),
	.w2(32'hba7f8b7c),
	.w3(32'h3b3bd45f),
	.w4(32'h3b680d85),
	.w5(32'h3bb87e15),
	.w6(32'hba67d909),
	.w7(32'h3b140c9e),
	.w8(32'hbb37f68d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002ba8),
	.w1(32'hbb9034d1),
	.w2(32'hbbf4d8f2),
	.w3(32'h3ca65ffe),
	.w4(32'hbc543f34),
	.w5(32'hba498855),
	.w6(32'h3c62316c),
	.w7(32'hba1664c3),
	.w8(32'hbbd847e4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ddf46),
	.w1(32'hbb74bbbd),
	.w2(32'hbaea10bc),
	.w3(32'hbbef7a78),
	.w4(32'hbb2802e4),
	.w5(32'h3ba68f30),
	.w6(32'hbb30cc11),
	.w7(32'hb9658e28),
	.w8(32'h3bd6223d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296500),
	.w1(32'hbbef5544),
	.w2(32'hbbe76038),
	.w3(32'hbb76f3f0),
	.w4(32'h3bb82dcd),
	.w5(32'h3aa5cae3),
	.w6(32'hbb938c66),
	.w7(32'h3afa0db9),
	.w8(32'hbb5dda9d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44846a),
	.w1(32'hb9b1241b),
	.w2(32'h3a0c4eb9),
	.w3(32'hbbd84eb8),
	.w4(32'hbaf0e908),
	.w5(32'hbb41059b),
	.w6(32'h3c4b54b7),
	.w7(32'h3ba39a2d),
	.w8(32'h3c764fad),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a56fad),
	.w1(32'hbb81eb31),
	.w2(32'hbaddcfe0),
	.w3(32'hbbd44f52),
	.w4(32'hb9081e57),
	.w5(32'h3ace2868),
	.w6(32'hbba055f8),
	.w7(32'hbb4624c1),
	.w8(32'hbbaa2697),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3973bb),
	.w1(32'hbbb8e3a8),
	.w2(32'h3c2cb824),
	.w3(32'h3baca9f6),
	.w4(32'hbad286e0),
	.w5(32'h3a5f8da2),
	.w6(32'h3afeb781),
	.w7(32'h3bd4649a),
	.w8(32'hbbbb784f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99bbbf),
	.w1(32'h3bf34365),
	.w2(32'h3c766857),
	.w3(32'hbb09f25b),
	.w4(32'hba805b98),
	.w5(32'hbb3c75b1),
	.w6(32'hbba1af6e),
	.w7(32'hbbd78cc5),
	.w8(32'h38d1a2a7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe1fd2),
	.w1(32'h39519ced),
	.w2(32'hbb9847c0),
	.w3(32'h3c02dae8),
	.w4(32'hbc0ba2de),
	.w5(32'hbbf764f7),
	.w6(32'hbc14189c),
	.w7(32'hbbb682db),
	.w8(32'h3c309c57),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56eef9),
	.w1(32'h3be84a6a),
	.w2(32'h3aa56f39),
	.w3(32'h3b9399d9),
	.w4(32'h3b643bfa),
	.w5(32'hbbc598d7),
	.w6(32'h3a4a4bc3),
	.w7(32'hbbad2e8c),
	.w8(32'hba84ffee),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d00fc),
	.w1(32'h3b57a264),
	.w2(32'hbc4fef72),
	.w3(32'hbad2fd5b),
	.w4(32'hbb872aa1),
	.w5(32'hba199612),
	.w6(32'h3a8eb1f8),
	.w7(32'hb9069e8b),
	.w8(32'hbb8a7d17),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00bb38),
	.w1(32'hbaed87ac),
	.w2(32'h3c14d6b0),
	.w3(32'h3c3e8add),
	.w4(32'hbc381b89),
	.w5(32'h39d51c63),
	.w6(32'h3be90772),
	.w7(32'hbb8e4ce4),
	.w8(32'hba9f7484),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be63b52),
	.w1(32'hbb93e498),
	.w2(32'h3b2813c2),
	.w3(32'hbbbeb506),
	.w4(32'hbbe7d32c),
	.w5(32'h39958fb8),
	.w6(32'hbbb3fb27),
	.w7(32'hb9d3cacb),
	.w8(32'h3a0b5022),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ef82c),
	.w1(32'h3930b1e0),
	.w2(32'h3c19d6d5),
	.w3(32'hbbf3df58),
	.w4(32'hbbd180dc),
	.w5(32'hbbedea5f),
	.w6(32'h3b3e9d5f),
	.w7(32'hbaa75c87),
	.w8(32'hba5131f5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806bba),
	.w1(32'h388653f1),
	.w2(32'hbb247d44),
	.w3(32'hbb454acb),
	.w4(32'h3be01328),
	.w5(32'h3b183836),
	.w6(32'hbc011a29),
	.w7(32'h3b02df2f),
	.w8(32'h3b2d7dfb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be31845),
	.w1(32'hbab785c5),
	.w2(32'hbbafca1b),
	.w3(32'h3b1bcd3c),
	.w4(32'hb803f210),
	.w5(32'hba4295fc),
	.w6(32'hba2fef6c),
	.w7(32'h3993e296),
	.w8(32'h3b269476),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee4113),
	.w1(32'hba114ba0),
	.w2(32'hbb4cd8fe),
	.w3(32'h383e748d),
	.w4(32'hbb40290f),
	.w5(32'h3aeb42aa),
	.w6(32'hbb819458),
	.w7(32'hbb54747a),
	.w8(32'hbb8a645c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081d5f),
	.w1(32'hbb613add),
	.w2(32'hba6ca93f),
	.w3(32'hbb9bd4e2),
	.w4(32'hbae5da23),
	.w5(32'hbc6bde52),
	.w6(32'h3a98e034),
	.w7(32'hb9b05824),
	.w8(32'hbbc975f9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f746d),
	.w1(32'h3bf63033),
	.w2(32'hbbb410b4),
	.w3(32'hbb94ab87),
	.w4(32'hbbbfe571),
	.w5(32'h3cf031ae),
	.w6(32'h3c233068),
	.w7(32'hbc00100d),
	.w8(32'hbaa68e07),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c5d78),
	.w1(32'h3c472376),
	.w2(32'h3afce895),
	.w3(32'hbb229739),
	.w4(32'hbb40f928),
	.w5(32'hbb926c54),
	.w6(32'hbb177be7),
	.w7(32'h3aabb4bc),
	.w8(32'hb9c9b512),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb575),
	.w1(32'h3c254d85),
	.w2(32'hbbd79632),
	.w3(32'hbb30364d),
	.w4(32'h3b5a6706),
	.w5(32'hbb6552f1),
	.w6(32'hbadab505),
	.w7(32'hb939f138),
	.w8(32'h3b98b6dd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab6d90),
	.w1(32'h3a51af69),
	.w2(32'h3bcbd6aa),
	.w3(32'hbb79dc14),
	.w4(32'hbad0f361),
	.w5(32'h3aa2c59e),
	.w6(32'h3b219562),
	.w7(32'h3b91ea8d),
	.w8(32'hbb081806),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b13b),
	.w1(32'h3b896c1a),
	.w2(32'hbbe8dcb1),
	.w3(32'hbba40d1f),
	.w4(32'hbc96eed6),
	.w5(32'h3b94a791),
	.w6(32'hbbe55f9d),
	.w7(32'h3c144c3d),
	.w8(32'h3b669b4e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40f4ce),
	.w1(32'hbc54905e),
	.w2(32'h3cccfc40),
	.w3(32'hbc0f4c83),
	.w4(32'h3b37a7a9),
	.w5(32'hbb81519f),
	.w6(32'hb9501c15),
	.w7(32'h3bb27f0c),
	.w8(32'hbbc41ff9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdc836),
	.w1(32'h3b100b79),
	.w2(32'h3ac05361),
	.w3(32'hbbdaf701),
	.w4(32'h3c42900d),
	.w5(32'hbb99e481),
	.w6(32'hb8e4a7fa),
	.w7(32'h3ba6b8eb),
	.w8(32'hbc761a5b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd5721),
	.w1(32'hb9e0f7d1),
	.w2(32'hba318d3c),
	.w3(32'hbad9ee55),
	.w4(32'hbac6b0cc),
	.w5(32'h3b1c7221),
	.w6(32'hbbec3908),
	.w7(32'hbbaa2fd3),
	.w8(32'h3a4c8221),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae66684),
	.w1(32'hbbb1d54b),
	.w2(32'h39831285),
	.w3(32'h3b1550d8),
	.w4(32'hbb50d512),
	.w5(32'h3ce55919),
	.w6(32'h3a928d95),
	.w7(32'hbbd59276),
	.w8(32'hba5316a5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983f1d8),
	.w1(32'h3b16318c),
	.w2(32'hbca791f6),
	.w3(32'hbb8cfb20),
	.w4(32'hb890edc6),
	.w5(32'h3a4b8152),
	.w6(32'hba83a425),
	.w7(32'hba54f5ef),
	.w8(32'h3aea37bd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9001c5),
	.w1(32'h3af0542b),
	.w2(32'hbaac422d),
	.w3(32'h3a828c3f),
	.w4(32'hbcb9eafc),
	.w5(32'hba2a3394),
	.w6(32'h3a0624f0),
	.w7(32'h38cfe798),
	.w8(32'h39fbf8db),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a981492),
	.w1(32'h3a1b5f9a),
	.w2(32'hbb3f632b),
	.w3(32'h3afdcd29),
	.w4(32'h3ba28df1),
	.w5(32'h3aaf14ba),
	.w6(32'h3a4ce913),
	.w7(32'h3ab1e706),
	.w8(32'hbb31254b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba094c99),
	.w1(32'hbb30d15f),
	.w2(32'h3a50845b),
	.w3(32'h3b12ca3f),
	.w4(32'h3809eba3),
	.w5(32'hba65d033),
	.w6(32'h3ae45bfb),
	.w7(32'hbab733a6),
	.w8(32'h3b3e4711),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f6f7),
	.w1(32'hba6cd0d3),
	.w2(32'h3ae939ca),
	.w3(32'h3a24f1d4),
	.w4(32'h3ac35889),
	.w5(32'h3a2118f3),
	.w6(32'h39af406a),
	.w7(32'h3aea6bcf),
	.w8(32'hbb128fb3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1b3e),
	.w1(32'h3b80730b),
	.w2(32'hbbcb0f73),
	.w3(32'h3ac36627),
	.w4(32'h3b17ab1f),
	.w5(32'hbb009a53),
	.w6(32'hb8a9be50),
	.w7(32'h3aa94bce),
	.w8(32'hba6e5b56),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ac279),
	.w1(32'h3a9322c4),
	.w2(32'hba59dbba),
	.w3(32'h3b7e155f),
	.w4(32'h3a7dd2f3),
	.w5(32'h39d03de8),
	.w6(32'h3b0fc508),
	.w7(32'h3aeebeba),
	.w8(32'hbbbc1c91),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaf4b6),
	.w1(32'h3bed1d1b),
	.w2(32'h3958404c),
	.w3(32'h3b29b038),
	.w4(32'hbb0f57bf),
	.w5(32'h3b2b2258),
	.w6(32'h3c73e459),
	.w7(32'hbad26c0f),
	.w8(32'hbb0384ff),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe876a),
	.w1(32'h3b3b0eee),
	.w2(32'hbb63a11c),
	.w3(32'hbb945569),
	.w4(32'hbbeba4d8),
	.w5(32'h3cb56064),
	.w6(32'h3a734157),
	.w7(32'h3aca778c),
	.w8(32'hba8107d3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd57f6),
	.w1(32'hb977db49),
	.w2(32'h39a5c292),
	.w3(32'hba1035e6),
	.w4(32'hbb0676a9),
	.w5(32'hba89871e),
	.w6(32'hbb1a7dfc),
	.w7(32'hbb1672a2),
	.w8(32'hb831c7ba),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13ac84),
	.w1(32'hbad79666),
	.w2(32'hbad09a9b),
	.w3(32'h3abfba05),
	.w4(32'h3a8a0f22),
	.w5(32'hba553d8d),
	.w6(32'hbaf1be15),
	.w7(32'h3a182579),
	.w8(32'h3b3067ce),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3ef5),
	.w1(32'h3965deb9),
	.w2(32'hba4b4fa2),
	.w3(32'h3a86a8b1),
	.w4(32'hbc8e6ec0),
	.w5(32'h3a5f0371),
	.w6(32'hbce6b41a),
	.w7(32'h3a161af0),
	.w8(32'h3b8057fb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354314a3),
	.w1(32'h3b0e8ae6),
	.w2(32'hb9a3eee5),
	.w3(32'h3b4ddbc3),
	.w4(32'h3b4c7408),
	.w5(32'hbaaa9c69),
	.w6(32'hb8bdc5eb),
	.w7(32'hba9dabfe),
	.w8(32'h3a042767),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25bc9d),
	.w1(32'h3a804142),
	.w2(32'h3b8b14ef),
	.w3(32'hba17d150),
	.w4(32'h3d120a00),
	.w5(32'hbaa9bb20),
	.w6(32'h3b9e7010),
	.w7(32'hbb4c6580),
	.w8(32'hbc1123b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c931438),
	.w1(32'h3712b845),
	.w2(32'h38305a81),
	.w3(32'hba3b0f29),
	.w4(32'hbb426d8f),
	.w5(32'hba19e58e),
	.w6(32'h39cbfe01),
	.w7(32'hbb48343b),
	.w8(32'h3b08d4dd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c802),
	.w1(32'h3a3f860e),
	.w2(32'h3a959aed),
	.w3(32'hbab76817),
	.w4(32'hbaac7001),
	.w5(32'hb876d018),
	.w6(32'h3b31c9b3),
	.w7(32'h3c098f87),
	.w8(32'h39637a48),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c35b5),
	.w1(32'h3cd1b09a),
	.w2(32'h3b1d1a63),
	.w3(32'h3af225a8),
	.w4(32'hb7caafcd),
	.w5(32'h3cf606de),
	.w6(32'hba06ba75),
	.w7(32'hbb098c31),
	.w8(32'hb99123b8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d10f1),
	.w1(32'h3accfb43),
	.w2(32'h39bb1f84),
	.w3(32'h3b3946b8),
	.w4(32'hbb37d238),
	.w5(32'hbcd2a542),
	.w6(32'hbc70e8f8),
	.w7(32'hba20bbf2),
	.w8(32'hbb0ada38),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a69f9),
	.w1(32'h3b02f018),
	.w2(32'h3a3287f9),
	.w3(32'hbc7803a6),
	.w4(32'h3b8f0d98),
	.w5(32'hbc5b7e8b),
	.w6(32'h38e77dd2),
	.w7(32'h3aa28dc6),
	.w8(32'h3aad7737),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961be8),
	.w1(32'h3a930c52),
	.w2(32'h3b0d006d),
	.w3(32'h395d1bf7),
	.w4(32'hbc5ebb66),
	.w5(32'h3b07a393),
	.w6(32'h39e07687),
	.w7(32'h3b54efeb),
	.w8(32'hb924bad8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbe2e),
	.w1(32'hb8d76cf0),
	.w2(32'hb9a1882d),
	.w3(32'h39645d1a),
	.w4(32'hbb78b785),
	.w5(32'h3b08783a),
	.w6(32'h397a8c9f),
	.w7(32'h3a905af3),
	.w8(32'h3a158eeb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4ee54),
	.w1(32'hba207ae9),
	.w2(32'hba4171c0),
	.w3(32'hbb1d2610),
	.w4(32'h3b9d6ea6),
	.w5(32'h3a544105),
	.w6(32'hba60edcf),
	.w7(32'h3a03ff74),
	.w8(32'hb9834bde),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956557f),
	.w1(32'h3a3d726a),
	.w2(32'hba6d1538),
	.w3(32'h3afd9838),
	.w4(32'h3a79f267),
	.w5(32'h3990850d),
	.w6(32'hb987b6bf),
	.w7(32'h3af3b7d1),
	.w8(32'h3948737f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ea20),
	.w1(32'h3a9a4ef0),
	.w2(32'h3ad143e6),
	.w3(32'hbb2244ec),
	.w4(32'hbaeec8f2),
	.w5(32'h3a1cdaa9),
	.w6(32'hbc95b118),
	.w7(32'h3aede8c4),
	.w8(32'h3921af82),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04736f),
	.w1(32'hbae4c278),
	.w2(32'h3ad946c3),
	.w3(32'h379ca87f),
	.w4(32'h398f0f6c),
	.w5(32'h3a7f478e),
	.w6(32'h3a529101),
	.w7(32'hbacc3aec),
	.w8(32'hbb43879f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08058d),
	.w1(32'h3aaaaec1),
	.w2(32'h3abcef6f),
	.w3(32'h3a89d5a1),
	.w4(32'h3b122055),
	.w5(32'hba3e8272),
	.w6(32'h3a6ec333),
	.w7(32'h3b91b905),
	.w8(32'hbb6b0ee9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996a41f),
	.w1(32'h3abd938d),
	.w2(32'h3aa0db04),
	.w3(32'h3adaca17),
	.w4(32'h3aff34bf),
	.w5(32'h3b239d0c),
	.w6(32'hb852a0cb),
	.w7(32'h3ad0385c),
	.w8(32'h3af9aa5e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45313c),
	.w1(32'h38bf0bc2),
	.w2(32'hbb75f63e),
	.w3(32'hbbd79266),
	.w4(32'hbc19be8a),
	.w5(32'h3af14bd0),
	.w6(32'hba5b50d4),
	.w7(32'h3a250727),
	.w8(32'h3ab15a71),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc95a),
	.w1(32'h3ac34872),
	.w2(32'hbb0f985b),
	.w3(32'hbc161198),
	.w4(32'h39d77562),
	.w5(32'hbb058ef3),
	.w6(32'hbafa877e),
	.w7(32'h3a6318c2),
	.w8(32'hba1c3819),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02149d),
	.w1(32'h3adcb149),
	.w2(32'hbb4b19d2),
	.w3(32'h3b8f4868),
	.w4(32'h3b27e35d),
	.w5(32'h3b6e2304),
	.w6(32'hbab80c32),
	.w7(32'h3a69a6e7),
	.w8(32'h3bfb7480),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c7121),
	.w1(32'h3a775c57),
	.w2(32'h39b506f5),
	.w3(32'hbb9c2226),
	.w4(32'hbb3963cf),
	.w5(32'h3b9402c0),
	.w6(32'hbb412f8c),
	.w7(32'hba97889c),
	.w8(32'hbc0d1006),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4526d1),
	.w1(32'h3b4e1533),
	.w2(32'h3b9f36d1),
	.w3(32'hbca2bccc),
	.w4(32'hb9edbc6f),
	.w5(32'hb99ac983),
	.w6(32'h3af04c59),
	.w7(32'hba50560b),
	.w8(32'h3b3a1a2f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9545),
	.w1(32'hbb4c4a9a),
	.w2(32'h3ba93c2a),
	.w3(32'h3a81ebb3),
	.w4(32'hba973a74),
	.w5(32'h3b8c572e),
	.w6(32'h3b01b821),
	.w7(32'h3b7880ab),
	.w8(32'h3b3f93c6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf93ab7),
	.w1(32'h3b603798),
	.w2(32'h397d1c88),
	.w3(32'hbae19d0a),
	.w4(32'hbb227bd6),
	.w5(32'h3bc01b0b),
	.w6(32'h3ba10358),
	.w7(32'hb9740228),
	.w8(32'hbba8a4ed),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a584790),
	.w1(32'hbb0e26fc),
	.w2(32'h3b020680),
	.w3(32'h3ccc71f0),
	.w4(32'hbb2e2e99),
	.w5(32'hba710279),
	.w6(32'hb90f1777),
	.w7(32'h3b3aadb1),
	.w8(32'hb9f335bc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db794),
	.w1(32'hbbcba338),
	.w2(32'h3c2040db),
	.w3(32'h3a32ca4b),
	.w4(32'h3ba381f0),
	.w5(32'hbbfffe66),
	.w6(32'hbaf0503b),
	.w7(32'hb998cefc),
	.w8(32'h3b36ed41),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc89e),
	.w1(32'hb9f6cda2),
	.w2(32'hb85b2a58),
	.w3(32'hbb3764da),
	.w4(32'hba52c8ee),
	.w5(32'hbb206473),
	.w6(32'hb9e01c8d),
	.w7(32'h3b1c0a84),
	.w8(32'h3b728648),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cbb3a),
	.w1(32'hbb1e799d),
	.w2(32'hba683e02),
	.w3(32'hba9e2be2),
	.w4(32'hbb096570),
	.w5(32'hb70b1d1b),
	.w6(32'hbbb57885),
	.w7(32'h3c4ef45a),
	.w8(32'h3c14bff8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c14b3),
	.w1(32'hba8f45fb),
	.w2(32'h3aa3e0f4),
	.w3(32'hbbf7fe87),
	.w4(32'hbb92181b),
	.w5(32'h3bd6d28c),
	.w6(32'h39017da4),
	.w7(32'h3c161794),
	.w8(32'h3ad21954),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b664d04),
	.w1(32'hbc1dbdb2),
	.w2(32'h3bcafbee),
	.w3(32'h3c2beb26),
	.w4(32'h3a510d99),
	.w5(32'hba34700a),
	.w6(32'h3aa32dc5),
	.w7(32'hba902d08),
	.w8(32'h3b733e5e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd985e),
	.w1(32'hbb66d9ae),
	.w2(32'h3aec9528),
	.w3(32'h3958b6ad),
	.w4(32'h3a5a268b),
	.w5(32'h3b9dcd37),
	.w6(32'hbba4031f),
	.w7(32'h3c3542f2),
	.w8(32'h3b09b2c8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414a5f),
	.w1(32'hbab47e8a),
	.w2(32'h3abb5a03),
	.w3(32'hbbacaf43),
	.w4(32'hb77829d5),
	.w5(32'hbb1a8efa),
	.w6(32'h39953768),
	.w7(32'hbba772a1),
	.w8(32'h3a3f25ec),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3616ee),
	.w1(32'hbc493fad),
	.w2(32'h3aafa052),
	.w3(32'hbbdc16d0),
	.w4(32'hbb9c01d9),
	.w5(32'h3bde75f1),
	.w6(32'h3a7c56c8),
	.w7(32'hb83823c3),
	.w8(32'hbb24a802),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb9de3),
	.w1(32'h3acf7ba4),
	.w2(32'h3b0db199),
	.w3(32'h3bd5ec90),
	.w4(32'hb960671c),
	.w5(32'h3b124ba2),
	.w6(32'hbae569d4),
	.w7(32'h39ffa78d),
	.w8(32'h38bdf832),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae51153),
	.w1(32'hb9d0dd05),
	.w2(32'hb7ba473c),
	.w3(32'hbb26018f),
	.w4(32'hbaae065e),
	.w5(32'h3a49f38b),
	.w6(32'hbb5f7d7c),
	.w7(32'h3a2ff5cd),
	.w8(32'hbabda6b3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba268481),
	.w1(32'h388e9b0f),
	.w2(32'hba196ba3),
	.w3(32'hbacdc723),
	.w4(32'hb991f282),
	.w5(32'hbb277841),
	.w6(32'hbb8fd9d6),
	.w7(32'hbb62bac5),
	.w8(32'hb8c78e27),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37b1ad),
	.w1(32'h38aa64bf),
	.w2(32'h3a6345e6),
	.w3(32'h3a92eb29),
	.w4(32'h3c34d184),
	.w5(32'hbb114744),
	.w6(32'h3bdeaeb2),
	.w7(32'h3c0d59c8),
	.w8(32'h3a4cd574),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b976a),
	.w1(32'hbbd99499),
	.w2(32'h3ae1786c),
	.w3(32'hba5d9fe9),
	.w4(32'h3b4ce441),
	.w5(32'h3b05f696),
	.w6(32'h3c612161),
	.w7(32'h3ac0e0f1),
	.w8(32'h3c343058),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9404),
	.w1(32'hbc0c3e84),
	.w2(32'hbb343aa3),
	.w3(32'h3a4059f7),
	.w4(32'hb91e47f7),
	.w5(32'hb8d564cf),
	.w6(32'hbb1918ab),
	.w7(32'hbb64c39e),
	.w8(32'h3bac4f62),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe89dd),
	.w1(32'h3af744f5),
	.w2(32'h3b31970f),
	.w3(32'h3c37a3af),
	.w4(32'hbb8f51a9),
	.w5(32'h3ab6937f),
	.w6(32'h3b9c0115),
	.w7(32'hbc507bb7),
	.w8(32'hbc5679bb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0efeed),
	.w1(32'h3a297690),
	.w2(32'hba2f1210),
	.w3(32'hba513d3e),
	.w4(32'h38c8d6ba),
	.w5(32'h34ba2e47),
	.w6(32'hb9ddfbaf),
	.w7(32'h3ac5c1a6),
	.w8(32'h3ab2816b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb605231),
	.w1(32'h3ad88f49),
	.w2(32'h3c9fa681),
	.w3(32'h3a1bae81),
	.w4(32'hbbdfd589),
	.w5(32'hba0c9e67),
	.w6(32'hb5a7a9ee),
	.w7(32'hba260bc9),
	.w8(32'hba2b77c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315d85),
	.w1(32'h3b2f0dc3),
	.w2(32'h3b494ffe),
	.w3(32'hbc09be4e),
	.w4(32'hbb5a001a),
	.w5(32'hba8591b7),
	.w6(32'hbae5dea2),
	.w7(32'h39d246c8),
	.w8(32'h3b170258),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66c326),
	.w1(32'h3bd7f722),
	.w2(32'h3b2ae782),
	.w3(32'h3a8fb6d5),
	.w4(32'hbbd6cc1e),
	.w5(32'h36289bf6),
	.w6(32'h3bd9554e),
	.w7(32'h3b03671f),
	.w8(32'h3b456c81),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a705556),
	.w1(32'h3b08acfe),
	.w2(32'hbb7d503f),
	.w3(32'hbc2e5745),
	.w4(32'h3b8b8d75),
	.w5(32'hbaf26943),
	.w6(32'h3a11eacc),
	.w7(32'h3b964280),
	.w8(32'h3b70da34),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978775),
	.w1(32'hbb33dffc),
	.w2(32'hb7f3327d),
	.w3(32'h3b29f2a7),
	.w4(32'hbac9d2ac),
	.w5(32'h3a109896),
	.w6(32'hba954a29),
	.w7(32'hbbb02d2b),
	.w8(32'hbbd84d0f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95246f),
	.w1(32'h3b519683),
	.w2(32'h3c35aa73),
	.w3(32'h3a814dd8),
	.w4(32'h3b85dc21),
	.w5(32'hba98f2ae),
	.w6(32'h3c0de616),
	.w7(32'hbc54132b),
	.w8(32'hba4da910),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb795a450),
	.w1(32'hbb75c2e9),
	.w2(32'hbbe8c30a),
	.w3(32'hbbebda2f),
	.w4(32'hbadeb9df),
	.w5(32'h3b8fc7db),
	.w6(32'hba371703),
	.w7(32'hbbbab43a),
	.w8(32'h3c0336e9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4b86),
	.w1(32'h3b9e3df0),
	.w2(32'hba256f2f),
	.w3(32'h3beb4952),
	.w4(32'hbb48f6b7),
	.w5(32'hbbf765aa),
	.w6(32'hbb481fba),
	.w7(32'hbb40d9e9),
	.w8(32'h3c49e104),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8ae6),
	.w1(32'hba27627c),
	.w2(32'h3b4e5ea8),
	.w3(32'h3b872356),
	.w4(32'hba8adfa6),
	.w5(32'hbc015127),
	.w6(32'h3b8327a1),
	.w7(32'h3c6b5fb9),
	.w8(32'hbb4207e3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0c30),
	.w1(32'hbb15c4a6),
	.w2(32'h3b5611bb),
	.w3(32'hbbbe015a),
	.w4(32'hbb8fb13b),
	.w5(32'hbbc597df),
	.w6(32'h3b8b7754),
	.w7(32'h3aadb454),
	.w8(32'hbb2f5f86),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cdc59),
	.w1(32'hbaebd2da),
	.w2(32'h3c02d6d4),
	.w3(32'h39f216bd),
	.w4(32'hb9e811da),
	.w5(32'h3b8ae247),
	.w6(32'hbab937f6),
	.w7(32'hbb9af8a9),
	.w8(32'hbb940868),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5ec20),
	.w1(32'hbb636409),
	.w2(32'hba9a6979),
	.w3(32'hba13e84e),
	.w4(32'hbbc80a19),
	.w5(32'hb957c3ce),
	.w6(32'h3ba503d0),
	.w7(32'h3bbf7bde),
	.w8(32'h3ac94810),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85be71),
	.w1(32'h3bad0049),
	.w2(32'h3a3dd598),
	.w3(32'h3b02ca23),
	.w4(32'h3b91f15e),
	.w5(32'hbb0c942f),
	.w6(32'hbc200c81),
	.w7(32'hbb857316),
	.w8(32'hb87e1d82),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5150f3),
	.w1(32'hbbb537eb),
	.w2(32'hba0830bd),
	.w3(32'h3a4037db),
	.w4(32'hbbb3dc01),
	.w5(32'hba32488d),
	.w6(32'h3cabec44),
	.w7(32'hb8819756),
	.w8(32'hbb0c9e0d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca436b1),
	.w1(32'hbacece8d),
	.w2(32'h3c296bdf),
	.w3(32'hbac9fcb2),
	.w4(32'h3b53f0e0),
	.w5(32'h3b329f97),
	.w6(32'h3c99e1a3),
	.w7(32'hbc15898e),
	.w8(32'hbba93cbe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cd7b2),
	.w1(32'h3c856622),
	.w2(32'h392b42b7),
	.w3(32'h3b6e2d02),
	.w4(32'h3bfeb41d),
	.w5(32'h3be236dc),
	.w6(32'h38ba1453),
	.w7(32'hba3fc71d),
	.w8(32'h3b2ea06f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc256a89),
	.w1(32'hba527595),
	.w2(32'h3ae1e131),
	.w3(32'h3ace7d43),
	.w4(32'h3bd10698),
	.w5(32'h3c548554),
	.w6(32'hbb4649b1),
	.w7(32'hbb31f383),
	.w8(32'hbb43d7d9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c69b4),
	.w1(32'hbbeda13a),
	.w2(32'hbb9ce111),
	.w3(32'hbc3b1b32),
	.w4(32'h3b0d1384),
	.w5(32'h3ccb5ddc),
	.w6(32'hbaac0344),
	.w7(32'h399647cb),
	.w8(32'h3853b4c6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3de11d),
	.w1(32'h3ac10da7),
	.w2(32'hbab0f6e9),
	.w3(32'hb9bf1edf),
	.w4(32'h3a93c816),
	.w5(32'hbba62c2c),
	.w6(32'hbb962e85),
	.w7(32'hbb989a60),
	.w8(32'h3b95b728),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d1eaf),
	.w1(32'hbbb6f863),
	.w2(32'hbb3e6a0d),
	.w3(32'h3b99ddba),
	.w4(32'hbaf35011),
	.w5(32'hbc45589e),
	.w6(32'h3b270c93),
	.w7(32'hbbae14c2),
	.w8(32'h3b194cdf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926d22e),
	.w1(32'h3b434327),
	.w2(32'h3ad4e440),
	.w3(32'hbb1ee4b8),
	.w4(32'hbbcdad92),
	.w5(32'h3c264c8b),
	.w6(32'hbb7b25ec),
	.w7(32'hbb33f79f),
	.w8(32'h3c006819),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4de4f3),
	.w1(32'hbb5a0b7b),
	.w2(32'hbb90e04e),
	.w3(32'hbb10e3c9),
	.w4(32'h3b19c7f5),
	.w5(32'hbb75934e),
	.w6(32'hbaa4e923),
	.w7(32'hb9890a40),
	.w8(32'h3b44af04),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2fd0),
	.w1(32'hbb18c342),
	.w2(32'h3b4c9567),
	.w3(32'hba3b4a62),
	.w4(32'hba4db220),
	.w5(32'hb9d8e3c4),
	.w6(32'hbafcdaec),
	.w7(32'hbb73acf6),
	.w8(32'hbb04c096),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ca40),
	.w1(32'hbb32273d),
	.w2(32'h3b83d47e),
	.w3(32'hbbdedfdd),
	.w4(32'hbb2fa243),
	.w5(32'h39ac44f5),
	.w6(32'hba9d5194),
	.w7(32'h3bc1358c),
	.w8(32'hbaa51ca3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad610d),
	.w1(32'hbc5d8eef),
	.w2(32'h3a998100),
	.w3(32'h3a09abcb),
	.w4(32'hbbce8e6b),
	.w5(32'hbae847d7),
	.w6(32'hbb13798e),
	.w7(32'hbb84f50b),
	.w8(32'hbbf11ff8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff543),
	.w1(32'hbc2ab565),
	.w2(32'h3ba641d5),
	.w3(32'h3c8342e3),
	.w4(32'h3b967a4b),
	.w5(32'h3bbb9593),
	.w6(32'hba756715),
	.w7(32'h3a04f1a0),
	.w8(32'hbb973c04),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a96d),
	.w1(32'hbbe5b496),
	.w2(32'h398f916a),
	.w3(32'hbbd774f4),
	.w4(32'hba8e9081),
	.w5(32'h3a5e7968),
	.w6(32'hbac434aa),
	.w7(32'hbaede51e),
	.w8(32'h3c58a6e3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb393f4),
	.w1(32'h3b2f5b0c),
	.w2(32'hbb68eb62),
	.w3(32'hbc080744),
	.w4(32'hba4397e4),
	.w5(32'h3b8749fc),
	.w6(32'h37baa5c1),
	.w7(32'h3aec340e),
	.w8(32'hb7ce12be),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b784dcb),
	.w1(32'h3b8fe5b0),
	.w2(32'h3a035ded),
	.w3(32'h3ad8f9b8),
	.w4(32'hba5a2eba),
	.w5(32'hba0bf18b),
	.w6(32'hbb4b6310),
	.w7(32'h3b0492f8),
	.w8(32'h3b7b61d8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd83438),
	.w1(32'h3b2993a9),
	.w2(32'hbbe116a9),
	.w3(32'hbb2ec599),
	.w4(32'h3ad71517),
	.w5(32'hbb675924),
	.w6(32'hba1a1f74),
	.w7(32'h3a66c04c),
	.w8(32'h3c977c3a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6ae0),
	.w1(32'h3b4fbf4a),
	.w2(32'h3a642ce3),
	.w3(32'hbb1ad389),
	.w4(32'hbb47b7de),
	.w5(32'h3c91a016),
	.w6(32'h3b2e2935),
	.w7(32'h3b769279),
	.w8(32'h3b62e830),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db971),
	.w1(32'h3bcd3208),
	.w2(32'hbb3fb92a),
	.w3(32'hba2e2140),
	.w4(32'hbaa7d88b),
	.w5(32'hbc771165),
	.w6(32'h3b814eb0),
	.w7(32'h3b0c2ad8),
	.w8(32'hbb8fd564),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2fe8a),
	.w1(32'hb944b207),
	.w2(32'h3aa9731d),
	.w3(32'h3b02afc8),
	.w4(32'hbb5cf9d8),
	.w5(32'hbbade640),
	.w6(32'h3bced739),
	.w7(32'hbb15a1b9),
	.w8(32'h399f70fa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88a772),
	.w1(32'h3b809d36),
	.w2(32'h399b0cb7),
	.w3(32'h3b510322),
	.w4(32'h3b871a7f),
	.w5(32'hbbbef01a),
	.w6(32'h3a531597),
	.w7(32'h3b26a14b),
	.w8(32'hbbdcf0c9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd5d14),
	.w1(32'h3a38f912),
	.w2(32'h3a52012f),
	.w3(32'h3c62aa32),
	.w4(32'hbb373fe1),
	.w5(32'h39849927),
	.w6(32'hbaa8e3a9),
	.w7(32'h3afadcb5),
	.w8(32'hb9d52c05),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1526),
	.w1(32'hb789c6c9),
	.w2(32'hba03d65e),
	.w3(32'hbb4b40dd),
	.w4(32'h39dc6193),
	.w5(32'hbb15cd17),
	.w6(32'h3a2794a3),
	.w7(32'h3b424311),
	.w8(32'hb9ce9b90),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c90f1),
	.w1(32'h3b886098),
	.w2(32'hb9d7f000),
	.w3(32'hba7dec9f),
	.w4(32'h3a61b0c3),
	.w5(32'hb81072db),
	.w6(32'h3b8d2c50),
	.w7(32'h3b65876c),
	.w8(32'hbabe204f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9583),
	.w1(32'h3b368faf),
	.w2(32'h3b7f4ffd),
	.w3(32'hba6baaf5),
	.w4(32'hba7cc48b),
	.w5(32'h3b0bb869),
	.w6(32'h3bb2b468),
	.w7(32'hba2cad29),
	.w8(32'hbbd7cca4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8c011),
	.w1(32'hba11a375),
	.w2(32'h3b9ab7d8),
	.w3(32'h3baf353c),
	.w4(32'hbb354d56),
	.w5(32'h3a3aecbf),
	.w6(32'hb9891173),
	.w7(32'hbaca4dfe),
	.w8(32'h3b904cb4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a61b1d),
	.w1(32'h3b3102bd),
	.w2(32'h3bbe7349),
	.w3(32'h3b227f40),
	.w4(32'h3b62de7e),
	.w5(32'h3a99e9b4),
	.w6(32'hbab3971c),
	.w7(32'h396920ba),
	.w8(32'h3aa7ed9a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96cdee),
	.w1(32'hbaf91139),
	.w2(32'h3acc3d62),
	.w3(32'hbad5fe0c),
	.w4(32'hba6213d7),
	.w5(32'h3b1175c8),
	.w6(32'h3a995556),
	.w7(32'hbadb6be8),
	.w8(32'hbbd25c5e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5bdf2),
	.w1(32'hbbd0ded9),
	.w2(32'h3bd69140),
	.w3(32'hbb72b3a3),
	.w4(32'h3bbaa7dc),
	.w5(32'hbc233ae0),
	.w6(32'hbbcbdb8f),
	.w7(32'h3c7a658d),
	.w8(32'hbb184845),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee796),
	.w1(32'hbb690371),
	.w2(32'h3b632b22),
	.w3(32'hb9f1d396),
	.w4(32'h3ac040a9),
	.w5(32'hbb0af6b0),
	.w6(32'h3a12f3b8),
	.w7(32'h3aab0951),
	.w8(32'hbb2d6dbd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39934fb2),
	.w1(32'h37f07703),
	.w2(32'hb9868c34),
	.w3(32'h3c408bad),
	.w4(32'h3c2a67a7),
	.w5(32'hbb259d86),
	.w6(32'h3ab275ab),
	.w7(32'hbaca901d),
	.w8(32'hbb93319a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b868dd6),
	.w1(32'hbb4c0084),
	.w2(32'h3b4f0499),
	.w3(32'h38a0f067),
	.w4(32'hbb2a9b68),
	.w5(32'hbacb60c2),
	.w6(32'hba8ae644),
	.w7(32'h3b68d870),
	.w8(32'hbb50506c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e523f),
	.w1(32'hb99f478e),
	.w2(32'hbb3640a4),
	.w3(32'hbaa98eca),
	.w4(32'h3adfccc5),
	.w5(32'hbb455a9e),
	.w6(32'hbb2b0d50),
	.w7(32'hbc0ae11b),
	.w8(32'hba8db9cd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75457),
	.w1(32'hb58c9842),
	.w2(32'hba98ac92),
	.w3(32'h39648cb5),
	.w4(32'h3b1d5389),
	.w5(32'hbb3d7e3f),
	.w6(32'h3b2353f9),
	.w7(32'hb83e496b),
	.w8(32'hb88c2d8e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b7f9),
	.w1(32'hb94737c1),
	.w2(32'h3a3e68b7),
	.w3(32'hbaddc503),
	.w4(32'h3b454e74),
	.w5(32'h3c8aa173),
	.w6(32'h3b3e0e9e),
	.w7(32'hbb886529),
	.w8(32'h3a6ed130),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb079d7),
	.w1(32'h3a3f99e6),
	.w2(32'hba38226d),
	.w3(32'hbbae9cd3),
	.w4(32'hbba464ba),
	.w5(32'hbb42515f),
	.w6(32'hbb79a03f),
	.w7(32'h3a48fc4b),
	.w8(32'h3b368b49),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba989f1d),
	.w1(32'h3b14595c),
	.w2(32'hb64e08f5),
	.w3(32'h3bb444bf),
	.w4(32'hbb733627),
	.w5(32'hb9c9cef3),
	.w6(32'h3af2f8f4),
	.w7(32'hba9ebeb5),
	.w8(32'h3c3106c2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900e281),
	.w1(32'h3a2f40f4),
	.w2(32'h3c49bfcd),
	.w3(32'hb9b6cdbb),
	.w4(32'h3a636e91),
	.w5(32'h3aee6bf9),
	.w6(32'h3aac9ac8),
	.w7(32'h3ab57029),
	.w8(32'hbac304a2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29a24d),
	.w1(32'h3b2096d7),
	.w2(32'hbb4e0d9b),
	.w3(32'h3c4d9946),
	.w4(32'h3a801dad),
	.w5(32'hbb93ca62),
	.w6(32'hb8a67bf3),
	.w7(32'hbc2b65ef),
	.w8(32'hbb3aa29e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba780b8b),
	.w1(32'h3b6079cc),
	.w2(32'h3abb4a0a),
	.w3(32'hbad88273),
	.w4(32'hbb8c4d78),
	.w5(32'h3b3ee499),
	.w6(32'h3b8326d1),
	.w7(32'h39fb6b05),
	.w8(32'h3a8e5c55),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa5af),
	.w1(32'h3b572c0f),
	.w2(32'h3add7c66),
	.w3(32'h3b48d0cc),
	.w4(32'h3b3f91f3),
	.w5(32'hba015ae8),
	.w6(32'hbb73f679),
	.w7(32'hbb63b8e1),
	.w8(32'hba33cd9c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28bca3),
	.w1(32'hba0808fb),
	.w2(32'h374c38e2),
	.w3(32'h3ac4cd04),
	.w4(32'hbac745de),
	.w5(32'hbb10eb12),
	.w6(32'h39c8d2dc),
	.w7(32'hbb1c41c2),
	.w8(32'hbae09dd2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe4a4c),
	.w1(32'h3aefade6),
	.w2(32'h3a29d60d),
	.w3(32'hba599d16),
	.w4(32'hbc13a17a),
	.w5(32'h3bcc7d3a),
	.w6(32'h3ac9deb7),
	.w7(32'hbb288e30),
	.w8(32'h3aafa4d1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95fdea4),
	.w1(32'hb9c318c9),
	.w2(32'h39bfc0a2),
	.w3(32'hbb883d41),
	.w4(32'hbab49bca),
	.w5(32'h3a8e24b5),
	.w6(32'h3a83ec9e),
	.w7(32'h3a859e76),
	.w8(32'h3b5cafbd),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08adc),
	.w1(32'h3aff5b64),
	.w2(32'h3b51685c),
	.w3(32'h38cb2f19),
	.w4(32'hbb373af9),
	.w5(32'h3aac9621),
	.w6(32'h3a203ab9),
	.w7(32'hbcb2a3f9),
	.w8(32'h3b29a94c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995a6b2),
	.w1(32'h3b1c1fce),
	.w2(32'h3aecb8c0),
	.w3(32'h3aa9a2b9),
	.w4(32'h3acf73b4),
	.w5(32'h3b674ce2),
	.w6(32'h3af7e7ff),
	.w7(32'h3ab74343),
	.w8(32'hba3d18ba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bebd),
	.w1(32'h3b2fe210),
	.w2(32'h3a813c72),
	.w3(32'h3a07cde8),
	.w4(32'h3b23e41d),
	.w5(32'h3b8c1458),
	.w6(32'h3b8af862),
	.w7(32'h3b60a122),
	.w8(32'hbaea1a2b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95719d),
	.w1(32'hba17a653),
	.w2(32'h3ab7def9),
	.w3(32'h3bb5d421),
	.w4(32'hbb9ec240),
	.w5(32'h3bc2450c),
	.w6(32'hbc9864c8),
	.w7(32'hba727339),
	.w8(32'hbb616a3e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906ed0a),
	.w1(32'hba912f1c),
	.w2(32'hbbd7285a),
	.w3(32'h3aae1fda),
	.w4(32'h3a7b0482),
	.w5(32'hbb684034),
	.w6(32'h3b752031),
	.w7(32'h3ba4c681),
	.w8(32'hbb2a3acf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30b40),
	.w1(32'hbc8a7b67),
	.w2(32'hbb7183a0),
	.w3(32'hba7b3fa2),
	.w4(32'hbbbf5be1),
	.w5(32'hbbab2a8f),
	.w6(32'hbc144cbe),
	.w7(32'h3b9b798a),
	.w8(32'hbb107fc9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f773a),
	.w1(32'h3b9b2c81),
	.w2(32'hbb1f6a14),
	.w3(32'hba45cd98),
	.w4(32'hbc2c68c7),
	.w5(32'hba852dfc),
	.w6(32'hbb2c4afe),
	.w7(32'h3bc0c32d),
	.w8(32'h3b7bcd23),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa588),
	.w1(32'hba8c7288),
	.w2(32'h3b8b1b77),
	.w3(32'h3bb76ca8),
	.w4(32'h3ba121b1),
	.w5(32'h3aec9270),
	.w6(32'h3c8d8581),
	.w7(32'hba740378),
	.w8(32'hb8695eae),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22c16b),
	.w1(32'hbbcbdee1),
	.w2(32'h3c5cabe0),
	.w3(32'h3a856589),
	.w4(32'hbc8e1af2),
	.w5(32'h3b821c22),
	.w6(32'h3a23dafe),
	.w7(32'h3b8794a7),
	.w8(32'h3b85ab44),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea3833),
	.w1(32'hbbdc4932),
	.w2(32'hbb2fbb56),
	.w3(32'h3aa97e16),
	.w4(32'h3b940768),
	.w5(32'h3b8c0c7d),
	.w6(32'h3bbc43d5),
	.w7(32'h39ec0b8d),
	.w8(32'h3bf13d36),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab115d),
	.w1(32'h3acfaa91),
	.w2(32'hb8d8313f),
	.w3(32'hbb37bd49),
	.w4(32'hbb60c6ff),
	.w5(32'h39225313),
	.w6(32'hb9c753b0),
	.w7(32'h3b1e0340),
	.w8(32'hbb5a4eb5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf1706),
	.w1(32'hbafc303d),
	.w2(32'h3bf4df1d),
	.w3(32'h3cb1b113),
	.w4(32'h3bc6ed4f),
	.w5(32'hbb3c6df1),
	.w6(32'h3b2ed21a),
	.w7(32'hb83ebc2d),
	.w8(32'hbb464f4b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1c79),
	.w1(32'hbaba7e53),
	.w2(32'hbb8abcb8),
	.w3(32'hba0cbf93),
	.w4(32'hbb26b2f3),
	.w5(32'hba7c76fa),
	.w6(32'hb9ab58dc),
	.w7(32'h3b676a73),
	.w8(32'h3b65a47e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c820c85),
	.w1(32'hb8002f17),
	.w2(32'h3a0d07ba),
	.w3(32'hbc3c0a1f),
	.w4(32'h3be224b9),
	.w5(32'hbc0c5677),
	.w6(32'hbbfa9620),
	.w7(32'hbb3fb34b),
	.w8(32'hba493270),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a4164),
	.w1(32'hbb9abff2),
	.w2(32'hbb0d1437),
	.w3(32'hbc001e38),
	.w4(32'hba028f4d),
	.w5(32'h3aebdcaa),
	.w6(32'h3c0f560b),
	.w7(32'hbbc36c4a),
	.w8(32'hbbfd6320),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac954b0),
	.w1(32'hbabdaa2b),
	.w2(32'h3c1307c0),
	.w3(32'hb8f47205),
	.w4(32'hbb1184a6),
	.w5(32'hbc1e89d3),
	.w6(32'h3c2f76e8),
	.w7(32'h397a6e11),
	.w8(32'h3c8a14d3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8f36),
	.w1(32'hbba9e3e8),
	.w2(32'hbc242b82),
	.w3(32'hbc1ff206),
	.w4(32'hba38518f),
	.w5(32'h3afba366),
	.w6(32'hbb39efcc),
	.w7(32'hbb294c65),
	.w8(32'h3a16a1ea),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee9c8),
	.w1(32'h3a776cfa),
	.w2(32'hbb3814a8),
	.w3(32'h3b2a55aa),
	.w4(32'hba9ea664),
	.w5(32'hb8d34b98),
	.w6(32'h3bb03f60),
	.w7(32'h3ad8a546),
	.w8(32'h3bd73028),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39928625),
	.w1(32'hbb4a691d),
	.w2(32'h3afadc8c),
	.w3(32'hbb9f9e42),
	.w4(32'hbc088537),
	.w5(32'h3be490f2),
	.w6(32'hbbc6069d),
	.w7(32'h3b904288),
	.w8(32'hbb29f91d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb544d08),
	.w1(32'h3c1b51aa),
	.w2(32'hbbf0c1da),
	.w3(32'hba876b16),
	.w4(32'h38083477),
	.w5(32'hbc0c5b97),
	.w6(32'hbc06507e),
	.w7(32'h3aa7c8c7),
	.w8(32'hbc3d4d3e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea1315),
	.w1(32'h3bcd1a6c),
	.w2(32'h3b83b3d4),
	.w3(32'hbb7fcd6f),
	.w4(32'hbb4eb1ea),
	.w5(32'h3ace31f9),
	.w6(32'hba0e0fb1),
	.w7(32'hba062301),
	.w8(32'hbbb301ce),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0bdd),
	.w1(32'h3c592205),
	.w2(32'hb94649da),
	.w3(32'h3bd0992a),
	.w4(32'hbbba76c1),
	.w5(32'hbb3d0e90),
	.w6(32'h3b8e5ae6),
	.w7(32'h3aea7b74),
	.w8(32'h3b718e32),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29372a),
	.w1(32'hb986e2cd),
	.w2(32'h39a8c508),
	.w3(32'hbc570d75),
	.w4(32'hbb2038c3),
	.w5(32'h3b39c4a8),
	.w6(32'hbbccfb28),
	.w7(32'hba6ac00b),
	.w8(32'hb9cba670),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905025),
	.w1(32'hb96cfaac),
	.w2(32'h3abd4773),
	.w3(32'hbafe1247),
	.w4(32'h3bd8ad34),
	.w5(32'h3c869082),
	.w6(32'h3b5ed6a4),
	.w7(32'h3c940cac),
	.w8(32'h3c21c876),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997465d),
	.w1(32'h3bd9ac1f),
	.w2(32'hba9dd4b0),
	.w3(32'h3b9b8c49),
	.w4(32'h3b5f4a8b),
	.w5(32'h3b8f071f),
	.w6(32'hbc3020a7),
	.w7(32'h3c944f49),
	.w8(32'hbb996c99),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2102),
	.w1(32'hbb193a17),
	.w2(32'hbc1ef009),
	.w3(32'h3bb4d03c),
	.w4(32'hbae9b194),
	.w5(32'h3b0aa322),
	.w6(32'h3b6ead1b),
	.w7(32'h35af6558),
	.w8(32'hbbb7d200),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a0e9),
	.w1(32'h3ac6561d),
	.w2(32'h3a335bee),
	.w3(32'h3b072bc2),
	.w4(32'h3c80e8b8),
	.w5(32'hbaf15ff8),
	.w6(32'hb9bad074),
	.w7(32'hbbaff868),
	.w8(32'hbc8d7b64),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaf033),
	.w1(32'h3a795533),
	.w2(32'hbb2081d5),
	.w3(32'h3b99ed75),
	.w4(32'h3b2dc93a),
	.w5(32'hb901f8e0),
	.w6(32'hbc0e3d77),
	.w7(32'hbc0eb3a2),
	.w8(32'h3af3277a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7ca0),
	.w1(32'hbb39f042),
	.w2(32'hbb594771),
	.w3(32'hbbadae48),
	.w4(32'hbae9ba37),
	.w5(32'hbae91498),
	.w6(32'h3af9e78c),
	.w7(32'hb978e77b),
	.w8(32'hbcb6241a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca68367),
	.w1(32'hba57ab8e),
	.w2(32'h3b16a0f2),
	.w3(32'h3a3e852a),
	.w4(32'h3bf4fd59),
	.w5(32'hbb364825),
	.w6(32'hbb9d6341),
	.w7(32'hb9e11d84),
	.w8(32'h39ce1bdd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d5b1),
	.w1(32'hbb919273),
	.w2(32'h3bf0a96f),
	.w3(32'hbb491ba7),
	.w4(32'h3b470e4f),
	.w5(32'hbb3c7302),
	.w6(32'h3af4b031),
	.w7(32'hbc3f08eb),
	.w8(32'hbc1be593),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b3f5),
	.w1(32'h3aa348a9),
	.w2(32'hbc102815),
	.w3(32'h3b323fd4),
	.w4(32'hbbebb892),
	.w5(32'hbb8ee1ac),
	.w6(32'h39aa36d7),
	.w7(32'hbbb5582b),
	.w8(32'h38a502dc),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c28ca),
	.w1(32'h3bc6c538),
	.w2(32'hbaf41324),
	.w3(32'h3b9ceb54),
	.w4(32'hbbe67ede),
	.w5(32'h3b6a94b9),
	.w6(32'h3bbff78b),
	.w7(32'h3a2fc628),
	.w8(32'hbc0a643e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e9698),
	.w1(32'h3b8b14ce),
	.w2(32'hbb9b23f1),
	.w3(32'hbaeeea2f),
	.w4(32'h3b82eace),
	.w5(32'h3c1f080f),
	.w6(32'h3b5f2564),
	.w7(32'h3c8ba30e),
	.w8(32'hbc9bbd88),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c5a16),
	.w1(32'h3c028565),
	.w2(32'hbacef92f),
	.w3(32'h3ab0a8e7),
	.w4(32'h3bd38683),
	.w5(32'hbbaa2dda),
	.w6(32'hbb88f4e7),
	.w7(32'hbb3b4e10),
	.w8(32'h3c031755),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a834937),
	.w1(32'hbaf9b161),
	.w2(32'hbc840c70),
	.w3(32'hbc0b3062),
	.w4(32'hbb56946b),
	.w5(32'hbb43dec7),
	.w6(32'hbbc4aff5),
	.w7(32'h3bad7ede),
	.w8(32'h3ade53da),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c99af),
	.w1(32'hba8d5fd6),
	.w2(32'h3a779060),
	.w3(32'h379d0074),
	.w4(32'hbb18ea02),
	.w5(32'h3b389db4),
	.w6(32'h3aa286d1),
	.w7(32'h3c73ecae),
	.w8(32'hbbc9051c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc5c90),
	.w1(32'hbbadef64),
	.w2(32'h3bb00199),
	.w3(32'hbbd05763),
	.w4(32'h3c0de19c),
	.w5(32'hbb3e7c2f),
	.w6(32'hbbcaf294),
	.w7(32'h3c82102b),
	.w8(32'h3a4b4741),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a9bf),
	.w1(32'hba7ec632),
	.w2(32'hbbccbae0),
	.w3(32'h3c584d90),
	.w4(32'h3ac354b2),
	.w5(32'hbb1b16c8),
	.w6(32'h3b7cbdf4),
	.w7(32'h3b92f019),
	.w8(32'hbb4efa99),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3e9d0),
	.w1(32'hbbec82dd),
	.w2(32'hbae59e7e),
	.w3(32'h3b3c461d),
	.w4(32'hb8a7c022),
	.w5(32'h3a93b3a1),
	.w6(32'hbb917651),
	.w7(32'h3cbb8bd2),
	.w8(32'h3cc8357e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33015b),
	.w1(32'hbb130f5b),
	.w2(32'h3bda1d9a),
	.w3(32'h3b37108a),
	.w4(32'hbc05a6da),
	.w5(32'hbc59d11f),
	.w6(32'hba5fdd52),
	.w7(32'hbc3613bf),
	.w8(32'hbb2ca357),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7992),
	.w1(32'hbbe4d16f),
	.w2(32'h3c3f709a),
	.w3(32'h3cf3ce91),
	.w4(32'h3c478cbc),
	.w5(32'h3ba1e858),
	.w6(32'hbb10a08c),
	.w7(32'h3ca39949),
	.w8(32'h3a86ff5a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24a674),
	.w1(32'h3c65a936),
	.w2(32'h3b264590),
	.w3(32'h3be96e5b),
	.w4(32'hba9a5021),
	.w5(32'h3bff2186),
	.w6(32'h3ba14c06),
	.w7(32'h3ac5ba0b),
	.w8(32'hbbb2b274),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c848b),
	.w1(32'h3c86a395),
	.w2(32'hbc081b90),
	.w3(32'h3c3c3eb1),
	.w4(32'hbb0e60c0),
	.w5(32'h3c04a6f5),
	.w6(32'h3c490219),
	.w7(32'hb7cf7740),
	.w8(32'hbc44ac07),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86038e6),
	.w1(32'h3c29a4a8),
	.w2(32'hbb9fc410),
	.w3(32'hbc0bfda9),
	.w4(32'h3ac3022f),
	.w5(32'h3c976197),
	.w6(32'h3bf48795),
	.w7(32'h3c8569c5),
	.w8(32'h3b84a448),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0f46),
	.w1(32'hbb4f5ac7),
	.w2(32'hba975ed4),
	.w3(32'h3c5dde4e),
	.w4(32'hbc348c74),
	.w5(32'h381e69f0),
	.w6(32'hbb910237),
	.w7(32'hbbac0246),
	.w8(32'h3c215327),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907bb64),
	.w1(32'h3c5259f4),
	.w2(32'h3a15ccd3),
	.w3(32'h3c67a55c),
	.w4(32'hb9a0a271),
	.w5(32'h3bddda35),
	.w6(32'hb4fd2fa2),
	.w7(32'h3a0265cd),
	.w8(32'hbbd7f7cf),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f1407),
	.w1(32'h38e5bcf0),
	.w2(32'h3c3cd8f9),
	.w3(32'h3a8bd409),
	.w4(32'hbb744796),
	.w5(32'h3a2ad760),
	.w6(32'h3aeaef46),
	.w7(32'h3b54c209),
	.w8(32'hbb8bb970),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb447cfa),
	.w1(32'h3bbf7767),
	.w2(32'hbb6b9a7f),
	.w3(32'h3adc0096),
	.w4(32'hba26b163),
	.w5(32'hbbc67415),
	.w6(32'h3b2cc281),
	.w7(32'h3a774231),
	.w8(32'hb9811477),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb325262),
	.w1(32'h3a41dc63),
	.w2(32'h3af63eeb),
	.w3(32'h3a9f50e8),
	.w4(32'hbb543ac5),
	.w5(32'h3bba2ce2),
	.w6(32'h3bcb4e63),
	.w7(32'hbb1ef71e),
	.w8(32'h3a379a5d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86afc5),
	.w1(32'hbba459cd),
	.w2(32'h3c34104b),
	.w3(32'h3c1a700b),
	.w4(32'h3a3ac3c1),
	.w5(32'h3aa8a32f),
	.w6(32'h3b808897),
	.w7(32'h3c713eb4),
	.w8(32'hbb2c9436),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23162),
	.w1(32'hba632b74),
	.w2(32'hbb4d0b76),
	.w3(32'hba49f7ba),
	.w4(32'h3c09e05e),
	.w5(32'h3ba50021),
	.w6(32'h3b5a74bf),
	.w7(32'hbb23894b),
	.w8(32'h3b5b0bc1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1851),
	.w1(32'h3cb49456),
	.w2(32'h3c8cd415),
	.w3(32'h3c28679c),
	.w4(32'h39591189),
	.w5(32'hbb9639f2),
	.w6(32'h3aaa4abd),
	.w7(32'h396d39c4),
	.w8(32'hbb5b25a9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6691ea),
	.w1(32'h3b4b1343),
	.w2(32'h3a4e1cfd),
	.w3(32'h3b46de13),
	.w4(32'hbc0d5e18),
	.w5(32'h3b16ee2c),
	.w6(32'h3c3b71bd),
	.w7(32'hbb8a2a6b),
	.w8(32'h3bf091fd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba979b4e),
	.w1(32'h3b12221a),
	.w2(32'h3a0ef8a2),
	.w3(32'h3c2de3a1),
	.w4(32'hbb30c9b0),
	.w5(32'hbaa763fb),
	.w6(32'hbc3e43d8),
	.w7(32'hbb1df18b),
	.w8(32'h3c44552c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0a4f8),
	.w1(32'h3ba9dea1),
	.w2(32'hb9aedcef),
	.w3(32'hbb4ed1bc),
	.w4(32'h3b8564e4),
	.w5(32'h38b646bd),
	.w6(32'hbb8e3bae),
	.w7(32'h3bf845df),
	.w8(32'h3b38b495),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82223b),
	.w1(32'hbb6e0045),
	.w2(32'h3bae1f0e),
	.w3(32'h3b927609),
	.w4(32'hba22bf95),
	.w5(32'h3c0cae7a),
	.w6(32'hb8ad45c0),
	.w7(32'h3b63d56a),
	.w8(32'h3c0718d7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906849d),
	.w1(32'h3c377d06),
	.w2(32'h3c87afa0),
	.w3(32'hbb00a1fc),
	.w4(32'h3d17cb70),
	.w5(32'hbb0cf936),
	.w6(32'hb9498b58),
	.w7(32'hbb0ded38),
	.w8(32'hbc2b832e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bf532),
	.w1(32'h3bb017d3),
	.w2(32'h38aa5d82),
	.w3(32'hbb304613),
	.w4(32'hbb1738df),
	.w5(32'h3b4ef0dd),
	.w6(32'h3c57eefb),
	.w7(32'h3bdb8726),
	.w8(32'h3bcba485),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8145ed),
	.w1(32'h3c68292a),
	.w2(32'hbb6b0cef),
	.w3(32'h3b7fec44),
	.w4(32'h3b8d79e2),
	.w5(32'h3a8955e5),
	.w6(32'hbbc11871),
	.w7(32'h3c687693),
	.w8(32'hb99e1dd0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0e619),
	.w1(32'h3ba86cfe),
	.w2(32'h3c04607b),
	.w3(32'h3b77f043),
	.w4(32'h3a227609),
	.w5(32'h3b7c4779),
	.w6(32'h3c1cb7bd),
	.w7(32'h3aba6a45),
	.w8(32'hbb91f645),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0555a1),
	.w1(32'hbb9ad654),
	.w2(32'h3b710ddc),
	.w3(32'hbbe52564),
	.w4(32'hba91caee),
	.w5(32'hbba584ab),
	.w6(32'hbb994cdc),
	.w7(32'h3b3077a1),
	.w8(32'hbab1f07d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4cbe8),
	.w1(32'hbbdddb3d),
	.w2(32'hbaf07697),
	.w3(32'h3bb6ac80),
	.w4(32'hbbb079f4),
	.w5(32'h3cd82dbb),
	.w6(32'hbb39171a),
	.w7(32'h3c057b06),
	.w8(32'hbbed0b63),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afa4d3),
	.w1(32'h3a27dc95),
	.w2(32'h3bfc6322),
	.w3(32'hbb866250),
	.w4(32'h3bbac1ad),
	.w5(32'hbb05bcfc),
	.w6(32'hbb83780f),
	.w7(32'hb97e3f96),
	.w8(32'hbb621971),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f3f8),
	.w1(32'hbbdf7d8c),
	.w2(32'hbad27ebd),
	.w3(32'h36136ec8),
	.w4(32'h3c16dedd),
	.w5(32'hbb1ac9b8),
	.w6(32'h3bf367a1),
	.w7(32'hbbb68243),
	.w8(32'hba25a019),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e910),
	.w1(32'h3b988ffd),
	.w2(32'hbb159a64),
	.w3(32'hbbffefd7),
	.w4(32'hba18e510),
	.w5(32'h3c03c2c5),
	.w6(32'h3c6c6d5f),
	.w7(32'hb9d6560a),
	.w8(32'hbbdf051e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7acac),
	.w1(32'hbb4ad785),
	.w2(32'h3a8d4ede),
	.w3(32'hbb3fca21),
	.w4(32'h3b78fde5),
	.w5(32'hba3f6194),
	.w6(32'hbb90e634),
	.w7(32'hbba358bc),
	.w8(32'hb9ae8a41),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dfba2),
	.w1(32'hbc0380f5),
	.w2(32'h3b740d1a),
	.w3(32'hba2ec0ea),
	.w4(32'h3b5df826),
	.w5(32'hbbbb7353),
	.w6(32'hbb29b1f8),
	.w7(32'hb9db7fa2),
	.w8(32'h3af6ec6c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0618b),
	.w1(32'hbb4eb305),
	.w2(32'hbb356a09),
	.w3(32'hbc2d07d5),
	.w4(32'h39f2aeb3),
	.w5(32'h3bf1d56a),
	.w6(32'h3b278408),
	.w7(32'hbabc7178),
	.w8(32'hba8a9b17),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc424ca4),
	.w1(32'h3be32f5d),
	.w2(32'h3c182001),
	.w3(32'hba832246),
	.w4(32'hbb46bdd6),
	.w5(32'hbb817e28),
	.w6(32'h3a5fe3dc),
	.w7(32'hbb2d662d),
	.w8(32'h3b0e4357),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6da48e),
	.w1(32'h3c110f4c),
	.w2(32'h3be77ac5),
	.w3(32'h3ce61cea),
	.w4(32'h3c49ff5c),
	.w5(32'h3c1e4644),
	.w6(32'hbbef44da),
	.w7(32'hbc4d8531),
	.w8(32'hbb19b7e5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbfc66),
	.w1(32'h398f2191),
	.w2(32'hbb9a836c),
	.w3(32'hbb16fb08),
	.w4(32'hbb394714),
	.w5(32'h3c45a5d6),
	.w6(32'h3bbcec58),
	.w7(32'hbc13c76c),
	.w8(32'hbb21e717),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4488b),
	.w1(32'hbb5d48f9),
	.w2(32'h3b9513e0),
	.w3(32'h3ba4b7e3),
	.w4(32'hb9ac82e8),
	.w5(32'h3c1a36d5),
	.w6(32'h3bcac2a4),
	.w7(32'h3b8ee326),
	.w8(32'hbc0449b9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144e1a),
	.w1(32'h3b61969b),
	.w2(32'hbaa0fa67),
	.w3(32'h3a685651),
	.w4(32'h3b7bd50f),
	.w5(32'hbb334e2e),
	.w6(32'h3c344c6d),
	.w7(32'h3b3e52b0),
	.w8(32'h3a8b3603),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbf741),
	.w1(32'hbb3d113f),
	.w2(32'h38adda0c),
	.w3(32'hbb3d45ce),
	.w4(32'h3bdd6f02),
	.w5(32'h3bb68584),
	.w6(32'hbb45a929),
	.w7(32'h3b811f8d),
	.w8(32'h38982860),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b742c3),
	.w1(32'hbb0aca30),
	.w2(32'hbb903a10),
	.w3(32'hbb9f31ce),
	.w4(32'hbb1fabc1),
	.w5(32'hb9b721c7),
	.w6(32'hbb20aea5),
	.w7(32'hba9fc8b8),
	.w8(32'h3b12cb69),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ade3e),
	.w1(32'hbba53da8),
	.w2(32'h3b82ca4e),
	.w3(32'hbc15c088),
	.w4(32'h3bb0aa1b),
	.w5(32'h3b567975),
	.w6(32'hba3df1f3),
	.w7(32'h3b912f55),
	.w8(32'hb9e93480),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c410dce),
	.w1(32'hbb923533),
	.w2(32'h3b6a410f),
	.w3(32'hbc1b1414),
	.w4(32'hbb38bf09),
	.w5(32'h39ee0621),
	.w6(32'h39245a2c),
	.w7(32'hbb65373d),
	.w8(32'hba19bd6b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c209),
	.w1(32'h3c9b87fe),
	.w2(32'h3b9bed47),
	.w3(32'hbab4e6aa),
	.w4(32'hbb0908e2),
	.w5(32'hbb6b6fe1),
	.w6(32'hbb4dee92),
	.w7(32'hb9b3a6ca),
	.w8(32'h3b2b8973),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976ee7f),
	.w1(32'h39b22a6f),
	.w2(32'hbb684366),
	.w3(32'hba69e392),
	.w4(32'hba9665ba),
	.w5(32'hbaa186fe),
	.w6(32'hbadc7cf0),
	.w7(32'h34c05a39),
	.w8(32'hba8647f6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7fa68),
	.w1(32'hbc156a72),
	.w2(32'hbbd078eb),
	.w3(32'hbb057ba3),
	.w4(32'hbbbec0d6),
	.w5(32'hbc12aac6),
	.w6(32'h3997b352),
	.w7(32'hbb678492),
	.w8(32'hb9dd1e75),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea4a15),
	.w1(32'hba814564),
	.w2(32'h3ba2b116),
	.w3(32'h3c8e6163),
	.w4(32'h3b8f2727),
	.w5(32'hbb2eba7c),
	.w6(32'h3b8d5ac4),
	.w7(32'h3b84dc74),
	.w8(32'hbbead192),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aca58),
	.w1(32'hbaa1d35b),
	.w2(32'hbaf1633a),
	.w3(32'hbb3c6cc8),
	.w4(32'h3c4f9f78),
	.w5(32'h3c0e1fbc),
	.w6(32'hbb831d6a),
	.w7(32'hbbab2992),
	.w8(32'hbbad2bfa),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32b60),
	.w1(32'hbb0c0930),
	.w2(32'hbb23b493),
	.w3(32'hbc294352),
	.w4(32'hbc571356),
	.w5(32'hbb5b9787),
	.w6(32'hbb4b7e94),
	.w7(32'hbb909e2d),
	.w8(32'h3c600fbc),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92be5bd),
	.w1(32'hba1b35dc),
	.w2(32'hb92b2652),
	.w3(32'hbb27cb3b),
	.w4(32'h3b9d2aca),
	.w5(32'hbb5fa60e),
	.w6(32'hbac396ec),
	.w7(32'h3c06d98e),
	.w8(32'hbbe73095),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13a8ba),
	.w1(32'h3c6dbbb4),
	.w2(32'h3b62dd8f),
	.w3(32'hbae7d7a4),
	.w4(32'hb995958b),
	.w5(32'h3a951b4b),
	.w6(32'hbb858f2b),
	.w7(32'hbac158b3),
	.w8(32'h3b30db82),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7b73),
	.w1(32'hbb8d5024),
	.w2(32'h3bbb9a49),
	.w3(32'h3be26cf0),
	.w4(32'hbbb1c2b2),
	.w5(32'h3b6c4637),
	.w6(32'hbb2c5293),
	.w7(32'h3b707df7),
	.w8(32'hbb87a801),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf729b),
	.w1(32'hbbc473ed),
	.w2(32'hbc335eab),
	.w3(32'h3b0d4d99),
	.w4(32'h3b3d8e65),
	.w5(32'h3be00c53),
	.w6(32'h3bed32f0),
	.w7(32'h3c0a90b1),
	.w8(32'hb8d50b7c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910482a),
	.w1(32'h3b7a1964),
	.w2(32'h3cb67afd),
	.w3(32'hbc77ada1),
	.w4(32'hba0e631b),
	.w5(32'h3ba10b84),
	.w6(32'hb9ac50f7),
	.w7(32'h3d0907f9),
	.w8(32'hbb4e8917),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db4fa),
	.w1(32'h3c4aa29e),
	.w2(32'h3bb61fe1),
	.w3(32'h3b89c58a),
	.w4(32'hbb1ddcd7),
	.w5(32'hbaa84e7c),
	.w6(32'h3a3c157c),
	.w7(32'h3b9951f2),
	.w8(32'h3b31ecdc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22c0ef),
	.w1(32'hb9fc5ae8),
	.w2(32'h39e940a4),
	.w3(32'hb981791d),
	.w4(32'hb9e4bc27),
	.w5(32'hb911dd6c),
	.w6(32'h38c8a7cb),
	.w7(32'hbac8aa21),
	.w8(32'h3c4bb45d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfc9fd),
	.w1(32'hbb7df311),
	.w2(32'hb9f43f61),
	.w3(32'h3b68e296),
	.w4(32'hb97a84a3),
	.w5(32'hbaad9521),
	.w6(32'hba621843),
	.w7(32'hba43f45c),
	.w8(32'h3a9f096d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18cdc3),
	.w1(32'h3b025d68),
	.w2(32'h39e5b5eb),
	.w3(32'hba85b444),
	.w4(32'hbac084c3),
	.w5(32'hbb396688),
	.w6(32'h3a867da8),
	.w7(32'hbbc298c6),
	.w8(32'hbadabf1f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ce95c),
	.w1(32'h3b455594),
	.w2(32'hba05b2bf),
	.w3(32'hbb16c0dc),
	.w4(32'hbb93a56e),
	.w5(32'hbbce5c22),
	.w6(32'h3a526cf2),
	.w7(32'hbaa4003b),
	.w8(32'h3b1f2737),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2ff53),
	.w1(32'hb98ca021),
	.w2(32'h39ce022b),
	.w3(32'hb893c717),
	.w4(32'hba199142),
	.w5(32'hbb019adc),
	.w6(32'hba4e5fe6),
	.w7(32'hb9ffac5a),
	.w8(32'h395ae2bb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81af5b),
	.w1(32'hbaf4aefa),
	.w2(32'h39a0142d),
	.w3(32'hba44b731),
	.w4(32'h3b14a545),
	.w5(32'h39c7f176),
	.w6(32'hbb117f5d),
	.w7(32'hbb94fbc2),
	.w8(32'hb8989eb5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e27eb),
	.w1(32'h391ccec2),
	.w2(32'hba9f3ab2),
	.w3(32'hbaf3d923),
	.w4(32'hbb8e0132),
	.w5(32'hbc366c7e),
	.w6(32'hbac97e84),
	.w7(32'hbb4ed39f),
	.w8(32'h3aae494f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23fd9b),
	.w1(32'h3a83ee6a),
	.w2(32'h39d14bad),
	.w3(32'hbb3e07c5),
	.w4(32'h3a7d3937),
	.w5(32'h3ad86298),
	.w6(32'h3a0b1dbd),
	.w7(32'h3a351c6a),
	.w8(32'hbb50b4d3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6f7fe),
	.w1(32'h3c79ad48),
	.w2(32'h398254b8),
	.w3(32'hb99e5999),
	.w4(32'h3bb8b9f5),
	.w5(32'hbb0712aa),
	.w6(32'hbab9a7a5),
	.w7(32'h3b181c5b),
	.w8(32'h3ab895de),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03d84),
	.w1(32'h3a736aa7),
	.w2(32'hbaa0f5d4),
	.w3(32'h3b679dbb),
	.w4(32'hbaf654c0),
	.w5(32'hbb0a56bf),
	.w6(32'hbb63e37c),
	.w7(32'hbb4f8608),
	.w8(32'h3c240c30),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bd38f),
	.w1(32'hbae606ec),
	.w2(32'h39f8fd7b),
	.w3(32'hbad6b7c2),
	.w4(32'hb55f2480),
	.w5(32'hbb280718),
	.w6(32'hbbbf4ec4),
	.w7(32'hbbb9f5b9),
	.w8(32'h37e7d561),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989ce0e),
	.w1(32'hba8d948f),
	.w2(32'h39b8a81c),
	.w3(32'hbbaaee0e),
	.w4(32'h3ab599a1),
	.w5(32'h3a9cb829),
	.w6(32'h3a477daf),
	.w7(32'hbb1d665f),
	.w8(32'hba6be948),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d2fe),
	.w1(32'hbbe7a4ff),
	.w2(32'h39df5424),
	.w3(32'hbb121ca2),
	.w4(32'hbae258f5),
	.w5(32'h3ac96e8e),
	.w6(32'h3a57a1eb),
	.w7(32'hbb206c62),
	.w8(32'h39a0da4b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99f2c7),
	.w1(32'h397bcb65),
	.w2(32'h3b36e83c),
	.w3(32'hb9602375),
	.w4(32'hbab24707),
	.w5(32'hba3b7a72),
	.w6(32'hbb9180af),
	.w7(32'hbb81ae1b),
	.w8(32'hbacb382e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a190c91),
	.w1(32'h3b3982cf),
	.w2(32'hbb14432b),
	.w3(32'hbb44ef10),
	.w4(32'hb9c191d5),
	.w5(32'hbb7367ec),
	.w6(32'hbaa4c6dd),
	.w7(32'h3cc3d775),
	.w8(32'hbb877ba2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eac8b9),
	.w1(32'hba4d150a),
	.w2(32'h3ac26899),
	.w3(32'h3be51a97),
	.w4(32'h3ad33b29),
	.w5(32'hba7bd4a3),
	.w6(32'hbc00905e),
	.w7(32'h3a41e35b),
	.w8(32'h3a0e18af),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb683b),
	.w1(32'hbb010070),
	.w2(32'h3b9211ac),
	.w3(32'hbae80ec9),
	.w4(32'hbaab5a2c),
	.w5(32'hb843c342),
	.w6(32'hbaeea151),
	.w7(32'hb82b60e9),
	.w8(32'h3a24dddb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30c9ce),
	.w1(32'h3aa2f531),
	.w2(32'hba3aeda0),
	.w3(32'hbb1350e7),
	.w4(32'h3c80ab50),
	.w5(32'h3a9a577e),
	.w6(32'hba7a2ab0),
	.w7(32'h3b59c571),
	.w8(32'h3c8aedcd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78fae68),
	.w1(32'hbc01caed),
	.w2(32'h3b86e193),
	.w3(32'h3a1d8aa8),
	.w4(32'hbb246c1f),
	.w5(32'hbacece2f),
	.w6(32'hbac60633),
	.w7(32'hbaf1b174),
	.w8(32'hbbe18912),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e99e21),
	.w1(32'h38560d06),
	.w2(32'hba840035),
	.w3(32'hb9cb8376),
	.w4(32'h3b1f09e2),
	.w5(32'hbaf211ba),
	.w6(32'h39e4f758),
	.w7(32'h3c5787bf),
	.w8(32'hba42bb04),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a534498),
	.w1(32'hbb10ab52),
	.w2(32'hba8003c6),
	.w3(32'hba8d609b),
	.w4(32'h3ac54fc2),
	.w5(32'hbaad42e0),
	.w6(32'h3a7f30b2),
	.w7(32'h3a7d3ff8),
	.w8(32'hba0521bd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e21dc),
	.w1(32'hba9ebae4),
	.w2(32'hbb384d60),
	.w3(32'hba86e017),
	.w4(32'hbb3dcc1a),
	.w5(32'hbacf909b),
	.w6(32'hbaefaa41),
	.w7(32'h3aa023a5),
	.w8(32'hb98af37b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0d5b2),
	.w1(32'h38a25cd3),
	.w2(32'hb920398b),
	.w3(32'hb904ae69),
	.w4(32'hba43ab34),
	.w5(32'hbab3caf4),
	.w6(32'hba05cabb),
	.w7(32'h3c155a6e),
	.w8(32'h396d0385),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a959b96),
	.w1(32'hba4abe3d),
	.w2(32'h3b0fdf0b),
	.w3(32'hb8efbd01),
	.w4(32'h3a3dd999),
	.w5(32'hba363483),
	.w6(32'hbae1c9cc),
	.w7(32'hbb287118),
	.w8(32'h370ada9c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989e405),
	.w1(32'hbc68e443),
	.w2(32'h3990c1fd),
	.w3(32'hbb13798e),
	.w4(32'hbb457fe8),
	.w5(32'h3b14add3),
	.w6(32'hbba2a78c),
	.w7(32'h3a15f363),
	.w8(32'h3abb5c2f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810b5d),
	.w1(32'h3993b1bf),
	.w2(32'hb9943ab0),
	.w3(32'hba55ddc0),
	.w4(32'h3a5a96d4),
	.w5(32'hbb53d131),
	.w6(32'hbaa9be9c),
	.w7(32'hb8f2db00),
	.w8(32'hbb3864d2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f0ff2),
	.w1(32'h3accc439),
	.w2(32'hbb9105ee),
	.w3(32'hbab99442),
	.w4(32'hba78cf63),
	.w5(32'hbb17f79a),
	.w6(32'h3be3415d),
	.w7(32'hbb3f0ba4),
	.w8(32'h39514127),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96ac43),
	.w1(32'hbb434e37),
	.w2(32'hbaab39ac),
	.w3(32'h3ab90613),
	.w4(32'h3b782b6a),
	.w5(32'h3a574f68),
	.w6(32'h3a2ff615),
	.w7(32'h3b88fe74),
	.w8(32'h3a274aa9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92564a),
	.w1(32'h3b33d2d5),
	.w2(32'h3aa86b4d),
	.w3(32'hb87359e1),
	.w4(32'h3ab9582e),
	.w5(32'h397d3434),
	.w6(32'hba734f2c),
	.w7(32'h3ae8b841),
	.w8(32'hba5b6c4c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ef01d),
	.w1(32'h3c7d3b89),
	.w2(32'hbb0d473a),
	.w3(32'hbae61c31),
	.w4(32'hbab52832),
	.w5(32'h391f650b),
	.w6(32'hbab4f0e0),
	.w7(32'hba2aaef1),
	.w8(32'h3b36c137),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule