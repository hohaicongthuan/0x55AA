module layer_10_featuremap_368(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc154c52),
	.w1(32'h3c0d6a59),
	.w2(32'h3c66094c),
	.w3(32'hbbb11b0d),
	.w4(32'hb99e8302),
	.w5(32'h3ca2367d),
	.w6(32'h3b807269),
	.w7(32'h3b1be681),
	.w8(32'hbb06c37f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce33c0a),
	.w1(32'hbb451a8c),
	.w2(32'hbcc2de36),
	.w3(32'h3b0fd063),
	.w4(32'h3bcaa474),
	.w5(32'hbbb910b6),
	.w6(32'h3b0bad50),
	.w7(32'hba9cadd7),
	.w8(32'hb96cc95a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cb469),
	.w1(32'hbab2e44b),
	.w2(32'hb933970d),
	.w3(32'hbc97ebc3),
	.w4(32'h3b64e6b9),
	.w5(32'h3a13bc89),
	.w6(32'h3d8e5145),
	.w7(32'h3b59fbef),
	.w8(32'hbb2570b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59cf20),
	.w1(32'hbc1ec571),
	.w2(32'hbb022559),
	.w3(32'hbd29186f),
	.w4(32'hbc14d75f),
	.w5(32'hbbda08c2),
	.w6(32'h3c3d6800),
	.w7(32'h3c645cce),
	.w8(32'hbb7c620f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50ca7),
	.w1(32'h3b38d073),
	.w2(32'hbbb518dc),
	.w3(32'hbc567268),
	.w4(32'h3bc2d5eb),
	.w5(32'hba072629),
	.w6(32'h392d687c),
	.w7(32'hbb5ba0eb),
	.w8(32'hbc87f270),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c83b),
	.w1(32'hbbffa38c),
	.w2(32'h3aa286fa),
	.w3(32'hba8f45b2),
	.w4(32'h3b2471b5),
	.w5(32'h3c737c4a),
	.w6(32'h3ad9d6df),
	.w7(32'hbbb19628),
	.w8(32'h3b97de1a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be20918),
	.w1(32'h3b4b35c0),
	.w2(32'h3b2f32d2),
	.w3(32'h3994ec15),
	.w4(32'h3c814aab),
	.w5(32'h3c510769),
	.w6(32'hbaadedcf),
	.w7(32'hbc455449),
	.w8(32'h3c9548e3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9c8e9),
	.w1(32'h388e635b),
	.w2(32'h3b82be76),
	.w3(32'hbc8504d8),
	.w4(32'hbb15340c),
	.w5(32'h3b944281),
	.w6(32'hbc033016),
	.w7(32'hbb99c1b1),
	.w8(32'h3c0ef8a4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdc82d),
	.w1(32'hbbc3d4fb),
	.w2(32'h3b833e01),
	.w3(32'hbbe0812a),
	.w4(32'hbc0c8557),
	.w5(32'h39e11902),
	.w6(32'h3a0b24ec),
	.w7(32'h3c1e42f4),
	.w8(32'h386ed418),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd11cb81),
	.w1(32'hbb7d1752),
	.w2(32'h3c00fb23),
	.w3(32'h3c38b482),
	.w4(32'h3b6c2458),
	.w5(32'hbc11bfa2),
	.w6(32'hbb83a4e9),
	.w7(32'hbc87b74a),
	.w8(32'hba9c371d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0422a7),
	.w1(32'hbbed755f),
	.w2(32'h3b8859d8),
	.w3(32'hbc35ad46),
	.w4(32'h3c60338e),
	.w5(32'h3c325e28),
	.w6(32'hbb37710c),
	.w7(32'hbb6f39f2),
	.w8(32'h3b46553f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6673a),
	.w1(32'hbab63fb0),
	.w2(32'hbd978884),
	.w3(32'hbad20db6),
	.w4(32'hbd48264a),
	.w5(32'hba5f36b7),
	.w6(32'hba95e2c1),
	.w7(32'hb82519d8),
	.w8(32'h3b820866),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1992c7),
	.w1(32'h3a942cae),
	.w2(32'h3c3e28cf),
	.w3(32'hba499e99),
	.w4(32'h3c034d50),
	.w5(32'h3c525b46),
	.w6(32'hb91d3708),
	.w7(32'h3bde586d),
	.w8(32'hbc75202b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a186bf4),
	.w1(32'hbd2e9767),
	.w2(32'h3b285bc4),
	.w3(32'hbc012f5d),
	.w4(32'h3c8b34da),
	.w5(32'hbadbb059),
	.w6(32'hbc8048e6),
	.w7(32'h3b88df4d),
	.w8(32'hbc3d9e46),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca299a2),
	.w1(32'h3c0e6c00),
	.w2(32'hba85efdb),
	.w3(32'h3a1a5381),
	.w4(32'hbc838866),
	.w5(32'h39cdaa79),
	.w6(32'hbb5c30eb),
	.w7(32'hbb4b3e78),
	.w8(32'h3a9dd04a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8204ea),
	.w1(32'h3b3301b6),
	.w2(32'h3c25c61c),
	.w3(32'h3c924b34),
	.w4(32'h39d96f4a),
	.w5(32'hbbdd9733),
	.w6(32'h3b68c61b),
	.w7(32'hbbe41088),
	.w8(32'hbb9534c3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdfa3a),
	.w1(32'h39ad12b9),
	.w2(32'h3b8a87e2),
	.w3(32'h3ab4eb43),
	.w4(32'h3a703d46),
	.w5(32'hbc29addc),
	.w6(32'hbb30c042),
	.w7(32'hbba5fd92),
	.w8(32'h3a90483d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a268),
	.w1(32'hbb8ef0a3),
	.w2(32'hbc448767),
	.w3(32'hbb6e8894),
	.w4(32'hba968058),
	.w5(32'hbb6b0fec),
	.w6(32'hbb71b17f),
	.w7(32'hbc99d2c6),
	.w8(32'hbb1ec13c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092ecf),
	.w1(32'hbb87eaaf),
	.w2(32'hb907d3da),
	.w3(32'hbb78aa35),
	.w4(32'hbbdaa431),
	.w5(32'h3c7f7d76),
	.w6(32'h3b16e746),
	.w7(32'hbacd9e86),
	.w8(32'hbbed59da),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc1762),
	.w1(32'hbc04e35b),
	.w2(32'h3b315b8f),
	.w3(32'h3b0c9bd6),
	.w4(32'h3c26f987),
	.w5(32'hbb5fc558),
	.w6(32'hbca8a8df),
	.w7(32'hbb8725d7),
	.w8(32'hba1a5abf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08b288),
	.w1(32'hba9f0b66),
	.w2(32'hb93da115),
	.w3(32'h3b62bb1e),
	.w4(32'hbbe65484),
	.w5(32'h3af44c28),
	.w6(32'h3b70e189),
	.w7(32'h3bcd0da2),
	.w8(32'hbc293fd0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd082829),
	.w1(32'hbc835d3d),
	.w2(32'h3b5f4191),
	.w3(32'h3b9ff633),
	.w4(32'h3ba0d63c),
	.w5(32'hbc5e9c10),
	.w6(32'hbc3dec44),
	.w7(32'h3b826a5f),
	.w8(32'hbbe30b32),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea3af5),
	.w1(32'h39dd0e9c),
	.w2(32'h3b8ad269),
	.w3(32'hba657850),
	.w4(32'h39086e56),
	.w5(32'h3c744e28),
	.w6(32'h3bd278f9),
	.w7(32'h3bcebc35),
	.w8(32'hbc84356a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38e6e),
	.w1(32'hbc4940e1),
	.w2(32'hbc00bbf4),
	.w3(32'h3bf3e807),
	.w4(32'hbbe10c4a),
	.w5(32'hb9892189),
	.w6(32'hbc0d065b),
	.w7(32'hbcc49f26),
	.w8(32'h3acaa766),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc019883),
	.w1(32'h3aad9f17),
	.w2(32'h3b72533c),
	.w3(32'h3b908314),
	.w4(32'hb91722c8),
	.w5(32'hbb63726a),
	.w6(32'hba2c5124),
	.w7(32'hbaa80992),
	.w8(32'hbb0faaca),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12fdcc),
	.w1(32'hbb347adc),
	.w2(32'h3c5604ad),
	.w3(32'hbc8bc3d2),
	.w4(32'hbc71feaa),
	.w5(32'h3aa4dbf8),
	.w6(32'h3a4c823a),
	.w7(32'hbc72b050),
	.w8(32'hb863de7f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15679d),
	.w1(32'hba780e4a),
	.w2(32'hb7dd3e5f),
	.w3(32'h3bce2ee5),
	.w4(32'hbbce214c),
	.w5(32'h3a501dda),
	.w6(32'hbb79c94d),
	.w7(32'hbb7cba46),
	.w8(32'hbaf1c032),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b9ed),
	.w1(32'h39cb811e),
	.w2(32'hbac4b02d),
	.w3(32'hbbddae4e),
	.w4(32'hbad1510d),
	.w5(32'hbb86a70d),
	.w6(32'h3a55f62f),
	.w7(32'h3b28ea31),
	.w8(32'h3a77ace7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c254e1c),
	.w1(32'hbc0d8ed0),
	.w2(32'h3b043028),
	.w3(32'hbc04ecd1),
	.w4(32'hbb1c8fda),
	.w5(32'h3b6aa475),
	.w6(32'h3b007984),
	.w7(32'hbb93dd37),
	.w8(32'hbb814fb2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0a1f),
	.w1(32'hbbbdb8a3),
	.w2(32'hbb1b421c),
	.w3(32'hbbf80477),
	.w4(32'h3b7b1181),
	.w5(32'hbb2e1294),
	.w6(32'h3b9e709f),
	.w7(32'hbb78d3f8),
	.w8(32'hbbd0f91d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc376a33),
	.w1(32'h3a5cb628),
	.w2(32'h3c4503bd),
	.w3(32'h3aff14d4),
	.w4(32'h3b1ef9dd),
	.w5(32'h3c1aaa09),
	.w6(32'hb9c8188e),
	.w7(32'hbc701d60),
	.w8(32'h3c2cb445),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78c730f),
	.w1(32'hb9c4143c),
	.w2(32'hba3aefa4),
	.w3(32'hbc7e086d),
	.w4(32'hbb767cc8),
	.w5(32'hbcbf055f),
	.w6(32'h3bf78d98),
	.w7(32'hbc904a48),
	.w8(32'hbc5178fe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0799df),
	.w1(32'h3be6ba4e),
	.w2(32'hbc36e20f),
	.w3(32'h3a1e9166),
	.w4(32'hbb6b7343),
	.w5(32'h3bda9cc2),
	.w6(32'h3be244c4),
	.w7(32'hbbc630d9),
	.w8(32'hbba4ed8b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06ac7a),
	.w1(32'h3b601274),
	.w2(32'h3c261eb9),
	.w3(32'hbb1f492c),
	.w4(32'hbb9d297a),
	.w5(32'h3bf963fc),
	.w6(32'h3989c2ca),
	.w7(32'hbad3f700),
	.w8(32'hbad47a86),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb680f),
	.w1(32'hbc19ac88),
	.w2(32'hbbafb5b0),
	.w3(32'h3b9c0bb0),
	.w4(32'h3b11d8a3),
	.w5(32'hbbdb1ef2),
	.w6(32'hbb4547a5),
	.w7(32'hbc5d35eb),
	.w8(32'hbc84407b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395669d8),
	.w1(32'h3ad680ac),
	.w2(32'hbbb3cf4a),
	.w3(32'hbab529ef),
	.w4(32'hbc0c488f),
	.w5(32'h3ab7845b),
	.w6(32'hbc122fa1),
	.w7(32'h3b093372),
	.w8(32'hbc0f2eff),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b5b7),
	.w1(32'h3c1e749e),
	.w2(32'hbbffd9fc),
	.w3(32'h3b319e4d),
	.w4(32'h3b229e27),
	.w5(32'hb9923497),
	.w6(32'hbb2ccdfc),
	.w7(32'hbb705330),
	.w8(32'hbc0c507f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54a768),
	.w1(32'hbb5b92a4),
	.w2(32'h3ae16451),
	.w3(32'h3d18fbe5),
	.w4(32'h3c10287a),
	.w5(32'hb981e7a6),
	.w6(32'h3ae89f04),
	.w7(32'h3b49f877),
	.w8(32'hbb8fafbb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39605c01),
	.w1(32'hbb0942f9),
	.w2(32'h3b9b30da),
	.w3(32'hbc6608f2),
	.w4(32'hbb4ba229),
	.w5(32'h3be5728c),
	.w6(32'hbb8a35e0),
	.w7(32'hba895036),
	.w8(32'h3b08ce53),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54ef29),
	.w1(32'hbc3d1d3d),
	.w2(32'hbb37f3e8),
	.w3(32'h3b27b669),
	.w4(32'h3b4c5029),
	.w5(32'hbb3caa36),
	.w6(32'hbb8e7348),
	.w7(32'hbb2910c3),
	.w8(32'hbb989272),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b02cd4),
	.w1(32'hbb2d2784),
	.w2(32'hbc421d2f),
	.w3(32'hbc87e4e1),
	.w4(32'hbc8d6fbb),
	.w5(32'hbc0541c3),
	.w6(32'hbb65bde7),
	.w7(32'hbc354243),
	.w8(32'hbafb4d77),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee49d),
	.w1(32'hbb17fefe),
	.w2(32'hbb5f89a6),
	.w3(32'hbb12010f),
	.w4(32'hbb13bf17),
	.w5(32'hbc985f0e),
	.w6(32'hbc155fa6),
	.w7(32'hbc379409),
	.w8(32'hbc1583e0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ad51b),
	.w1(32'h3c10841b),
	.w2(32'h3b784279),
	.w3(32'h3c0c5256),
	.w4(32'hbc20fff5),
	.w5(32'h3b445c7f),
	.w6(32'h3b85dff5),
	.w7(32'hbad58f37),
	.w8(32'hbc00f5d0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b3f2),
	.w1(32'h3a0e1abb),
	.w2(32'h3c35a1e9),
	.w3(32'hbb03e64e),
	.w4(32'h3a16c5ba),
	.w5(32'hbb08a74e),
	.w6(32'hbaa93865),
	.w7(32'h3bc964ec),
	.w8(32'hba76c4c3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1de6f4),
	.w1(32'hb9ef3018),
	.w2(32'h3c241a00),
	.w3(32'h3b316ed2),
	.w4(32'h3c1b5514),
	.w5(32'hbcbf07c6),
	.w6(32'h39ce5d23),
	.w7(32'hbb1da81e),
	.w8(32'h3a192e6f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5e12b),
	.w1(32'hbbd084b8),
	.w2(32'h3bd5b450),
	.w3(32'hbc397e91),
	.w4(32'hbbeb58fa),
	.w5(32'hbb89e888),
	.w6(32'h3a6ec9d6),
	.w7(32'h3b8968b0),
	.w8(32'h3b1c027a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86b4cf),
	.w1(32'h3b1020da),
	.w2(32'hbc1a7ed2),
	.w3(32'h3b7c6c31),
	.w4(32'h3a49ff2e),
	.w5(32'hbc422b21),
	.w6(32'h3bb6ff80),
	.w7(32'h3ac500b1),
	.w8(32'h3949cea7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39888208),
	.w1(32'hbaebaf45),
	.w2(32'h3bd8c90c),
	.w3(32'hbac67a61),
	.w4(32'hbbb237f3),
	.w5(32'h3b471699),
	.w6(32'hbbd0277d),
	.w7(32'h3b9dd170),
	.w8(32'h3b2064aa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d98cd9),
	.w1(32'hba989444),
	.w2(32'h3c1e0606),
	.w3(32'hbbc5b2de),
	.w4(32'h3aa039fc),
	.w5(32'h3b571476),
	.w6(32'hbb0812c9),
	.w7(32'hba7ca43d),
	.w8(32'h3bb22f72),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d119f),
	.w1(32'h3b97ff53),
	.w2(32'hbc0aedde),
	.w3(32'h3a154bb8),
	.w4(32'h3b7963a4),
	.w5(32'h3c2a9149),
	.w6(32'h3bd91595),
	.w7(32'h3b5b7abf),
	.w8(32'hbab44363),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b66ff),
	.w1(32'hba98fde5),
	.w2(32'hbb0e54b9),
	.w3(32'h3bb407be),
	.w4(32'h3b448413),
	.w5(32'h3a323330),
	.w6(32'hbc03b1f7),
	.w7(32'h3b2cbeb4),
	.w8(32'hbacaec43),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a354292),
	.w1(32'hba97e478),
	.w2(32'h3ba76cbf),
	.w3(32'hbaf96fc9),
	.w4(32'h387c7694),
	.w5(32'h3afc582f),
	.w6(32'hbc062d05),
	.w7(32'hbb675206),
	.w8(32'hbbfab010),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7972f),
	.w1(32'h3c59c358),
	.w2(32'h3b384860),
	.w3(32'hbbab72e5),
	.w4(32'h39d8481a),
	.w5(32'hbca152fe),
	.w6(32'hba456b68),
	.w7(32'hbbcc45a0),
	.w8(32'hba5f7c07),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa81f0d),
	.w1(32'hbc1b336a),
	.w2(32'hbb43ce24),
	.w3(32'hbb52864d),
	.w4(32'hbbd6a365),
	.w5(32'hbac8125c),
	.w6(32'hbb162e1c),
	.w7(32'hbc81ed6f),
	.w8(32'hbaf2e4c4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6ee4),
	.w1(32'h3c69e16e),
	.w2(32'hbb4f1cfa),
	.w3(32'h3b40b80d),
	.w4(32'h3aa37e43),
	.w5(32'h3bc0b0b4),
	.w6(32'hbbdec060),
	.w7(32'h398d7dfc),
	.w8(32'h3bb80e17),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cf86d),
	.w1(32'hbb45ffa0),
	.w2(32'h3a3b722e),
	.w3(32'hbb14578a),
	.w4(32'h3b059dce),
	.w5(32'hbc069b14),
	.w6(32'hbb101461),
	.w7(32'hb900bc3d),
	.w8(32'h3c29591a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54efe8),
	.w1(32'h3bca88c1),
	.w2(32'hbb4e8f09),
	.w3(32'h3c68e98c),
	.w4(32'hbb59ae30),
	.w5(32'hbb9783ca),
	.w6(32'hbc8bc898),
	.w7(32'hbbbf79f1),
	.w8(32'h3b42bf0b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb0ee),
	.w1(32'hbbc88afe),
	.w2(32'hba664b85),
	.w3(32'h3d24de9a),
	.w4(32'hbb1bebb0),
	.w5(32'h3b6d7563),
	.w6(32'h3b852806),
	.w7(32'h3a1da667),
	.w8(32'h3be95345),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc897cf),
	.w1(32'hbb66a14c),
	.w2(32'h3a22b8f2),
	.w3(32'h393eb6d7),
	.w4(32'hbb8ebfc7),
	.w5(32'h3b872509),
	.w6(32'hbb83fd15),
	.w7(32'hbc8f3b1a),
	.w8(32'h3951a849),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77964f),
	.w1(32'hbc25282f),
	.w2(32'h3be9e62f),
	.w3(32'hbbda404b),
	.w4(32'hb7d21610),
	.w5(32'h3a97e6fc),
	.w6(32'hbba1a3f4),
	.w7(32'h3c03d46b),
	.w8(32'hbc039741),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280813),
	.w1(32'h3bec7b61),
	.w2(32'hba02a7d1),
	.w3(32'hbc237a65),
	.w4(32'h3bf80f8c),
	.w5(32'h3b31d59b),
	.w6(32'hbd080f13),
	.w7(32'hba8700dd),
	.w8(32'hb9dea9e8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce12da0),
	.w1(32'hbc21ea3b),
	.w2(32'hb858b7a0),
	.w3(32'hbc326bc1),
	.w4(32'hbb01d005),
	.w5(32'hbd3c4ceb),
	.w6(32'hbc4d53b8),
	.w7(32'h3be10bf3),
	.w8(32'hbb7b14cf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8119fc),
	.w1(32'h3b5f998b),
	.w2(32'h3c1b5ccb),
	.w3(32'h3b9a42d5),
	.w4(32'hba1a35ef),
	.w5(32'hbbebc20f),
	.w6(32'hbbf534c0),
	.w7(32'h3baf9f2d),
	.w8(32'hbbacb5ce),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21823d),
	.w1(32'h3c1b89d9),
	.w2(32'h3c607ab2),
	.w3(32'hbbae0a08),
	.w4(32'h3bf7ee30),
	.w5(32'hbd069512),
	.w6(32'hba46419c),
	.w7(32'hbb407371),
	.w8(32'h3c0e7a4a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc301f),
	.w1(32'h3b12b5e0),
	.w2(32'h3b62dbbf),
	.w3(32'h3b9c08bf),
	.w4(32'h3bfc3a38),
	.w5(32'hbc621518),
	.w6(32'hb9a47a09),
	.w7(32'h3ba09718),
	.w8(32'hbcbb4af5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7596a4),
	.w1(32'hbc44464f),
	.w2(32'hbbd13d61),
	.w3(32'hbb0a4a7a),
	.w4(32'h3aac5d7c),
	.w5(32'hb9295c9d),
	.w6(32'hbc7c7b9c),
	.w7(32'hbc48aa32),
	.w8(32'h3acaae2e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bbc3a),
	.w1(32'hbbb0e180),
	.w2(32'h3ba6277a),
	.w3(32'hbc88f1d9),
	.w4(32'hbb4421e4),
	.w5(32'h3add204d),
	.w6(32'hbab25908),
	.w7(32'hba5e017c),
	.w8(32'hbc19e326),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2177e),
	.w1(32'hbcd733d0),
	.w2(32'h3cad80f4),
	.w3(32'hbb9ed235),
	.w4(32'hbba59d39),
	.w5(32'h3c288b84),
	.w6(32'hbba8f3a5),
	.w7(32'hba93ead0),
	.w8(32'h3c24c2c4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b933e),
	.w1(32'h3bee9226),
	.w2(32'h3bb4da32),
	.w3(32'hbb1dea5d),
	.w4(32'hb73e9451),
	.w5(32'h3b7e9a8f),
	.w6(32'hbbda1eb1),
	.w7(32'hbc0d1cb6),
	.w8(32'h3ac8e8f0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1bb76),
	.w1(32'hbae3bfa5),
	.w2(32'h3b5f0cd5),
	.w3(32'h3ba0db10),
	.w4(32'hbbacccf0),
	.w5(32'hbc7d9028),
	.w6(32'h3ba54427),
	.w7(32'h3b3b7cdf),
	.w8(32'hbc724d11),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610ec0),
	.w1(32'h3c02256f),
	.w2(32'hbc55257a),
	.w3(32'hbca24065),
	.w4(32'h3b6676d9),
	.w5(32'h3bc8c466),
	.w6(32'hbbf45e80),
	.w7(32'hbc2b685e),
	.w8(32'hbb886dff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b9733),
	.w1(32'hbb12ee5a),
	.w2(32'h3ba21434),
	.w3(32'h3bf1d0b5),
	.w4(32'h3b86f042),
	.w5(32'h3b134a86),
	.w6(32'h3ae3e69b),
	.w7(32'h3bcefeeb),
	.w8(32'h3c27368e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f419c),
	.w1(32'h3b31efac),
	.w2(32'h3a7ffd7c),
	.w3(32'h3ad0eaed),
	.w4(32'hbc0001a4),
	.w5(32'hbcd6b85c),
	.w6(32'h3ba9b8a1),
	.w7(32'h3b684e64),
	.w8(32'hbc3c6782),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510927),
	.w1(32'h39bc3984),
	.w2(32'h3a90f5bd),
	.w3(32'hba7b6909),
	.w4(32'h3abe5eb5),
	.w5(32'hba7c1bc4),
	.w6(32'h3c3e5b64),
	.w7(32'h3bbb1d09),
	.w8(32'h3c8ff899),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f9a0a),
	.w1(32'h3b89fb8d),
	.w2(32'h3887bff3),
	.w3(32'h3a970f52),
	.w4(32'hbcd3bc81),
	.w5(32'hbb839cca),
	.w6(32'hbbbc3a24),
	.w7(32'hbc09b6bf),
	.w8(32'h3c4307f5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883dee),
	.w1(32'h3ab7be15),
	.w2(32'h39cbcbb0),
	.w3(32'h3c3c02cd),
	.w4(32'hbb3b87a2),
	.w5(32'hbb29e228),
	.w6(32'h3c9a7c79),
	.w7(32'hbba6003d),
	.w8(32'h3c32810f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881c2b),
	.w1(32'h3c18db1e),
	.w2(32'h3ba8c9ee),
	.w3(32'h3bacc3eb),
	.w4(32'hbaeab30c),
	.w5(32'h3bb1d2c4),
	.w6(32'hba7ad083),
	.w7(32'h3c6dff9f),
	.w8(32'h3b31d8d8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eedcdf),
	.w1(32'h3b9f8893),
	.w2(32'h3c6265e4),
	.w3(32'h3b9ce0bd),
	.w4(32'h3b976207),
	.w5(32'h3ba8b1b0),
	.w6(32'hbb3de7e2),
	.w7(32'h3c3f9bc5),
	.w8(32'hbb9021ea),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5ac8),
	.w1(32'h3b2d7ff2),
	.w2(32'hbc238fee),
	.w3(32'h3b8ec546),
	.w4(32'hba4236ac),
	.w5(32'h39ec8857),
	.w6(32'h3b965999),
	.w7(32'h3b2efa99),
	.w8(32'hbc03f341),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3b5d6),
	.w1(32'h3b5a3c40),
	.w2(32'h3cc5ef96),
	.w3(32'h3bae7597),
	.w4(32'hbb998807),
	.w5(32'hbb8c82d8),
	.w6(32'hba4ccb3a),
	.w7(32'h3c7d5864),
	.w8(32'hbc92c9a4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb40d3),
	.w1(32'h3b6ca95a),
	.w2(32'hbaba8309),
	.w3(32'hbbf8cb6d),
	.w4(32'hbb53aea2),
	.w5(32'hbbba5591),
	.w6(32'hba8a92ad),
	.w7(32'h3ba91a63),
	.w8(32'h3bb2abdd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1cfc5),
	.w1(32'h3c288221),
	.w2(32'h3b4061c5),
	.w3(32'h3b6dbfb5),
	.w4(32'h3b0088f1),
	.w5(32'h3c77c8d7),
	.w6(32'hbbcc2009),
	.w7(32'h3b42c593),
	.w8(32'h3c805d90),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ed965),
	.w1(32'h3c077984),
	.w2(32'h3b54810c),
	.w3(32'hbb2cbf73),
	.w4(32'h3b0377ea),
	.w5(32'hbbdfa29f),
	.w6(32'hbbce2d05),
	.w7(32'hbad4950e),
	.w8(32'hba9732d5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24830b),
	.w1(32'hbb739a75),
	.w2(32'hbbd94517),
	.w3(32'hba6ab05e),
	.w4(32'hbba3ba6b),
	.w5(32'h3b5d249e),
	.w6(32'hbc7be58c),
	.w7(32'hbc36040b),
	.w8(32'h3bfd2ba1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b16aa),
	.w1(32'h3b44b24c),
	.w2(32'hbb6e8295),
	.w3(32'hbc3d644c),
	.w4(32'hbc4a4321),
	.w5(32'h3b83cdbc),
	.w6(32'hbb866c20),
	.w7(32'hbccd26ad),
	.w8(32'h3956ff25),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d003),
	.w1(32'h3c40ff34),
	.w2(32'h3c37be26),
	.w3(32'hba526983),
	.w4(32'hbb1c8b9e),
	.w5(32'hbba53e18),
	.w6(32'h3c48d405),
	.w7(32'hbcc3a06c),
	.w8(32'hbc18e832),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c541d07),
	.w1(32'hbb4441e3),
	.w2(32'hbc69bfbc),
	.w3(32'h3bbf7917),
	.w4(32'h3ba322b2),
	.w5(32'h3c021d0b),
	.w6(32'h3b5ad633),
	.w7(32'hbbbb5ae1),
	.w8(32'hbad3860f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5652c),
	.w1(32'hbc985aeb),
	.w2(32'hbb0de8ed),
	.w3(32'hbab2c3a3),
	.w4(32'h3b8124b8),
	.w5(32'hb8398444),
	.w6(32'hb9e9e135),
	.w7(32'h3c939d06),
	.w8(32'h3ca9dfe5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e0bc9),
	.w1(32'h3cfe6f31),
	.w2(32'h3cb9aa93),
	.w3(32'h3a3ba507),
	.w4(32'hbc1b9300),
	.w5(32'hbcc260c1),
	.w6(32'h3b592c75),
	.w7(32'hbc5c105f),
	.w8(32'hbc3699fd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967426),
	.w1(32'h3c61bfa8),
	.w2(32'hbcb90339),
	.w3(32'hbc23e6f7),
	.w4(32'hb9e83f97),
	.w5(32'hbbd8a644),
	.w6(32'hbaf91635),
	.w7(32'h3c9d1dea),
	.w8(32'hbc4f1f8d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86bd21),
	.w1(32'h3bb7bb42),
	.w2(32'hbc91dd4f),
	.w3(32'h3ac9bc82),
	.w4(32'hbbd851ff),
	.w5(32'h3a912e08),
	.w6(32'h3cf58ea9),
	.w7(32'hbba9d2b0),
	.w8(32'h3c095eaf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4df7c),
	.w1(32'h3b773c84),
	.w2(32'h3c5ae88b),
	.w3(32'hbb9d4701),
	.w4(32'h3c8ade2a),
	.w5(32'hbb1e1e25),
	.w6(32'hbbaf653c),
	.w7(32'hbc630ace),
	.w8(32'hbb227c92),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3a746),
	.w1(32'h3c56e258),
	.w2(32'hbc215d02),
	.w3(32'hbbd78366),
	.w4(32'h3ab9a4e7),
	.w5(32'hbb930b5b),
	.w6(32'hbb9fe06e),
	.w7(32'hbc84cc5d),
	.w8(32'h3c027eb8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a3a4d),
	.w1(32'h3bb00485),
	.w2(32'h3c8345d8),
	.w3(32'hbbe040cd),
	.w4(32'h3c1d3542),
	.w5(32'h3bb1f4ae),
	.w6(32'h3b1d721c),
	.w7(32'hbb0580f5),
	.w8(32'hbb56e639),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc942a01),
	.w1(32'hbc28ecc7),
	.w2(32'h3b3fbc55),
	.w3(32'hbb5952c7),
	.w4(32'hbc1049cb),
	.w5(32'hbc36c262),
	.w6(32'hbb4c5f50),
	.w7(32'hbc823e36),
	.w8(32'hbbb23be6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2beba4),
	.w1(32'hbb03a85a),
	.w2(32'hbb562c77),
	.w3(32'hbacf8a27),
	.w4(32'hbaa4c908),
	.w5(32'hbc13c5e2),
	.w6(32'h3b904f86),
	.w7(32'h3c402dec),
	.w8(32'h3b1c3b34),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee23cf),
	.w1(32'h3bc7289b),
	.w2(32'hba035097),
	.w3(32'h3bc10548),
	.w4(32'hbae2478c),
	.w5(32'hbcae32d3),
	.w6(32'h3b949868),
	.w7(32'hbb05aea3),
	.w8(32'hb8055acb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892701),
	.w1(32'hbbf2ab92),
	.w2(32'hbb002a8a),
	.w3(32'h3953f55f),
	.w4(32'h3b82d621),
	.w5(32'h3bbbc450),
	.w6(32'h3b5d0440),
	.w7(32'h3c79e2dc),
	.w8(32'hbb5b4e47),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a250c),
	.w1(32'hbb5a78f2),
	.w2(32'hbc097bf6),
	.w3(32'hbc0f0cc4),
	.w4(32'h3aba47d5),
	.w5(32'h3ab09ab2),
	.w6(32'h3a91f0d2),
	.w7(32'h3b1d0873),
	.w8(32'h39fcad3f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf619cb),
	.w1(32'hbb86bbee),
	.w2(32'h3b9cb891),
	.w3(32'h3ab6a3f5),
	.w4(32'h3b5e4a19),
	.w5(32'h3b48bf5e),
	.w6(32'hbab311ad),
	.w7(32'hbc283f23),
	.w8(32'h3b5c07f0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762dfa),
	.w1(32'h3bfb320c),
	.w2(32'hbb5c367d),
	.w3(32'h3b0e5f77),
	.w4(32'hbbad827f),
	.w5(32'h3934bf97),
	.w6(32'h3b19a059),
	.w7(32'hbc820a99),
	.w8(32'hbafbb892),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baedfd0),
	.w1(32'h3bdc7fce),
	.w2(32'h3bdcf79b),
	.w3(32'hbb0bbab4),
	.w4(32'hbaca286a),
	.w5(32'h396ffb28),
	.w6(32'h3c0326b5),
	.w7(32'hbc201e76),
	.w8(32'h3afbbbcf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eb727),
	.w1(32'h39c712d1),
	.w2(32'hbc83b20d),
	.w3(32'hbb1271ec),
	.w4(32'hbbd667d9),
	.w5(32'h3d2885f1),
	.w6(32'h3a89ebee),
	.w7(32'hbc85569f),
	.w8(32'h3c01fe73),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81e9d4),
	.w1(32'h39e7e13c),
	.w2(32'hb9a9f3c5),
	.w3(32'h3bdd8a6d),
	.w4(32'hbb417800),
	.w5(32'hbbb54b81),
	.w6(32'h3bab128b),
	.w7(32'h3b3a636f),
	.w8(32'h3c29566f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7cfac),
	.w1(32'h3b85918f),
	.w2(32'hbb9be6a3),
	.w3(32'h3b143c47),
	.w4(32'hbc82efdc),
	.w5(32'hbcba95b9),
	.w6(32'h3c034e73),
	.w7(32'hbb35792f),
	.w8(32'h3930d1ff),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3ada9),
	.w1(32'hbb3319ca),
	.w2(32'h3b4f4ea0),
	.w3(32'h3b8eef66),
	.w4(32'hbb2c62fa),
	.w5(32'hbc4715c0),
	.w6(32'h3a208a4b),
	.w7(32'hbb8920de),
	.w8(32'hbbab1d75),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce190d6),
	.w1(32'hbc824405),
	.w2(32'hb9b6a8c8),
	.w3(32'hbbdc7ea8),
	.w4(32'h3b46d71d),
	.w5(32'h3a4050cb),
	.w6(32'hbc3d0f3d),
	.w7(32'hbc8b7eaf),
	.w8(32'h39f90286),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac62664),
	.w1(32'h3b26fd42),
	.w2(32'hb9e5ef3e),
	.w3(32'h3b3d55a0),
	.w4(32'hbbd430e1),
	.w5(32'h3c091262),
	.w6(32'h3bf6bb24),
	.w7(32'h3b68f01f),
	.w8(32'hba936630),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f61e),
	.w1(32'hbb8d0470),
	.w2(32'hbb253806),
	.w3(32'h3c2a9baa),
	.w4(32'hba880daa),
	.w5(32'hbb36b9c2),
	.w6(32'h3b317c12),
	.w7(32'h3b80a38f),
	.w8(32'h3c303dd3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28c5d5),
	.w1(32'h3baa5f7a),
	.w2(32'h3ac8327d),
	.w3(32'hbb019668),
	.w4(32'h3b6b64a8),
	.w5(32'h3b969f5f),
	.w6(32'hbbc3bf37),
	.w7(32'hbb9dd180),
	.w8(32'hba9a901a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3628),
	.w1(32'hbbd078f9),
	.w2(32'hba68078f),
	.w3(32'h3af62528),
	.w4(32'hbca9b9dc),
	.w5(32'h3c12d279),
	.w6(32'hbbe8b111),
	.w7(32'h3aeb3c8d),
	.w8(32'h3c0c42b0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a0b81),
	.w1(32'hbbd72296),
	.w2(32'hbc17e77e),
	.w3(32'h3b03aee4),
	.w4(32'hbbe923c8),
	.w5(32'h3ac87be9),
	.w6(32'hbb8f6ff7),
	.w7(32'hbbd08aa4),
	.w8(32'h3bdf2bbc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b926),
	.w1(32'hbbae5ccd),
	.w2(32'h3b0bce91),
	.w3(32'h3beb01e4),
	.w4(32'hbbbc8422),
	.w5(32'hbc899eee),
	.w6(32'hbb800c03),
	.w7(32'hbbf9bb74),
	.w8(32'hbb4f74df),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c717ba5),
	.w1(32'hbb8c5757),
	.w2(32'h3ae88652),
	.w3(32'h3c001ed6),
	.w4(32'hbbcc1fda),
	.w5(32'hbbbf34d0),
	.w6(32'hbb996103),
	.w7(32'h39ea0b51),
	.w8(32'hbb6f7c3f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00f3f),
	.w1(32'hbc1b6e80),
	.w2(32'h3c2539fd),
	.w3(32'h3c274592),
	.w4(32'h3bbbcc91),
	.w5(32'hbc888c88),
	.w6(32'h3c21be20),
	.w7(32'h3d01683c),
	.w8(32'h3b204552),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322e6b),
	.w1(32'h3a8b87ac),
	.w2(32'hbc25aade),
	.w3(32'hbc0334c6),
	.w4(32'hba5309f4),
	.w5(32'hbc828b46),
	.w6(32'hbc15f12a),
	.w7(32'hbb9c6afd),
	.w8(32'h3bc3c2ff),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c4261),
	.w1(32'h3b2a359b),
	.w2(32'hbb275896),
	.w3(32'hbae23f1f),
	.w4(32'hbc61552f),
	.w5(32'hbcb11493),
	.w6(32'h3c69ee96),
	.w7(32'hbab30256),
	.w8(32'hbbe40f82),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41cca6),
	.w1(32'h3c298511),
	.w2(32'hbb46812f),
	.w3(32'h3b8ab644),
	.w4(32'hbb8e1edd),
	.w5(32'hbc24c344),
	.w6(32'hb9fda5f7),
	.w7(32'hbb55aa72),
	.w8(32'hbbebfef8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a937565),
	.w1(32'hbb8fd2f2),
	.w2(32'h3c07d119),
	.w3(32'hbaf12206),
	.w4(32'hba8dabf7),
	.w5(32'hbc368790),
	.w6(32'hbc417df1),
	.w7(32'h3b3f066e),
	.w8(32'hbbe572f9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0896bb),
	.w1(32'hbc0654b0),
	.w2(32'h3b307c23),
	.w3(32'h3c6fffd8),
	.w4(32'hbc0ecbd7),
	.w5(32'hba8303c0),
	.w6(32'h3acc2c96),
	.w7(32'h3c71258d),
	.w8(32'h3bc31101),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec8487),
	.w1(32'hbb8988b6),
	.w2(32'h3c375981),
	.w3(32'h3b5052be),
	.w4(32'hbb4bd91f),
	.w5(32'hbbf0859d),
	.w6(32'hbc19c4b2),
	.w7(32'hbbf2e12c),
	.w8(32'hbb5775ab),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446fda),
	.w1(32'hba3030f9),
	.w2(32'h3c829ac9),
	.w3(32'h39dd9a47),
	.w4(32'h3a72bbe6),
	.w5(32'h3b07a98a),
	.w6(32'h3c0e02c1),
	.w7(32'h3a0fc23d),
	.w8(32'hbbefc324),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8277c),
	.w1(32'h3b970937),
	.w2(32'hbb0f1e60),
	.w3(32'hbb12cc20),
	.w4(32'hb9ffa403),
	.w5(32'hbd0aefaf),
	.w6(32'hbc72c294),
	.w7(32'hbc857d1d),
	.w8(32'hbc13c441),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaaedb),
	.w1(32'h3b62bb64),
	.w2(32'h3aca2871),
	.w3(32'hbbbe86c7),
	.w4(32'h3ba0e72f),
	.w5(32'h3b46bbbf),
	.w6(32'h3b167c41),
	.w7(32'h3bc8ab17),
	.w8(32'hbb807ae3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f4b6),
	.w1(32'hbc21c3fa),
	.w2(32'h3bdd6da2),
	.w3(32'hbc8563ad),
	.w4(32'hbb3ff352),
	.w5(32'hbbdf9961),
	.w6(32'h3b095f60),
	.w7(32'h3c67898b),
	.w8(32'h3ae6d6bd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55570b),
	.w1(32'h38bbf9f3),
	.w2(32'hbb802f7d),
	.w3(32'hbb23f9ea),
	.w4(32'hbd09b383),
	.w5(32'hbb92020c),
	.w6(32'hbd32e374),
	.w7(32'h3a4263bb),
	.w8(32'hbb6e1f30),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f18b9),
	.w1(32'hbc1e6b06),
	.w2(32'hbc4da804),
	.w3(32'hbc1124df),
	.w4(32'h398c9e9e),
	.w5(32'h3c31c028),
	.w6(32'hbafb2c3a),
	.w7(32'h3c8e5496),
	.w8(32'hbc58c4a6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139668),
	.w1(32'hb946aff1),
	.w2(32'h3c1928e4),
	.w3(32'hbd06dbc4),
	.w4(32'hbb82f3b4),
	.w5(32'h3b9901cd),
	.w6(32'h3cee3668),
	.w7(32'h3a467abd),
	.w8(32'h3c312838),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3789fb),
	.w1(32'hbc28e351),
	.w2(32'hbbbe7240),
	.w3(32'h3c49d4b2),
	.w4(32'h3aaecab7),
	.w5(32'h3bbae8dc),
	.w6(32'hbbe76f2b),
	.w7(32'hbbe3c15c),
	.w8(32'hbc34de90),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba560412),
	.w1(32'hbc804ec6),
	.w2(32'hbb7cbc82),
	.w3(32'hba6cb3cf),
	.w4(32'hba8b8b09),
	.w5(32'h3b7f86c6),
	.w6(32'hbad0f5bd),
	.w7(32'hb93d1e8a),
	.w8(32'hbb22b5dc),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b47a),
	.w1(32'hbbc04b19),
	.w2(32'hbbb0bcc5),
	.w3(32'h3c47b674),
	.w4(32'hbc1a5a5e),
	.w5(32'h3bf02a49),
	.w6(32'h3a5a130a),
	.w7(32'hbbf8b66b),
	.w8(32'hbc285245),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a0c02),
	.w1(32'hba5f063c),
	.w2(32'hbaeadadd),
	.w3(32'hbbc991bd),
	.w4(32'hbb8b6a27),
	.w5(32'hb8901e7d),
	.w6(32'hbc87a372),
	.w7(32'hba4e2c22),
	.w8(32'h396a6201),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b8728),
	.w1(32'hbb8031ef),
	.w2(32'hba947772),
	.w3(32'h3ae2281a),
	.w4(32'h3b68c2ea),
	.w5(32'hbbebb6f5),
	.w6(32'hbb61c028),
	.w7(32'hbd051561),
	.w8(32'h3c1661b2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc347a7d),
	.w1(32'hbbac17e4),
	.w2(32'h3c033c0f),
	.w3(32'hbc43a327),
	.w4(32'hbc710cf3),
	.w5(32'hbc80c996),
	.w6(32'hbb9ef17d),
	.w7(32'h3aadf3d1),
	.w8(32'hbc19b4f2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb3d24),
	.w1(32'hbc7be0fb),
	.w2(32'h3b3f1c2e),
	.w3(32'hbbb6882a),
	.w4(32'hbcd3b866),
	.w5(32'h3c3d144d),
	.w6(32'h3bc4c6e6),
	.w7(32'hbbac24a8),
	.w8(32'h3b2bb5da),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1606ad),
	.w1(32'h3b802251),
	.w2(32'h3ab24579),
	.w3(32'hbbf6fa0f),
	.w4(32'h3b73f543),
	.w5(32'h3ac91dc2),
	.w6(32'h3bca6815),
	.w7(32'hbc6d70e2),
	.w8(32'hb81bd218),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ae5e0),
	.w1(32'hbbf4fe5a),
	.w2(32'h3b8cee22),
	.w3(32'h39b96707),
	.w4(32'h3c9a21bc),
	.w5(32'hbba4b5b0),
	.w6(32'hb8b7d85f),
	.w7(32'hbc0bf99d),
	.w8(32'h3b9fadc3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc5128),
	.w1(32'hbc6c1ad6),
	.w2(32'hbb9b1432),
	.w3(32'hbcb2ea05),
	.w4(32'hbc640c5b),
	.w5(32'hbbcae458),
	.w6(32'hbbc30090),
	.w7(32'h3befe53e),
	.w8(32'h3b7769a8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ed76),
	.w1(32'hba04f2db),
	.w2(32'h3c1005ab),
	.w3(32'h3bb530e1),
	.w4(32'h38cdf4b3),
	.w5(32'hbadd01c1),
	.w6(32'hba480ca2),
	.w7(32'h3b671002),
	.w8(32'h3b1c0b70),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d4d0e),
	.w1(32'h3a5fcc74),
	.w2(32'h3b4d79ad),
	.w3(32'hbababf89),
	.w4(32'h3c3176e2),
	.w5(32'hbc50d075),
	.w6(32'hbcb6921b),
	.w7(32'h3ac17982),
	.w8(32'h3ca5c8a5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37587f),
	.w1(32'hbb91bd21),
	.w2(32'h3bcc0aef),
	.w3(32'h3cc97b67),
	.w4(32'h3c445ba6),
	.w5(32'hbbb922e1),
	.w6(32'hbbe48acb),
	.w7(32'hb90d50f1),
	.w8(32'hbb9ec78a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86651e),
	.w1(32'h3cc685bf),
	.w2(32'hbb30fb8e),
	.w3(32'h3babd9c8),
	.w4(32'hbb1bb4ee),
	.w5(32'hbb1f3e77),
	.w6(32'hbc122a8c),
	.w7(32'h3b689eb6),
	.w8(32'h3bcbd034),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64ebec),
	.w1(32'hbb005ccf),
	.w2(32'h3b23cff3),
	.w3(32'h3bec08fa),
	.w4(32'hb7f166d2),
	.w5(32'hbc4e7bf4),
	.w6(32'hbb30fc73),
	.w7(32'h3b3787e3),
	.w8(32'h3c0477b4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4df1c),
	.w1(32'h3aa10cf4),
	.w2(32'hbb397cb7),
	.w3(32'h3bc5b563),
	.w4(32'h3af91cac),
	.w5(32'h3bb4e481),
	.w6(32'h3cde5c6f),
	.w7(32'hb9b895fb),
	.w8(32'hbcf805a6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d7a86),
	.w1(32'h3b72cc58),
	.w2(32'h3c78432a),
	.w3(32'h3be25f5e),
	.w4(32'h3d394fd5),
	.w5(32'hbc785ca1),
	.w6(32'h3c365f18),
	.w7(32'hb9ee4f9b),
	.w8(32'hbc1f54e9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6621),
	.w1(32'hbd06b3de),
	.w2(32'hbc6349cb),
	.w3(32'hbb577799),
	.w4(32'h3c87efa3),
	.w5(32'h3b15264d),
	.w6(32'h3c1da8eb),
	.w7(32'h3cc05947),
	.w8(32'hbbb3d229),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be402fc),
	.w1(32'hbb24dd64),
	.w2(32'h3b8a4021),
	.w3(32'hbba007d6),
	.w4(32'h3c0dcb97),
	.w5(32'hbb94e741),
	.w6(32'h3b51462c),
	.w7(32'h3c8c09ba),
	.w8(32'hbc0ccfa0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a07f),
	.w1(32'h398024cc),
	.w2(32'hbafd1ccd),
	.w3(32'h3d2f8ed5),
	.w4(32'h3b2e589a),
	.w5(32'h3b1a4012),
	.w6(32'h3c1c51e4),
	.w7(32'h3bc6fe24),
	.w8(32'hbb95cf99),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca87301),
	.w1(32'hbc091b04),
	.w2(32'hbc7cf30e),
	.w3(32'h3ba21ddf),
	.w4(32'hba305f6c),
	.w5(32'hba894fcd),
	.w6(32'h3aad8a5f),
	.w7(32'hba291c6f),
	.w8(32'h3b1616ef),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd70d4a),
	.w1(32'hbb03a654),
	.w2(32'h39a32545),
	.w3(32'h3c97ac4e),
	.w4(32'h3bd90b69),
	.w5(32'hbc36552d),
	.w6(32'h3a2c4001),
	.w7(32'h3c814477),
	.w8(32'h39b6f9eb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97f267),
	.w1(32'h3b9ffa8a),
	.w2(32'hbc3f795e),
	.w3(32'h3afac065),
	.w4(32'h3b0979a8),
	.w5(32'h3a4cd4d8),
	.w6(32'hb97c6ae0),
	.w7(32'hbd072ea3),
	.w8(32'hbc05ddca),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7cd2e),
	.w1(32'h3c852828),
	.w2(32'h3ba4c6f1),
	.w3(32'hb90fccf2),
	.w4(32'hbc26ee29),
	.w5(32'h3a39ecc6),
	.w6(32'hbd565325),
	.w7(32'hbbb3ab8d),
	.w8(32'h3b9878f4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aab64),
	.w1(32'hb9069761),
	.w2(32'h3c623357),
	.w3(32'h3cb90277),
	.w4(32'hbbe15ca9),
	.w5(32'h3b156f52),
	.w6(32'h3a53abaf),
	.w7(32'hbc4f5e2d),
	.w8(32'hbbc041b4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06a7e9),
	.w1(32'hbbc8581d),
	.w2(32'hbd3d6e90),
	.w3(32'hbb5fa042),
	.w4(32'hbb3d8187),
	.w5(32'hba386653),
	.w6(32'hbb739eca),
	.w7(32'h3c3bbdeb),
	.w8(32'hbd44cf9f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd565),
	.w1(32'hbb037d67),
	.w2(32'hb9638cba),
	.w3(32'h3a3723da),
	.w4(32'h3baea2bf),
	.w5(32'h3c847b99),
	.w6(32'hbb3fb6fe),
	.w7(32'h3bae914e),
	.w8(32'hbba4af3d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64df15),
	.w1(32'hbb74ea0a),
	.w2(32'h3d6d32cf),
	.w3(32'hbc723991),
	.w4(32'hbaa221df),
	.w5(32'h3bb79198),
	.w6(32'hbb8b76ec),
	.w7(32'hbd10c976),
	.w8(32'hbbec616e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1832ba),
	.w1(32'hbbcc7f6d),
	.w2(32'h3bda68c8),
	.w3(32'hbb927a4e),
	.w4(32'hbb01625a),
	.w5(32'hbbc080b3),
	.w6(32'hbb826dc0),
	.w7(32'hbbb11297),
	.w8(32'h3bc8675d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5013a),
	.w1(32'h3bd46238),
	.w2(32'hbb9fe7a7),
	.w3(32'hbbae0ab1),
	.w4(32'h3c57a507),
	.w5(32'hbc7e58b4),
	.w6(32'h3ac2f8cb),
	.w7(32'h3bae5a40),
	.w8(32'hbb47dadd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8dcb),
	.w1(32'hbbb7908b),
	.w2(32'h39880144),
	.w3(32'h3ad94508),
	.w4(32'h3bdaac4b),
	.w5(32'h3b815397),
	.w6(32'hbbeabcff),
	.w7(32'hbc127da9),
	.w8(32'h3b4463d6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094c19),
	.w1(32'h3c097c35),
	.w2(32'h3b387ba0),
	.w3(32'h3bb5a6b1),
	.w4(32'h3c7731b3),
	.w5(32'h3c956d7a),
	.w6(32'h3b9d5b34),
	.w7(32'hbce0e03c),
	.w8(32'h3b3330cb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fad78),
	.w1(32'h3b4469b2),
	.w2(32'hbaad4105),
	.w3(32'hba904892),
	.w4(32'h3a72c35c),
	.w5(32'h3c4906cb),
	.w6(32'h3c375991),
	.w7(32'hbc13b3cd),
	.w8(32'hba3d0010),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3707),
	.w1(32'hbb84c1b7),
	.w2(32'hbd28ee96),
	.w3(32'hba4fd8e6),
	.w4(32'hbb65ecc2),
	.w5(32'hbb3d9966),
	.w6(32'hbc9694a9),
	.w7(32'hbc445bce),
	.w8(32'hbacc84d3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a501de8),
	.w1(32'hb8d91a2c),
	.w2(32'hbb7fb09b),
	.w3(32'h395fdd45),
	.w4(32'hbc62d649),
	.w5(32'h38d40bc3),
	.w6(32'h3ad7ad5c),
	.w7(32'hbbfaa038),
	.w8(32'hbd08e2d0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd117c7),
	.w1(32'hbb8ecafb),
	.w2(32'h3b08c661),
	.w3(32'h3c9e0bad),
	.w4(32'hb9f62154),
	.w5(32'h3b42e44b),
	.w6(32'hbc57039b),
	.w7(32'hbd1b2bca),
	.w8(32'hbbcceb01),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6948c7),
	.w1(32'h3ad616b6),
	.w2(32'hbb6e9328),
	.w3(32'hbc5ff94e),
	.w4(32'h3b5513cb),
	.w5(32'hbb43fb0f),
	.w6(32'hb8df3242),
	.w7(32'h3a1a7eac),
	.w8(32'h3d4d56d2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a1cb9),
	.w1(32'h3adf1c8c),
	.w2(32'h3b57761f),
	.w3(32'h3b3eaeff),
	.w4(32'h3afe9a11),
	.w5(32'hbbf33ef5),
	.w6(32'hbbf885be),
	.w7(32'hb92074e3),
	.w8(32'hbbdf81fd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60d7a9),
	.w1(32'h3c47bcdf),
	.w2(32'h3c911b90),
	.w3(32'hbbc99b75),
	.w4(32'h3b8156c9),
	.w5(32'h3c776c32),
	.w6(32'hb9cb12d9),
	.w7(32'h3a1d54ce),
	.w8(32'h3c66cf62),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dbe63),
	.w1(32'hbca8d11b),
	.w2(32'hbb979dba),
	.w3(32'hbc39a0ba),
	.w4(32'hbb6d824b),
	.w5(32'h3ae64b3a),
	.w6(32'h3c656f12),
	.w7(32'h3b4cf3b3),
	.w8(32'h3c400f37),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60c8b),
	.w1(32'h3bcd22dd),
	.w2(32'h3be80994),
	.w3(32'hbbd2da53),
	.w4(32'h3b735ffe),
	.w5(32'h3b84830b),
	.w6(32'hbb946a8a),
	.w7(32'h3a8bbf69),
	.w8(32'hbc5c3bea),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6809b1),
	.w1(32'h3cfcfcf2),
	.w2(32'hbc3ad6d0),
	.w3(32'hbb2ea7d7),
	.w4(32'hbb7c0bf5),
	.w5(32'h3a00c200),
	.w6(32'h3a8b9ab8),
	.w7(32'hbc51ab86),
	.w8(32'h3c80d331),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ceaae),
	.w1(32'h3d273999),
	.w2(32'h3d0062f8),
	.w3(32'h3ac60c38),
	.w4(32'hbc25bc3b),
	.w5(32'hbb2057dd),
	.w6(32'hbc384e2f),
	.w7(32'hb8077536),
	.w8(32'hbcadcbd5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe18436),
	.w1(32'hbc23d736),
	.w2(32'h3c6ff6fe),
	.w3(32'hbb82311c),
	.w4(32'h3bdd8576),
	.w5(32'hba45adf4),
	.w6(32'hbc2ea3f2),
	.w7(32'hbab96b6c),
	.w8(32'hbbd1aac8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a434c),
	.w1(32'hbc083dcb),
	.w2(32'h3bdab678),
	.w3(32'hbc10b33d),
	.w4(32'hbc3c82f4),
	.w5(32'h3c59f61a),
	.w6(32'hbc152691),
	.w7(32'hbb2a0f70),
	.w8(32'h3c4838a6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac099b9),
	.w1(32'h3c1cc185),
	.w2(32'h3c650872),
	.w3(32'hbba048f4),
	.w4(32'h3be63e9f),
	.w5(32'hbce13dbf),
	.w6(32'h3a8fce21),
	.w7(32'h3a98b653),
	.w8(32'hbc9a070d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b609),
	.w1(32'hbc58bd6c),
	.w2(32'hbbaf31f7),
	.w3(32'hbbc004d8),
	.w4(32'hbad06402),
	.w5(32'hbcc240d1),
	.w6(32'h3bd80334),
	.w7(32'h3aaf74f9),
	.w8(32'h38709b16),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ab430),
	.w1(32'hbbc86abc),
	.w2(32'hbce04a63),
	.w3(32'hbb87f5fa),
	.w4(32'h3ac05085),
	.w5(32'h3b3c93e8),
	.w6(32'hbb734218),
	.w7(32'h3aad47c5),
	.w8(32'hbc8b9a7c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4de4a8),
	.w1(32'h3a4a7803),
	.w2(32'hba558731),
	.w3(32'h3b231fd3),
	.w4(32'h3c1b706c),
	.w5(32'h3a15c7dc),
	.w6(32'h3bed6462),
	.w7(32'h3b0c92fa),
	.w8(32'hbbcd0457),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0a6be),
	.w1(32'hbc6c14bd),
	.w2(32'hbc1ba371),
	.w3(32'hbc5b8f2c),
	.w4(32'hbb514765),
	.w5(32'h3b566ac8),
	.w6(32'h3a09d116),
	.w7(32'h398bac34),
	.w8(32'hbb5e1113),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e29a),
	.w1(32'hba97b672),
	.w2(32'h3c3b2b9f),
	.w3(32'h3b325582),
	.w4(32'hbba71458),
	.w5(32'hbc0bc63e),
	.w6(32'h3c819f2a),
	.w7(32'h3b148998),
	.w8(32'hbb8bb65a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a827b2e),
	.w1(32'hbc838e54),
	.w2(32'h3a094888),
	.w3(32'hbbb9ebfe),
	.w4(32'h3b297898),
	.w5(32'h3bf464b5),
	.w6(32'hbbd83be2),
	.w7(32'hbb23539a),
	.w8(32'hbc84bb8e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39799385),
	.w1(32'h3c3eb833),
	.w2(32'h3b8689a0),
	.w3(32'hbbee53c4),
	.w4(32'hbb204391),
	.w5(32'h3b144ecf),
	.w6(32'h3a4dd13c),
	.w7(32'hbb3e4dc9),
	.w8(32'h3bc37f9e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cacd4f2),
	.w1(32'hba20ee94),
	.w2(32'hbb1c9a89),
	.w3(32'h3a926053),
	.w4(32'hbcae9d12),
	.w5(32'hbc51f0f7),
	.w6(32'hbb67d7bb),
	.w7(32'hbbf71e01),
	.w8(32'hbb3c7c6f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608362),
	.w1(32'h3bfeca0a),
	.w2(32'hbc1adfb7),
	.w3(32'hbcb3c861),
	.w4(32'h3add8fca),
	.w5(32'h394737b2),
	.w6(32'hb8ba19e7),
	.w7(32'hbb9adf95),
	.w8(32'h3c07a662),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39268751),
	.w1(32'h3c077be2),
	.w2(32'h3caf9807),
	.w3(32'h3c4d45d7),
	.w4(32'h3c304db1),
	.w5(32'hbca5909d),
	.w6(32'hbb20c7ea),
	.w7(32'h3b3cbe19),
	.w8(32'hbc76f6c2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128a0d),
	.w1(32'hbbf6040c),
	.w2(32'hbca4f7b1),
	.w3(32'h3ba77b2b),
	.w4(32'hbab88205),
	.w5(32'h39602126),
	.w6(32'h3ba5b88e),
	.w7(32'h3b5ff0d3),
	.w8(32'hbc911d3e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf945c5),
	.w1(32'h3a039dca),
	.w2(32'h3ce7eac9),
	.w3(32'h3a07ac47),
	.w4(32'h3badaed8),
	.w5(32'h3c1c9acc),
	.w6(32'hba906ee3),
	.w7(32'h3aac8357),
	.w8(32'h3bba2873),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1363ab),
	.w1(32'hbc81a228),
	.w2(32'hbc19e629),
	.w3(32'hba70669b),
	.w4(32'h3a293c28),
	.w5(32'h3c91d0fc),
	.w6(32'hbb2f8c09),
	.w7(32'h3ada5f71),
	.w8(32'h3b0d50a1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5dec0),
	.w1(32'hbc1c0abe),
	.w2(32'h3b5aab2c),
	.w3(32'hb98226e5),
	.w4(32'hbbc82e98),
	.w5(32'hbb486cab),
	.w6(32'hbbe237a5),
	.w7(32'hbb9aa168),
	.w8(32'h3abcd67f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b521dc6),
	.w1(32'h3ac85935),
	.w2(32'hb85dc199),
	.w3(32'hbc2bdd77),
	.w4(32'h3ba8d099),
	.w5(32'hbb532f59),
	.w6(32'hbc22e52f),
	.w7(32'h3aef3af8),
	.w8(32'hbc22a70e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74cf81),
	.w1(32'h3b2fd39b),
	.w2(32'h3aba993b),
	.w3(32'h3c15ba1b),
	.w4(32'h3c59cef2),
	.w5(32'hbbf843a0),
	.w6(32'hbb44cbf3),
	.w7(32'hbc881532),
	.w8(32'h3c358237),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceed968),
	.w1(32'hba73085d),
	.w2(32'h3b57d003),
	.w3(32'h3be768de),
	.w4(32'h3bb731a3),
	.w5(32'h3ba3c1ac),
	.w6(32'hbbbd71c4),
	.w7(32'hba9e5df5),
	.w8(32'h3aec22aa),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6af78),
	.w1(32'h3c4adaab),
	.w2(32'hba7984b3),
	.w3(32'hbbb02dab),
	.w4(32'hbb18656b),
	.w5(32'h3bf8e454),
	.w6(32'hbc381f9d),
	.w7(32'h3c8186cd),
	.w8(32'h3c1f083c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9b22),
	.w1(32'hbaeb71e5),
	.w2(32'hbad6d040),
	.w3(32'hba965c72),
	.w4(32'hbc79a423),
	.w5(32'hbb8ae3b9),
	.w6(32'h3a85c754),
	.w7(32'h3bec116c),
	.w8(32'h3a0c842a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f0963),
	.w1(32'hbaa5ed45),
	.w2(32'hbb19cb07),
	.w3(32'hbbc9571c),
	.w4(32'h3b381212),
	.w5(32'h3b3ece45),
	.w6(32'hbc23b62e),
	.w7(32'hbc475b58),
	.w8(32'hbc038f86),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf211f7),
	.w1(32'hbb5e792a),
	.w2(32'h3a670edb),
	.w3(32'hbbaec63d),
	.w4(32'h3ba4193c),
	.w5(32'hbc674fa1),
	.w6(32'h3b2ea45d),
	.w7(32'h3b2b93f2),
	.w8(32'hbb2a7f9e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4e621),
	.w1(32'hbbc5bb80),
	.w2(32'h3bff3778),
	.w3(32'hbc595be4),
	.w4(32'hbab9c3c6),
	.w5(32'hbbba1c98),
	.w6(32'h3c799f67),
	.w7(32'hbc38ff82),
	.w8(32'hba015516),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e42c0),
	.w1(32'h3c4c1287),
	.w2(32'h3b28f3bb),
	.w3(32'h3b907def),
	.w4(32'hb76e3269),
	.w5(32'hbaa77c9e),
	.w6(32'hbba44aa5),
	.w7(32'hbbac3c45),
	.w8(32'hbc35f678),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a93c4),
	.w1(32'hbaa1eca3),
	.w2(32'hbb72ebaa),
	.w3(32'h3a8c5458),
	.w4(32'h3b18509c),
	.w5(32'h3cc8c454),
	.w6(32'h3afa629c),
	.w7(32'h3b46a9e9),
	.w8(32'h3aceb8c9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43425a),
	.w1(32'h3cae6c62),
	.w2(32'hbc121002),
	.w3(32'hbb193226),
	.w4(32'hbc6f3d7a),
	.w5(32'h3c4050fe),
	.w6(32'h3b73513c),
	.w7(32'h3a54dda4),
	.w8(32'hbbfe6745),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f3dcc),
	.w1(32'hbca1192d),
	.w2(32'h3c58fad4),
	.w3(32'h3a5db053),
	.w4(32'hbb848735),
	.w5(32'h3c255e2c),
	.w6(32'h3b2dccec),
	.w7(32'h3be101c7),
	.w8(32'h3b6e8676),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bdd1),
	.w1(32'hbbf01bab),
	.w2(32'hba3c9ca8),
	.w3(32'hb9efffd0),
	.w4(32'h3b8444fd),
	.w5(32'hbc6724c7),
	.w6(32'hbb6ebd40),
	.w7(32'hbbef1157),
	.w8(32'hbb2499fc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae4ff1),
	.w1(32'hbb77a07d),
	.w2(32'hbc0638bf),
	.w3(32'hbc032eb8),
	.w4(32'h3a047ea7),
	.w5(32'hbc7a0c63),
	.w6(32'h3b3a0b39),
	.w7(32'h3c3df837),
	.w8(32'hbb9f2849),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2350),
	.w1(32'h3c21a58e),
	.w2(32'hb9c61efe),
	.w3(32'h3bbe4921),
	.w4(32'hbd07ba6c),
	.w5(32'h3b8bb299),
	.w6(32'h3c7a9183),
	.w7(32'h3ca4aa10),
	.w8(32'h3c0e5e6d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c3ba),
	.w1(32'hbcfb5173),
	.w2(32'h3c9b36a4),
	.w3(32'h3c071844),
	.w4(32'h3b88eb99),
	.w5(32'hbb5af02a),
	.w6(32'h3956ccb4),
	.w7(32'hba5f95d5),
	.w8(32'h3abeee96),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e36a8),
	.w1(32'hbc3664ec),
	.w2(32'hbc257413),
	.w3(32'h3c33a996),
	.w4(32'h3b95254e),
	.w5(32'h3a7b6181),
	.w6(32'h3b0c4cf5),
	.w7(32'h3a4e1f03),
	.w8(32'hbc24edda),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912400),
	.w1(32'hbc574519),
	.w2(32'h3bbdb47c),
	.w3(32'h3c7909ba),
	.w4(32'hbbff91d0),
	.w5(32'hbb17d00b),
	.w6(32'hbce9ebab),
	.w7(32'hbcaefdfa),
	.w8(32'hbb4cfb08),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4da0e4),
	.w1(32'hbbe6ebf0),
	.w2(32'hbb948a3a),
	.w3(32'hbc45fcb5),
	.w4(32'h3a83c84e),
	.w5(32'h3c3621d1),
	.w6(32'h3a70a2e6),
	.w7(32'hbb1e4d7c),
	.w8(32'hbaa0198f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd491a4),
	.w1(32'h3a8fc948),
	.w2(32'h3b941028),
	.w3(32'h3b6a470d),
	.w4(32'h3c365154),
	.w5(32'h3d22ddfa),
	.w6(32'hba66c05a),
	.w7(32'h3c226740),
	.w8(32'hbab6128e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15816c),
	.w1(32'hbbb468a1),
	.w2(32'h3bbc9353),
	.w3(32'hbbbef27b),
	.w4(32'hbaa5d650),
	.w5(32'h3bff5bf9),
	.w6(32'h3b219306),
	.w7(32'hbc29980c),
	.w8(32'hbc9d9707),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc99b5),
	.w1(32'h3be0b0c5),
	.w2(32'h3a7b83ea),
	.w3(32'h3b7e52d7),
	.w4(32'h3ca6b022),
	.w5(32'hbb24e085),
	.w6(32'h3aa023d7),
	.w7(32'h3a697a60),
	.w8(32'h3bb90cd9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac91ac),
	.w1(32'hbc148dee),
	.w2(32'h36b0a0f5),
	.w3(32'h3c15f0a8),
	.w4(32'h3bc11f59),
	.w5(32'hbb758d7c),
	.w6(32'hb997d2ec),
	.w7(32'hbbc612f6),
	.w8(32'hbad6f544),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fb7c8),
	.w1(32'hbc9bad68),
	.w2(32'hba92880f),
	.w3(32'hbc204786),
	.w4(32'h3c787f03),
	.w5(32'hbc2e37bc),
	.w6(32'hbbe93293),
	.w7(32'hbb930a8b),
	.w8(32'h3bc549e4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8df86e),
	.w1(32'h3b9078ee),
	.w2(32'hbc83c998),
	.w3(32'h3a308642),
	.w4(32'hbb71125f),
	.w5(32'hbd0c0ae1),
	.w6(32'h3bfc8174),
	.w7(32'h3c000e99),
	.w8(32'h3a81fc08),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b3bf5),
	.w1(32'h3ad4f2b8),
	.w2(32'h3b35ec5b),
	.w3(32'hbb8cc481),
	.w4(32'hbc855f24),
	.w5(32'hbab151ca),
	.w6(32'hbbe18dcf),
	.w7(32'h3b056ab0),
	.w8(32'hbabce62d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cc5d3),
	.w1(32'hbb9bad96),
	.w2(32'hbbdbf596),
	.w3(32'h3b5a451f),
	.w4(32'hbae738c6),
	.w5(32'hbc8688a2),
	.w6(32'h3c17b2b2),
	.w7(32'hbbefa822),
	.w8(32'hbb6c6bc2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27886),
	.w1(32'h3a9202a5),
	.w2(32'h3b3d26b1),
	.w3(32'hbc65616e),
	.w4(32'hbc866ae7),
	.w5(32'hbb5d2f4b),
	.w6(32'hbaba5502),
	.w7(32'h39aa11bb),
	.w8(32'hb9b47614),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d7647),
	.w1(32'h3be72077),
	.w2(32'h3c4800df),
	.w3(32'h3bf4eb15),
	.w4(32'h3b4de229),
	.w5(32'h3c995cf9),
	.w6(32'hba90a595),
	.w7(32'hbb8895de),
	.w8(32'h3bc602df),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc680e28),
	.w1(32'hbb34a7c9),
	.w2(32'h3c8259fd),
	.w3(32'h3bc6b61c),
	.w4(32'h3bb699c1),
	.w5(32'hbb6f0bcd),
	.w6(32'hbb833c33),
	.w7(32'hbbe75945),
	.w8(32'hbc04462b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9adb0),
	.w1(32'hbbf1cabb),
	.w2(32'hbb0b8ef9),
	.w3(32'h3c0d785a),
	.w4(32'hbb2da068),
	.w5(32'h3c41ac16),
	.w6(32'hbcd16f35),
	.w7(32'h3b133433),
	.w8(32'hbac515ec),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac485),
	.w1(32'h3c41e2eb),
	.w2(32'hbb237a46),
	.w3(32'h39e94ae7),
	.w4(32'h3b900b0c),
	.w5(32'h3bcafdd6),
	.w6(32'h3ae2cd58),
	.w7(32'hbcb1dda6),
	.w8(32'h3bb2232f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c6be),
	.w1(32'hbc8ca6f2),
	.w2(32'h3b946489),
	.w3(32'hbb8bdd74),
	.w4(32'hbc1cbc8e),
	.w5(32'hba4b1d67),
	.w6(32'h3b90ff75),
	.w7(32'hbb89e9f9),
	.w8(32'hbcd477a6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec81e),
	.w1(32'h3a686355),
	.w2(32'h3a56229a),
	.w3(32'h39802df7),
	.w4(32'h3a8e5868),
	.w5(32'h3b617917),
	.w6(32'hb7e9a3ed),
	.w7(32'h3aaf4ab8),
	.w8(32'hbc8b3f8a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8f7d),
	.w1(32'hbc3314aa),
	.w2(32'hbb3aacb9),
	.w3(32'hbb6d1873),
	.w4(32'hbbf02a56),
	.w5(32'hbc76f489),
	.w6(32'h3bc7f9b0),
	.w7(32'hbc0daf2d),
	.w8(32'h3beec4e0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e0ba),
	.w1(32'hba2781fd),
	.w2(32'h3c451cb6),
	.w3(32'hbc677618),
	.w4(32'hbc3a3978),
	.w5(32'hbb7429f4),
	.w6(32'hbbeba5fc),
	.w7(32'hbb6bd0db),
	.w8(32'h3bd01124),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc404980),
	.w1(32'hbba47624),
	.w2(32'hbbf31cb4),
	.w3(32'h3c80cfe9),
	.w4(32'h39fd60fd),
	.w5(32'h3ba1da0c),
	.w6(32'h3bc99e1f),
	.w7(32'hbb8d65ab),
	.w8(32'h3c13e346),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8794b2),
	.w1(32'h3bcae754),
	.w2(32'h3ac586c7),
	.w3(32'h3ad1c7c9),
	.w4(32'hbc19f900),
	.w5(32'hbc41d0d4),
	.w6(32'hbb578fce),
	.w7(32'h3b774d8d),
	.w8(32'hbb956d7c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46e894),
	.w1(32'h3b78d654),
	.w2(32'h3b398cce),
	.w3(32'h3bee9ea8),
	.w4(32'h3c1e5933),
	.w5(32'h3c49386d),
	.w6(32'h3a1e02af),
	.w7(32'h3bafa14c),
	.w8(32'h389bc875),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c683),
	.w1(32'h3bb2b91a),
	.w2(32'hbc45e5d4),
	.w3(32'hbbc48ad9),
	.w4(32'hbc6513ea),
	.w5(32'hbc03247b),
	.w6(32'hbbb2985a),
	.w7(32'hba95e586),
	.w8(32'hbae4d5cb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0220f5),
	.w1(32'h3c9a6566),
	.w2(32'hbb0144cc),
	.w3(32'h3a729b14),
	.w4(32'h3b39adf9),
	.w5(32'h3b8a681c),
	.w6(32'h3a971165),
	.w7(32'h3b985da6),
	.w8(32'h3c833548),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b167036),
	.w1(32'hbbc11c13),
	.w2(32'hbb7c3589),
	.w3(32'hbc804217),
	.w4(32'hbb8edbb0),
	.w5(32'hbc44a0bb),
	.w6(32'h3a8b2e9f),
	.w7(32'h3b217a11),
	.w8(32'hbc15e803),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1d1f0),
	.w1(32'h3b0caeb5),
	.w2(32'h389345e5),
	.w3(32'hb9f36874),
	.w4(32'hbc34aef6),
	.w5(32'h3c683d2b),
	.w6(32'h38b42582),
	.w7(32'hbc17423b),
	.w8(32'hb9bddf83),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b52d8),
	.w1(32'hbc44d6b8),
	.w2(32'hbafbc3ec),
	.w3(32'h38da80d6),
	.w4(32'hbb822e1e),
	.w5(32'hbc6c5f96),
	.w6(32'hbb6d32f0),
	.w7(32'h3b2d8536),
	.w8(32'hbc83a1b7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb5046),
	.w1(32'h3b4d69c7),
	.w2(32'h3a27f5a5),
	.w3(32'h3a2ef701),
	.w4(32'h3d2ad9c0),
	.w5(32'hbc1d1d58),
	.w6(32'hbb46ad84),
	.w7(32'hbb38cad9),
	.w8(32'hbc37ec60),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a382f),
	.w1(32'h3ae31f0d),
	.w2(32'hb9e07287),
	.w3(32'h3bd3959a),
	.w4(32'h3bd25e72),
	.w5(32'hbbc146ae),
	.w6(32'h3ace855c),
	.w7(32'hba98cc06),
	.w8(32'h3c16fbbe),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd53c4a9),
	.w1(32'hbc1e7243),
	.w2(32'hbbee5790),
	.w3(32'hbc166bb4),
	.w4(32'hb9d7a7d5),
	.w5(32'hbc35eeef),
	.w6(32'hbae7e57c),
	.w7(32'hbc0151a0),
	.w8(32'hbbb9cde5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec949f),
	.w1(32'hbbd09058),
	.w2(32'h3b3cef78),
	.w3(32'h395b2f54),
	.w4(32'h3bd43869),
	.w5(32'hba38131e),
	.w6(32'h3b9c72d0),
	.w7(32'hbbe4e07a),
	.w8(32'hbc258dd5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55288a),
	.w1(32'hba7a178a),
	.w2(32'hba2e9ea9),
	.w3(32'h3ac1ec3a),
	.w4(32'h3b81c4f4),
	.w5(32'h3c8fc1d2),
	.w6(32'h3b9a7568),
	.w7(32'h3cee2e79),
	.w8(32'hbc1cd68d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94a29f),
	.w1(32'hbbaddb21),
	.w2(32'hbc183268),
	.w3(32'hbbe05e0f),
	.w4(32'hbbf3ef46),
	.w5(32'hba83da5a),
	.w6(32'hbc06b51f),
	.w7(32'h3a893e94),
	.w8(32'hbbbfe882),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84a735),
	.w1(32'hbb6a279f),
	.w2(32'h3b881e8f),
	.w3(32'hbbb90f2d),
	.w4(32'h3c680351),
	.w5(32'hba90322c),
	.w6(32'hbb57b084),
	.w7(32'hbbeb1086),
	.w8(32'hbb85c9e6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8507dd),
	.w1(32'h3acaa617),
	.w2(32'hba96e8b4),
	.w3(32'hba1eae62),
	.w4(32'h3bb2577e),
	.w5(32'h3b8a511e),
	.w6(32'h3d13c435),
	.w7(32'hbaa8462c),
	.w8(32'h3bec2130),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca696),
	.w1(32'h3b16a200),
	.w2(32'hbbd56f0b),
	.w3(32'hbb105a88),
	.w4(32'hbd108e56),
	.w5(32'hbc3fd083),
	.w6(32'hbbcfa632),
	.w7(32'h3be588d1),
	.w8(32'h3c3eed4a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7e9b2f),
	.w1(32'hbd4631de),
	.w2(32'h3b0c2732),
	.w3(32'hba780943),
	.w4(32'hbc39fc62),
	.w5(32'hb98d33f9),
	.w6(32'hbc240407),
	.w7(32'h3c36e779),
	.w8(32'h3c0498f2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6325f6),
	.w1(32'h3bd74d61),
	.w2(32'hbab19330),
	.w3(32'hbb7f04fc),
	.w4(32'h3ae14f94),
	.w5(32'hbac7fd3d),
	.w6(32'hbb508976),
	.w7(32'h3bc6b2c1),
	.w8(32'h3b432483),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a23e),
	.w1(32'h3b22365f),
	.w2(32'hbb8f2b2f),
	.w3(32'h3b045ac2),
	.w4(32'h3c7d3753),
	.w5(32'h3a6a1960),
	.w6(32'h3c06dee7),
	.w7(32'h3af79bd0),
	.w8(32'h3b5870a7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39765b83),
	.w1(32'hbcb5e2ed),
	.w2(32'h3b52c0c2),
	.w3(32'hba7f7056),
	.w4(32'h3b9e54cf),
	.w5(32'h3b5b067a),
	.w6(32'hba5de01f),
	.w7(32'h3b82fff2),
	.w8(32'hbd14f2af),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f744d),
	.w1(32'hbb929794),
	.w2(32'hbbd3723e),
	.w3(32'h3cbd4b93),
	.w4(32'hbae86a16),
	.w5(32'hbb6755bd),
	.w6(32'hbc482ecd),
	.w7(32'hbab2ecb2),
	.w8(32'h3c8e7016),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fd178),
	.w1(32'h3c1dc417),
	.w2(32'h3a3c656a),
	.w3(32'hbbb4a92b),
	.w4(32'h3b1b4b3c),
	.w5(32'h3afbe5c4),
	.w6(32'h3b860d8b),
	.w7(32'h3cff1f16),
	.w8(32'hbaab2a53),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72a6a1),
	.w1(32'hbba97771),
	.w2(32'hb99b4c2b),
	.w3(32'hbc1dbf4f),
	.w4(32'hbc01edef),
	.w5(32'h3a8507a4),
	.w6(32'h3c1be220),
	.w7(32'h3ac752c2),
	.w8(32'hba356dc6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1059d),
	.w1(32'h39256236),
	.w2(32'hbb650ed3),
	.w3(32'h3bf471da),
	.w4(32'hbbd54529),
	.w5(32'hbcaf1388),
	.w6(32'hbd326bea),
	.w7(32'hbbfd8b9e),
	.w8(32'h3c5e542a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40d288),
	.w1(32'hbb4b025e),
	.w2(32'hbb355884),
	.w3(32'h3b814110),
	.w4(32'h3bfd3927),
	.w5(32'h3a5130cd),
	.w6(32'hbaabbd7d),
	.w7(32'hbbe46541),
	.w8(32'h38cf4e74),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22a7a4),
	.w1(32'hbcd19d68),
	.w2(32'h3ba3ff6b),
	.w3(32'hba42d9dd),
	.w4(32'hbd0a3906),
	.w5(32'hbc8321e0),
	.w6(32'h3d0095e6),
	.w7(32'h3c97ebef),
	.w8(32'h3bb3974a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12a293),
	.w1(32'hbb9ce918),
	.w2(32'h3b1c6e04),
	.w3(32'h3cc06f06),
	.w4(32'h3b03242d),
	.w5(32'h3a1bc35d),
	.w6(32'hbc0b2574),
	.w7(32'hbaceb871),
	.w8(32'hbcdd87ae),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14e981),
	.w1(32'hba900385),
	.w2(32'hbc0d033f),
	.w3(32'hb922119f),
	.w4(32'hbca0d692),
	.w5(32'hbbcaacec),
	.w6(32'hbc215e26),
	.w7(32'h3c2743ff),
	.w8(32'hbc5fbf29),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87e20d),
	.w1(32'hbb1018b9),
	.w2(32'hbb69504e),
	.w3(32'h3c212f17),
	.w4(32'hba2ec40d),
	.w5(32'hbb6e25e5),
	.w6(32'h3c7450d3),
	.w7(32'hbc5b741d),
	.w8(32'hbd6ef56c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2bf0),
	.w1(32'hbc9506b3),
	.w2(32'hbc7863fb),
	.w3(32'hbb5740ba),
	.w4(32'hbb8ab7c0),
	.w5(32'h3b1be17d),
	.w6(32'h3ab6f656),
	.w7(32'hba48ad5e),
	.w8(32'hbb8e5211),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cc9ab),
	.w1(32'hbca98046),
	.w2(32'hbbd708fc),
	.w3(32'h3d0ce9de),
	.w4(32'hbb9f5d2a),
	.w5(32'hbc025e81),
	.w6(32'hbc5d1515),
	.w7(32'hbb062c7f),
	.w8(32'hba5c29a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule