module layer_8_featuremap_93(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b2aa),
	.w1(32'h3dfc41f1),
	.w2(32'h3d2e57cf),
	.w3(32'h3d563d94),
	.w4(32'h3d89786b),
	.w5(32'h3dd44e3a),
	.w6(32'h3d92f14c),
	.w7(32'hbbdd8b4d),
	.w8(32'h3d9c3422),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9d204c),
	.w1(32'h3d9feda5),
	.w2(32'h3c26c180),
	.w3(32'h3cf7fed4),
	.w4(32'h3d83c719),
	.w5(32'h3cff4bd1),
	.w6(32'h3d2a9d5f),
	.w7(32'hbb450dd5),
	.w8(32'h3cb85ac5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d287b30),
	.w1(32'h3d4d5647),
	.w2(32'h3d71a2fa),
	.w3(32'h3cc60df9),
	.w4(32'h3d15904f),
	.w5(32'h3c45b332),
	.w6(32'h3da6e9be),
	.w7(32'h3b35b3cd),
	.w8(32'h3d34afb4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1190a1),
	.w1(32'h3d70a0c1),
	.w2(32'h3dc5d18e),
	.w3(32'h3ca019f5),
	.w4(32'h3c2caa8e),
	.w5(32'h3e19d6e1),
	.w6(32'h3dadebeb),
	.w7(32'h3cd9a16c),
	.w8(32'h3d7e431c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed7c36),
	.w1(32'h3d7dc3bf),
	.w2(32'h3d981903),
	.w3(32'h3c97862e),
	.w4(32'h3db6ee4d),
	.w5(32'h3c5f3a82),
	.w6(32'hbbac94bc),
	.w7(32'h3d9d6b90),
	.w8(32'hbb5dd528),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da93595),
	.w1(32'h3c124d83),
	.w2(32'hbba516db),
	.w3(32'h3d120cf4),
	.w4(32'h39b0259c),
	.w5(32'h3d503d66),
	.w6(32'h3c164e35),
	.w7(32'hbb554dc2),
	.w8(32'h3cb793a4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dcc3889),
	.w1(32'h3dd744aa),
	.w2(32'h3d102429),
	.w3(32'h3deef8d1),
	.w4(32'h3dd60d84),
	.w5(32'h3dbdfde3),
	.w6(32'hb8f45631),
	.w7(32'h3c91b5b2),
	.w8(32'h3c6deeda),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c628715),
	.w1(32'h3d900e48),
	.w2(32'h3d7605c2),
	.w3(32'h3cedd291),
	.w4(32'h3dbcf295),
	.w5(32'h3de09dcb),
	.w6(32'h3d6772e5),
	.w7(32'h3d8f2382),
	.w8(32'h3d5bf4de),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d104b0e),
	.w1(32'h3e0013fd),
	.w2(32'h3b8ab8fb),
	.w3(32'h3c15c85d),
	.w4(32'h3da4d6e7),
	.w5(32'h3bb0fa7e),
	.w6(32'h3caa1f6c),
	.w7(32'h3b975cd9),
	.w8(32'h3d993756),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee7348),
	.w1(32'h3dc54601),
	.w2(32'h3d2ab738),
	.w3(32'h3e0e9615),
	.w4(32'h3d8f3bec),
	.w5(32'h3db21a78),
	.w6(32'h3de4759a),
	.w7(32'h3d62e800),
	.w8(32'h3d99cf52),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8e9e51),
	.w1(32'h3d066b1b),
	.w2(32'h3d4f8f3e),
	.w3(32'h39065232),
	.w4(32'h3adf8268),
	.w5(32'h3bf8632c),
	.w6(32'h3cad79da),
	.w7(32'hbb1b65cd),
	.w8(32'h3d131314),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8178c6),
	.w1(32'h3d9eb3df),
	.w2(32'h3ca27de6),
	.w3(32'h3c90f8ce),
	.w4(32'h3ccb8dc3),
	.w5(32'h3db405f1),
	.w6(32'hba94b0b4),
	.w7(32'h3d9f6bcb),
	.w8(32'h3c093b3b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930db6),
	.w1(32'h3da8688b),
	.w2(32'h3b83ab1c),
	.w3(32'h3d0098de),
	.w4(32'h3bc5980c),
	.w5(32'h3b921428),
	.w6(32'h3d9947f3),
	.w7(32'h3bb7c388),
	.w8(32'h3b61ee8b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf91e),
	.w1(32'hbaa79786),
	.w2(32'hba963441),
	.w3(32'hba1e0612),
	.w4(32'hba538f7d),
	.w5(32'hba55648a),
	.w6(32'hba4ec250),
	.w7(32'hba7a3931),
	.w8(32'hba8e343f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aea5d7),
	.w1(32'h381b1cfa),
	.w2(32'h3883f36e),
	.w3(32'hb80769c6),
	.w4(32'h37c0f192),
	.w5(32'h38422724),
	.w6(32'hb7ca6ebb),
	.w7(32'h37137be9),
	.w8(32'h381cbed8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08351d),
	.w1(32'h39e75901),
	.w2(32'h39e54497),
	.w3(32'h39d38ec2),
	.w4(32'h39cdc36f),
	.w5(32'h39c00b15),
	.w6(32'h3962a70e),
	.w7(32'h39b49405),
	.w8(32'h39ecda24),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae770fc),
	.w1(32'hbb077145),
	.w2(32'h39672e64),
	.w3(32'hb9abb567),
	.w4(32'hb9acb739),
	.w5(32'h3ad8c56f),
	.w6(32'h39c59533),
	.w7(32'hba57945b),
	.w8(32'h3b2d54d0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2dc07),
	.w1(32'h3c20a64d),
	.w2(32'h3bfb4dd5),
	.w3(32'h3b988ad5),
	.w4(32'h3be7790c),
	.w5(32'h3c195a4d),
	.w6(32'h3b0d151d),
	.w7(32'hba79bebe),
	.w8(32'hbaeaf962),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c721353),
	.w1(32'h3cce50aa),
	.w2(32'h3cea8b23),
	.w3(32'h3bcfbd79),
	.w4(32'h3ca72589),
	.w5(32'h3d2f1282),
	.w6(32'hbc9c59c9),
	.w7(32'hbc2cda83),
	.w8(32'h3cb86d7f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c0b24),
	.w1(32'h3af15753),
	.w2(32'h3bd7280c),
	.w3(32'hbc318a90),
	.w4(32'hbc2289a2),
	.w5(32'hbbb9165f),
	.w6(32'hbc1778f3),
	.w7(32'hbbb7fdb4),
	.w8(32'hba7b4d0f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a6d3),
	.w1(32'hbbb51e61),
	.w2(32'hbbc38ea2),
	.w3(32'hbb5ccbea),
	.w4(32'hbc41f783),
	.w5(32'hbbde648f),
	.w6(32'hb720cd18),
	.w7(32'hbc1b6140),
	.w8(32'hbb566d9b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6620e9),
	.w1(32'hbc889be2),
	.w2(32'hbc32b4cc),
	.w3(32'hbc45a966),
	.w4(32'hbc50423f),
	.w5(32'hbbfc2886),
	.w6(32'hbc576bac),
	.w7(32'hbc59b057),
	.w8(32'hbc032337),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a0ac0),
	.w1(32'h3b32c691),
	.w2(32'h3c839b87),
	.w3(32'hbc8db525),
	.w4(32'hbbc1d182),
	.w5(32'h3c890170),
	.w6(32'hbcafc780),
	.w7(32'hbc82cb8e),
	.w8(32'h3c5ba3da),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e8e86),
	.w1(32'h3b80055c),
	.w2(32'hb952f885),
	.w3(32'h3ad0038d),
	.w4(32'h3aa15d99),
	.w5(32'hbb46b36e),
	.w6(32'h3ae908e0),
	.w7(32'hba0139f1),
	.w8(32'hbb398000),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12daf8),
	.w1(32'h3ac8d6b7),
	.w2(32'h3aa64454),
	.w3(32'h3ae7f1d2),
	.w4(32'h3b01374d),
	.w5(32'h3ad56459),
	.w6(32'h3b0bc370),
	.w7(32'h3b1abd85),
	.w8(32'h3b143d00),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6aeb),
	.w1(32'h3b60e7d9),
	.w2(32'h3c5370e9),
	.w3(32'hbb7610ef),
	.w4(32'h3b25b0f0),
	.w5(32'h3c60f558),
	.w6(32'hbbfd91fa),
	.w7(32'hbc073905),
	.w8(32'h3b5604f3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9003967),
	.w1(32'h3a276dd2),
	.w2(32'h39fce993),
	.w3(32'hb9475345),
	.w4(32'h39a4ed3d),
	.w5(32'h397c9774),
	.w6(32'hb9d8dfd8),
	.w7(32'h390c6c7e),
	.w8(32'h39441895),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde0d40),
	.w1(32'hbc7e942a),
	.w2(32'hbb44c0e5),
	.w3(32'hbc680782),
	.w4(32'hbc7a8071),
	.w5(32'h3b160e33),
	.w6(32'hbc6fe10a),
	.w7(32'hbd567bed),
	.w8(32'hbbca30ec),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2712d),
	.w1(32'h3bdc307e),
	.w2(32'h3c4680b1),
	.w3(32'h3b42dfc1),
	.w4(32'h3baac713),
	.w5(32'h3c453e7c),
	.w6(32'hbaa24bc5),
	.w7(32'hba8ce4a5),
	.w8(32'h3ba1d1f6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a301973),
	.w1(32'h3839f644),
	.w2(32'hba5290f7),
	.w3(32'h3b08df99),
	.w4(32'h3ac71b7e),
	.w5(32'h3a253933),
	.w6(32'h3ace913a),
	.w7(32'h3a85569d),
	.w8(32'h39c2603b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39a89),
	.w1(32'h3a61ece4),
	.w2(32'h3ae9b9f2),
	.w3(32'hb825a7dc),
	.w4(32'h3acd0cb0),
	.w5(32'h3b2d203f),
	.w6(32'h3a8102d0),
	.w7(32'h3b27e824),
	.w8(32'h3b3f8172),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcaab3),
	.w1(32'hba399c77),
	.w2(32'hba9a1527),
	.w3(32'h3890f474),
	.w4(32'hb98b7261),
	.w5(32'hba90c973),
	.w6(32'hbb4ec5aa),
	.w7(32'hbb4df04b),
	.w8(32'hbb1c9bb8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb18ce),
	.w1(32'h39640734),
	.w2(32'h3956a947),
	.w3(32'h37176a07),
	.w4(32'h38fe8b2e),
	.w5(32'h395007f7),
	.w6(32'h381b9582),
	.w7(32'h39116cd1),
	.w8(32'h3980a440),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afdd37),
	.w1(32'h39046af7),
	.w2(32'h38bdb81b),
	.w3(32'hb6bd9050),
	.w4(32'h3853d750),
	.w5(32'h38322106),
	.w6(32'hb7cb1d21),
	.w7(32'h38a8613e),
	.w8(32'h382f7aad),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305548),
	.w1(32'hbc3bf96e),
	.w2(32'hbc52523c),
	.w3(32'hbc58498a),
	.w4(32'hbc63b9b1),
	.w5(32'hbc794480),
	.w6(32'hbbf29534),
	.w7(32'hbbb5b396),
	.w8(32'hbc059786),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716c12c),
	.w1(32'h3b6b74c5),
	.w2(32'h3bfab828),
	.w3(32'h3b469993),
	.w4(32'h3b5a4b96),
	.w5(32'h3c225092),
	.w6(32'hbb03c2b6),
	.w7(32'hbbd5df02),
	.w8(32'h3b6e5ca4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e9c19),
	.w1(32'h36065fdf),
	.w2(32'h37eb8bfe),
	.w3(32'hb88d8cf8),
	.w4(32'h36c6db47),
	.w5(32'hb7da50f2),
	.w6(32'hb8a1de44),
	.w7(32'h37a797ea),
	.w8(32'hb86c52b5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2751f),
	.w1(32'hb6ca5dde),
	.w2(32'h3a86f999),
	.w3(32'hbb1071aa),
	.w4(32'hbae5af37),
	.w5(32'hba1d0263),
	.w6(32'hbbc59737),
	.w7(32'hbbeacd24),
	.w8(32'hbb96b17f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869311),
	.w1(32'hbadb3dd6),
	.w2(32'hbac59ddd),
	.w3(32'hba9d0ad6),
	.w4(32'hbae58848),
	.w5(32'hbaa4e290),
	.w6(32'hba8b0fab),
	.w7(32'hbac1bccb),
	.w8(32'hba82ba54),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba640ff3),
	.w1(32'hb9e939fd),
	.w2(32'hba216e4e),
	.w3(32'hbb03989b),
	.w4(32'hba8fa81f),
	.w5(32'hba71b4ea),
	.w6(32'hbac8b25f),
	.w7(32'hba4e619a),
	.w8(32'hba6490cc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c163778),
	.w1(32'h3d02f74b),
	.w2(32'h3d284887),
	.w3(32'h3c6b9c54),
	.w4(32'h3cbff452),
	.w5(32'h3d0bb4e1),
	.w6(32'hbae10022),
	.w7(32'h3c0228d2),
	.w8(32'h3cc491b1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e6cc4),
	.w1(32'h3ab345bb),
	.w2(32'h3a2fa5ab),
	.w3(32'h3a6ec106),
	.w4(32'h3b04ea41),
	.w5(32'h3b70f4e4),
	.w6(32'hba4a4497),
	.w7(32'hba9b2252),
	.w8(32'h3b208975),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfa68d),
	.w1(32'hbad23b11),
	.w2(32'hbb034dc9),
	.w3(32'hb8e05781),
	.w4(32'hba7d5fc6),
	.w5(32'hbaea51b7),
	.w6(32'hb944989d),
	.w7(32'hba87f352),
	.w8(32'hbaef0b0d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1317d2),
	.w1(32'h3b5f0495),
	.w2(32'h3b7eb31e),
	.w3(32'h3b80fdf4),
	.w4(32'h3b3f8599),
	.w5(32'h3baa57ba),
	.w6(32'hb9b30c54),
	.w7(32'hbae73fd2),
	.w8(32'h3b65406d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51db64),
	.w1(32'h3c958abe),
	.w2(32'h3c9e7bef),
	.w3(32'h3c456192),
	.w4(32'h3c502568),
	.w5(32'h3ca167f2),
	.w6(32'h3b0e9b72),
	.w7(32'h3b17a534),
	.w8(32'h3c8335fc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39325a81),
	.w1(32'h3b86e114),
	.w2(32'h3b9a32fc),
	.w3(32'h3aceaa9f),
	.w4(32'h3b400363),
	.w5(32'h3bc8b1dd),
	.w6(32'hbbb7a9f6),
	.w7(32'hbb4748ac),
	.w8(32'h3b19309e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37774e25),
	.w1(32'h37ce28c7),
	.w2(32'h377e9259),
	.w3(32'hb74c804a),
	.w4(32'h37925530),
	.w5(32'h3637ee70),
	.w6(32'hb8630df4),
	.w7(32'h35e10b30),
	.w8(32'h36ed5f48),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dca4f),
	.w1(32'hbb81763c),
	.w2(32'h3b8e56e2),
	.w3(32'hbc24f630),
	.w4(32'hbb95d9e8),
	.w5(32'h3c129435),
	.w6(32'hbc93028d),
	.w7(32'hbc5e5137),
	.w8(32'h3b8e06c5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b057532),
	.w1(32'h3b57d67b),
	.w2(32'h3b1f59bc),
	.w3(32'h3b952a4c),
	.w4(32'h3b70ffea),
	.w5(32'h3b653584),
	.w6(32'h3b3ba03d),
	.w7(32'h3aa5c701),
	.w8(32'h3b240e0a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a151af1),
	.w1(32'h3c192d80),
	.w2(32'h3c8de6aa),
	.w3(32'h3bcbd178),
	.w4(32'h3c0ec264),
	.w5(32'h3c7bbe3e),
	.w6(32'h3b017f88),
	.w7(32'h3b5b12f4),
	.w8(32'h3c5ba305),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ae5ba),
	.w1(32'hba9989ca),
	.w2(32'h3b971d65),
	.w3(32'hbb6e2336),
	.w4(32'hbb514b46),
	.w5(32'hbb63f1ad),
	.w6(32'hbbf0dce6),
	.w7(32'hbc40b219),
	.w8(32'hbc6e26d9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8e4a),
	.w1(32'h3c0ca321),
	.w2(32'h3c9acc05),
	.w3(32'hbbad9f11),
	.w4(32'h3c977752),
	.w5(32'h3cfce4f5),
	.w6(32'hbc8ac763),
	.w7(32'hbab17b95),
	.w8(32'h3c8e7964),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996a810),
	.w1(32'h3b265e94),
	.w2(32'h3ba24068),
	.w3(32'h3b199702),
	.w4(32'h3b8d6025),
	.w5(32'h3bca214b),
	.w6(32'hbb245c74),
	.w7(32'hbac30a3b),
	.w8(32'h3b30d7d6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5e137),
	.w1(32'h3c782689),
	.w2(32'h3cb51871),
	.w3(32'h3be17c84),
	.w4(32'h3badc177),
	.w5(32'h3c7cebd8),
	.w6(32'h3bc2f5e1),
	.w7(32'h3bbb1afa),
	.w8(32'h3c209525),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382b51fa),
	.w1(32'h39165adc),
	.w2(32'h3951a672),
	.w3(32'hb85d4ec7),
	.w4(32'h387c2e5c),
	.w5(32'h39069bac),
	.w6(32'hb8d9e7b0),
	.w7(32'hb7056c0c),
	.w8(32'h38cf4137),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1193),
	.w1(32'h3c7b012d),
	.w2(32'h3cf10940),
	.w3(32'hbb7bd412),
	.w4(32'h3b8f0fe2),
	.w5(32'h3cd68f02),
	.w6(32'hbbdaa1bc),
	.w7(32'hbbc59102),
	.w8(32'h3c11314e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28f350),
	.w1(32'h39a979f2),
	.w2(32'h39c03014),
	.w3(32'hbb38ebd1),
	.w4(32'hbb524ba8),
	.w5(32'hbaa034a1),
	.w6(32'hbb15bfcd),
	.w7(32'h39b0ed62),
	.w8(32'h3ad9603b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fbc6c),
	.w1(32'hbad6058f),
	.w2(32'hb87e0ae6),
	.w3(32'h3b58119d),
	.w4(32'h3bf48ae5),
	.w5(32'h3c1a4c43),
	.w6(32'hba8253e9),
	.w7(32'hbb4e23a6),
	.w8(32'h3b53da29),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0301d),
	.w1(32'hbb6852f6),
	.w2(32'hb9ed4c08),
	.w3(32'hbba18199),
	.w4(32'hbbbb4950),
	.w5(32'hba397d36),
	.w6(32'hbb800751),
	.w7(32'hbbecbf61),
	.w8(32'h3a35afb6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb439c2),
	.w1(32'h3c108613),
	.w2(32'h3c297193),
	.w3(32'h3ae8310c),
	.w4(32'h3b9d49cd),
	.w5(32'h3bc89628),
	.w6(32'h3b49bfd8),
	.w7(32'h3b9a899e),
	.w8(32'h3c180a5b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31e797),
	.w1(32'h3a1d154e),
	.w2(32'h39eb2de3),
	.w3(32'h3a26b55f),
	.w4(32'h3a1bdbd1),
	.w5(32'h3a1e5058),
	.w6(32'h3a3290ca),
	.w7(32'h3a6e5a06),
	.w8(32'h3a5850e0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ca4b5),
	.w1(32'hba619c81),
	.w2(32'h388a7618),
	.w3(32'hbac4239c),
	.w4(32'hba2ad02b),
	.w5(32'h38bb917a),
	.w6(32'hba9a5cca),
	.w7(32'hba358e0d),
	.w8(32'hb99e51d6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d022e),
	.w1(32'h3cd7b303),
	.w2(32'h3cf2f906),
	.w3(32'h3c72f141),
	.w4(32'h3cbce26b),
	.w5(32'h3d07696c),
	.w6(32'hba4a2614),
	.w7(32'h3bad5b31),
	.w8(32'h3c59f9d4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4921cc),
	.w1(32'hba4e3ef9),
	.w2(32'hbad232a3),
	.w3(32'h3b8258c1),
	.w4(32'h3bc7d666),
	.w5(32'h3b92c9f8),
	.w6(32'h3b79b7b7),
	.w7(32'h3b8af005),
	.w8(32'h3b424c24),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a193c8a),
	.w1(32'hba8ac348),
	.w2(32'hbac2e029),
	.w3(32'h3b1cbfcd),
	.w4(32'hb930cd70),
	.w5(32'hba204606),
	.w6(32'h3b261fb3),
	.w7(32'h3928d896),
	.w8(32'hbacdd1f9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e78c2b),
	.w1(32'h3b4e8997),
	.w2(32'h3b25ecf3),
	.w3(32'h3b63180f),
	.w4(32'h3b9489ce),
	.w5(32'h3ba465aa),
	.w6(32'h3ad2d393),
	.w7(32'h3a3961fb),
	.w8(32'h3b835c5f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b9bbc),
	.w1(32'h3b878954),
	.w2(32'h3bbc050e),
	.w3(32'h3bb377c2),
	.w4(32'h3b900947),
	.w5(32'h3bb1bc10),
	.w6(32'h3b9ba990),
	.w7(32'h3b22a5a0),
	.w8(32'h3b84b4c3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98145c),
	.w1(32'h397116b4),
	.w2(32'h3b81b617),
	.w3(32'h39fa79d3),
	.w4(32'h3a7f758a),
	.w5(32'h3ba9432a),
	.w6(32'hbb905446),
	.w7(32'hbbb7cc89),
	.w8(32'hbb0ab015),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922e404),
	.w1(32'hb9b3af2e),
	.w2(32'hb99e66c7),
	.w3(32'hb96b2479),
	.w4(32'hb98e7a29),
	.w5(32'hb950bab0),
	.w6(32'hb9a5bbb1),
	.w7(32'hb982212a),
	.w8(32'hb989c6e4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb60e),
	.w1(32'hbc3df821),
	.w2(32'hbbb9e3e1),
	.w3(32'h3bead536),
	.w4(32'hbb1580a9),
	.w5(32'h3bcdf275),
	.w6(32'h3c248b01),
	.w7(32'hbc507eb4),
	.w8(32'h3c47aaf8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984563e),
	.w1(32'hb90b33f2),
	.w2(32'hb9c491bc),
	.w3(32'hb787884d),
	.w4(32'h38ed34ba),
	.w5(32'hb92213bb),
	.w6(32'h3908b0f0),
	.w7(32'h396592a5),
	.w8(32'hb8d127ba),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06894),
	.w1(32'h3ae57f86),
	.w2(32'h3aa9047f),
	.w3(32'hba3fbc5a),
	.w4(32'hb96eb672),
	.w5(32'h3aed2d45),
	.w6(32'hbb5d35e0),
	.w7(32'hbaea8860),
	.w8(32'h3b625fb6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d384b0),
	.w1(32'h39882b1e),
	.w2(32'hb7ca4b4d),
	.w3(32'h38e10c61),
	.w4(32'h3a1e076e),
	.w5(32'h396998c2),
	.w6(32'h394b32e3),
	.w7(32'h39d11880),
	.w8(32'h39136d5c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c022b95),
	.w1(32'h3c756289),
	.w2(32'h3c224bcc),
	.w3(32'h3c46c33a),
	.w4(32'h3c4b8e7d),
	.w5(32'h3c1c6862),
	.w6(32'h3bc498e8),
	.w7(32'hba32e75d),
	.w8(32'hbaf50312),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cf07b),
	.w1(32'h3896d632),
	.w2(32'h38abd7ee),
	.w3(32'hb4cf7ec4),
	.w4(32'hb761fe54),
	.w5(32'h37854d5e),
	.w6(32'hb7c04ceb),
	.w7(32'hb8547b22),
	.w8(32'hb771d7a6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e20b9b),
	.w1(32'hb9cfea86),
	.w2(32'h3a1fafca),
	.w3(32'hbb329ca9),
	.w4(32'hb9d3fd05),
	.w5(32'h3b2749ba),
	.w6(32'hbbb739b4),
	.w7(32'hbb7ad3f1),
	.w8(32'h3b079830),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38625c0f),
	.w1(32'h38f1a1b6),
	.w2(32'h3a0d2f52),
	.w3(32'h383308a3),
	.w4(32'h3b1eb732),
	.w5(32'h3999c868),
	.w6(32'h36e28a3c),
	.w7(32'hbb05cb75),
	.w8(32'hbaadec05),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec80ae),
	.w1(32'h3c185e36),
	.w2(32'h3c737f6e),
	.w3(32'hb9719e31),
	.w4(32'h3c133aeb),
	.w5(32'h3c25b4a4),
	.w6(32'hbc005cb1),
	.w7(32'hbb341660),
	.w8(32'h3a253b7f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f0d2e),
	.w1(32'h3b7c3d8f),
	.w2(32'h3c989391),
	.w3(32'hbb2d5744),
	.w4(32'h3c6e1560),
	.w5(32'h3c643062),
	.w6(32'hbba6c148),
	.w7(32'h3bd756f3),
	.w8(32'h3bd35396),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8247ac),
	.w1(32'h3b1df844),
	.w2(32'h3c3ba588),
	.w3(32'hba4b6b4f),
	.w4(32'h3bb17969),
	.w5(32'h3b04b30c),
	.w6(32'hba506f6b),
	.w7(32'h3be0fc90),
	.w8(32'h3b703461),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b906f78),
	.w1(32'h3b4e39b9),
	.w2(32'h3b32a129),
	.w3(32'h3b17ff92),
	.w4(32'h3b6ab5bf),
	.w5(32'h3cab11e1),
	.w6(32'h3b2bbfdf),
	.w7(32'hbbcc6e2d),
	.w8(32'h3c4ec59e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbf52e),
	.w1(32'h3ccf64ad),
	.w2(32'h3bd9b1d3),
	.w3(32'h3b6fd8e7),
	.w4(32'h3bba45b7),
	.w5(32'h3c4e9cb2),
	.w6(32'h3c1071df),
	.w7(32'h3c341744),
	.w8(32'h3cc8fb98),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53ae73),
	.w1(32'h3c9a6737),
	.w2(32'h3bfdaffe),
	.w3(32'h3c53b71e),
	.w4(32'h3c194c9b),
	.w5(32'h3c556f4b),
	.w6(32'h3b7bd72e),
	.w7(32'hbbfd29a9),
	.w8(32'h3bf0b3ba),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1b866),
	.w1(32'h3d312f1c),
	.w2(32'h3d5b43c2),
	.w3(32'h3d2ab1c6),
	.w4(32'h3d0511af),
	.w5(32'h3ce9e29e),
	.w6(32'h3c0866de),
	.w7(32'h3b9cfc79),
	.w8(32'h3c69fa57),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa9f3b),
	.w1(32'h3c1a1d5a),
	.w2(32'h3c81c40e),
	.w3(32'h3b85d20d),
	.w4(32'h3b5ec4b2),
	.w5(32'h3c2bb722),
	.w6(32'hbc0f2dc5),
	.w7(32'hbc87b3a2),
	.w8(32'h3b4b95b6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69c55c),
	.w1(32'h3b0702b0),
	.w2(32'h3c3c45b5),
	.w3(32'hbbd2b0ba),
	.w4(32'h3b3feaca),
	.w5(32'h3bba5402),
	.w6(32'hbbcf28f7),
	.w7(32'h3bc4cd45),
	.w8(32'h3bffdc68),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b95e6),
	.w1(32'hbb9cb5bd),
	.w2(32'hbbea8b15),
	.w3(32'hbaddf93a),
	.w4(32'hbbd8dae9),
	.w5(32'hbbee471f),
	.w6(32'hbb598b3e),
	.w7(32'hbbd67c96),
	.w8(32'hbba95d67),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb694e5),
	.w1(32'hbc3435ed),
	.w2(32'h3b936315),
	.w3(32'hbbdddb4d),
	.w4(32'h3ba423bb),
	.w5(32'h3c267a87),
	.w6(32'hbc0da250),
	.w7(32'h3b8e070c),
	.w8(32'h3ba6aa9a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b7c3),
	.w1(32'h3ba39797),
	.w2(32'h3b8f59b6),
	.w3(32'h3b08aecf),
	.w4(32'h36742c2b),
	.w5(32'hbbe46144),
	.w6(32'hb998e262),
	.w7(32'hb7196ae9),
	.w8(32'hbbca58be),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b3b0),
	.w1(32'hbb57f1f0),
	.w2(32'h3bb0a228),
	.w3(32'hbb6d47dd),
	.w4(32'hbbadcdde),
	.w5(32'h3a8f5d3a),
	.w6(32'hbbab6c05),
	.w7(32'hbbdb9925),
	.w8(32'hbb9a0c79),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb689217),
	.w1(32'h3b931ff8),
	.w2(32'h3bf03ab6),
	.w3(32'h3a8019da),
	.w4(32'hb9a34cf2),
	.w5(32'h3ac74b27),
	.w6(32'hbbc9f3fa),
	.w7(32'h3a907de8),
	.w8(32'hbb447777),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9a55),
	.w1(32'h3a078736),
	.w2(32'hbb82ef91),
	.w3(32'hb930bd04),
	.w4(32'hbacd06c1),
	.w5(32'hbbab51de),
	.w6(32'h3c09b8be),
	.w7(32'hbaa2d278),
	.w8(32'hbb8273b9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c66c),
	.w1(32'hbc786859),
	.w2(32'hbb900f82),
	.w3(32'hbc4f7aa9),
	.w4(32'hba862c0b),
	.w5(32'hbb1ed83b),
	.w6(32'hbc377b03),
	.w7(32'h3b89255d),
	.w8(32'hbb2af0b2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa87019),
	.w1(32'h3c09bc5e),
	.w2(32'h3c88cfc2),
	.w3(32'h3b43b13a),
	.w4(32'h3c2becab),
	.w5(32'h3ba076ad),
	.w6(32'hbaac130e),
	.w7(32'hbb936898),
	.w8(32'hbb84999c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde1ddd),
	.w1(32'h3c8ab546),
	.w2(32'h3c1d06a1),
	.w3(32'h3a073087),
	.w4(32'h3b8f5dc8),
	.w5(32'h3b9b7136),
	.w6(32'h3bd793e5),
	.w7(32'h3b4b020a),
	.w8(32'h3b76443e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c4c17),
	.w1(32'h3bd7617c),
	.w2(32'h3c7525f5),
	.w3(32'h3bdaba73),
	.w4(32'h3c19b444),
	.w5(32'h3c1c5085),
	.w6(32'h3b321298),
	.w7(32'h3b4c2f50),
	.w8(32'h3bbb85a7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d157),
	.w1(32'hbc38cf54),
	.w2(32'h3bf9bb78),
	.w3(32'hbc406159),
	.w4(32'h3988a209),
	.w5(32'hbb619550),
	.w6(32'hbcd0b4ad),
	.w7(32'hbc5b35a5),
	.w8(32'hbb81ec06),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f6cb6),
	.w1(32'hbc3be5d2),
	.w2(32'hb97a7d1d),
	.w3(32'hbc390114),
	.w4(32'h3bc76bf0),
	.w5(32'h3c698838),
	.w6(32'hbc872590),
	.w7(32'h3a8f1981),
	.w8(32'h3c3cf2d0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51459),
	.w1(32'h3c985a06),
	.w2(32'h3c0f7c1c),
	.w3(32'h3c720926),
	.w4(32'h3c34f2fa),
	.w5(32'hb9122233),
	.w6(32'h3c90ea54),
	.w7(32'h3c06ec26),
	.w8(32'hba6fe8c8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08ea0a),
	.w1(32'h3bba631a),
	.w2(32'hbc641662),
	.w3(32'h3b987229),
	.w4(32'hbc17046e),
	.w5(32'hbc880dfd),
	.w6(32'h3b3ccca5),
	.w7(32'hbc133d19),
	.w8(32'hbbcbd96a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5025c5),
	.w1(32'hbc0a1892),
	.w2(32'hbbc4d668),
	.w3(32'hbc89fdbf),
	.w4(32'hba4b86e0),
	.w5(32'h3a55e519),
	.w6(32'hbc364fe5),
	.w7(32'hbb49af76),
	.w8(32'hbb1f5ee0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a8de),
	.w1(32'hbbfed940),
	.w2(32'h3c7020ed),
	.w3(32'hbab95549),
	.w4(32'h3be38960),
	.w5(32'h3a69a0d9),
	.w6(32'hbbe5ed1f),
	.w7(32'h3c219b3d),
	.w8(32'hbb16cef5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7882),
	.w1(32'hbc160709),
	.w2(32'h3b2afcf6),
	.w3(32'hbc134773),
	.w4(32'h3c1768ba),
	.w5(32'h3a8c1370),
	.w6(32'hbc3a4989),
	.w7(32'h3c0c831e),
	.w8(32'h3acda6f1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c358efe),
	.w1(32'h3bc9f134),
	.w2(32'hbb807802),
	.w3(32'h3a1a2055),
	.w4(32'h39eec588),
	.w5(32'hbbf5d439),
	.w6(32'h3b54e0ac),
	.w7(32'h3c216f71),
	.w8(32'h3bf1509d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79b9f5),
	.w1(32'hb8f636e6),
	.w2(32'h3b3219c1),
	.w3(32'h3b7050f2),
	.w4(32'hbb8fbb8c),
	.w5(32'hbc2d8752),
	.w6(32'h3b9eb88c),
	.w7(32'hbbf352d9),
	.w8(32'hba6645d6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d1f2),
	.w1(32'hbc38ba24),
	.w2(32'hbb0ae8b1),
	.w3(32'h3af93b9e),
	.w4(32'hbb0abf58),
	.w5(32'hbbfffc76),
	.w6(32'h3b5f9001),
	.w7(32'hbc22095a),
	.w8(32'h3a222599),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55ffeb),
	.w1(32'hbbc1b8be),
	.w2(32'hba6fcd62),
	.w3(32'hba3bec68),
	.w4(32'h3c34c498),
	.w5(32'hba3a1038),
	.w6(32'hbb97c4ec),
	.w7(32'h3c14bc2b),
	.w8(32'hba3f6197),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea8771),
	.w1(32'h3c230e3d),
	.w2(32'hbb5d2077),
	.w3(32'h3b4ba800),
	.w4(32'hb9768106),
	.w5(32'hbb4f9187),
	.w6(32'h3ad63746),
	.w7(32'hbb8887ff),
	.w8(32'hbb1c5805),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b035c4b),
	.w1(32'hbb27a2d0),
	.w2(32'hbb4ecc97),
	.w3(32'hbba77623),
	.w4(32'hbb9f213e),
	.w5(32'hbc3057ed),
	.w6(32'hbaea69a7),
	.w7(32'hba82c572),
	.w8(32'hbc450ead),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6643d),
	.w1(32'h3a0cdc5a),
	.w2(32'h3c6555f5),
	.w3(32'hbc0e238f),
	.w4(32'h3c96c54e),
	.w5(32'h3aa48355),
	.w6(32'hbc242c98),
	.w7(32'h3c080762),
	.w8(32'hbc08c4e4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2129c),
	.w1(32'h3c1b0446),
	.w2(32'hbb9e5fcd),
	.w3(32'h3bbd2c47),
	.w4(32'hbb170f0a),
	.w5(32'hbbc2c08c),
	.w6(32'h3ba5bf17),
	.w7(32'hbb926b4b),
	.w8(32'hbc75fefb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24f354),
	.w1(32'hbb8e94cf),
	.w2(32'hbc1b8ad4),
	.w3(32'h3b56a67b),
	.w4(32'hbb4b4c63),
	.w5(32'hbb81ab3d),
	.w6(32'hbbe2b578),
	.w7(32'hbc02d8d2),
	.w8(32'hbc534cff),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc804705),
	.w1(32'hbc88274f),
	.w2(32'h3a60ca0a),
	.w3(32'hbc958586),
	.w4(32'h3bcd58ac),
	.w5(32'hb8cd3df3),
	.w6(32'hbc642556),
	.w7(32'h3c198941),
	.w8(32'hbb0f1b4d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be072),
	.w1(32'h3b7e44f8),
	.w2(32'h3c27142a),
	.w3(32'h3bb03544),
	.w4(32'h3bc861a6),
	.w5(32'h3c411737),
	.w6(32'h3be62491),
	.w7(32'h3ba3bf3b),
	.w8(32'h3c0e9628),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c471b5e),
	.w1(32'hbbc53dc4),
	.w2(32'h3c5603c8),
	.w3(32'h3b53e97a),
	.w4(32'hba705735),
	.w5(32'h3c5960e7),
	.w6(32'hbb8cb48d),
	.w7(32'hbb8bf8b6),
	.w8(32'h3b8d0b49),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3589e),
	.w1(32'h3bcb7718),
	.w2(32'h3c6d1987),
	.w3(32'h3c79b553),
	.w4(32'h3c918371),
	.w5(32'h3c846488),
	.w6(32'h3a52fe5f),
	.w7(32'h3c2f7369),
	.w8(32'h3bcbe468),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d797f),
	.w1(32'h3c53fc7c),
	.w2(32'hbbd62c31),
	.w3(32'h3c63774d),
	.w4(32'hbc074451),
	.w5(32'h3ad78c6e),
	.w6(32'h3c15eb9c),
	.w7(32'hbbf71f9e),
	.w8(32'h3bff7cef),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc62f56),
	.w1(32'hbca583f8),
	.w2(32'h3b68a77c),
	.w3(32'hbc274e91),
	.w4(32'h3b6bbae1),
	.w5(32'h3ba47db9),
	.w6(32'hbc777b25),
	.w7(32'hbb9eabed),
	.w8(32'hba080ef9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b55dd),
	.w1(32'hba9ef519),
	.w2(32'hb91df7cc),
	.w3(32'hbb5b1273),
	.w4(32'h3bf02efd),
	.w5(32'h3b502ea9),
	.w6(32'hbb24445f),
	.w7(32'h3b3efd8d),
	.w8(32'hba9eda31),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4e80),
	.w1(32'hba9a4642),
	.w2(32'hbb8a75e3),
	.w3(32'hbbaa63d8),
	.w4(32'hbb1148fb),
	.w5(32'h3adbf2d5),
	.w6(32'hbb34b641),
	.w7(32'hbbebf59c),
	.w8(32'hba03d40a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a42a9),
	.w1(32'hbb8e3711),
	.w2(32'h3cb156ae),
	.w3(32'hbc223f28),
	.w4(32'h3c11f3e5),
	.w5(32'h3c6f6658),
	.w6(32'hbc41e6b3),
	.w7(32'h3c91d9f7),
	.w8(32'h3c98dd77),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ce365),
	.w1(32'h3b63bb3c),
	.w2(32'hbbdf6cfd),
	.w3(32'h3c335a1d),
	.w4(32'hbba425ae),
	.w5(32'hbbd1ac86),
	.w6(32'h3be64bc6),
	.w7(32'hbc5cbe39),
	.w8(32'hbc235a3e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46586f),
	.w1(32'hbad5ca9d),
	.w2(32'h3b5da3e0),
	.w3(32'hbb619d1d),
	.w4(32'h3b11724d),
	.w5(32'h390c16b3),
	.w6(32'hbbe547f0),
	.w7(32'hba49a5ba),
	.w8(32'h39853812),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a204f7),
	.w1(32'hbb724d0e),
	.w2(32'h3a2be155),
	.w3(32'hbbe1880a),
	.w4(32'hb9c15e4a),
	.w5(32'h3a84d80e),
	.w6(32'hbb61fcd2),
	.w7(32'h3c172e90),
	.w8(32'h3b4eb7e5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc89e),
	.w1(32'hbc4731b5),
	.w2(32'h39722323),
	.w3(32'hbabf8dcb),
	.w4(32'hbc656741),
	.w5(32'hbc3b9953),
	.w6(32'hbc7e7d45),
	.w7(32'hbbea6176),
	.w8(32'hbb7dccd1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b418bb7),
	.w1(32'hbb813e0e),
	.w2(32'h3b00491f),
	.w3(32'h3c2befba),
	.w4(32'hbb479162),
	.w5(32'h3b77ad33),
	.w6(32'hb99af9c0),
	.w7(32'hbb85ac98),
	.w8(32'h3b35e195),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b104f18),
	.w1(32'h3bea8a4a),
	.w2(32'hbc26d2c6),
	.w3(32'hbb90811f),
	.w4(32'hbbec1ec0),
	.w5(32'hb9e27338),
	.w6(32'hba6cc980),
	.w7(32'hbc396a59),
	.w8(32'hbabc9175),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3f72),
	.w1(32'hbca34065),
	.w2(32'hba3c3060),
	.w3(32'hbc48352c),
	.w4(32'hbbbd5226),
	.w5(32'h3acb14a1),
	.w6(32'hbc92e86a),
	.w7(32'hbc14bdb3),
	.w8(32'hbbae28cd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule