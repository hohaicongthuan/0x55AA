module layer_10_featuremap_435(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74baf8),
	.w1(32'h3b08669f),
	.w2(32'h3abfc129),
	.w3(32'hb98632e9),
	.w4(32'h3b1a5cbb),
	.w5(32'h3a7650b7),
	.w6(32'hbaffc0bf),
	.w7(32'h3b10c245),
	.w8(32'h3af2728a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a342),
	.w1(32'h3b1b5a93),
	.w2(32'hb9d72cce),
	.w3(32'h3a54e190),
	.w4(32'hbb4c8cf9),
	.w5(32'hbb667add),
	.w6(32'hb98430e8),
	.w7(32'hbbd0f966),
	.w8(32'hbbced164),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a1d9d),
	.w1(32'h38a74069),
	.w2(32'h391b6bca),
	.w3(32'hba8dffe1),
	.w4(32'h3a72f558),
	.w5(32'h3a472b95),
	.w6(32'hbaf880fe),
	.w7(32'h398c795b),
	.w8(32'h3aa5fcfc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3a7f9),
	.w1(32'hbac75c23),
	.w2(32'hb9edd27d),
	.w3(32'h3b1a7588),
	.w4(32'hbb18916a),
	.w5(32'h3ab00f55),
	.w6(32'h3b055212),
	.w7(32'hbabd3c08),
	.w8(32'h3a803916),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393343a9),
	.w1(32'h3a72a98c),
	.w2(32'h39e964b6),
	.w3(32'h3ad4a419),
	.w4(32'hb90f5708),
	.w5(32'h3a39a655),
	.w6(32'h3a1bb211),
	.w7(32'hba353232),
	.w8(32'h3a77a66a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a059937),
	.w1(32'h3a266151),
	.w2(32'hbaa0a334),
	.w3(32'h3a1a0eb0),
	.w4(32'h3a8f6a6a),
	.w5(32'hb8ad1f1d),
	.w6(32'h3a9ad141),
	.w7(32'h39ff42ba),
	.w8(32'hba1d8592),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5692c8),
	.w1(32'h38fc5fce),
	.w2(32'hbbaea325),
	.w3(32'h3bcafa8f),
	.w4(32'h379917bc),
	.w5(32'hbc11efa5),
	.w6(32'hbb6266c6),
	.w7(32'hbb6c38b3),
	.w8(32'hbb4007dc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc804bfc),
	.w1(32'hbc633012),
	.w2(32'hbc42d4c7),
	.w3(32'hbc90c2de),
	.w4(32'h3be6d87c),
	.w5(32'h3bfabfc8),
	.w6(32'hbc31ce36),
	.w7(32'hbc0a26d7),
	.w8(32'h3bff0d39),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaee75),
	.w1(32'hbb06cee8),
	.w2(32'hb93a8409),
	.w3(32'hbb17a50d),
	.w4(32'hbb02652f),
	.w5(32'hb971ff73),
	.w6(32'hbaf5c3b9),
	.w7(32'hbb40b8ed),
	.w8(32'hba9fa10e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d2e2),
	.w1(32'h3b99ea0c),
	.w2(32'h3ba68b57),
	.w3(32'h3a9e6c9f),
	.w4(32'h3b638604),
	.w5(32'hba85e2d9),
	.w6(32'hbba3c693),
	.w7(32'hbb0073e0),
	.w8(32'hbac585e0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17551f),
	.w1(32'hba629847),
	.w2(32'hbb03db5c),
	.w3(32'h3a5e887e),
	.w4(32'hb9d2ee24),
	.w5(32'h374e6004),
	.w6(32'h3a2639c5),
	.w7(32'h3a01e24b),
	.w8(32'hb9df041f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cbc36),
	.w1(32'h3b84057c),
	.w2(32'h3ab38861),
	.w3(32'h3bdef726),
	.w4(32'h3b98cd62),
	.w5(32'hbb3a7266),
	.w6(32'hbb598c93),
	.w7(32'h3a36e7c7),
	.w8(32'h3b47a942),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8892fe),
	.w1(32'h3a19bc08),
	.w2(32'hbb4ba63d),
	.w3(32'hb9edf246),
	.w4(32'hb98424ed),
	.w5(32'hbbdf90af),
	.w6(32'hba9ecf3b),
	.w7(32'hbb48e632),
	.w8(32'hbb8f86de),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872263),
	.w1(32'hbb8236dd),
	.w2(32'hbb9b2e1a),
	.w3(32'hba9b6578),
	.w4(32'hbb87d7fe),
	.w5(32'hbb9a6d1d),
	.w6(32'hbb008bd8),
	.w7(32'hbbdfcdd0),
	.w8(32'hbb2a2c9e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed4bb0),
	.w1(32'h3af4e420),
	.w2(32'hbab9da6c),
	.w3(32'h3b7debc4),
	.w4(32'hbb98bf4a),
	.w5(32'hbaff8057),
	.w6(32'h397910bb),
	.w7(32'hbbb4b244),
	.w8(32'hbb7b8150),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90d85),
	.w1(32'h38e77f8e),
	.w2(32'hb8b96cfe),
	.w3(32'hbaf75ad5),
	.w4(32'hbc013b11),
	.w5(32'hbb796a2d),
	.w6(32'hbb95b8f8),
	.w7(32'hbb94d929),
	.w8(32'hba923360),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59355),
	.w1(32'h39d721bf),
	.w2(32'h3a98f462),
	.w3(32'hba9a5c85),
	.w4(32'h3a43bb21),
	.w5(32'h3ab28491),
	.w6(32'hb9775151),
	.w7(32'h3aeb1118),
	.w8(32'h3b06449d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c43d6),
	.w1(32'hbc490d67),
	.w2(32'hbc18b3ab),
	.w3(32'hbc91bd7d),
	.w4(32'hbbdfe41e),
	.w5(32'hbaf70dba),
	.w6(32'hbc40e897),
	.w7(32'h3be399f1),
	.w8(32'h3c4a513c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb739db4),
	.w1(32'hbb6aca6f),
	.w2(32'hba9b5da2),
	.w3(32'hbbd8798e),
	.w4(32'hbb50ed4f),
	.w5(32'h3adb8e46),
	.w6(32'hbbc99506),
	.w7(32'hba669dbd),
	.w8(32'h3b8671e6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d929),
	.w1(32'h3a14be88),
	.w2(32'hbb2ef501),
	.w3(32'hbadf536b),
	.w4(32'hb9d487e3),
	.w5(32'hbabc4fe1),
	.w6(32'hba5b9737),
	.w7(32'h3ad12515),
	.w8(32'hba5fa72d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb132394),
	.w1(32'h39fbfc54),
	.w2(32'hba941fad),
	.w3(32'hbb8d3e46),
	.w4(32'hb94d3888),
	.w5(32'hba0deccf),
	.w6(32'hbb4026ac),
	.w7(32'hba3fa8d5),
	.w8(32'hb9c1327e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2922a),
	.w1(32'h3a9fd49c),
	.w2(32'hbb463c7b),
	.w3(32'h3acecd8e),
	.w4(32'h39edaccc),
	.w5(32'hb9f06484),
	.w6(32'h3b77a57f),
	.w7(32'hb949e746),
	.w8(32'hbb62946e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98fecd),
	.w1(32'hbca8e4e6),
	.w2(32'hbb988a7f),
	.w3(32'hbcc6c342),
	.w4(32'hbb88268a),
	.w5(32'hbaad1aa5),
	.w6(32'hbc9a3d1e),
	.w7(32'h3bf6655f),
	.w8(32'h3c12c895),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acea736),
	.w1(32'h3b886baf),
	.w2(32'h3b5988b9),
	.w3(32'h3b87f15b),
	.w4(32'h39880e0b),
	.w5(32'hbbad7655),
	.w6(32'hba3a1daf),
	.w7(32'hbb8d25a8),
	.w8(32'hbbfb7cf4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0e01e),
	.w1(32'h3b5a0f79),
	.w2(32'h3bd32c1e),
	.w3(32'h3a1c5d1b),
	.w4(32'hbb82639d),
	.w5(32'hbb5e26be),
	.w6(32'hbb463ae3),
	.w7(32'hbc78bce3),
	.w8(32'hbc4db9aa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc6e2),
	.w1(32'h39bc253d),
	.w2(32'hbab7d630),
	.w3(32'hbadc367c),
	.w4(32'h38feeb18),
	.w5(32'hbab30eb7),
	.w6(32'hba5b6084),
	.w7(32'hb9ffaa10),
	.w8(32'hba8eb70e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace1f3e),
	.w1(32'h3abed0c7),
	.w2(32'h3a118874),
	.w3(32'hba74f1b2),
	.w4(32'h3a86f74e),
	.w5(32'h3a377213),
	.w6(32'hba6d147d),
	.w7(32'hba84518e),
	.w8(32'hbaa2b453),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c6f4),
	.w1(32'hb9663b75),
	.w2(32'hbb4fafba),
	.w3(32'h3b30c4fb),
	.w4(32'hbb62a957),
	.w5(32'hbc936f49),
	.w6(32'h3b9067bd),
	.w7(32'h3ab457ad),
	.w8(32'hbbb7b934),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e18444),
	.w1(32'h3a4d9d94),
	.w2(32'h39269a53),
	.w3(32'h393cf454),
	.w4(32'hb961f82f),
	.w5(32'hb9895c1e),
	.w6(32'h396c9e54),
	.w7(32'hb95e6f0b),
	.w8(32'h3aa77022),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a5eb),
	.w1(32'h3be3d577),
	.w2(32'h3bcce17f),
	.w3(32'h3c15298d),
	.w4(32'hbba482d4),
	.w5(32'hbc25dae1),
	.w6(32'h3c46c405),
	.w7(32'hbba1ef92),
	.w8(32'hbc346d05),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75f810),
	.w1(32'h3ad15a2c),
	.w2(32'h3b04be8f),
	.w3(32'h3aee1d80),
	.w4(32'hb90c19c2),
	.w5(32'hb98cacce),
	.w6(32'h3b63e67d),
	.w7(32'h3abcd7b1),
	.w8(32'h3a4fb1ea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6fa3),
	.w1(32'hbb462e69),
	.w2(32'hbaf460c2),
	.w3(32'hbaa560d1),
	.w4(32'hbafa9569),
	.w5(32'hbae1814b),
	.w6(32'h39d6d241),
	.w7(32'hbab061ac),
	.w8(32'hb7abb068),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c7bc),
	.w1(32'h3b22d9e0),
	.w2(32'h3afc267f),
	.w3(32'h3abb3ca5),
	.w4(32'h3b522da9),
	.w5(32'h3a39281e),
	.w6(32'hb8d943ad),
	.w7(32'h3a822edd),
	.w8(32'h3b2a6f76),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9643),
	.w1(32'hba12489d),
	.w2(32'h3acc764e),
	.w3(32'hba66fcf3),
	.w4(32'hbb22af81),
	.w5(32'hbacd0aa3),
	.w6(32'hbb07eec0),
	.w7(32'hbbb6aeb6),
	.w8(32'hbbaefce2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ad3f4),
	.w1(32'hba2c232c),
	.w2(32'h3a640152),
	.w3(32'hba15ffb1),
	.w4(32'hbb44fbd6),
	.w5(32'hbaaa0c08),
	.w6(32'hbac76738),
	.w7(32'hbb463754),
	.w8(32'h3a8bf72c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee5f0),
	.w1(32'h3ab2e610),
	.w2(32'h3b11473b),
	.w3(32'hbb7c5f68),
	.w4(32'h3b0a1eb1),
	.w5(32'h3b4832ef),
	.w6(32'hbb78b94d),
	.w7(32'h3a04e6d3),
	.w8(32'h3ad7b8e4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0044),
	.w1(32'hbb267e12),
	.w2(32'hb9bd6e3d),
	.w3(32'hbab4d97a),
	.w4(32'hba7847e3),
	.w5(32'hbae50a6f),
	.w6(32'hbc465eba),
	.w7(32'hbc69e22f),
	.w8(32'hba906442),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13a925),
	.w1(32'h3b447be2),
	.w2(32'hbb3cc98c),
	.w3(32'h3b9f7868),
	.w4(32'hbc191db4),
	.w5(32'hbc6c138d),
	.w6(32'hbb5aaf1d),
	.w7(32'hbc82271b),
	.w8(32'hbc8b863f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d1130),
	.w1(32'h3b74ee5f),
	.w2(32'hbc0750a8),
	.w3(32'h3c8b5ae9),
	.w4(32'hbbc75e61),
	.w5(32'hbc9f7300),
	.w6(32'h3c586640),
	.w7(32'hbbd66ff0),
	.w8(32'hbc81b2f4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf5f87),
	.w1(32'hba87a886),
	.w2(32'h39d2c279),
	.w3(32'hbb0fce4d),
	.w4(32'hbb30f39b),
	.w5(32'hbabbc9e6),
	.w6(32'hbb5f1734),
	.w7(32'hbb96cfbf),
	.w8(32'hbada265b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a4322),
	.w1(32'hbac94d53),
	.w2(32'hbadf66ad),
	.w3(32'hb89dbc0a),
	.w4(32'hbb96d223),
	.w5(32'hbb458b14),
	.w6(32'hbaacb3be),
	.w7(32'hbb6bbd40),
	.w8(32'hbb2f5b3a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cc57e),
	.w1(32'h3a0f197a),
	.w2(32'hbaaaa205),
	.w3(32'hbb41fef0),
	.w4(32'hbae433f0),
	.w5(32'hbaac65fc),
	.w6(32'hbb8bc1b7),
	.w7(32'hbaa97f65),
	.w8(32'hbb124455),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7edf58),
	.w1(32'hbac4a37d),
	.w2(32'h3af2a65f),
	.w3(32'hbad99c6c),
	.w4(32'hba30b5f5),
	.w5(32'h3abd1fff),
	.w6(32'hbacb0c11),
	.w7(32'hb9918969),
	.w8(32'hb8adda6f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92546b),
	.w1(32'h3b31ba7a),
	.w2(32'hbb86433f),
	.w3(32'hb9582376),
	.w4(32'h39688954),
	.w5(32'hbb60dc80),
	.w6(32'hbb6216c7),
	.w7(32'h3bec983d),
	.w8(32'h3b9a692b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77c6714),
	.w1(32'h3b5647a1),
	.w2(32'h3b6430ca),
	.w3(32'h3b72593a),
	.w4(32'hba1760e9),
	.w5(32'hbb36f4ad),
	.w6(32'h3b3cb2d8),
	.w7(32'hbbc35d91),
	.w8(32'hbbc1c979),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f645),
	.w1(32'h3bdfdc19),
	.w2(32'h3be48e17),
	.w3(32'h3b00f9d7),
	.w4(32'h3abb69fe),
	.w5(32'h3b50f148),
	.w6(32'hbb09d31d),
	.w7(32'hbbe1a58c),
	.w8(32'hbbd14819),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95ecbd),
	.w1(32'hbb44d2e5),
	.w2(32'h3a668a12),
	.w3(32'hbbb0fd3b),
	.w4(32'hbb05f6a7),
	.w5(32'h396ffcd6),
	.w6(32'hbc1cd00f),
	.w7(32'hbb9a3602),
	.w8(32'hbb0c9eae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8def61),
	.w1(32'hbc8e23d1),
	.w2(32'hbc2ee677),
	.w3(32'hbcb5750c),
	.w4(32'hbba34f50),
	.w5(32'h3b6d4f48),
	.w6(32'hbcbad60b),
	.w7(32'h3b218854),
	.w8(32'h3c45c849),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43b420),
	.w1(32'h3a814c7c),
	.w2(32'h3a324dc8),
	.w3(32'hbb3b6abb),
	.w4(32'h387301f7),
	.w5(32'h3ab21bc2),
	.w6(32'hbb1737af),
	.w7(32'h3a2cb97e),
	.w8(32'h3a5eeb40),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c79a29),
	.w1(32'h394884c2),
	.w2(32'hb97e62c4),
	.w3(32'hbadc4620),
	.w4(32'hb9d5aae3),
	.w5(32'h3a00bc3a),
	.w6(32'hbae830a3),
	.w7(32'hb9cb18bc),
	.w8(32'h3a25770a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac56d3b),
	.w1(32'hbaad15ec),
	.w2(32'hba5df9cd),
	.w3(32'h3ab40ff7),
	.w4(32'hba6342c0),
	.w5(32'hbab2db4d),
	.w6(32'hb884cedc),
	.w7(32'hbae7cb1e),
	.w8(32'hba86a8c6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b111),
	.w1(32'hba8c0154),
	.w2(32'hbbe55f84),
	.w3(32'hbb08f460),
	.w4(32'hba98b876),
	.w5(32'hbb95b3c7),
	.w6(32'hbb2c82c4),
	.w7(32'h3a02836a),
	.w8(32'hbbba2615),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ceb5),
	.w1(32'hba849031),
	.w2(32'h389f0edc),
	.w3(32'hbbb78784),
	.w4(32'h39ff35c6),
	.w5(32'h3b0cc243),
	.w6(32'hbbbd9419),
	.w7(32'h3a1a5458),
	.w8(32'h39abb184),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f78af),
	.w1(32'hbc44819b),
	.w2(32'hbb9ebfad),
	.w3(32'hbc505b79),
	.w4(32'hbb4632db),
	.w5(32'h3b02ed5b),
	.w6(32'hbc4bf072),
	.w7(32'h3a23a05c),
	.w8(32'h3c203284),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0216f),
	.w1(32'hbba2e6b1),
	.w2(32'hbb10d40f),
	.w3(32'hbaed8390),
	.w4(32'hb9fc0a92),
	.w5(32'h3ad01067),
	.w6(32'h3962fc33),
	.w7(32'hb90c8dac),
	.w8(32'h39a3b77b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c37d0),
	.w1(32'hbaf3dee5),
	.w2(32'h39e4b477),
	.w3(32'hba5ba965),
	.w4(32'hbab2c4b3),
	.w5(32'h3a95d01f),
	.w6(32'hb9ed47d8),
	.w7(32'hbae6c050),
	.w8(32'h3882a7f6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a970),
	.w1(32'h3ac2e217),
	.w2(32'h3b1dbaaf),
	.w3(32'hb9804e1f),
	.w4(32'h3a413065),
	.w5(32'h3a8ce081),
	.w6(32'h39bcab8e),
	.w7(32'h39907a4c),
	.w8(32'h3adc2dac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d54ed),
	.w1(32'hbaf17283),
	.w2(32'hbb905182),
	.w3(32'h3b29e63d),
	.w4(32'hba0ba329),
	.w5(32'hbb55a981),
	.w6(32'h3b478ace),
	.w7(32'hba48e4be),
	.w8(32'hbbb10171),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad5e59),
	.w1(32'hbb0382a7),
	.w2(32'hbb255924),
	.w3(32'hba6c8120),
	.w4(32'hba46f54d),
	.w5(32'hba82c7a8),
	.w6(32'hbb004c31),
	.w7(32'hbadde4c6),
	.w8(32'hbabe5ec5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a277),
	.w1(32'hbac88e4d),
	.w2(32'h390d6bb8),
	.w3(32'hba91f65c),
	.w4(32'hba476736),
	.w5(32'hba257cf9),
	.w6(32'hb9f63cee),
	.w7(32'hbab13dbf),
	.w8(32'hba67adcc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd7ea9),
	.w1(32'hbb54ff13),
	.w2(32'hbb29cee6),
	.w3(32'hbba5d308),
	.w4(32'hba8bf58f),
	.w5(32'h3a845abb),
	.w6(32'hbba1557f),
	.w7(32'h39bbfd58),
	.w8(32'h3ac1ee28),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc532549),
	.w1(32'hbb8c481c),
	.w2(32'hbba48864),
	.w3(32'hbc2d7843),
	.w4(32'hbaf24851),
	.w5(32'hbc0293d1),
	.w6(32'hba290801),
	.w7(32'h3b95e91d),
	.w8(32'hba88f11e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b48885),
	.w1(32'hbb27e139),
	.w2(32'hba8f55f2),
	.w3(32'h39ec42ec),
	.w4(32'hbb63e2b7),
	.w5(32'hbac6443f),
	.w6(32'hba0e7d43),
	.w7(32'hba96a0b2),
	.w8(32'hb683d826),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0151e9),
	.w1(32'h3a734fa8),
	.w2(32'h3a225d70),
	.w3(32'h38879711),
	.w4(32'h39bc380d),
	.w5(32'h3aaeb59c),
	.w6(32'hb7a4a405),
	.w7(32'hb8b20a6e),
	.w8(32'h3b046199),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b6b0d),
	.w1(32'h3b1b3202),
	.w2(32'h3b560727),
	.w3(32'h3a3a4adf),
	.w4(32'h3b118626),
	.w5(32'h3ad69a95),
	.w6(32'h3a77aaf2),
	.w7(32'h3b2edfcb),
	.w8(32'h3b6d8c23),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463d50),
	.w1(32'h3b57959e),
	.w2(32'h3b055429),
	.w3(32'h3b4ddc88),
	.w4(32'h3a6f4298),
	.w5(32'h39af112f),
	.w6(32'h3b583024),
	.w7(32'h3a6eae51),
	.w8(32'hba82723d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c051b),
	.w1(32'h3be737c0),
	.w2(32'h3c13596d),
	.w3(32'h3c013da4),
	.w4(32'h3ba3afa5),
	.w5(32'hbb7185f4),
	.w6(32'hbc1c4a1f),
	.w7(32'h3c0653a3),
	.w8(32'h3c52d49e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96ac11),
	.w1(32'h3b66e4d0),
	.w2(32'h3b6c0237),
	.w3(32'hb81c4ad0),
	.w4(32'h393109a6),
	.w5(32'h3b9c4d92),
	.w6(32'hbba04f4d),
	.w7(32'hbbb071ab),
	.w8(32'hbbf4f3fb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c5b4e),
	.w1(32'hbc0f0c07),
	.w2(32'hbb1996b4),
	.w3(32'hbb3cffbd),
	.w4(32'h3a8f1af2),
	.w5(32'h3ae355be),
	.w6(32'hbaaa4a4e),
	.w7(32'h3b71d750),
	.w8(32'h3b694c88),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a0d9),
	.w1(32'h3c052f4a),
	.w2(32'h3b4ac411),
	.w3(32'h3b2ba700),
	.w4(32'hbb7cc390),
	.w5(32'hbc5f046a),
	.w6(32'hbb11335c),
	.w7(32'hbc837474),
	.w8(32'hbc813ed2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1185f),
	.w1(32'h3b31aa66),
	.w2(32'h3b2c603b),
	.w3(32'hbba68f87),
	.w4(32'h3b41dd1f),
	.w5(32'h3bb34382),
	.w6(32'hbbdfc9e4),
	.w7(32'h3b261ac6),
	.w8(32'h3ba5d148),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f349ef),
	.w1(32'h3b9e84cf),
	.w2(32'hba9cd617),
	.w3(32'h3b1cfb91),
	.w4(32'h3a555e60),
	.w5(32'h3ae0d782),
	.w6(32'hb9a43a94),
	.w7(32'hb8ca8f70),
	.w8(32'h3b968a2c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8eb5),
	.w1(32'h3bc5720b),
	.w2(32'h39bfb53c),
	.w3(32'h3b541798),
	.w4(32'h3b8f9355),
	.w5(32'h3b183340),
	.w6(32'hbaafdf46),
	.w7(32'h3ba288f4),
	.w8(32'h3b1aa760),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72cad3),
	.w1(32'hbc6b0d90),
	.w2(32'hbc52181b),
	.w3(32'hb97f434a),
	.w4(32'hbbe91c14),
	.w5(32'hbbfd19ae),
	.w6(32'h3a50b87b),
	.w7(32'hbc1e427d),
	.w8(32'hbc236e84),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136fae),
	.w1(32'h3afa1977),
	.w2(32'h3b0384b9),
	.w3(32'hbc1f4876),
	.w4(32'hbc1bed5a),
	.w5(32'hbb4fec35),
	.w6(32'hbc848e82),
	.w7(32'hbbef25f8),
	.w8(32'hbab753f3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f33b),
	.w1(32'hbc938470),
	.w2(32'hbbd5a5c1),
	.w3(32'hbc4d104e),
	.w4(32'hbc39601a),
	.w5(32'hbac473ec),
	.w6(32'hbaa53cb9),
	.w7(32'hbbae57cf),
	.w8(32'h3bba51de),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fd469),
	.w1(32'hbc47e42e),
	.w2(32'hbbb2b53d),
	.w3(32'hbc22ac90),
	.w4(32'hbc4574a7),
	.w5(32'h3c02702b),
	.w6(32'hbc97a34a),
	.w7(32'hbb7817e7),
	.w8(32'h3c39dcd3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d79a3),
	.w1(32'h3b9975f0),
	.w2(32'h3b4feab3),
	.w3(32'h3bcf93dd),
	.w4(32'hbb4fb2a6),
	.w5(32'hbbfba607),
	.w6(32'h3b8631c4),
	.w7(32'hbc07f757),
	.w8(32'hbc3745bc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cfe70),
	.w1(32'h3bcd6ed4),
	.w2(32'h3c178cf2),
	.w3(32'hbb8fe7b2),
	.w4(32'h3c277db7),
	.w5(32'h3c1f44bf),
	.w6(32'h3b576276),
	.w7(32'h3c157b1d),
	.w8(32'h3ba1c543),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc29696),
	.w1(32'hbc1bbf31),
	.w2(32'h39a0450a),
	.w3(32'h3c2c9cb8),
	.w4(32'hb9f42f24),
	.w5(32'hbc173e92),
	.w6(32'hbaac0afe),
	.w7(32'hba99c637),
	.w8(32'h3b8017d3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aa7f6),
	.w1(32'h3aa8ccb0),
	.w2(32'h3c011006),
	.w3(32'h3b81df29),
	.w4(32'h39831814),
	.w5(32'h3b003c20),
	.w6(32'hbb0d0c90),
	.w7(32'hbb2c9574),
	.w8(32'hbb932817),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3830f2),
	.w1(32'hbc8a73f9),
	.w2(32'hbc50c656),
	.w3(32'hbb52ce5e),
	.w4(32'hbc2becb1),
	.w5(32'hbbce0c0b),
	.w6(32'hbbe6daba),
	.w7(32'hbb0a54e4),
	.w8(32'h39bde650),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ddfe),
	.w1(32'hb902f962),
	.w2(32'h3a94dfda),
	.w3(32'hbb832cd3),
	.w4(32'hbaa9e77a),
	.w5(32'hb9d5c1a8),
	.w6(32'h373663f1),
	.w7(32'h39416703),
	.w8(32'hbb27a66f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc584),
	.w1(32'h3b01d35d),
	.w2(32'hba82fc8e),
	.w3(32'h3ab00549),
	.w4(32'h3a6459c6),
	.w5(32'hbb8d68e0),
	.w6(32'hb9b84bff),
	.w7(32'hbba6051e),
	.w8(32'hbbcc9ce6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f6fb),
	.w1(32'hbbe8197f),
	.w2(32'hbc004d78),
	.w3(32'hba409c09),
	.w4(32'hbbfb0ebb),
	.w5(32'hbc508e3c),
	.w6(32'hb931b9ee),
	.w7(32'h3a9b3a42),
	.w8(32'hbb79ef21),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d18a),
	.w1(32'h3ae4e96d),
	.w2(32'hbb583280),
	.w3(32'hbc0afc2b),
	.w4(32'h3c10211c),
	.w5(32'hbb0abbda),
	.w6(32'hbb8e3cd1),
	.w7(32'hbb65c2b2),
	.w8(32'hbb493459),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb018162),
	.w1(32'h3b6894ba),
	.w2(32'h3b17a10d),
	.w3(32'hb9a81b28),
	.w4(32'hbba9748e),
	.w5(32'hbc557d02),
	.w6(32'hbb64d45f),
	.w7(32'hbbe9bc42),
	.w8(32'hbc4e35b7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151db3),
	.w1(32'hbb785f4e),
	.w2(32'hbb2ce0fe),
	.w3(32'hbbe2f66e),
	.w4(32'hbba69a72),
	.w5(32'hbbaa457a),
	.w6(32'hbb280a90),
	.w7(32'hbb9b30c1),
	.w8(32'h3af740db),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e1a86),
	.w1(32'h3ae0cf13),
	.w2(32'h3b32bbc9),
	.w3(32'hbbc20711),
	.w4(32'hbaa04086),
	.w5(32'h3b6405ed),
	.w6(32'hba380ccb),
	.w7(32'hbbef66c5),
	.w8(32'hbc001ebf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc831bf3),
	.w1(32'hbc2ca2d4),
	.w2(32'hbad0f5bf),
	.w3(32'hbc98a8c7),
	.w4(32'hbb5bf597),
	.w5(32'h3c0654b7),
	.w6(32'hbc6b7283),
	.w7(32'h3abe5afe),
	.w8(32'h3c24ece3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56ae1c),
	.w1(32'h3c08a657),
	.w2(32'hbb6b2879),
	.w3(32'h3c00ab28),
	.w4(32'h3a8057f6),
	.w5(32'hbc0de9db),
	.w6(32'h3b84a99f),
	.w7(32'h3a2ee4ee),
	.w8(32'hbbf6132a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbced29e),
	.w1(32'h3b36b3af),
	.w2(32'h3b2d68c1),
	.w3(32'hbb3a660b),
	.w4(32'hb79765f2),
	.w5(32'hbc16cc47),
	.w6(32'hbbb57bb6),
	.w7(32'hba6c00f8),
	.w8(32'h3b720d3d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2509e4),
	.w1(32'h3b1e44fc),
	.w2(32'hbb01deaf),
	.w3(32'hb95e12db),
	.w4(32'h3b94be71),
	.w5(32'h3afdf62e),
	.w6(32'h3b372aa4),
	.w7(32'hbb7cd7c5),
	.w8(32'hbbc57001),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b1f6),
	.w1(32'h3ae04de8),
	.w2(32'h3be7f449),
	.w3(32'h3bae5ac5),
	.w4(32'h3c049d86),
	.w5(32'h3c2d8dec),
	.w6(32'hbb8c83d3),
	.w7(32'hbaba919f),
	.w8(32'h3bee9815),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a396e7f),
	.w1(32'h3b642c0f),
	.w2(32'h3bb9c22c),
	.w3(32'h3c22851f),
	.w4(32'hbad6b05f),
	.w5(32'hbb4b1f22),
	.w6(32'h38fa7f1f),
	.w7(32'hbb9ca697),
	.w8(32'h3a1e56cc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e0e4),
	.w1(32'h3bcb8519),
	.w2(32'hbb868c7e),
	.w3(32'h3bec8a67),
	.w4(32'hbaf40c6b),
	.w5(32'hbc148c42),
	.w6(32'h3b767379),
	.w7(32'hba0c3794),
	.w8(32'hbb9c4e26),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059ed7),
	.w1(32'h3a01d442),
	.w2(32'hbc159ff8),
	.w3(32'h3b3cc81e),
	.w4(32'hbb896d48),
	.w5(32'hbbc6866d),
	.w6(32'hbb66fc41),
	.w7(32'hbbd0004a),
	.w8(32'hbb971466),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f2b31),
	.w1(32'hbbf316d0),
	.w2(32'hbb95619f),
	.w3(32'hbc12efb0),
	.w4(32'hbb07b369),
	.w5(32'hbb076e82),
	.w6(32'hbc5237e7),
	.w7(32'hbab7fb01),
	.w8(32'hbb701aeb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9edf),
	.w1(32'h3b798e9b),
	.w2(32'h3bc28b50),
	.w3(32'h3c9d986d),
	.w4(32'h3b91b09a),
	.w5(32'hbc63be4b),
	.w6(32'h3bc2e352),
	.w7(32'h3b904d3b),
	.w8(32'h3b73deed),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc590498),
	.w1(32'hbc85efef),
	.w2(32'hbc047491),
	.w3(32'hbd182081),
	.w4(32'hbc8a192a),
	.w5(32'h3a94b47a),
	.w6(32'hbce6990a),
	.w7(32'hbc4182db),
	.w8(32'h3b885075),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06ce6a),
	.w1(32'hbbf6c460),
	.w2(32'hbc98df10),
	.w3(32'h3ac8310e),
	.w4(32'hbbe052bb),
	.w5(32'hbc8a1dd0),
	.w6(32'hba506185),
	.w7(32'hbc6da306),
	.w8(32'hbc962c89),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36f197),
	.w1(32'hbb848b45),
	.w2(32'h381dbf5d),
	.w3(32'hbac91a94),
	.w4(32'hbc0c3b13),
	.w5(32'hbc58bd04),
	.w6(32'hbc2e61d6),
	.w7(32'hbc8be223),
	.w8(32'hbc9770ec),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f019e),
	.w1(32'h3c1d5867),
	.w2(32'h3b3a8ac8),
	.w3(32'hbb5c72ab),
	.w4(32'h3bd4307f),
	.w5(32'h3b78aa08),
	.w6(32'hbc70c207),
	.w7(32'h3c5bd017),
	.w8(32'h3c563104),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0493),
	.w1(32'hbc7e092e),
	.w2(32'hbc4da5f6),
	.w3(32'h3b54b744),
	.w4(32'hbc2912a1),
	.w5(32'hbc5af2b1),
	.w6(32'h3c3ae689),
	.w7(32'hbbbf718b),
	.w8(32'hbc2d4e98),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd099380),
	.w1(32'hbd14b839),
	.w2(32'hbcf2c8d8),
	.w3(32'hbd0961b3),
	.w4(32'hbc349ee8),
	.w5(32'hbb5ea72b),
	.w6(32'hbd278769),
	.w7(32'hbbeec727),
	.w8(32'h3beb52af),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b923ad1),
	.w1(32'h3a6e98c0),
	.w2(32'hbc0757b2),
	.w3(32'h3c13fd83),
	.w4(32'hbb2f6c39),
	.w5(32'hbc69b7e8),
	.w6(32'h3bd24ebd),
	.w7(32'h3a8b296e),
	.w8(32'hbbc95410),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d1718),
	.w1(32'hbbdb6a33),
	.w2(32'hbba02392),
	.w3(32'h3b116add),
	.w4(32'hbb6a9a01),
	.w5(32'hbb5d34c9),
	.w6(32'h3ad7f9f3),
	.w7(32'h3b815940),
	.w8(32'h3a9ea146),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70f7b8),
	.w1(32'h3b43e9e9),
	.w2(32'hba600ecb),
	.w3(32'hbb2eee92),
	.w4(32'hb99b2764),
	.w5(32'hbb49598c),
	.w6(32'hbb3a52df),
	.w7(32'h3b717b45),
	.w8(32'h3b3b32a1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b309117),
	.w1(32'h3c0878fa),
	.w2(32'h3b7b0c0a),
	.w3(32'h3b114c34),
	.w4(32'h3abb79aa),
	.w5(32'hbbadb4b2),
	.w6(32'h3b0fd817),
	.w7(32'hba2de2b1),
	.w8(32'hbad8491c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ca928),
	.w1(32'h3bd92781),
	.w2(32'h3baed440),
	.w3(32'hb92fc1c0),
	.w4(32'h3b8d0e4d),
	.w5(32'hbbbc15a6),
	.w6(32'h3b21fc84),
	.w7(32'hbbdf0cbd),
	.w8(32'hbbbd9153),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4cf47),
	.w1(32'h3bec44d2),
	.w2(32'h39f1551b),
	.w3(32'h3c6a62d9),
	.w4(32'hba4dece5),
	.w5(32'hbc0f712e),
	.w6(32'h3c957745),
	.w7(32'hbb77faa7),
	.w8(32'hbbb8bfb6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8813),
	.w1(32'h3c426af8),
	.w2(32'h3bc090e4),
	.w3(32'h3b9f1900),
	.w4(32'h3b9477e2),
	.w5(32'hba14d7e6),
	.w6(32'h3b636849),
	.w7(32'hbbc39f17),
	.w8(32'hbbbeeb60),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52fd86),
	.w1(32'h3be504c4),
	.w2(32'h3c20bedb),
	.w3(32'hbb40b82d),
	.w4(32'h3b974816),
	.w5(32'h3c67474b),
	.w6(32'hbab468a2),
	.w7(32'h3b32298a),
	.w8(32'h3c022b99),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf12d),
	.w1(32'hbbe0a72b),
	.w2(32'hb8d81238),
	.w3(32'h3b1bbd71),
	.w4(32'hbbd6169f),
	.w5(32'hbbd6e356),
	.w6(32'h3a56fbfe),
	.w7(32'hb93f61b2),
	.w8(32'h3c026c61),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e00dd),
	.w1(32'h3b4adba8),
	.w2(32'h3b89eacf),
	.w3(32'h3bf2bcc2),
	.w4(32'h3b2966c1),
	.w5(32'hbb60378b),
	.w6(32'h3be10102),
	.w7(32'hbb91db7b),
	.w8(32'hbc0a8387),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6b48),
	.w1(32'h3b5a7997),
	.w2(32'h39b42fae),
	.w3(32'h3b2ae7f5),
	.w4(32'h3a82401e),
	.w5(32'h3b01eafe),
	.w6(32'hbbcb7226),
	.w7(32'hba3b1247),
	.w8(32'h3abf8937),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189274),
	.w1(32'h3c04e458),
	.w2(32'h3c0617b5),
	.w3(32'hba3eff1c),
	.w4(32'h3bb8c02c),
	.w5(32'h3c024a93),
	.w6(32'hba596ba4),
	.w7(32'h3b988440),
	.w8(32'h3ba053be),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122c31),
	.w1(32'h3ade90c3),
	.w2(32'h3b85b0b0),
	.w3(32'h3c4c03ec),
	.w4(32'h3c8c9e6e),
	.w5(32'h3ca398ff),
	.w6(32'h3c009103),
	.w7(32'h3c47940d),
	.w8(32'h3c58fdc0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24bbba),
	.w1(32'hbb03acfd),
	.w2(32'hbbd5e429),
	.w3(32'h3cb9d8e8),
	.w4(32'hb9da2da7),
	.w5(32'hbae108e1),
	.w6(32'h3c7a3e6a),
	.w7(32'h3b2285c7),
	.w8(32'h3b2bc077),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39017efc),
	.w1(32'hbc2c5d05),
	.w2(32'hbc28a923),
	.w3(32'h3ac8a14e),
	.w4(32'hbbf36c74),
	.w5(32'hbc798101),
	.w6(32'h3af730e9),
	.w7(32'hbc369b31),
	.w8(32'hbc5e5399),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ab37),
	.w1(32'h38fff3c6),
	.w2(32'h3b6216bb),
	.w3(32'hbc6966fd),
	.w4(32'hbaf6bdc3),
	.w5(32'h3bbaf49a),
	.w6(32'hbc8859bb),
	.w7(32'h3a53ef71),
	.w8(32'h3a409e2f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8e56),
	.w1(32'h3b9836d7),
	.w2(32'hba94143b),
	.w3(32'h39f9e637),
	.w4(32'hbae32c3a),
	.w5(32'hbb7e25a7),
	.w6(32'hbb8a6697),
	.w7(32'hba8409ac),
	.w8(32'hbb7bed32),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c2b88),
	.w1(32'h3c22df85),
	.w2(32'h3b1c01a1),
	.w3(32'hba20a135),
	.w4(32'hbb8dd6ac),
	.w5(32'hbb6b83e8),
	.w6(32'h3aadb365),
	.w7(32'hbc1699f1),
	.w8(32'hbbd39f6e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97c04f),
	.w1(32'h3b6d0731),
	.w2(32'h3a9ffcc9),
	.w3(32'h3bd55e62),
	.w4(32'h3b6f555c),
	.w5(32'hbb976ce0),
	.w6(32'h3c4b4d75),
	.w7(32'hba268bfd),
	.w8(32'hbbbfff76),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab449ff),
	.w1(32'h3c2f53b7),
	.w2(32'h3b680f5a),
	.w3(32'hbba264f0),
	.w4(32'h3c4ec7f5),
	.w5(32'h3c036f7c),
	.w6(32'h39d15d6b),
	.w7(32'h3c4e8817),
	.w8(32'h3c29f849),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b895f0d),
	.w1(32'h3c814f1f),
	.w2(32'h3c5b3073),
	.w3(32'h3c3bf5c9),
	.w4(32'h3c968d4c),
	.w5(32'h3c9e648d),
	.w6(32'h3c62fd39),
	.w7(32'h3c6abc0f),
	.w8(32'h3c7fb8ce),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c804d75),
	.w1(32'h3b12bd08),
	.w2(32'h3b69b317),
	.w3(32'h3cc14e62),
	.w4(32'hbb28a8b1),
	.w5(32'hbb92b4fa),
	.w6(32'h3c5bcd62),
	.w7(32'hbb36ee5e),
	.w8(32'hba879b40),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31ae7d),
	.w1(32'h3c22e06b),
	.w2(32'h3af85b52),
	.w3(32'hbbcc9d94),
	.w4(32'h3b949302),
	.w5(32'hbb4ac061),
	.w6(32'hbbb50f9f),
	.w7(32'h3b4d35c4),
	.w8(32'hbafe2583),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcc40a),
	.w1(32'hbb20bee6),
	.w2(32'h3afba34d),
	.w3(32'hbb9ece4e),
	.w4(32'hbb9e13cb),
	.w5(32'hbbc09106),
	.w6(32'hbb8b0a92),
	.w7(32'hbb8d0121),
	.w8(32'h3acdb1b5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb731152),
	.w1(32'hb91a1146),
	.w2(32'h3c259191),
	.w3(32'hbbd9832a),
	.w4(32'h3ba2f47c),
	.w5(32'h3bf80fe9),
	.w6(32'hbb96dfed),
	.w7(32'h3be7fee8),
	.w8(32'h3c43814b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c300cd0),
	.w1(32'hbc81ad83),
	.w2(32'hbc78c2c4),
	.w3(32'h3c293500),
	.w4(32'hbc266a9b),
	.w5(32'hbc715305),
	.w6(32'h3c00ea8c),
	.w7(32'hbc2fffb4),
	.w8(32'hbc0e1b9f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57368d),
	.w1(32'h3a87aa85),
	.w2(32'hbb35d6b4),
	.w3(32'hbc0ff5ce),
	.w4(32'h3bbf8d2c),
	.w5(32'h3c078e70),
	.w6(32'hb9e7ff6b),
	.w7(32'h39b2e2f3),
	.w8(32'h3bb77c78),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282708),
	.w1(32'hbabfab5a),
	.w2(32'hba118302),
	.w3(32'h3c08084a),
	.w4(32'hb89bea01),
	.w5(32'hbb55266c),
	.w6(32'h3a735197),
	.w7(32'hbb0227f9),
	.w8(32'hbb882009),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb038449),
	.w1(32'h3b9985ba),
	.w2(32'h3c0ed5b0),
	.w3(32'h3a25c7c4),
	.w4(32'h3b1b1eb2),
	.w5(32'h3b3d38e2),
	.w6(32'h3823106a),
	.w7(32'hba83216e),
	.w8(32'hbae46214),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58f134),
	.w1(32'hbc62b578),
	.w2(32'hbc1528ad),
	.w3(32'hbc0a1d00),
	.w4(32'hbbc3034b),
	.w5(32'hbbed886c),
	.w6(32'hbc7794c1),
	.w7(32'hbad9d912),
	.w8(32'h3bce1a68),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00604a),
	.w1(32'h3c1e7173),
	.w2(32'h3c018c57),
	.w3(32'hbba6d498),
	.w4(32'hbb26c8b3),
	.w5(32'hbb78bb43),
	.w6(32'hbbb2829f),
	.w7(32'hbc87188c),
	.w8(32'hbc335087),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd03b58),
	.w1(32'hbcaa3100),
	.w2(32'hbca3195e),
	.w3(32'hbbb2c48b),
	.w4(32'hbc61c37d),
	.w5(32'hbc8c5a52),
	.w6(32'hbc864889),
	.w7(32'hbc3c571c),
	.w8(32'hbbcb7882),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc5f82),
	.w1(32'h3a831825),
	.w2(32'h3b0456a7),
	.w3(32'hbca57506),
	.w4(32'h3be9d67f),
	.w5(32'h3baec4d7),
	.w6(32'hbc97145d),
	.w7(32'hb83711ab),
	.w8(32'h3a8abeed),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0c952),
	.w1(32'h3ae1283f),
	.w2(32'h3bd1bd2e),
	.w3(32'hbb7baa72),
	.w4(32'hbb877c2e),
	.w5(32'h3aa2fc41),
	.w6(32'hba58ef99),
	.w7(32'hbb34f885),
	.w8(32'h3ac7fd86),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb28b6),
	.w1(32'hba32e842),
	.w2(32'h3b008bea),
	.w3(32'hbb696516),
	.w4(32'hbb1f1ad5),
	.w5(32'hbb513fc0),
	.w6(32'h3b1ef132),
	.w7(32'hbb2ac439),
	.w8(32'hba36c24c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60852),
	.w1(32'h39e20da2),
	.w2(32'hb9a5a266),
	.w3(32'h3b2ea03b),
	.w4(32'h3b97b63d),
	.w5(32'h3ab6f875),
	.w6(32'h3ae845b3),
	.w7(32'hba63fec5),
	.w8(32'h3a475828),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade4821),
	.w1(32'hbbdf6bcc),
	.w2(32'hbc267484),
	.w3(32'h3c10b950),
	.w4(32'hbc7ac2c4),
	.w5(32'hbc9d2f14),
	.w6(32'h3c2b625a),
	.w7(32'hbc57b262),
	.w8(32'hbc741c5d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1418ae),
	.w1(32'hbaeb902a),
	.w2(32'hbb0a98df),
	.w3(32'hbc46868a),
	.w4(32'h3b911d2c),
	.w5(32'h3aa18440),
	.w6(32'hbc1183db),
	.w7(32'h3bf2db58),
	.w8(32'h3c019042),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad96a),
	.w1(32'hb7d84b6d),
	.w2(32'h3b832c2d),
	.w3(32'h3bbfb05b),
	.w4(32'h39a25f27),
	.w5(32'h39f76ee7),
	.w6(32'h3c1a3695),
	.w7(32'hb90cb2da),
	.w8(32'h3b1a399c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af956fe),
	.w1(32'h3b4c5295),
	.w2(32'h3b950c5a),
	.w3(32'h3bb7c225),
	.w4(32'h3bd849b1),
	.w5(32'h3bf3337d),
	.w6(32'h3b23a92a),
	.w7(32'h3c4c8322),
	.w8(32'h3bf2529a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d195),
	.w1(32'hb94b19e0),
	.w2(32'h3b9ebe7e),
	.w3(32'h3b787dcc),
	.w4(32'hbbed12c4),
	.w5(32'hbb4188e8),
	.w6(32'h3b862caa),
	.w7(32'hbb98efed),
	.w8(32'hba44a1f3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd530),
	.w1(32'h3b79729f),
	.w2(32'hbbb0cd3e),
	.w3(32'h3b43072b),
	.w4(32'hbbc6edc6),
	.w5(32'hbc39d554),
	.w6(32'hba5909fa),
	.w7(32'hbb91c570),
	.w8(32'hbb5d9243),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196a9e),
	.w1(32'h3c1f4b36),
	.w2(32'hb989dba4),
	.w3(32'hbbf614c5),
	.w4(32'hb905177f),
	.w5(32'h3a04b96f),
	.w6(32'hbb82beac),
	.w7(32'h3a233e71),
	.w8(32'hbbbba3d3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067480),
	.w1(32'hbbb2ed22),
	.w2(32'hbb503a1c),
	.w3(32'hbb1efc62),
	.w4(32'h39b89a22),
	.w5(32'hbad7d6d9),
	.w6(32'hbbcb03e5),
	.w7(32'hbb0bc924),
	.w8(32'hbb951689),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba297d6),
	.w1(32'h3abe3c32),
	.w2(32'h3a608d37),
	.w3(32'h3acb1381),
	.w4(32'h3a7469df),
	.w5(32'hbb6ae386),
	.w6(32'hbc3a2b31),
	.w7(32'hbc06cf1a),
	.w8(32'hbac423a2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e4e5),
	.w1(32'h3b9e9ae9),
	.w2(32'hbad17fd9),
	.w3(32'h3b524d06),
	.w4(32'hbaa63532),
	.w5(32'hbc02d882),
	.w6(32'hbb81842a),
	.w7(32'hbbb8d2bd),
	.w8(32'hbbdd4ab8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287346),
	.w1(32'h3b7343a1),
	.w2(32'h3c0c050e),
	.w3(32'hbc1190c5),
	.w4(32'h3c3a19b1),
	.w5(32'h3c6af6de),
	.w6(32'hbbe16158),
	.w7(32'hbb1d8338),
	.w8(32'hb930f691),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e7f7),
	.w1(32'h3b3791e5),
	.w2(32'hba8df351),
	.w3(32'h3bd86f95),
	.w4(32'hbb2b3f5f),
	.w5(32'hbbabe8bc),
	.w6(32'hbadfb20c),
	.w7(32'hbaf82743),
	.w8(32'hbc4d67ec),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d9ce),
	.w1(32'h3b4de9a9),
	.w2(32'h3af75ee5),
	.w3(32'h3aa0f624),
	.w4(32'hbaac84b1),
	.w5(32'hbb49da9c),
	.w6(32'hbb530cb7),
	.w7(32'hbbb7b5c6),
	.w8(32'hbbef198a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822683),
	.w1(32'h3b9809a9),
	.w2(32'h3b80bfea),
	.w3(32'hb9b7c1c9),
	.w4(32'h3af3358e),
	.w5(32'h3b875b95),
	.w6(32'hba829b46),
	.w7(32'h3ac431c0),
	.w8(32'h3b2aa257),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac84f31),
	.w1(32'h3bcaa531),
	.w2(32'h3b94e78c),
	.w3(32'h3b1e2947),
	.w4(32'h3b06edd9),
	.w5(32'hbb59fe7d),
	.w6(32'h3b93bc89),
	.w7(32'hba83952b),
	.w8(32'hbb95dd2b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aad04),
	.w1(32'h3bbc52cc),
	.w2(32'h3c08c041),
	.w3(32'hbb1754a2),
	.w4(32'h3acf3b8e),
	.w5(32'h3bbe10e7),
	.w6(32'h38a15081),
	.w7(32'hba8c3a99),
	.w8(32'h3ad871dd),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cdc24),
	.w1(32'hbba2dcb2),
	.w2(32'hbb5c738b),
	.w3(32'h3bc8da99),
	.w4(32'hbbd4f9b3),
	.w5(32'hbb9a4a63),
	.w6(32'h3be70d32),
	.w7(32'hbbd0dcef),
	.w8(32'hbba08f65),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6ddaf),
	.w1(32'hbbc3d43f),
	.w2(32'hbb1c78d3),
	.w3(32'hbb45a8cc),
	.w4(32'hbbbc94ab),
	.w5(32'hbb4bedaa),
	.w6(32'hbb50d9b7),
	.w7(32'hb9799402),
	.w8(32'h3b0e9114),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a25c3),
	.w1(32'hbca27077),
	.w2(32'hbc8edba4),
	.w3(32'hbad0e579),
	.w4(32'hbc8fe0c7),
	.w5(32'hbc8f6764),
	.w6(32'h3abe9e38),
	.w7(32'hbc7a1066),
	.w8(32'hbc3dbcde),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad5f57),
	.w1(32'h3b18ff3b),
	.w2(32'h3bde6a0b),
	.w3(32'hbc8a9ac6),
	.w4(32'h3a9a5778),
	.w5(32'h3bc3cdfb),
	.w6(32'hbc7d404b),
	.w7(32'hbbb29fbd),
	.w8(32'h3b760fae),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8472e0),
	.w1(32'h3b3e73ea),
	.w2(32'h39638dce),
	.w3(32'h39fe1ad0),
	.w4(32'h3b81c3cf),
	.w5(32'hba8b097a),
	.w6(32'hbab8802f),
	.w7(32'h3abcc660),
	.w8(32'h3ad77462),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4223f3),
	.w1(32'h3bcac691),
	.w2(32'h3bb3ff57),
	.w3(32'h3b609a56),
	.w4(32'hbc3efff4),
	.w5(32'hbc199ffa),
	.w6(32'h3c175a30),
	.w7(32'hbc08cba2),
	.w8(32'hbc2b96a4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba984b9),
	.w1(32'hbb3e9555),
	.w2(32'h3af4b9bf),
	.w3(32'hbb81f406),
	.w4(32'h3b18cd81),
	.w5(32'h3bbc42a4),
	.w6(32'hbbf436f7),
	.w7(32'h3a847160),
	.w8(32'h3a89d8ca),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c834613),
	.w1(32'hbb43d0f4),
	.w2(32'hbbfef7a8),
	.w3(32'h3c80aaba),
	.w4(32'hbbfd60a2),
	.w5(32'hbc0554ab),
	.w6(32'h3a920647),
	.w7(32'hbbfa799c),
	.w8(32'hbae9dfbf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc819),
	.w1(32'hbc2dc3be),
	.w2(32'hbb5eaf0e),
	.w3(32'hbbee95b7),
	.w4(32'hbc06b396),
	.w5(32'hbb6c6fda),
	.w6(32'hbb89f297),
	.w7(32'hbbb82046),
	.w8(32'hbb1abe72),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a520),
	.w1(32'h39feaf53),
	.w2(32'hbbac777d),
	.w3(32'h390014b2),
	.w4(32'h3a015994),
	.w5(32'hbbdcb848),
	.w6(32'h3af7be98),
	.w7(32'hbb28fc3b),
	.w8(32'hbb23d39b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bebb91),
	.w1(32'h3b41f109),
	.w2(32'h3b3b8a14),
	.w3(32'h3b5b9b9e),
	.w4(32'h38991137),
	.w5(32'hbb71ae16),
	.w6(32'h3b965687),
	.w7(32'hba72c923),
	.w8(32'hba5a6f42),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a099b),
	.w1(32'hbc15c7d1),
	.w2(32'hbc0e08f6),
	.w3(32'hbbceac58),
	.w4(32'hbc398c1b),
	.w5(32'hbb6da423),
	.w6(32'hbc164388),
	.w7(32'hbc63463f),
	.w8(32'hbab35454),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc872980),
	.w1(32'hbb97ad32),
	.w2(32'hbbb88149),
	.w3(32'hbbbcc3ae),
	.w4(32'hb99155c3),
	.w5(32'hbabdfb68),
	.w6(32'hbb70f979),
	.w7(32'h3a785317),
	.w8(32'h3b296c22),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a361ad0),
	.w1(32'h3ad9531e),
	.w2(32'hba52e4fc),
	.w3(32'h3be72fef),
	.w4(32'hb9a65590),
	.w5(32'hbc1e4bb5),
	.w6(32'h3c1f4c64),
	.w7(32'hbb5a8d22),
	.w8(32'hbbe9c1e3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44d299),
	.w1(32'hbb17db00),
	.w2(32'hba909d55),
	.w3(32'hbad6f420),
	.w4(32'hbc0158e7),
	.w5(32'hbab1d2ce),
	.w6(32'hbb81f8dc),
	.w7(32'hbb6c1ee2),
	.w8(32'h38fcfd51),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88cd2b),
	.w1(32'h3a8abf9b),
	.w2(32'hbc0c86bf),
	.w3(32'h3b345a02),
	.w4(32'h3ab2153f),
	.w5(32'hbbf40820),
	.w6(32'h3b5022a7),
	.w7(32'h3bb9ba1a),
	.w8(32'hba643252),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7684c),
	.w1(32'hbade5bc1),
	.w2(32'h3ba9ec23),
	.w3(32'hbb1165c9),
	.w4(32'h3a48aa20),
	.w5(32'hb919f0fd),
	.w6(32'hbb9aae0c),
	.w7(32'hbb5699d3),
	.w8(32'h3ba5b227),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9017b6a),
	.w1(32'h3b6e9750),
	.w2(32'h3bce9cdc),
	.w3(32'h3ace94d9),
	.w4(32'h3c34c134),
	.w5(32'h3c2e6a15),
	.w6(32'hbb3f4636),
	.w7(32'h3c283cbd),
	.w8(32'h3c6f5541),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b921fa1),
	.w1(32'hbbad6f0e),
	.w2(32'hbb74262e),
	.w3(32'h3c10cdb5),
	.w4(32'hbb82cb32),
	.w5(32'hba0b6f18),
	.w6(32'h3c2f6f88),
	.w7(32'hbae11963),
	.w8(32'h3b0cc817),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc998c),
	.w1(32'h3bb2129a),
	.w2(32'h3c126d2d),
	.w3(32'hbacd5f2c),
	.w4(32'h3a82a5de),
	.w5(32'h3b527ab7),
	.w6(32'hbbdd3a01),
	.w7(32'h3b57692a),
	.w8(32'h3a95ad7b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99bdb3),
	.w1(32'h3b3c5906),
	.w2(32'h3bb6afc0),
	.w3(32'h3b986439),
	.w4(32'hbb0316e6),
	.w5(32'h3b03c1b0),
	.w6(32'hba1a1132),
	.w7(32'hbad6f0fd),
	.w8(32'h3ae886ae),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb1a4),
	.w1(32'h3a9362c9),
	.w2(32'h382118bc),
	.w3(32'h3b66fdac),
	.w4(32'h37eb21a4),
	.w5(32'hbb4d764b),
	.w6(32'h386d0901),
	.w7(32'h3a224325),
	.w8(32'hbb222d23),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51cd89),
	.w1(32'hba2edb91),
	.w2(32'hbac36312),
	.w3(32'h39dfb23b),
	.w4(32'h3abd2056),
	.w5(32'hba65b202),
	.w6(32'hbb32f4f0),
	.w7(32'hbb0775cd),
	.w8(32'hbb328c5f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cd023),
	.w1(32'hbb599c03),
	.w2(32'h3a1012bb),
	.w3(32'h3ba56822),
	.w4(32'hbc116075),
	.w5(32'hbbd7471a),
	.w6(32'hbbf359b2),
	.w7(32'hbc097b5d),
	.w8(32'hbc1efc7e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5032f1),
	.w1(32'h3c05fb32),
	.w2(32'h3be9373d),
	.w3(32'hbb839415),
	.w4(32'hba7f7cb2),
	.w5(32'hbb8475cc),
	.w6(32'hbb801765),
	.w7(32'h3a9cedd0),
	.w8(32'hba189a4b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ddd0a),
	.w1(32'hbc0d3170),
	.w2(32'hbb7ae9e9),
	.w3(32'hbb76c3c1),
	.w4(32'hbbef3145),
	.w5(32'hbbc00d47),
	.w6(32'h3a8cc0cb),
	.w7(32'hbbaa93b9),
	.w8(32'hbb676737),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6865de),
	.w1(32'h3c946a6f),
	.w2(32'h3cdbd8c5),
	.w3(32'hbbfd1bde),
	.w4(32'h3c961384),
	.w5(32'h3c46f5e1),
	.w6(32'hbabdc66d),
	.w7(32'h3c9422c1),
	.w8(32'h3c516d8f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd61123),
	.w1(32'hbc4e3278),
	.w2(32'hbbf94c2b),
	.w3(32'h3cb94217),
	.w4(32'hbc163337),
	.w5(32'hbc7afe61),
	.w6(32'h3ca7f79b),
	.w7(32'hbc2e1691),
	.w8(32'hbc3fe8b3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78152d),
	.w1(32'hbc00e776),
	.w2(32'hbb9c23ad),
	.w3(32'hbc2a6e07),
	.w4(32'hb8024f11),
	.w5(32'hbab50728),
	.w6(32'hbbed0ba4),
	.w7(32'hbc46dc00),
	.w8(32'hbbc29f4c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a33f0),
	.w1(32'hbc227879),
	.w2(32'hbbad3d87),
	.w3(32'hbb361cf9),
	.w4(32'hbb5e36bd),
	.w5(32'hbbc41990),
	.w6(32'hba620e30),
	.w7(32'h393a1464),
	.w8(32'h3b18f21b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc632729),
	.w1(32'hbbf14913),
	.w2(32'hbb0fc21b),
	.w3(32'hbc062777),
	.w4(32'h39e90f91),
	.w5(32'h3baa3783),
	.w6(32'hb97bd68f),
	.w7(32'h3c1a8cc3),
	.w8(32'h3c49f880),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bc7b8),
	.w1(32'h3c673c86),
	.w2(32'h3beafff0),
	.w3(32'h3c7ce8b5),
	.w4(32'hb97b5794),
	.w5(32'hbc9e1029),
	.w6(32'h3c399d97),
	.w7(32'hba53fa47),
	.w8(32'hbbf6a7e0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3790a),
	.w1(32'h3c5d9942),
	.w2(32'h3c079dec),
	.w3(32'hba49d0e1),
	.w4(32'h3c826a7e),
	.w5(32'h3b184c8c),
	.w6(32'hba579db6),
	.w7(32'h3bfb198c),
	.w8(32'h3b8b9f02),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c063839),
	.w1(32'h3b2ac0eb),
	.w2(32'h3ac01e56),
	.w3(32'h3bf33a43),
	.w4(32'hbb1d5b8d),
	.w5(32'hbba52dac),
	.w6(32'h3c203262),
	.w7(32'hbbf51d1a),
	.w8(32'hbc35fad0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a239c),
	.w1(32'h3b5c8009),
	.w2(32'hba91e870),
	.w3(32'hbc23cc0c),
	.w4(32'hbb13cac9),
	.w5(32'hbb330892),
	.w6(32'hbc008357),
	.w7(32'hb8f95819),
	.w8(32'h3b121114),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aadc2),
	.w1(32'h396407e1),
	.w2(32'h3bd56f7c),
	.w3(32'h3ab66a17),
	.w4(32'h3a9e4779),
	.w5(32'h3c081a7d),
	.w6(32'h3bc733eb),
	.w7(32'h3af495d8),
	.w8(32'h3bbb0ef7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badcf96),
	.w1(32'hbc08065e),
	.w2(32'hbc2de29a),
	.w3(32'h3c17eac1),
	.w4(32'hbbfb00d8),
	.w5(32'hbc66a1bb),
	.w6(32'h3bc75b32),
	.w7(32'hbbfa641f),
	.w8(32'hbba40640),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af5dd),
	.w1(32'hbb787347),
	.w2(32'h3b5204f7),
	.w3(32'hbc1b63f4),
	.w4(32'h38b29427),
	.w5(32'h3b9f723b),
	.w6(32'hbbf93d4f),
	.w7(32'hbb80c4dc),
	.w8(32'h3b43f439),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfea427),
	.w1(32'h3c56366a),
	.w2(32'h3cb4b2b1),
	.w3(32'h3ba4414a),
	.w4(32'hbad372d0),
	.w5(32'hba8cc089),
	.w6(32'hbb8c2d6b),
	.w7(32'hbc3bd345),
	.w8(32'hbbcc42bb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34fcf9),
	.w1(32'hb953b3c5),
	.w2(32'h3b2bbda0),
	.w3(32'h3a288bac),
	.w4(32'hbb1cb470),
	.w5(32'hbb423855),
	.w6(32'h3b349b5d),
	.w7(32'hb9c43ad4),
	.w8(32'hbae7e7bc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55a6e4),
	.w1(32'h3b469533),
	.w2(32'h39687c06),
	.w3(32'hb911eaed),
	.w4(32'hbac98cfb),
	.w5(32'hbb6be111),
	.w6(32'h3795b114),
	.w7(32'hbb645c89),
	.w8(32'hbb6de387),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878fe7),
	.w1(32'hbba77223),
	.w2(32'hbbc6466c),
	.w3(32'hbb5bdd46),
	.w4(32'hbb59de9a),
	.w5(32'hbb15a5d0),
	.w6(32'hbba4f3f5),
	.w7(32'hbb56f840),
	.w8(32'hbb146cca),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e7290),
	.w1(32'h3a5f7eb9),
	.w2(32'h3ac12b12),
	.w3(32'h39c3b49a),
	.w4(32'h3a10657a),
	.w5(32'hbb0520ea),
	.w6(32'hbafbdfcc),
	.w7(32'h3ba6d88c),
	.w8(32'hba9b0481),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90737),
	.w1(32'hbb8b52bb),
	.w2(32'hbc1c61f3),
	.w3(32'hbbf04bef),
	.w4(32'h3b0dcb09),
	.w5(32'hbbc23e60),
	.w6(32'hbb08074c),
	.w7(32'h3bca5b37),
	.w8(32'hbb5e5c11),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07aadd),
	.w1(32'h3a4427ac),
	.w2(32'h3946ee74),
	.w3(32'hbacb4aa6),
	.w4(32'h3b211055),
	.w5(32'h397a572d),
	.w6(32'h3a85a56e),
	.w7(32'h3a9e0f3d),
	.w8(32'hb9bdff31),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a2a9d),
	.w1(32'h3aa9b7b2),
	.w2(32'h3afbdf63),
	.w3(32'hba83f06b),
	.w4(32'hba0cb464),
	.w5(32'h38a95069),
	.w6(32'hb9b26b46),
	.w7(32'h3aeb0f2f),
	.w8(32'h3b294a14),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b090e01),
	.w1(32'h3b8a49ee),
	.w2(32'h3a9f3399),
	.w3(32'h3b840d99),
	.w4(32'hba71d18e),
	.w5(32'hba4c6bb9),
	.w6(32'h3a741416),
	.w7(32'hbb296d94),
	.w8(32'hbb857085),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200e10),
	.w1(32'h3b2a29a8),
	.w2(32'hba60b9b7),
	.w3(32'h39a50393),
	.w4(32'hbb0caad0),
	.w5(32'hbbc19bde),
	.w6(32'h3a9b54b0),
	.w7(32'hbb81a140),
	.w8(32'hbbc4fda0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba38de4),
	.w1(32'hb9e3abb5),
	.w2(32'hbb21365d),
	.w3(32'hbb5ded16),
	.w4(32'hbb6acebe),
	.w5(32'hba240afc),
	.w6(32'hba633d27),
	.w7(32'hbb82c579),
	.w8(32'hbab47995),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b614381),
	.w1(32'h3b931dcb),
	.w2(32'hbb3849fd),
	.w3(32'h3b8a2f9f),
	.w4(32'hbb44c8b1),
	.w5(32'hbc02211c),
	.w6(32'h3ad9425a),
	.w7(32'hbbc77fc9),
	.w8(32'hbbca7d84),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e13c),
	.w1(32'h3a8fc814),
	.w2(32'h3ae23d46),
	.w3(32'hba9c8452),
	.w4(32'hb6a60b6b),
	.w5(32'h3a90d50c),
	.w6(32'hbb45ab8e),
	.w7(32'hb91babee),
	.w8(32'hba911b4d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939d74),
	.w1(32'h3c650246),
	.w2(32'h3c20403c),
	.w3(32'hbaff76e5),
	.w4(32'h3c00c814),
	.w5(32'h3b31f267),
	.w6(32'hbb6ac5f6),
	.w7(32'h3bcc8855),
	.w8(32'h3b956525),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cc3c7),
	.w1(32'h3990dd59),
	.w2(32'hb936c53b),
	.w3(32'h3b511324),
	.w4(32'h3902834b),
	.w5(32'hba07553b),
	.w6(32'h3bdae262),
	.w7(32'hbb03f262),
	.w8(32'h39bfa927),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905c114),
	.w1(32'hbac55907),
	.w2(32'h39643cec),
	.w3(32'hba6f23f6),
	.w4(32'hb9406317),
	.w5(32'hba06770d),
	.w6(32'hb788441c),
	.w7(32'h38e4bfd3),
	.w8(32'hbb139b52),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3389cd),
	.w1(32'h3bce849f),
	.w2(32'hba7994ed),
	.w3(32'hba2cb787),
	.w4(32'h3bb58bf4),
	.w5(32'h3bb1a9af),
	.w6(32'hbc11fa45),
	.w7(32'h3a6c4f02),
	.w8(32'hb9d79835),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4cf40),
	.w1(32'hba97f479),
	.w2(32'h3adb5f9a),
	.w3(32'hbbc59796),
	.w4(32'h3c0509f9),
	.w5(32'h3bc03f62),
	.w6(32'hbc151efe),
	.w7(32'h3b805375),
	.w8(32'h3b017ddf),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75141b),
	.w1(32'h3b91cd75),
	.w2(32'h3bdb6d69),
	.w3(32'h3b3e9138),
	.w4(32'hb8b5095d),
	.w5(32'hb994259c),
	.w6(32'h3a6b5b4c),
	.w7(32'hbc050a66),
	.w8(32'hbc081d5c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45bc87),
	.w1(32'h3a7363c6),
	.w2(32'h3bb89628),
	.w3(32'h3c08501b),
	.w4(32'h3ab93189),
	.w5(32'hbb597274),
	.w6(32'hbab8261e),
	.w7(32'h3b378cf1),
	.w8(32'h3b5aea90),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320819),
	.w1(32'h3acffff9),
	.w2(32'hbab665b0),
	.w3(32'hba39e78d),
	.w4(32'h3aaa57cc),
	.w5(32'h3a44f1a0),
	.w6(32'hbb603a19),
	.w7(32'hbacb43a2),
	.w8(32'hba35f36d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f5501),
	.w1(32'hbb47823d),
	.w2(32'hb91b085f),
	.w3(32'hba803b89),
	.w4(32'hbb235347),
	.w5(32'h3a0d94f6),
	.w6(32'hbaab1583),
	.w7(32'hbb6fe0f5),
	.w8(32'h3a643ba1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7985c5),
	.w1(32'h3b26711c),
	.w2(32'hbb95d628),
	.w3(32'hbb81ebd2),
	.w4(32'h38f25510),
	.w5(32'h3a82f825),
	.w6(32'hbc7a1111),
	.w7(32'hbba0c846),
	.w8(32'hb9a895fa),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5896),
	.w1(32'hbc40d752),
	.w2(32'hbb22a73f),
	.w3(32'hbc1bf0d0),
	.w4(32'hbb71fd48),
	.w5(32'h3baab7c8),
	.w6(32'hbbdd2bb0),
	.w7(32'hbab8dc6a),
	.w8(32'h3c310ffd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc217746),
	.w1(32'hbbd27fd3),
	.w2(32'hbade6ec1),
	.w3(32'hbc44509e),
	.w4(32'hbbc59256),
	.w5(32'h3bd165d7),
	.w6(32'hbcaf45f3),
	.w7(32'hbbca5415),
	.w8(32'h3beb9538),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e13f0),
	.w1(32'h3b80b7bf),
	.w2(32'h3b3aeac1),
	.w3(32'h3a37a3e0),
	.w4(32'h3a83b507),
	.w5(32'h3a97f521),
	.w6(32'hbacbf7ab),
	.w7(32'h3b14b00d),
	.w8(32'hb984b978),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab39696),
	.w1(32'h3bcc021d),
	.w2(32'h3b249a8b),
	.w3(32'h3bbce39a),
	.w4(32'h3b14e346),
	.w5(32'h39d764bd),
	.w6(32'h3bc9c4b2),
	.w7(32'hbb3ce7c2),
	.w8(32'hbaee45cd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4492e6),
	.w1(32'hb8596423),
	.w2(32'hba61e4db),
	.w3(32'h3b48ac49),
	.w4(32'h3a8241cd),
	.w5(32'h3b21c790),
	.w6(32'h3b70cc71),
	.w7(32'hba8a22c6),
	.w8(32'hba5c1a55),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66cc99),
	.w1(32'hbb3e9883),
	.w2(32'h3a74e6d6),
	.w3(32'h391bd5c0),
	.w4(32'hbb8770ff),
	.w5(32'hba845985),
	.w6(32'h39349c6f),
	.w7(32'hbb58f5da),
	.w8(32'hbb029931),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808ce5),
	.w1(32'h3bba2de0),
	.w2(32'h3a93fa8b),
	.w3(32'h391d64ba),
	.w4(32'h3a9876d8),
	.w5(32'hba8ddb01),
	.w6(32'hbabec5ab),
	.w7(32'h3aa09068),
	.w8(32'h3b0b5bf9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a757291),
	.w1(32'hbb3bfef2),
	.w2(32'hbb81c61b),
	.w3(32'h3ac2ed0a),
	.w4(32'hbace378e),
	.w5(32'hbb877594),
	.w6(32'h3a460cf1),
	.w7(32'hbb8fa41d),
	.w8(32'hbbdc9bae),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc1fb),
	.w1(32'h3ae10471),
	.w2(32'hbba368d6),
	.w3(32'hbc026e0e),
	.w4(32'h3b02a60d),
	.w5(32'hbba82a58),
	.w6(32'hbc3bc023),
	.w7(32'h3b343902),
	.w8(32'hba849116),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae94a8d),
	.w1(32'hbb2f57c9),
	.w2(32'hb9387ab0),
	.w3(32'hbba2a076),
	.w4(32'hba6e85ff),
	.w5(32'h3b8cc94b),
	.w6(32'hbbc24c2f),
	.w7(32'hbafb8e27),
	.w8(32'hbac71c7a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af820ee),
	.w1(32'h3b7bf8c4),
	.w2(32'hbb715e85),
	.w3(32'h3b337501),
	.w4(32'h3ad485bf),
	.w5(32'hbb18c706),
	.w6(32'hbb37a536),
	.w7(32'hbafd1112),
	.w8(32'hbbc2ad5c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf092a8),
	.w1(32'hba86e8c1),
	.w2(32'hbaead8d8),
	.w3(32'hba0f3e29),
	.w4(32'hbaba0a45),
	.w5(32'hbb43aec5),
	.w6(32'hba4b5130),
	.w7(32'hbb06b5c2),
	.w8(32'hbae2a889),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedaea4),
	.w1(32'hbc2194b8),
	.w2(32'hbbde7ebd),
	.w3(32'hbc933e9f),
	.w4(32'hbc378ad9),
	.w5(32'hbb8f9d24),
	.w6(32'hbcc6ac79),
	.w7(32'hbbab1f33),
	.w8(32'h3b42495f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5068f8),
	.w1(32'h3adaa964),
	.w2(32'hb956f12a),
	.w3(32'hbbbc64e3),
	.w4(32'hba6cfbbf),
	.w5(32'hbab86741),
	.w6(32'hbc0c1287),
	.w7(32'hba28360a),
	.w8(32'h3a69be39),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18a047),
	.w1(32'hbb38d21f),
	.w2(32'hb9997f8a),
	.w3(32'hbb822211),
	.w4(32'hb83c30e2),
	.w5(32'hba477d8b),
	.w6(32'hbb0aab46),
	.w7(32'h3a8adf74),
	.w8(32'hb9c4a34b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0333),
	.w1(32'h3a6aeea5),
	.w2(32'hba3b4a32),
	.w3(32'h395663c5),
	.w4(32'h3b30e855),
	.w5(32'h3ad14a03),
	.w6(32'hbb4917c4),
	.w7(32'h3b05539a),
	.w8(32'h3bbfd793),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d963),
	.w1(32'h3bb28f26),
	.w2(32'h3a9fa1ab),
	.w3(32'hb9527ca9),
	.w4(32'h3bb97880),
	.w5(32'h3b4dbec6),
	.w6(32'hba49f7db),
	.w7(32'h3b90b36d),
	.w8(32'h3a8d4e62),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947855),
	.w1(32'h3acfe4c2),
	.w2(32'hb98a076d),
	.w3(32'h3b7c2301),
	.w4(32'h3a4ae37a),
	.w5(32'hba84b213),
	.w6(32'h3b73d4e4),
	.w7(32'h3a3fa1e5),
	.w8(32'hbad052c0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b3cc8),
	.w1(32'hba987913),
	.w2(32'h3a3c73d5),
	.w3(32'h38c9bccb),
	.w4(32'hb9a46a92),
	.w5(32'hbb3a61ab),
	.w6(32'hbaf32d37),
	.w7(32'h3ad300c0),
	.w8(32'hba5564a4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee420f),
	.w1(32'hba02560e),
	.w2(32'h3ad30b23),
	.w3(32'hba0ebc80),
	.w4(32'hbb223cfe),
	.w5(32'h3910ffb3),
	.w6(32'hb9ac2772),
	.w7(32'h3ac5c4b7),
	.w8(32'h398c786c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7ab6e),
	.w1(32'h3b5441ae),
	.w2(32'h3acde9ec),
	.w3(32'h3af49e9b),
	.w4(32'h387ac32f),
	.w5(32'h3a821f73),
	.w6(32'h3a0670eb),
	.w7(32'hbae1a41c),
	.w8(32'hbad78cad),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba177132),
	.w1(32'h3b77fbeb),
	.w2(32'hb990da0f),
	.w3(32'h3bf3b44e),
	.w4(32'h3a2172ae),
	.w5(32'hbbfcd876),
	.w6(32'h3a87af4e),
	.w7(32'h3ad7b42f),
	.w8(32'hb9e138c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a71b2),
	.w1(32'h3aea4c0e),
	.w2(32'h38b7db8c),
	.w3(32'hba712d68),
	.w4(32'h3b93da53),
	.w5(32'hba0012f6),
	.w6(32'hbaf62274),
	.w7(32'h3b4ddc03),
	.w8(32'h3afa965b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79d518),
	.w1(32'hb90f55fe),
	.w2(32'h3b14025b),
	.w3(32'h3aa71695),
	.w4(32'hb89b7ec1),
	.w5(32'hbb0525dd),
	.w6(32'hbb5791c0),
	.w7(32'h3c018b96),
	.w8(32'h3baed2f8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6ea60),
	.w1(32'hbb45c4b5),
	.w2(32'hb98dc78e),
	.w3(32'hba7ecf85),
	.w4(32'hba5c318e),
	.w5(32'h3aaf3a88),
	.w6(32'hb95ebd6e),
	.w7(32'h3a83f5bc),
	.w8(32'h3a176817),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837101),
	.w1(32'hbae0340c),
	.w2(32'hbb01451d),
	.w3(32'hbb19a889),
	.w4(32'hbb5bd05b),
	.w5(32'hbb058e7c),
	.w6(32'hbae96826),
	.w7(32'hbb0b6c92),
	.w8(32'hba859837),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2834a),
	.w1(32'h3b23a966),
	.w2(32'h39af216e),
	.w3(32'h3b3849d2),
	.w4(32'h3b1b8e3f),
	.w5(32'h3a1931ae),
	.w6(32'h399c2ad7),
	.w7(32'h3b373ab1),
	.w8(32'hb976d114),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125606),
	.w1(32'hb9dc5dce),
	.w2(32'h3a4af498),
	.w3(32'hbaedfbc3),
	.w4(32'h3b98ac7e),
	.w5(32'h3b6e4a01),
	.w6(32'hba7e74aa),
	.w7(32'h3ba98984),
	.w8(32'h3b6e4298),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b16e6),
	.w1(32'hbb9c03ae),
	.w2(32'hbac68f06),
	.w3(32'hbb90c46c),
	.w4(32'hbbca85ce),
	.w5(32'hbb2ab6a5),
	.w6(32'hba327d33),
	.w7(32'hbb6ef2ba),
	.w8(32'hbaea4af5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b150fdb),
	.w1(32'hbae34783),
	.w2(32'hba3605bc),
	.w3(32'h3a095769),
	.w4(32'hbbbdc40c),
	.w5(32'hba92a8ea),
	.w6(32'hbac7b412),
	.w7(32'hbb2d09f8),
	.w8(32'hbb4c05f5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb49f07),
	.w1(32'h3c1620fc),
	.w2(32'h3bd253f2),
	.w3(32'hbbc76d57),
	.w4(32'h3c40a67f),
	.w5(32'h3c070ddc),
	.w6(32'hbbb73f52),
	.w7(32'h3c2df919),
	.w8(32'h3c1501b4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba945636),
	.w1(32'hbb4d55dd),
	.w2(32'hbb730f0a),
	.w3(32'h3adb176e),
	.w4(32'hbb83709c),
	.w5(32'hbb770cad),
	.w6(32'h3be2b553),
	.w7(32'hbb787813),
	.w8(32'hbb1f6d8b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68a074),
	.w1(32'h39df8c61),
	.w2(32'h3a11e4ab),
	.w3(32'hbb09ba79),
	.w4(32'hba9414f5),
	.w5(32'h3a1e4688),
	.w6(32'hba8a562a),
	.w7(32'hbab1c3c1),
	.w8(32'h3ab1921a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8509c4),
	.w1(32'h3af52c24),
	.w2(32'h3a560d07),
	.w3(32'h3af132bb),
	.w4(32'hbb09a3f0),
	.w5(32'hbb1cdb83),
	.w6(32'hba005058),
	.w7(32'hbacfeac0),
	.w8(32'h3b1832fd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2daac7),
	.w1(32'h3af4b977),
	.w2(32'h3b730627),
	.w3(32'h3ae6d48d),
	.w4(32'hb9ea53af),
	.w5(32'hba5a9d26),
	.w6(32'h3b3c4112),
	.w7(32'h3b9d83f9),
	.w8(32'h3b56b7e8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48244),
	.w1(32'hbb865b31),
	.w2(32'h3a691b40),
	.w3(32'hbb2e3155),
	.w4(32'hba661490),
	.w5(32'hbbadedfa),
	.w6(32'hbb0d85a6),
	.w7(32'h3bcad11c),
	.w8(32'h3c13a625),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dfdb4),
	.w1(32'hbb593244),
	.w2(32'hba902d92),
	.w3(32'h3a60a9f1),
	.w4(32'hbb60cec1),
	.w5(32'hb8dfcba6),
	.w6(32'h3b135f41),
	.w7(32'hbb4347a3),
	.w8(32'hba963880),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd22198),
	.w1(32'h36fa8b12),
	.w2(32'h3b847b3b),
	.w3(32'hbb0cec94),
	.w4(32'h3b8810ef),
	.w5(32'h3bd78589),
	.w6(32'hbbc28927),
	.w7(32'hbaaf2a3d),
	.w8(32'hbb964f19),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule