module upsampling2d2x2(data_in, data_out, valid_in, valid_out);
    parameter DATA_WIDTH = 32;
    parameter IMG_WIDTH = 13;
    parameter IMG_HEIGHT = 13;
endmodule