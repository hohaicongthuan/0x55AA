module layer_8_featuremap_239(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcc1c2),
	.w1(32'hbbd76747),
	.w2(32'h3b9e7d73),
	.w3(32'hbbf53f71),
	.w4(32'hbc989ec0),
	.w5(32'hbc0d0147),
	.w6(32'hbc9c969e),
	.w7(32'h3aa184c8),
	.w8(32'h3b725909),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb49125),
	.w1(32'h3be7215e),
	.w2(32'h3b0a991e),
	.w3(32'hbbc42254),
	.w4(32'h3be8ae24),
	.w5(32'h3b051bac),
	.w6(32'h3becfa7e),
	.w7(32'h3b8a153b),
	.w8(32'h3ba26bf5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06e964),
	.w1(32'hbbc6954c),
	.w2(32'hb952e102),
	.w3(32'h3ba77da1),
	.w4(32'h3a10b3d2),
	.w5(32'h3b2e4cbd),
	.w6(32'h3c54b678),
	.w7(32'h3ca5c972),
	.w8(32'h3bd936c0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd9784),
	.w1(32'h3c283e30),
	.w2(32'h3c12bb50),
	.w3(32'hba61f156),
	.w4(32'h3a29f110),
	.w5(32'h3bcd73e0),
	.w6(32'h3bd884c4),
	.w7(32'h3c59eeec),
	.w8(32'h3c13472f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03df6c),
	.w1(32'h3c11dd71),
	.w2(32'hba8551d1),
	.w3(32'h3b31d8ae),
	.w4(32'h3ba81b57),
	.w5(32'hb936aae8),
	.w6(32'h3bd3e218),
	.w7(32'h3928927a),
	.w8(32'h3a97b47d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e9679),
	.w1(32'h3c1ced30),
	.w2(32'h3c427c5d),
	.w3(32'h3b89c371),
	.w4(32'h3c8b233e),
	.w5(32'h3cb0d672),
	.w6(32'h3c4fae29),
	.w7(32'h3c506a8c),
	.w8(32'hb9a81413),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c89d4),
	.w1(32'hbb84a53a),
	.w2(32'hbbd553d7),
	.w3(32'h3c85c3bf),
	.w4(32'hbb27000a),
	.w5(32'hbb46825b),
	.w6(32'h3a84eba3),
	.w7(32'hbb8181dc),
	.w8(32'hbb255f76),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7ab98),
	.w1(32'h3ce80fb6),
	.w2(32'h3ca32bd2),
	.w3(32'h3b24d5a1),
	.w4(32'h3cdbd274),
	.w5(32'h3b95dbc4),
	.w6(32'h3c9471be),
	.w7(32'h3c932a53),
	.w8(32'h3c0b5c32),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b871f97),
	.w1(32'h3c289b81),
	.w2(32'hbc5ce833),
	.w3(32'hbc959329),
	.w4(32'h3c195291),
	.w5(32'hbc79b269),
	.w6(32'h3c17ad32),
	.w7(32'hbbbbfdd1),
	.w8(32'hbbfc8074),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1740ac),
	.w1(32'h3a36de46),
	.w2(32'h3b83e653),
	.w3(32'hbc8301f7),
	.w4(32'hbb6101d9),
	.w5(32'hbb91b33a),
	.w6(32'hbc2f8422),
	.w7(32'h3c00938f),
	.w8(32'h3ac9a0a9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90e3f4),
	.w1(32'h3bdecc99),
	.w2(32'h39b7ee95),
	.w3(32'hbc168952),
	.w4(32'hbb108449),
	.w5(32'h3b805fef),
	.w6(32'hbc0c2b63),
	.w7(32'hbc29d3a9),
	.w8(32'hbba62687),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91cdc0),
	.w1(32'hbba8eb96),
	.w2(32'hba744b75),
	.w3(32'hbc3089a8),
	.w4(32'hbc2e204f),
	.w5(32'hbc0ffb06),
	.w6(32'hbc323719),
	.w7(32'hbbe1f153),
	.w8(32'hbb9bca9e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c17e1),
	.w1(32'hbc17fe4d),
	.w2(32'hbc59c215),
	.w3(32'h3bac7a66),
	.w4(32'hbb83be3b),
	.w5(32'hbc67704d),
	.w6(32'h3bae58b0),
	.w7(32'hbadecd5f),
	.w8(32'hbb95dea6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea9d6d),
	.w1(32'h3ba3b829),
	.w2(32'h3cd42549),
	.w3(32'h3ac0427b),
	.w4(32'h3c0c9601),
	.w5(32'h3c55da26),
	.w6(32'hbaf463cf),
	.w7(32'h3ca9720d),
	.w8(32'h3c937d35),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda800c),
	.w1(32'hbc06e5b6),
	.w2(32'hbb36cb64),
	.w3(32'h3c45436f),
	.w4(32'hbc01e6b3),
	.w5(32'hbb6f452a),
	.w6(32'hbbd0f82c),
	.w7(32'hbb83d47a),
	.w8(32'hbb66bb8d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff05db),
	.w1(32'hbbf682d7),
	.w2(32'hbc4eed2c),
	.w3(32'hbb422fca),
	.w4(32'hbcb3b8c0),
	.w5(32'hbc57c947),
	.w6(32'hbb8c2edb),
	.w7(32'hbbfb9606),
	.w8(32'h3ae9ce61),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac17293),
	.w1(32'hbbed1a47),
	.w2(32'h396d5574),
	.w3(32'hbaacf42d),
	.w4(32'hbb86d2f5),
	.w5(32'h3b6ad6c8),
	.w6(32'h3aedcdfc),
	.w7(32'h3b64ab12),
	.w8(32'h3b0bf83e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4152a),
	.w1(32'hbb96ca70),
	.w2(32'h3bc791e1),
	.w3(32'hbb1175a8),
	.w4(32'hbc4d4d56),
	.w5(32'hbb585ed7),
	.w6(32'hbc2e9575),
	.w7(32'hbb4891e9),
	.w8(32'hbb0c7419),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002b6a),
	.w1(32'h3c563a29),
	.w2(32'h3cac0290),
	.w3(32'hbbb17821),
	.w4(32'hbc635f42),
	.w5(32'h3b453433),
	.w6(32'hbd21655e),
	.w7(32'hbcbac015),
	.w8(32'hbca3b415),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd2215),
	.w1(32'h3b299c44),
	.w2(32'h3bf84445),
	.w3(32'hbbec1fb1),
	.w4(32'hbbe5b613),
	.w5(32'hbc06de5c),
	.w6(32'hbc2d72df),
	.w7(32'hbc30229f),
	.w8(32'hbc00f41c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e0223),
	.w1(32'h3b8e4514),
	.w2(32'h3c6d940e),
	.w3(32'hbbb898b9),
	.w4(32'hbbbbc271),
	.w5(32'h3b83a6de),
	.w6(32'h3c9f2da3),
	.w7(32'h3c506c6e),
	.w8(32'h38a96790),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a1b4),
	.w1(32'h3c9ceaf5),
	.w2(32'h3cf78e94),
	.w3(32'h3c64ee09),
	.w4(32'h3cbf0b52),
	.w5(32'h3ca52f37),
	.w6(32'h3c4627e6),
	.w7(32'h3c8aa102),
	.w8(32'h3c5d58ee),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6af0),
	.w1(32'h3c138faf),
	.w2(32'h3cf750a0),
	.w3(32'hbc8c3ab0),
	.w4(32'hbba359ae),
	.w5(32'h3bf1d910),
	.w6(32'hbc4e63f9),
	.w7(32'h3bfa8496),
	.w8(32'hbc5c1bcf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dae67),
	.w1(32'h3c81cb1d),
	.w2(32'h3cd3b7f2),
	.w3(32'hba8a68c1),
	.w4(32'h3c8525ac),
	.w5(32'h3ca8c968),
	.w6(32'h3b3777b1),
	.w7(32'h3c219d9a),
	.w8(32'h3c62c42c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bcf6e),
	.w1(32'h3c36f91d),
	.w2(32'h3bc6a176),
	.w3(32'h39324760),
	.w4(32'h3c3b4abd),
	.w5(32'h3bf8c829),
	.w6(32'h3c0b4cbb),
	.w7(32'h3c2b04d6),
	.w8(32'hba87bbcc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b822f),
	.w1(32'h3be74381),
	.w2(32'h3cb4e0ae),
	.w3(32'hbb267fbe),
	.w4(32'h3be73561),
	.w5(32'h3a45721b),
	.w6(32'hbc1685cc),
	.w7(32'h3c874255),
	.w8(32'h3bbf14e6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92f2ad),
	.w1(32'hbb450a5e),
	.w2(32'hbc88aa16),
	.w3(32'hbc024da6),
	.w4(32'hbb8bb1be),
	.w5(32'hbc690bc2),
	.w6(32'h3bf64dcd),
	.w7(32'h3c1b7cdf),
	.w8(32'h3c4f3c27),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183be6),
	.w1(32'h3d059b20),
	.w2(32'h3e114e9c),
	.w3(32'hbcb204b4),
	.w4(32'hbb554f34),
	.w5(32'h3d91f7f5),
	.w6(32'h3b39b5e4),
	.w7(32'hbc40b392),
	.w8(32'h3c820df5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cceb997),
	.w1(32'h3c1b0c7d),
	.w2(32'h3b678266),
	.w3(32'h3c6d1ebc),
	.w4(32'hbae4b7ec),
	.w5(32'hbb4bce5a),
	.w6(32'hbba0b4cf),
	.w7(32'hbbf46e48),
	.w8(32'hbb1057b7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0e2c3),
	.w1(32'h3a8e6365),
	.w2(32'hbb535660),
	.w3(32'hbb9cd2e1),
	.w4(32'hbbc196d6),
	.w5(32'hbc3c8e59),
	.w6(32'h3a212ff8),
	.w7(32'hbaa649bf),
	.w8(32'hbc0fd122),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc811e4b),
	.w1(32'h3b530d29),
	.w2(32'h3bce2ba7),
	.w3(32'hbcbc3610),
	.w4(32'hb95ba7e5),
	.w5(32'h39dbb9b8),
	.w6(32'h3c01ccd7),
	.w7(32'h3c4e4a3e),
	.w8(32'h3c1c7b92),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b092b81),
	.w1(32'h3c26d6be),
	.w2(32'h3a6db4e1),
	.w3(32'hba426819),
	.w4(32'h3bff08c7),
	.w5(32'h3b702c03),
	.w6(32'h3c3eab6d),
	.w7(32'h39c210cc),
	.w8(32'hbc1610d7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ee4bf),
	.w1(32'hbb590be1),
	.w2(32'h3cb0f224),
	.w3(32'hbb758b6a),
	.w4(32'hbc1e2a64),
	.w5(32'h3c3ce3de),
	.w6(32'hbb8bf5db),
	.w7(32'h3be24ac3),
	.w8(32'h3c8001c2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb0515),
	.w1(32'h3cb5dafe),
	.w2(32'h3cc034e9),
	.w3(32'h3c38a5b1),
	.w4(32'h3cbf4967),
	.w5(32'h3cc2ebac),
	.w6(32'h3c09c912),
	.w7(32'h3c06d0eb),
	.w8(32'h3c221e85),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca17f5f),
	.w1(32'hbc50eaa3),
	.w2(32'hbc8cefe7),
	.w3(32'h3c9bbe55),
	.w4(32'hbc652134),
	.w5(32'hbca3ac53),
	.w6(32'hb9a46a36),
	.w7(32'hbb09493b),
	.w8(32'hbbe339f2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1f25b),
	.w1(32'h3c8639a9),
	.w2(32'h3cb6e488),
	.w3(32'hbc838dd8),
	.w4(32'hbc25c546),
	.w5(32'hbb59f154),
	.w6(32'h3c0f4165),
	.w7(32'h3c944641),
	.w8(32'h3c0966f3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9989090),
	.w1(32'h3b99197a),
	.w2(32'h3ba5d0d9),
	.w3(32'hbb003de7),
	.w4(32'hba77200a),
	.w5(32'h3a97d06e),
	.w6(32'h3b519078),
	.w7(32'h3b2ad7e1),
	.w8(32'hbad5db2a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd0e5),
	.w1(32'h3c0384bf),
	.w2(32'h3c54e419),
	.w3(32'h3ace55e2),
	.w4(32'h3bcd4a3e),
	.w5(32'h3c13ed2e),
	.w6(32'hbab938d0),
	.w7(32'h3b1df805),
	.w8(32'h3ab007b2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e10c8),
	.w1(32'hbba45c00),
	.w2(32'hbbf6ae96),
	.w3(32'h3ba6d308),
	.w4(32'hbc2fb9df),
	.w5(32'hba8bd135),
	.w6(32'h3bfbedb9),
	.w7(32'hbb6cbcc1),
	.w8(32'h3966dd5b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec8977),
	.w1(32'h3cf73237),
	.w2(32'h3d237a7f),
	.w3(32'h3c386f2b),
	.w4(32'h3cb5d862),
	.w5(32'h3ce59b4c),
	.w6(32'h3c422fbc),
	.w7(32'h3c8c883e),
	.w8(32'h3c356d97),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cecf8a5),
	.w1(32'hb98dded9),
	.w2(32'h3b0ab66f),
	.w3(32'h3c0edc25),
	.w4(32'hbca0364b),
	.w5(32'hbca005ba),
	.w6(32'hbceb6d7e),
	.w7(32'hbcf8756e),
	.w8(32'hbc9a491f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eb92f),
	.w1(32'hbb866fa0),
	.w2(32'h3b824328),
	.w3(32'hbc458611),
	.w4(32'hbc333c7d),
	.w5(32'h3b0a00a2),
	.w6(32'h3b1ab5db),
	.w7(32'h3b5b80e1),
	.w8(32'h3b67e178),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f467),
	.w1(32'hbb0dc623),
	.w2(32'h3bd09dae),
	.w3(32'hbb89df6a),
	.w4(32'h39bf1eaa),
	.w5(32'h3c4c56de),
	.w6(32'h3abd107a),
	.w7(32'h3b2252e0),
	.w8(32'h3b356d4a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f53e),
	.w1(32'hbc549867),
	.w2(32'hbc98d2fa),
	.w3(32'hbaeed2e6),
	.w4(32'hbc957166),
	.w5(32'hbc52ec27),
	.w6(32'hbc882ac7),
	.w7(32'hbc767195),
	.w8(32'hbbe86f4b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd94121),
	.w1(32'h3c8cd2e1),
	.w2(32'h3cf8e36b),
	.w3(32'hbc0b29ca),
	.w4(32'hbbbc2879),
	.w5(32'h3c385e0d),
	.w6(32'hbbcc5bed),
	.w7(32'h3c078ce5),
	.w8(32'hbb2ed0a2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd7ef0),
	.w1(32'h3c34951b),
	.w2(32'h3aa737bd),
	.w3(32'hbbc48233),
	.w4(32'h3bc38bca),
	.w5(32'h3ae6892b),
	.w6(32'h3c0f7125),
	.w7(32'h3a433bad),
	.w8(32'h3b81be5a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c24f),
	.w1(32'hbca0fd7d),
	.w2(32'hbcb88830),
	.w3(32'hbb114081),
	.w4(32'hbc8e9168),
	.w5(32'hbca207ad),
	.w6(32'hbc05d5a7),
	.w7(32'hbc71f64b),
	.w8(32'hbc35af55),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd47b92),
	.w1(32'h3d04fb77),
	.w2(32'h3d569855),
	.w3(32'hbc39089f),
	.w4(32'h3c24dd37),
	.w5(32'h3c862a49),
	.w6(32'h3b64ec12),
	.w7(32'h3c7cf240),
	.w8(32'h3b1fe2f1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c558724),
	.w1(32'h3cc43939),
	.w2(32'h3cf84fce),
	.w3(32'h3c3dbd4f),
	.w4(32'h3b0a76b0),
	.w5(32'h3bcafbb8),
	.w6(32'h3c3f1f78),
	.w7(32'h3ca19a4a),
	.w8(32'h3c245bd4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f9080),
	.w1(32'h3c4aa827),
	.w2(32'h3c9b8e85),
	.w3(32'hba88b10b),
	.w4(32'hbc1db6af),
	.w5(32'h3bb7ca85),
	.w6(32'h3bc3aab8),
	.w7(32'h3bc417d4),
	.w8(32'h3bef9520),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2056f2),
	.w1(32'h3bdcc167),
	.w2(32'h3bb9cd37),
	.w3(32'h3cd3a7a0),
	.w4(32'h3b6a52c7),
	.w5(32'hbaa8de06),
	.w6(32'h3bb355fe),
	.w7(32'hbad00279),
	.w8(32'h3aa275f0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adb153),
	.w1(32'h3ca524b5),
	.w2(32'h3c8add7a),
	.w3(32'hbbdfe6b9),
	.w4(32'h3c11f56f),
	.w5(32'h3c69a80c),
	.w6(32'hbc7759ea),
	.w7(32'hbc4846a2),
	.w8(32'hbb8c488f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e553),
	.w1(32'h3adf3ef7),
	.w2(32'hbc17fd73),
	.w3(32'hbb29c409),
	.w4(32'h3aaa279a),
	.w5(32'hbc0bfdfe),
	.w6(32'hbc2496ba),
	.w7(32'hbc540722),
	.w8(32'hbbc51518),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52ff32),
	.w1(32'hbbb7bb65),
	.w2(32'hbbda5a94),
	.w3(32'hbc10cdbf),
	.w4(32'hbc91a361),
	.w5(32'hbc79b3a5),
	.w6(32'hbc85811e),
	.w7(32'hbcb0640c),
	.w8(32'hbc2b4456),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d60e),
	.w1(32'h3b2877fd),
	.w2(32'h3c82e9f1),
	.w3(32'hbbf2795f),
	.w4(32'h3bccfd1b),
	.w5(32'h3c181ae5),
	.w6(32'hbb18c5ed),
	.w7(32'h3c072e73),
	.w8(32'h3cb44d79),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3f371),
	.w1(32'h3bc861f5),
	.w2(32'h3d1d4bb7),
	.w3(32'h3cdb2e2f),
	.w4(32'hbc4f0f65),
	.w5(32'h3b1c66e9),
	.w6(32'hbbf5d0a8),
	.w7(32'hbb145862),
	.w8(32'h3b4c6934),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e75ea),
	.w1(32'hbbd76b12),
	.w2(32'h3bfba978),
	.w3(32'hb992afee),
	.w4(32'hbba76c1a),
	.w5(32'h3aa4edde),
	.w6(32'h3b8d4c04),
	.w7(32'h3bcc4602),
	.w8(32'h3c58dbe7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e1688),
	.w1(32'h3c3e12af),
	.w2(32'h3c25dfe5),
	.w3(32'h3c6d94fd),
	.w4(32'h3a10291c),
	.w5(32'h3c2bbaa7),
	.w6(32'h3b8b9672),
	.w7(32'hba12447d),
	.w8(32'h3bbbc2c9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445634),
	.w1(32'hbbabd44e),
	.w2(32'h3af1b022),
	.w3(32'h3aab689b),
	.w4(32'h39d4351d),
	.w5(32'h3aea63be),
	.w6(32'h39f87e19),
	.w7(32'hbae69972),
	.w8(32'h3b18a6a9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137ce0),
	.w1(32'h3c985346),
	.w2(32'h3cc420ee),
	.w3(32'h3b09b481),
	.w4(32'h3cabd65a),
	.w5(32'h3c655149),
	.w6(32'h3bf8dbb8),
	.w7(32'h3c5bfc77),
	.w8(32'h3be0129e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c62a7),
	.w1(32'hbb41065e),
	.w2(32'hbc2beebe),
	.w3(32'h3be677ba),
	.w4(32'h3c43dda9),
	.w5(32'h3a283161),
	.w6(32'hba939b0b),
	.w7(32'hbc112eaa),
	.w8(32'hb9ff61a7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dc2a0),
	.w1(32'h3ae2127f),
	.w2(32'hba0b67a5),
	.w3(32'hb9eceff9),
	.w4(32'hbb65851e),
	.w5(32'hbbdbdde6),
	.w6(32'h3b0f7891),
	.w7(32'h3b1aed6b),
	.w8(32'hbac69f08),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b185cca),
	.w1(32'h3d145baf),
	.w2(32'h3cac263d),
	.w3(32'hbc435aeb),
	.w4(32'h3c873459),
	.w5(32'h3b9e1104),
	.w6(32'hbb6caf3e),
	.w7(32'hbc306e50),
	.w8(32'hbc82b06e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc504d0c),
	.w1(32'hbc39b758),
	.w2(32'hbbf66201),
	.w3(32'hbb5adfff),
	.w4(32'hbb3903fb),
	.w5(32'hbb0fcc40),
	.w6(32'hbc03a68b),
	.w7(32'hba57b40f),
	.w8(32'h3ba88bf2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e449d),
	.w1(32'hbbf17a77),
	.w2(32'hbbd12ab3),
	.w3(32'hbb0e0b61),
	.w4(32'hbb5fe039),
	.w5(32'hbba1a857),
	.w6(32'hbbca2167),
	.w7(32'hbc07f3fe),
	.w8(32'hbc09c7bc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9d695),
	.w1(32'h3cd7e514),
	.w2(32'h3d321ca7),
	.w3(32'hbbb76fc1),
	.w4(32'h3cbc0eac),
	.w5(32'h3cec3e5b),
	.w6(32'h3b37c785),
	.w7(32'h3c3af067),
	.w8(32'h3c2418dd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd95d9d),
	.w1(32'h3c1da2aa),
	.w2(32'h38dcdb89),
	.w3(32'h3c70c47e),
	.w4(32'h3bf5b8a3),
	.w5(32'h3c2c769e),
	.w6(32'h3ca6d151),
	.w7(32'h3c0cf42d),
	.w8(32'hbb852136),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55357d),
	.w1(32'hbb285635),
	.w2(32'hbb820b85),
	.w3(32'h3c2c8001),
	.w4(32'hba9944d1),
	.w5(32'h3bbeabfa),
	.w6(32'h3b4a633a),
	.w7(32'h3b6bcae8),
	.w8(32'h3bd7660d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb696eb4),
	.w1(32'h3ab548f4),
	.w2(32'h3c7d5399),
	.w3(32'hbb455e36),
	.w4(32'hbb5b8f4e),
	.w5(32'h3c834687),
	.w6(32'hbb0cd98d),
	.w7(32'h3b98b9fd),
	.w8(32'hbb8e0734),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82fd51),
	.w1(32'h3b8050fa),
	.w2(32'h3c89d3ea),
	.w3(32'h3bf33529),
	.w4(32'hbaa394d5),
	.w5(32'h3c273ca3),
	.w6(32'h3b2861a8),
	.w7(32'h3b8d8208),
	.w8(32'hbc44bd2c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b229a31),
	.w1(32'h3bdbbf06),
	.w2(32'hbb1bb215),
	.w3(32'hbac52ce8),
	.w4(32'h3c2120ce),
	.w5(32'h3af01036),
	.w6(32'h3b66ab90),
	.w7(32'hbbbcf65c),
	.w8(32'hbb6a5daf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989d7d),
	.w1(32'h3b889d01),
	.w2(32'h3c43d24e),
	.w3(32'hbbdabce7),
	.w4(32'h3bd4df4c),
	.w5(32'h3c12ea6b),
	.w6(32'h3c0a6bc2),
	.w7(32'h3cafa8c4),
	.w8(32'h3c8970d1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92c8de),
	.w1(32'h3c814f45),
	.w2(32'h3c4a3855),
	.w3(32'h3c56d609),
	.w4(32'h3ae1e927),
	.w5(32'h3b94a05b),
	.w6(32'h3cc5ff82),
	.w7(32'h3ce5131c),
	.w8(32'h3caffa2e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb70df7),
	.w1(32'h3ba14228),
	.w2(32'h3bc654ff),
	.w3(32'h3c739865),
	.w4(32'hbad88b94),
	.w5(32'hbc243ff7),
	.w6(32'hbbc36301),
	.w7(32'hbb3034bc),
	.w8(32'hbb0ef58d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518e1a),
	.w1(32'h3c1c958b),
	.w2(32'h3c05c1f1),
	.w3(32'hbbb9b320),
	.w4(32'h3baf39f0),
	.w5(32'h3bfa2133),
	.w6(32'h3c3cb338),
	.w7(32'h3be3ae7f),
	.w8(32'h3bf00b92),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5adec5),
	.w1(32'h3ca969c0),
	.w2(32'h3d13f86a),
	.w3(32'h3b4c4ffd),
	.w4(32'hbb167748),
	.w5(32'h3cad010f),
	.w6(32'h3b2177fa),
	.w7(32'h3be809e7),
	.w8(32'h3c99be17),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd014f4),
	.w1(32'h3b966297),
	.w2(32'h3c4c0962),
	.w3(32'h3c654a0c),
	.w4(32'h3b342bc8),
	.w5(32'h3b885582),
	.w6(32'h3c1edf7c),
	.w7(32'h3c3fcfab),
	.w8(32'h3c2eb39a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0156dc),
	.w1(32'hba62dbd3),
	.w2(32'h3c4e51bd),
	.w3(32'hbb98b72a),
	.w4(32'hbc54ca21),
	.w5(32'h3abb3e01),
	.w6(32'hbc839dee),
	.w7(32'hbbed2e5c),
	.w8(32'hbaa7e1a0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88be97),
	.w1(32'h3c018eab),
	.w2(32'h3cfb61b5),
	.w3(32'h3bdf4bd0),
	.w4(32'h3b9f8c32),
	.w5(32'h3c94270a),
	.w6(32'h3acd1e47),
	.w7(32'h3c01c2c5),
	.w8(32'h3c18dae4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf708a3),
	.w1(32'hbba7e759),
	.w2(32'h3bf1835f),
	.w3(32'h3a0d1c5d),
	.w4(32'hbb6b3070),
	.w5(32'h3c3a0cad),
	.w6(32'hbbfa5460),
	.w7(32'h3a97a283),
	.w8(32'h3be24545),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1b3e5),
	.w1(32'hbbad217f),
	.w2(32'h3bd29302),
	.w3(32'h3bd37121),
	.w4(32'hbc7261cd),
	.w5(32'hbc0f693b),
	.w6(32'h3c4b5b20),
	.w7(32'h3c658514),
	.w8(32'h3c13a049),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac3ff2),
	.w1(32'h3b4ac1d5),
	.w2(32'h3cccb044),
	.w3(32'hbc1b064f),
	.w4(32'hbb01c042),
	.w5(32'h3c685f1c),
	.w6(32'h3beb6d11),
	.w7(32'h3c43c6a2),
	.w8(32'h3c5ba11b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7db0e0),
	.w1(32'hbbb671fc),
	.w2(32'h3cc21d9a),
	.w3(32'h3a38e09b),
	.w4(32'hbc70e59d),
	.w5(32'h3c35d0ca),
	.w6(32'hbc802e08),
	.w7(32'hbc03522b),
	.w8(32'hbbe715cc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e0f95),
	.w1(32'h3cb6cf97),
	.w2(32'h3bf1cf6b),
	.w3(32'h3b5a8514),
	.w4(32'h3aed8f8c),
	.w5(32'h3c2b1c4a),
	.w6(32'hbc5664cd),
	.w7(32'hbc98e268),
	.w8(32'hbc684b56),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46294e),
	.w1(32'h3c985b1f),
	.w2(32'h3d14ffec),
	.w3(32'hba3fb092),
	.w4(32'hbbe7cb97),
	.w5(32'h3c73a693),
	.w6(32'hbcdd271c),
	.w7(32'hbc59e973),
	.w8(32'hbc5ba48d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c835f7c),
	.w1(32'h3b26532b),
	.w2(32'h3ba5c5c6),
	.w3(32'hb98b29ae),
	.w4(32'hbb3c7bcc),
	.w5(32'h3a0b892a),
	.w6(32'h391e36a3),
	.w7(32'h3bb91030),
	.w8(32'h3bebee04),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4044f),
	.w1(32'hbb83ffa0),
	.w2(32'hbb22d1fe),
	.w3(32'h3a7a3a3a),
	.w4(32'h3a9b4dcc),
	.w5(32'h3b67dea5),
	.w6(32'hbba740ef),
	.w7(32'hbb870f10),
	.w8(32'hbc208069),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf728b),
	.w1(32'h39b69e90),
	.w2(32'hbb59f52d),
	.w3(32'hba401535),
	.w4(32'h3b803eba),
	.w5(32'h3b0d8643),
	.w6(32'hbbf10833),
	.w7(32'hbc85506c),
	.w8(32'hbc960b82),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc219aa6),
	.w1(32'h3aedaebd),
	.w2(32'h3b49ecd9),
	.w3(32'hbb51f955),
	.w4(32'h3b2382ea),
	.w5(32'h3b6090e7),
	.w6(32'hbb045595),
	.w7(32'hba64abfa),
	.w8(32'hbaf33d93),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c641),
	.w1(32'h3c56a879),
	.w2(32'h3c4693fa),
	.w3(32'h3b18e1ec),
	.w4(32'h3b18c985),
	.w5(32'hb9c61bb9),
	.w6(32'h3ba2099f),
	.w7(32'h3c343e17),
	.w8(32'hbbf95b53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b875e),
	.w1(32'h3bb11957),
	.w2(32'h3c3845f0),
	.w3(32'h3aef1beb),
	.w4(32'hbb41754f),
	.w5(32'h3b95ab11),
	.w6(32'h3c863033),
	.w7(32'h3ce8f77e),
	.w8(32'h3cdc19e0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c558d4c),
	.w1(32'h3c7309a6),
	.w2(32'h3cb94e37),
	.w3(32'h3c54b522),
	.w4(32'h3c8ee723),
	.w5(32'h3cf50ef3),
	.w6(32'h3c1e5495),
	.w7(32'h3c2f585c),
	.w8(32'h3c41b7f7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb54a4),
	.w1(32'h392f8f69),
	.w2(32'hbc4e7281),
	.w3(32'h3cd795d1),
	.w4(32'hbac5835e),
	.w5(32'hbc1c64cd),
	.w6(32'h3bfb9043),
	.w7(32'h3aabe907),
	.w8(32'hbad7230c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf78e7d),
	.w1(32'hbaa26448),
	.w2(32'hbb192397),
	.w3(32'hbc07db00),
	.w4(32'hbb63413f),
	.w5(32'hbb4dbd90),
	.w6(32'hbbb6d965),
	.w7(32'hbbf5617e),
	.w8(32'hbb5158fc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f705),
	.w1(32'hbbb0f626),
	.w2(32'hbca1f811),
	.w3(32'h3a1d3934),
	.w4(32'hbbddccad),
	.w5(32'hbc6d5561),
	.w6(32'hbc05b760),
	.w7(32'h3a91898e),
	.w8(32'h3be70d82),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952af8a),
	.w1(32'h3b086ab8),
	.w2(32'h3c0dc082),
	.w3(32'hbbe5ab66),
	.w4(32'hba614d5d),
	.w5(32'h3bf49fc2),
	.w6(32'hbbc044dc),
	.w7(32'h3a8b4c06),
	.w8(32'h3c19a11c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09a98d),
	.w1(32'h3cab00d0),
	.w2(32'h3d0861fd),
	.w3(32'hbae105b5),
	.w4(32'h3bdfb166),
	.w5(32'h3cac2448),
	.w6(32'hbb7ea3eb),
	.w7(32'h3ba054a5),
	.w8(32'h3b895c0c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd63ffe),
	.w1(32'hba89e205),
	.w2(32'h3c25187c),
	.w3(32'h3c8f7183),
	.w4(32'hbbfab8e1),
	.w5(32'hbb931549),
	.w6(32'h3bdfe14f),
	.w7(32'hbb9c2e9e),
	.w8(32'h3b351e0f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99888d),
	.w1(32'hbc645d85),
	.w2(32'hbc7fe476),
	.w3(32'h3c24f919),
	.w4(32'hbcae09c2),
	.w5(32'hbc793588),
	.w6(32'h3b8de0d8),
	.w7(32'hbbe13aa5),
	.w8(32'h3b3fe3fa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37544d),
	.w1(32'h3b8243d9),
	.w2(32'h3c300bb8),
	.w3(32'h3ba60316),
	.w4(32'h3ba89acd),
	.w5(32'h3c75c6fc),
	.w6(32'h3b0541fd),
	.w7(32'h3beb9106),
	.w8(32'h3c0d7c87),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65d9bb),
	.w1(32'h3c1b4f8a),
	.w2(32'h3c0be5cd),
	.w3(32'h3c81441b),
	.w4(32'h3b6bd1e7),
	.w5(32'h3c8d1856),
	.w6(32'h3b8d12d5),
	.w7(32'h39bbebaa),
	.w8(32'hba0b1f0b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcab22),
	.w1(32'h3b0e3964),
	.w2(32'hbcdce778),
	.w3(32'h3c43d939),
	.w4(32'h3c01929f),
	.w5(32'hbb92e2ea),
	.w6(32'h3953c6d8),
	.w7(32'hbc5a186a),
	.w8(32'hbc8c33ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc53c13),
	.w1(32'h3c044f82),
	.w2(32'h3cac4e33),
	.w3(32'hbc3ec9fe),
	.w4(32'h3beb70b5),
	.w5(32'h3c7a4412),
	.w6(32'hbab4a2f3),
	.w7(32'h3bf8eaab),
	.w8(32'h3bc3a7f9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf6741e),
	.w1(32'h3c2785f3),
	.w2(32'h3ba9beaa),
	.w3(32'h3c511c2c),
	.w4(32'h3bd08fa0),
	.w5(32'hba8ee0ff),
	.w6(32'h3c829799),
	.w7(32'h3c233c26),
	.w8(32'hbb070c5f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0900c),
	.w1(32'hbd0db4d4),
	.w2(32'hbd07aaf1),
	.w3(32'hbb20d181),
	.w4(32'hbcca895c),
	.w5(32'hbc9ab763),
	.w6(32'hbca04bd1),
	.w7(32'hbc7e5123),
	.w8(32'h396514b4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5e6bb),
	.w1(32'h3ae3224a),
	.w2(32'hbb873e1c),
	.w3(32'hbbdf982a),
	.w4(32'hbb9dc903),
	.w5(32'hbbbb4599),
	.w6(32'h3a25a649),
	.w7(32'hbc201f68),
	.w8(32'hba80ba9a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be589c3),
	.w1(32'h3bcfe9c1),
	.w2(32'hba6b245b),
	.w3(32'h3b126e03),
	.w4(32'h3bdc55f6),
	.w5(32'hba8f39f9),
	.w6(32'hbbb599d8),
	.w7(32'hbbcaa31a),
	.w8(32'hbbe5eef8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82288b),
	.w1(32'hba079158),
	.w2(32'h3c00d1c5),
	.w3(32'h39c74ba3),
	.w4(32'hbbbb33ba),
	.w5(32'h3bed74ae),
	.w6(32'h3c3664cc),
	.w7(32'h3c5d5479),
	.w8(32'h3c33f78e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b832d),
	.w1(32'hbbc5fbd8),
	.w2(32'hbccb0b12),
	.w3(32'h3be70807),
	.w4(32'h3bc42059),
	.w5(32'hbc36e32d),
	.w6(32'h3b3a88a9),
	.w7(32'hbb8dbc24),
	.w8(32'hbc26073a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5046a),
	.w1(32'h3c0c4ed2),
	.w2(32'h3b070288),
	.w3(32'hbc6e0eea),
	.w4(32'h3be0eb67),
	.w5(32'h3a51521d),
	.w6(32'h3abde35a),
	.w7(32'hba7f1fb9),
	.w8(32'hba293f10),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ca42),
	.w1(32'h3b9e3737),
	.w2(32'h3cb2a0e5),
	.w3(32'h3b9620bc),
	.w4(32'h3c55c96d),
	.w5(32'h3c9e0f05),
	.w6(32'h3a06de68),
	.w7(32'h3c58bfa1),
	.w8(32'h3c475db8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee705a),
	.w1(32'hbb49de7d),
	.w2(32'hbc0e10e2),
	.w3(32'h3c7844a7),
	.w4(32'hbb4faaae),
	.w5(32'hbc02593d),
	.w6(32'h3a559c88),
	.w7(32'hbbe3ab60),
	.w8(32'hbb112004),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc640916),
	.w1(32'h3ca70bb6),
	.w2(32'h3ce5396c),
	.w3(32'hbc1315a4),
	.w4(32'h3c9880ff),
	.w5(32'h3ca412e6),
	.w6(32'h3cb3f32e),
	.w7(32'h3cd3c6bc),
	.w8(32'h3c9a8f70),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb581d7),
	.w1(32'hbc1401d1),
	.w2(32'hbcc7ae50),
	.w3(32'h3c8ac028),
	.w4(32'h39691e7a),
	.w5(32'hbc2fbf75),
	.w6(32'h3bfad62b),
	.w7(32'h3b6c13bc),
	.w8(32'hbc494d3a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbd0a2),
	.w1(32'h3c0cdddc),
	.w2(32'h3c0c3413),
	.w3(32'hbc092a5c),
	.w4(32'h3bb06b1f),
	.w5(32'h3bc7eb53),
	.w6(32'h3bc92338),
	.w7(32'h3be7750c),
	.w8(32'h3b1f4416),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7e1a6),
	.w1(32'h3a8c2f39),
	.w2(32'hba956245),
	.w3(32'hbaa3765e),
	.w4(32'h3aa6c06b),
	.w5(32'hbae1db57),
	.w6(32'hbb8debea),
	.w7(32'hbbdea83a),
	.w8(32'hbb948197),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0169cc),
	.w1(32'hbbd5faf3),
	.w2(32'hbc4b5370),
	.w3(32'hba25e9b3),
	.w4(32'hbc2153cc),
	.w5(32'hbc00bab6),
	.w6(32'hbc2f29dc),
	.w7(32'hbc81c850),
	.w8(32'hbc57d31e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94a765),
	.w1(32'h3c6da26c),
	.w2(32'h3cdb8e20),
	.w3(32'hbc88b25c),
	.w4(32'h3c3566e5),
	.w5(32'h3cade4cd),
	.w6(32'h3b3a6fc2),
	.w7(32'h3c62fb24),
	.w8(32'h3c1592fe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c409239),
	.w1(32'h3c29800a),
	.w2(32'h3cd5faf5),
	.w3(32'h3c2b19d1),
	.w4(32'h3a486aaf),
	.w5(32'h3c18e44c),
	.w6(32'h3c114337),
	.w7(32'h3c74f55e),
	.w8(32'h3c1fdee6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98d40e),
	.w1(32'h3b4a52c1),
	.w2(32'h3bf44057),
	.w3(32'h3bb2654f),
	.w4(32'hba05d6e1),
	.w5(32'h3af29dfd),
	.w6(32'h3b495f19),
	.w7(32'h3b2d347f),
	.w8(32'hbaf34420),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50deab),
	.w1(32'h3bb75b7c),
	.w2(32'h3c8caf92),
	.w3(32'hbad98edc),
	.w4(32'hbb9bf227),
	.w5(32'h3c4f561a),
	.w6(32'h3ba8cb0c),
	.w7(32'h3c063759),
	.w8(32'h3c0eb566),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c029943),
	.w1(32'h3b0baf8a),
	.w2(32'h3bc534ee),
	.w3(32'h3bdf52f7),
	.w4(32'hbc227125),
	.w5(32'h3bc83179),
	.w6(32'hbc1bc5aa),
	.w7(32'hbbb35057),
	.w8(32'h3b62d7bf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0c24),
	.w1(32'hbb0c1a32),
	.w2(32'hbc4449ce),
	.w3(32'h3a967a52),
	.w4(32'h3b03124c),
	.w5(32'hbbbebf85),
	.w6(32'h3b78d04f),
	.w7(32'hbac8ba36),
	.w8(32'h3ade66e6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc345009),
	.w1(32'h3ca04e07),
	.w2(32'h3cce39f6),
	.w3(32'hbb5efe8f),
	.w4(32'h3c6b71a7),
	.w5(32'h3c73ee37),
	.w6(32'h3c5595aa),
	.w7(32'h3c92143a),
	.w8(32'h3c32dabe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca32dcb),
	.w1(32'hb9faad9f),
	.w2(32'h3b79ea2c),
	.w3(32'h3c038add),
	.w4(32'h3c5101da),
	.w5(32'h3c4744b3),
	.w6(32'hbbf40817),
	.w7(32'h38589e52),
	.w8(32'hba438d3c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c180370),
	.w1(32'h3ce50577),
	.w2(32'h3d0bf48d),
	.w3(32'h3c1e13d1),
	.w4(32'h3c9ba6a8),
	.w5(32'h3c9a309c),
	.w6(32'h3c4edb81),
	.w7(32'h3c40b640),
	.w8(32'h3b2b6845),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca52349),
	.w1(32'h3b3e7aa7),
	.w2(32'h3c2806be),
	.w3(32'h3bd98532),
	.w4(32'h3a90d594),
	.w5(32'h3b2f8360),
	.w6(32'hb927a2cd),
	.w7(32'h3ac30c51),
	.w8(32'h3a89eb95),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fe053),
	.w1(32'hbc04a4b2),
	.w2(32'hba2f2fe5),
	.w3(32'h39b71d13),
	.w4(32'hbc1781fc),
	.w5(32'h3b7b9331),
	.w6(32'hbaacdd2f),
	.w7(32'h3b64151e),
	.w8(32'h3ba9c3dd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule