module layer_10_featuremap_472(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33cbff4d),
	.w1(32'hb317b577),
	.w2(32'hb494ff4e),
	.w3(32'h330e5cb1),
	.w4(32'h34ab884d),
	.w5(32'h343af5d5),
	.w6(32'h33ab9a33),
	.w7(32'h341feb24),
	.w8(32'h349c6a2b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900c78a),
	.w1(32'h38b584d8),
	.w2(32'h385276c5),
	.w3(32'hb95cd509),
	.w4(32'h38111284),
	.w5(32'h38baaa13),
	.w6(32'hb9e53f54),
	.w7(32'hb98c913b),
	.w8(32'hb87685bd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4376f6c),
	.w1(32'hb42009c8),
	.w2(32'hb408eae0),
	.w3(32'hb383a6d9),
	.w4(32'h341b90f4),
	.w5(32'hb47bee40),
	.w6(32'h3446da72),
	.w7(32'hb5400e69),
	.w8(32'hb469098e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca0c9d),
	.w1(32'h39176cf3),
	.w2(32'hb4e5fee6),
	.w3(32'h378880b9),
	.w4(32'h36268aec),
	.w5(32'h35e5620e),
	.w6(32'h3754b8da),
	.w7(32'hb8836cdb),
	.w8(32'hb7ad6533),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f4683),
	.w1(32'hb626f436),
	.w2(32'hb59855f6),
	.w3(32'hb5b1eeb9),
	.w4(32'h35502702),
	.w5(32'hb49afc47),
	.w6(32'h35293cee),
	.w7(32'h360038f8),
	.w8(32'h346e5ab0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34bcf29b),
	.w1(32'h3508ce6b),
	.w2(32'h341f1774),
	.w3(32'h33dc9d93),
	.w4(32'h33ef7c24),
	.w5(32'h3416f243),
	.w6(32'h3495fc47),
	.w7(32'h34bb8231),
	.w8(32'hb404dfd7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1e002),
	.w1(32'hb93eab98),
	.w2(32'hbac49ce4),
	.w3(32'h39b82c72),
	.w4(32'hbaa22010),
	.w5(32'hba9c0577),
	.w6(32'hb8eeb835),
	.w7(32'hba5a1a4d),
	.w8(32'hb9edebf9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef58a1),
	.w1(32'h3a4aa57f),
	.w2(32'h3aaeafda),
	.w3(32'hb935d481),
	.w4(32'h3a660a68),
	.w5(32'hb8d8d144),
	.w6(32'hba6f2c8d),
	.w7(32'hba356c5a),
	.w8(32'hb925cae0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb52b967f),
	.w1(32'h366019c4),
	.w2(32'h355b12f1),
	.w3(32'hb3ba5ad6),
	.w4(32'h3681716e),
	.w5(32'hb5f6da67),
	.w6(32'h33822fe7),
	.w7(32'h3624e56e),
	.w8(32'hb6a9dd2c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02c3d9),
	.w1(32'h3902626f),
	.w2(32'h39517457),
	.w3(32'hb7eb49cf),
	.w4(32'hb9a4912c),
	.w5(32'hb923f9c0),
	.w6(32'hb9097328),
	.w7(32'hb92ca8b2),
	.w8(32'h38ca4d7c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b77a74),
	.w1(32'hb6b01d56),
	.w2(32'hb6a809e7),
	.w3(32'hb6ce0622),
	.w4(32'hb6f95442),
	.w5(32'hb629cabd),
	.w6(32'hb5cccf6c),
	.w7(32'hb6d9280f),
	.w8(32'hb687a720),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbebf2),
	.w1(32'h3a10d241),
	.w2(32'hba338b91),
	.w3(32'h3a0308fb),
	.w4(32'hba7af341),
	.w5(32'hba845df0),
	.w6(32'h37ab75ef),
	.w7(32'hbacbdb4d),
	.w8(32'hba0b9be3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989af2f),
	.w1(32'hb94ac47a),
	.w2(32'h3784b470),
	.w3(32'hb81179ef),
	.w4(32'hb9d555d2),
	.w5(32'hb94e9394),
	.w6(32'hb74ef756),
	.w7(32'hb8622c7b),
	.w8(32'h39b73049),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e0f78),
	.w1(32'hba7cf506),
	.w2(32'hb9921ffb),
	.w3(32'hba0f64f8),
	.w4(32'hba0756c5),
	.w5(32'h376cd35c),
	.w6(32'hb8af5b38),
	.w7(32'hb92d918c),
	.w8(32'h399e6b2d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ab3e29),
	.w1(32'h387b8fb8),
	.w2(32'h37be9f7b),
	.w3(32'hb856ad6a),
	.w4(32'hb72830b5),
	.w5(32'h38179319),
	.w6(32'hb931c9e8),
	.w7(32'hb92d1626),
	.w8(32'hb8c76f3a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d0b61),
	.w1(32'hb9607db6),
	.w2(32'h3a34cf07),
	.w3(32'hba3200e7),
	.w4(32'h39e4287e),
	.w5(32'h3a4aafd5),
	.w6(32'hba6d7ba6),
	.w7(32'h39eba2ed),
	.w8(32'h3a7559c3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3659e1d3),
	.w1(32'h377cb287),
	.w2(32'h36c1af2e),
	.w3(32'h3630455b),
	.w4(32'h37275a89),
	.w5(32'h36e18228),
	.w6(32'h37a11b59),
	.w7(32'h3673c827),
	.w8(32'h35c63533),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899ff6b),
	.w1(32'hb9927b08),
	.w2(32'h38cb1aa0),
	.w3(32'hb971d744),
	.w4(32'hb994fab2),
	.w5(32'h39a383d1),
	.w6(32'hba0ebab8),
	.w7(32'hb796d7a2),
	.w8(32'h3a793613),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b071ec),
	.w1(32'hb8b8124c),
	.w2(32'hb8a209a8),
	.w3(32'h38965b11),
	.w4(32'hb8f831a4),
	.w5(32'h3775ee46),
	.w6(32'hb78dec86),
	.w7(32'h380cc4ef),
	.w8(32'h39b6b3bb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3641b6c1),
	.w1(32'hb71719af),
	.w2(32'hb57d173f),
	.w3(32'h36b8f8cc),
	.w4(32'hb6910004),
	.w5(32'hb6b67d4e),
	.w6(32'h36177a4a),
	.w7(32'hb6fbc68c),
	.w8(32'hb6a63fef),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3654027e),
	.w1(32'h34ba63a6),
	.w2(32'hb6450d36),
	.w3(32'hb61453f2),
	.w4(32'hb68b8c05),
	.w5(32'h35ba47f3),
	.w6(32'h364c932a),
	.w7(32'hb5cf7027),
	.w8(32'h369a1bfc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d8f5d5),
	.w1(32'h38ff0c80),
	.w2(32'h38bb4ecc),
	.w3(32'hb8131c56),
	.w4(32'h38944946),
	.w5(32'h389101fa),
	.w6(32'hb8e4772e),
	.w7(32'hb857cf7a),
	.w8(32'hb8065cff),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a626a0f),
	.w1(32'hb9e95172),
	.w2(32'hb9cd4900),
	.w3(32'h39d25487),
	.w4(32'hba5cd609),
	.w5(32'h39f4592c),
	.w6(32'hba8a71f3),
	.w7(32'hba365700),
	.w8(32'h3918778a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0aa8d),
	.w1(32'h383a6966),
	.w2(32'hb7ed683d),
	.w3(32'h392a0302),
	.w4(32'h3843860e),
	.w5(32'hb792fc79),
	.w6(32'h38c7403e),
	.w7(32'h37911b44),
	.w8(32'hb7c74fc1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9149857),
	.w1(32'h3896d1a3),
	.w2(32'h39067c26),
	.w3(32'hb989c2c3),
	.w4(32'h399dda51),
	.w5(32'h388ec9e8),
	.w6(32'hba0bc757),
	.w7(32'hb9de6483),
	.w8(32'hb9dd3b57),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376bb28b),
	.w1(32'h378470ab),
	.w2(32'h361b84fd),
	.w3(32'h38000554),
	.w4(32'h3798fca6),
	.w5(32'h36a963cb),
	.w6(32'h37f08549),
	.w7(32'h375cca4f),
	.w8(32'h366c753b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b21fb9),
	.w1(32'h3669b020),
	.w2(32'h36893131),
	.w3(32'h366e677b),
	.w4(32'h371be412),
	.w5(32'h3635a1d1),
	.w6(32'h34bd4f90),
	.w7(32'h367ee9e0),
	.w8(32'hb58b1be6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c568c),
	.w1(32'h3ad53d14),
	.w2(32'h398a1bc5),
	.w3(32'hba878c65),
	.w4(32'h3aa03634),
	.w5(32'hba161bff),
	.w6(32'hbb017438),
	.w7(32'h3a3937a1),
	.w8(32'h388a4870),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h340c2848),
	.w1(32'h374588c0),
	.w2(32'h373af26c),
	.w3(32'hb5970b28),
	.w4(32'h3690b185),
	.w5(32'h370949d6),
	.w6(32'hb5f8db08),
	.w7(32'h35be56ca),
	.w8(32'h36ccc421),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996c41f),
	.w1(32'h399faf4f),
	.w2(32'h3985722a),
	.w3(32'hb9ff1747),
	.w4(32'h39983955),
	.w5(32'hb8bd5f41),
	.w6(32'hba7e3a33),
	.w7(32'h38b0f8cb),
	.w8(32'hb9c61480),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h331ecf8d),
	.w1(32'h33b3f2ef),
	.w2(32'h3375457d),
	.w3(32'h34ecfe7f),
	.w4(32'h330ede5a),
	.w5(32'hb3cde2b7),
	.w6(32'h358456b6),
	.w7(32'h3468c1cf),
	.w8(32'hb4bb86be),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35be83d2),
	.w1(32'h36963630),
	.w2(32'hb4e94264),
	.w3(32'h35809d0e),
	.w4(32'h360cb662),
	.w5(32'hb5e3964d),
	.w6(32'h3573c16b),
	.w7(32'hb64ef92a),
	.w8(32'hb6544ce1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f4e3a),
	.w1(32'hb8378556),
	.w2(32'hb8b44a3d),
	.w3(32'h390d1e70),
	.w4(32'hb8f357b3),
	.w5(32'hb81e9014),
	.w6(32'hb70925a1),
	.w7(32'hb8fbf012),
	.w8(32'h391d00c2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acd309),
	.w1(32'hb86f35ba),
	.w2(32'h37b5cb25),
	.w3(32'hb96ae7a3),
	.w4(32'h38b2023f),
	.w5(32'h37dbc2f1),
	.w6(32'hb9966eb6),
	.w7(32'hb91f1fb2),
	.w8(32'hb840573f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a228d6),
	.w1(32'h3963c033),
	.w2(32'h38855a10),
	.w3(32'h383fba59),
	.w4(32'hb7c6dfe8),
	.w5(32'hb89571bf),
	.w6(32'hb8c89501),
	.w7(32'hb93b34f7),
	.w8(32'hb808faa2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4e7a2),
	.w1(32'h38b696f1),
	.w2(32'hb9d23589),
	.w3(32'h39c74009),
	.w4(32'hb9079e13),
	.w5(32'hb89a2795),
	.w6(32'h3910e14e),
	.w7(32'hb928b8b6),
	.w8(32'h390702ec),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34dd34d0),
	.w1(32'h3aa3c1f0),
	.w2(32'hba9bebe9),
	.w3(32'h3af9a09a),
	.w4(32'hba6ec336),
	.w5(32'hbada7bc1),
	.w6(32'hba80fc30),
	.w7(32'hbb384071),
	.w8(32'hb9fb28cf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f2b7),
	.w1(32'h3995da71),
	.w2(32'h3960b3f0),
	.w3(32'hb9ded47a),
	.w4(32'h3998f113),
	.w5(32'h39bac084),
	.w6(32'hba2156df),
	.w7(32'hb9a0f265),
	.w8(32'hb9e6e639),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb2d14),
	.w1(32'hb99013c0),
	.w2(32'h38acf243),
	.w3(32'hb9faa58f),
	.w4(32'h38a0ef57),
	.w5(32'hb7f46bd4),
	.w6(32'hb9fa9f7a),
	.w7(32'hb97facf0),
	.w8(32'hba12838b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d241a6),
	.w1(32'h37716364),
	.w2(32'h3721fa88),
	.w3(32'h3734d141),
	.w4(32'hb72d5667),
	.w5(32'h3813a56e),
	.w6(32'hb8f28253),
	.w7(32'hb901d770),
	.w8(32'hb7f2c793),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3657fc86),
	.w1(32'h366df87a),
	.w2(32'hb4a967e6),
	.w3(32'h3540de1f),
	.w4(32'h350554a2),
	.w5(32'hb60c0acb),
	.w6(32'h35cd8b89),
	.w7(32'hb617f240),
	.w8(32'hb62c1504),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb651b212),
	.w1(32'h366bcf07),
	.w2(32'h3539ff11),
	.w3(32'hb666c82d),
	.w4(32'h3720e253),
	.w5(32'h36125b97),
	.w6(32'hb623ba41),
	.w7(32'h362da26f),
	.w8(32'hb6ba80fe),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5ea1c),
	.w1(32'h386718f1),
	.w2(32'h37b26622),
	.w3(32'h38161774),
	.w4(32'h38943aba),
	.w5(32'h38344c37),
	.w6(32'h38860039),
	.w7(32'h38c41d5f),
	.w8(32'h3848698b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9970541),
	.w1(32'hba154b7e),
	.w2(32'h39003491),
	.w3(32'hba81c896),
	.w4(32'hba054175),
	.w5(32'hb8af0c59),
	.w6(32'hba1e9a47),
	.w7(32'h3a359dd5),
	.w8(32'h3a17be99),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8befb0a),
	.w1(32'h39195f0e),
	.w2(32'h370e6874),
	.w3(32'hb87a4cb4),
	.w4(32'h39a4ec76),
	.w5(32'hb71592d9),
	.w6(32'hb89f6e0f),
	.w7(32'h388c946d),
	.w8(32'hb9c00a7f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890e86a),
	.w1(32'hb9097e6f),
	.w2(32'hb94c1f2b),
	.w3(32'h3a04bd5f),
	.w4(32'h39e62f25),
	.w5(32'h39596ad7),
	.w6(32'h3a07f03a),
	.w7(32'h392f80f3),
	.w8(32'hb9a2a560),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1e910),
	.w1(32'h3951bc30),
	.w2(32'h39752f2e),
	.w3(32'hb8b00b3e),
	.w4(32'h3931cbda),
	.w5(32'h37d6c3a3),
	.w6(32'hb9040106),
	.w7(32'hb7f5cfcd),
	.w8(32'hb8e09001),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a586ab8),
	.w1(32'hb7befcab),
	.w2(32'hb8271471),
	.w3(32'h3a0507bd),
	.w4(32'hb99de263),
	.w5(32'hb76112c2),
	.w6(32'h39a883ff),
	.w7(32'hb990827a),
	.w8(32'h3a2e0610),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3552c40e),
	.w1(32'h35d5f0ee),
	.w2(32'hb577ff98),
	.w3(32'h35a7dec7),
	.w4(32'hb3d12066),
	.w5(32'hb62458ed),
	.w6(32'h354f0191),
	.w7(32'hb5b647fb),
	.w8(32'hb62dc283),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369dbb33),
	.w1(32'h36ea3030),
	.w2(32'hb50d2431),
	.w3(32'h3707b0b1),
	.w4(32'h36a3697f),
	.w5(32'hb67c6611),
	.w6(32'h36f4c124),
	.w7(32'h3574b4e2),
	.w8(32'hb68cd53a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4aeb11f),
	.w1(32'hb6794112),
	.w2(32'h36010756),
	.w3(32'hb6bd3547),
	.w4(32'hb6b26e9e),
	.w5(32'h34c2b355),
	.w6(32'hb621f4a3),
	.w7(32'hb6f8eebd),
	.w8(32'h3617c8a2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c4d5c),
	.w1(32'hb9f668fb),
	.w2(32'hb98ff152),
	.w3(32'hb9a03bd5),
	.w4(32'hb9960e9d),
	.w5(32'h392e54fb),
	.w6(32'hb9ed6610),
	.w7(32'h388942f3),
	.w8(32'h38ca5ead),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb10a3),
	.w1(32'h3908a7c7),
	.w2(32'h396570a0),
	.w3(32'h37c4df51),
	.w4(32'h388d8f9f),
	.w5(32'h396df271),
	.w6(32'hb89a968f),
	.w7(32'h38d5be11),
	.w8(32'h39670d8f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09390f),
	.w1(32'hb790f078),
	.w2(32'h386b601a),
	.w3(32'h3958bba4),
	.w4(32'hb9944ed9),
	.w5(32'hb913a599),
	.w6(32'hb7cde295),
	.w7(32'hb9a521e7),
	.w8(32'h3a103d1e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983455d),
	.w1(32'hb92b6827),
	.w2(32'h36cf4658),
	.w3(32'hb99f2362),
	.w4(32'h38cc073b),
	.w5(32'h38782011),
	.w6(32'hb8a0fa51),
	.w7(32'h39229da4),
	.w8(32'h39370148),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70f0d73),
	.w1(32'h37cd91e8),
	.w2(32'hb761ce2c),
	.w3(32'hb79f9c8d),
	.w4(32'h36634923),
	.w5(32'hb6b2c1da),
	.w6(32'hb8209711),
	.w7(32'hb8083e19),
	.w8(32'hb7c64680),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a55d40),
	.w1(32'hb41e221a),
	.w2(32'h3685230c),
	.w3(32'hb55cab40),
	.w4(32'h3692ac09),
	.w5(32'h3682ec58),
	.w6(32'hb596d854),
	.w7(32'h361e31d7),
	.w8(32'h368d902e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f5766),
	.w1(32'hb7701f8e),
	.w2(32'h35af63d2),
	.w3(32'hb76e2313),
	.w4(32'h381de434),
	.w5(32'h3682a5a5),
	.w6(32'hb87fbf02),
	.w7(32'h3691775e),
	.w8(32'hb873c398),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37267258),
	.w1(32'h380f45a5),
	.w2(32'h38074959),
	.w3(32'h370a1c17),
	.w4(32'h37e61b84),
	.w5(32'h37e6b18a),
	.w6(32'hb6f32e27),
	.w7(32'h35821ff7),
	.w8(32'h3768c2bf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d4f78),
	.w1(32'h37ecc13b),
	.w2(32'h378c6c15),
	.w3(32'h381e1991),
	.w4(32'h37ff4e28),
	.w5(32'hb763e30f),
	.w6(32'h361be918),
	.w7(32'h379e84f4),
	.w8(32'h379bc9a6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6894574),
	.w1(32'hb9500a68),
	.w2(32'h385aa351),
	.w3(32'hb94f73e8),
	.w4(32'hb9595662),
	.w5(32'h38d264bf),
	.w6(32'hb9a559f8),
	.w7(32'hb8730be1),
	.w8(32'h39b71ab8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6a986),
	.w1(32'hb9b1028f),
	.w2(32'h3840dc0a),
	.w3(32'hba78ac06),
	.w4(32'hb8e8a306),
	.w5(32'h38c76404),
	.w6(32'hba8aae62),
	.w7(32'h399d646b),
	.w8(32'h39e8895b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb34df6b6),
	.w1(32'h35c358a9),
	.w2(32'h35ac4b19),
	.w3(32'h35132a3b),
	.w4(32'h362df1bd),
	.w5(32'h35b4860c),
	.w6(32'h34d1b1c5),
	.w7(32'h359336c1),
	.w8(32'hb592964a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d6be1e),
	.w1(32'h36086cf0),
	.w2(32'h3230af78),
	.w3(32'h359219c1),
	.w4(32'h36240fc1),
	.w5(32'h3411178e),
	.w6(32'h3534b611),
	.w7(32'h35c62f67),
	.w8(32'hb61f2160),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h347a8601),
	.w1(32'h34db8dfb),
	.w2(32'h3445949c),
	.w3(32'h34d17b16),
	.w4(32'h3481a7d8),
	.w5(32'hb4098bb1),
	.w6(32'h34a30fab),
	.w7(32'h328e1ce3),
	.w8(32'hb48986eb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33b0b99a),
	.w1(32'h35758dc1),
	.w2(32'hb53fb196),
	.w3(32'h35a1b529),
	.w4(32'h3609577c),
	.w5(32'h35d0b9b0),
	.w6(32'h35d12c79),
	.w7(32'h35e1220d),
	.w8(32'h34c6fecc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6620c),
	.w1(32'h3a90a057),
	.w2(32'h3b075d45),
	.w3(32'hb7b21722),
	.w4(32'hb93e1b6e),
	.w5(32'hb91b992d),
	.w6(32'hba19c5de),
	.w7(32'hba56b4cb),
	.w8(32'h3a2a25d8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d46394),
	.w1(32'hba213625),
	.w2(32'hb99740bd),
	.w3(32'h39935cf9),
	.w4(32'h39dda168),
	.w5(32'h3a2ad64b),
	.w6(32'h39672141),
	.w7(32'h390323a7),
	.w8(32'h3a1aca17),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12de1d),
	.w1(32'hba007b91),
	.w2(32'h38a9d138),
	.w3(32'hba5bf353),
	.w4(32'hb9bcaf12),
	.w5(32'h39fcafb1),
	.w6(32'hba383689),
	.w7(32'h39f16687),
	.w8(32'h39d79ad7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9378caf),
	.w1(32'h3acb5dc4),
	.w2(32'h3a997f37),
	.w3(32'hb990190a),
	.w4(32'h3becd5c8),
	.w5(32'h3a94e195),
	.w6(32'hb9c67f90),
	.w7(32'h3b1dd6c0),
	.w8(32'h3a915196),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40bb7f),
	.w1(32'hbbe5cb52),
	.w2(32'hbbbe324b),
	.w3(32'h3b86d241),
	.w4(32'hbba6bb81),
	.w5(32'hbb3bb6e9),
	.w6(32'hba0721a1),
	.w7(32'hbc238719),
	.w8(32'hbbda5108),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280c8b),
	.w1(32'h3c1384e0),
	.w2(32'h3ad7ef5a),
	.w3(32'hba2ecece),
	.w4(32'h3c0a4e9d),
	.w5(32'h3bf44633),
	.w6(32'hb9530778),
	.w7(32'h3bc901e7),
	.w8(32'h3c516f67),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af43ffa),
	.w1(32'h3b57a894),
	.w2(32'hb98df1d2),
	.w3(32'hba83d459),
	.w4(32'h3b3770e2),
	.w5(32'hbb448bbd),
	.w6(32'h3c1e86ca),
	.w7(32'hb9243a9d),
	.w8(32'hbbd1fd9f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1503a4),
	.w1(32'h3c12bc75),
	.w2(32'h3b7e26c6),
	.w3(32'hbaf97155),
	.w4(32'h3c55d7b3),
	.w5(32'h3c3715df),
	.w6(32'hba4903ca),
	.w7(32'h3c0db15d),
	.w8(32'h3c0a0b7b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc508dd),
	.w1(32'h39c5140b),
	.w2(32'hba83d5b9),
	.w3(32'h3c6fc314),
	.w4(32'hbc003cdc),
	.w5(32'hbb836d7b),
	.w6(32'h3c255f75),
	.w7(32'hbb167ba2),
	.w8(32'hbb8e2891),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c2502),
	.w1(32'hbc0aafc8),
	.w2(32'hbc1c91aa),
	.w3(32'hbba2b48c),
	.w4(32'hbbaaf598),
	.w5(32'hbbe139bb),
	.w6(32'hbb205ccb),
	.w7(32'hbb12c943),
	.w8(32'hbb50946d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d46ac),
	.w1(32'hbba6d3a8),
	.w2(32'hbb8f8453),
	.w3(32'hbbde6a59),
	.w4(32'hbb3c8392),
	.w5(32'hbabdb9ce),
	.w6(32'hbbcc2e54),
	.w7(32'hb9adf3f6),
	.w8(32'h3b4fa175),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a5962),
	.w1(32'h3ad27049),
	.w2(32'h3b4ab3cc),
	.w3(32'h3b676653),
	.w4(32'h3bdbf22b),
	.w5(32'h3c03bf2a),
	.w6(32'h3b1a956d),
	.w7(32'hb941b3b1),
	.w8(32'h3ab3dbe7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc0416),
	.w1(32'h3b4d0f3a),
	.w2(32'h3b29c98c),
	.w3(32'h3c0cb9e4),
	.w4(32'h3a49b7d3),
	.w5(32'hb996b744),
	.w6(32'h3c04c402),
	.w7(32'h3bd02cea),
	.w8(32'h3b601e06),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af40a53),
	.w1(32'hbb616043),
	.w2(32'hba16a7b3),
	.w3(32'h3b2bff6d),
	.w4(32'h3b4f63c0),
	.w5(32'h3a84edd5),
	.w6(32'h3bbf6543),
	.w7(32'h3a597cb9),
	.w8(32'h3b91be28),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4305ef),
	.w1(32'h3bb4524f),
	.w2(32'h3b5aacfb),
	.w3(32'h3b888ac9),
	.w4(32'h3b963831),
	.w5(32'h3baade37),
	.w6(32'h3b063651),
	.w7(32'hba70ba83),
	.w8(32'hba99863b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1314a),
	.w1(32'hba1c6983),
	.w2(32'h39fc71c2),
	.w3(32'h3b67c579),
	.w4(32'h39aafb90),
	.w5(32'h3b3cc47a),
	.w6(32'hba0a7ced),
	.w7(32'hb90d0718),
	.w8(32'h3b2ca02b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be044),
	.w1(32'h3c2c9052),
	.w2(32'h3c4b52af),
	.w3(32'hba0308e5),
	.w4(32'h3b50402e),
	.w5(32'h3bb9acf0),
	.w6(32'h3993851d),
	.w7(32'h3b0a5605),
	.w8(32'h3b306ea6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b004f),
	.w1(32'hbb1032ed),
	.w2(32'hbbbc560e),
	.w3(32'h3b0acdd9),
	.w4(32'h3a98656b),
	.w5(32'hbac20699),
	.w6(32'h3bb02cbc),
	.w7(32'h3ade9e0d),
	.w8(32'hbb227a9f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875bc5),
	.w1(32'h3b55505b),
	.w2(32'hbb3d9e80),
	.w3(32'hbb8304b5),
	.w4(32'h3c18728b),
	.w5(32'h3bbc0a74),
	.w6(32'hbb4c46cb),
	.w7(32'h3cbd9c24),
	.w8(32'h3c880940),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e35c5),
	.w1(32'hbb5c2de2),
	.w2(32'hbb8fc143),
	.w3(32'h3b167881),
	.w4(32'hbb146653),
	.w5(32'hbad388f3),
	.w6(32'h3c58f0ce),
	.w7(32'hb953a077),
	.w8(32'hbad0f94f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2568d5),
	.w1(32'h3b1773a2),
	.w2(32'hbb4c9e9e),
	.w3(32'h3a1b9875),
	.w4(32'h3b03cbd0),
	.w5(32'h3aabfd77),
	.w6(32'hba9ba9f1),
	.w7(32'h3b02edcc),
	.w8(32'h3c055268),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411b25),
	.w1(32'hbb95c5c5),
	.w2(32'hbc8903c6),
	.w3(32'h3b48934d),
	.w4(32'hb9697272),
	.w5(32'hbbab6cb0),
	.w6(32'h3b6a9860),
	.w7(32'hb99beb2a),
	.w8(32'hbaa81ca6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb336852),
	.w1(32'hbb519898),
	.w2(32'hbb853c17),
	.w3(32'hbaee10d0),
	.w4(32'hbba97459),
	.w5(32'h3b59e938),
	.w6(32'h3b5fa5ae),
	.w7(32'h3aee4d67),
	.w8(32'h3a96976b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9328fa),
	.w1(32'hbb84c281),
	.w2(32'hbb4b4657),
	.w3(32'h3ae094ad),
	.w4(32'hbbab9e03),
	.w5(32'h3b6ba63b),
	.w6(32'h3a9c76b0),
	.w7(32'h3a8d856c),
	.w8(32'h3bafbd53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e9d3),
	.w1(32'hbac678af),
	.w2(32'hba2da16c),
	.w3(32'h3ab58e51),
	.w4(32'hbb276256),
	.w5(32'hba4609f2),
	.w6(32'h3bbeaf64),
	.w7(32'hb9b99966),
	.w8(32'h396938f4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e92c7),
	.w1(32'hbaf238f2),
	.w2(32'hbb388ac8),
	.w3(32'h3b3f1cfc),
	.w4(32'h3b239ebf),
	.w5(32'h3b81657f),
	.w6(32'h3a8115e6),
	.w7(32'h3b282d90),
	.w8(32'h3b670991),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e17a),
	.w1(32'h3ab2c336),
	.w2(32'h3b92c9ba),
	.w3(32'h3b3dae50),
	.w4(32'h3b01098b),
	.w5(32'h3ada1063),
	.w6(32'h3b2a7ee7),
	.w7(32'hbacbdec9),
	.w8(32'h3bb63257),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c8754),
	.w1(32'hbbb8f295),
	.w2(32'hbbcee94c),
	.w3(32'hbacb3bbc),
	.w4(32'hba14b22c),
	.w5(32'hbbca5a93),
	.w6(32'h3b5830c7),
	.w7(32'hbbf54617),
	.w8(32'hbc1c4652),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9fc82),
	.w1(32'hbadf994c),
	.w2(32'hbb35d419),
	.w3(32'hbb8cff45),
	.w4(32'hba826b45),
	.w5(32'hb9d698e4),
	.w6(32'hbc327db4),
	.w7(32'h3b28ad37),
	.w8(32'h3b332ec4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab99be2),
	.w1(32'h3c361577),
	.w2(32'h3aa3bad2),
	.w3(32'h3b839869),
	.w4(32'h3c05940c),
	.w5(32'h39c72d01),
	.w6(32'h3b074ebd),
	.w7(32'h3b47b834),
	.w8(32'hbbc97c74),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39576ab1),
	.w1(32'h3be92c20),
	.w2(32'h3b26e733),
	.w3(32'h3b7cd46e),
	.w4(32'h3c4a3b59),
	.w5(32'h3c1b35b9),
	.w6(32'hbb16b240),
	.w7(32'h3c1741d1),
	.w8(32'h3bcd508f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bb289),
	.w1(32'hba4def94),
	.w2(32'hbb8d7888),
	.w3(32'h3bdef383),
	.w4(32'h3a2749bb),
	.w5(32'h3b4eccc4),
	.w6(32'h3b95a8e0),
	.w7(32'h3bd44d21),
	.w8(32'h3bb686fb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e004ac),
	.w1(32'hbabeef39),
	.w2(32'h3a5a9bca),
	.w3(32'h3b52a1ec),
	.w4(32'hbac302a3),
	.w5(32'hba8683ab),
	.w6(32'h3b8e4a8f),
	.w7(32'h3b5309a7),
	.w8(32'hb7aa9408),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb7fd9),
	.w1(32'hba38c0b1),
	.w2(32'hb9812f71),
	.w3(32'h3ad3d3bd),
	.w4(32'hbbce427c),
	.w5(32'hbba1dcd3),
	.w6(32'hb8d1a1f9),
	.w7(32'h3b3b0337),
	.w8(32'h3adcbd78),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dfd03),
	.w1(32'h3bb5cf2f),
	.w2(32'h3a832db9),
	.w3(32'h3b1a195f),
	.w4(32'h3c75da71),
	.w5(32'h3c4b28da),
	.w6(32'h3bc6078a),
	.w7(32'h3c45bec8),
	.w8(32'h3c61bbdc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe1ee5),
	.w1(32'h3b8d2921),
	.w2(32'hbab799b0),
	.w3(32'h3c2dbac9),
	.w4(32'h3bb37482),
	.w5(32'hbadda473),
	.w6(32'h3c43be2b),
	.w7(32'h3c76f331),
	.w8(32'h387f06be),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a654c70),
	.w1(32'hbc18ad24),
	.w2(32'hbc22e73e),
	.w3(32'h3b294588),
	.w4(32'hbc603188),
	.w5(32'hbc11ede1),
	.w6(32'hba7ae668),
	.w7(32'hbb80b4ed),
	.w8(32'hba8b44d5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1fda),
	.w1(32'hbc337643),
	.w2(32'hbc6b2465),
	.w3(32'hbc38db52),
	.w4(32'hba8df805),
	.w5(32'hbbd4297b),
	.w6(32'hbb5483c9),
	.w7(32'h3be238df),
	.w8(32'hbb5ab4db),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78cf92),
	.w1(32'h3c231c5a),
	.w2(32'h3c5e5399),
	.w3(32'hbbf1ed42),
	.w4(32'h3b523540),
	.w5(32'hb8a9ee3f),
	.w6(32'h3a8ddc1b),
	.w7(32'hbbd8f1db),
	.w8(32'hbbfc4ddf),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd325dd),
	.w1(32'h3af4532e),
	.w2(32'h3b05346f),
	.w3(32'h3add2e8a),
	.w4(32'hbb14ab45),
	.w5(32'hbaf96ac5),
	.w6(32'hba8dd92e),
	.w7(32'hb9fda705),
	.w8(32'hba9393f1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe38c7),
	.w1(32'h3b17af6f),
	.w2(32'h3b71399a),
	.w3(32'h3a933abb),
	.w4(32'hba1a5329),
	.w5(32'hba447f35),
	.w6(32'h3a658f7c),
	.w7(32'h397d879e),
	.w8(32'hbacec8ab),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc0e1),
	.w1(32'h3a5c81f9),
	.w2(32'hb8ab847c),
	.w3(32'hbaa96712),
	.w4(32'h3b7c09c9),
	.w5(32'h3b88d67f),
	.w6(32'hbb9c2054),
	.w7(32'h3b28ac68),
	.w8(32'h3b02edd0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977ba1d),
	.w1(32'h3b54534c),
	.w2(32'h3b0f6d93),
	.w3(32'h3b80e5de),
	.w4(32'hbb202e2d),
	.w5(32'hb8de5e2e),
	.w6(32'h3b91459e),
	.w7(32'h3b3aacab),
	.w8(32'h3ad627be),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7adb4b),
	.w1(32'hbb8513d0),
	.w2(32'hbb6e0556),
	.w3(32'hbbb1218f),
	.w4(32'h3a8421c9),
	.w5(32'hbb856434),
	.w6(32'hba2a47b4),
	.w7(32'hbbe0e517),
	.w8(32'hbbdc932c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a71ab),
	.w1(32'hbbd66fa0),
	.w2(32'hbb2630b3),
	.w3(32'h3b3224bb),
	.w4(32'hbb47b35c),
	.w5(32'hbb332f60),
	.w6(32'hbb99151c),
	.w7(32'hbbadd73a),
	.w8(32'hbb0173d6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35f00c),
	.w1(32'h3aee76e9),
	.w2(32'h3b3bedbf),
	.w3(32'hba133810),
	.w4(32'h3af2f52d),
	.w5(32'h3c1099a1),
	.w6(32'hbb29e4b9),
	.w7(32'h3a8bf909),
	.w8(32'h3a573be1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b87d3),
	.w1(32'hbb94b467),
	.w2(32'hbc2109fc),
	.w3(32'h3b342c19),
	.w4(32'hbbbd5e36),
	.w5(32'hbbee501b),
	.w6(32'h3af65324),
	.w7(32'h3a47ba12),
	.w8(32'hb86fde65),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3268e),
	.w1(32'hbbb39b3f),
	.w2(32'hbc0eacd5),
	.w3(32'hbbbcc380),
	.w4(32'h3c05544b),
	.w5(32'hba2ea2aa),
	.w6(32'hba80e8ab),
	.w7(32'h3c1e4fcf),
	.w8(32'h3898b3ed),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df9e3),
	.w1(32'h39c84a2b),
	.w2(32'h3a59ea49),
	.w3(32'hbc04214c),
	.w4(32'h3b0ad718),
	.w5(32'h39585d28),
	.w6(32'hbbf24a11),
	.w7(32'h3b312de0),
	.w8(32'h3bb7ab95),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47ee2b),
	.w1(32'h399ba85d),
	.w2(32'hbb1fa0bd),
	.w3(32'hbb25851a),
	.w4(32'h3af84125),
	.w5(32'h3ac2d3b5),
	.w6(32'h3b8f1d59),
	.w7(32'h3b108b06),
	.w8(32'h3b79fbca),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec16a),
	.w1(32'hbb47846f),
	.w2(32'hbbd2d427),
	.w3(32'h3b0763a6),
	.w4(32'hbb4b24d5),
	.w5(32'hbbb4c03a),
	.w6(32'h3b626565),
	.w7(32'hbad34948),
	.w8(32'hbb4355f1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80250e),
	.w1(32'hbb8d1889),
	.w2(32'hbb6524f3),
	.w3(32'hbb14677a),
	.w4(32'h3b18d12d),
	.w5(32'hba83939d),
	.w6(32'hbb5de229),
	.w7(32'h3ae2932f),
	.w8(32'h3b079d44),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1d356),
	.w1(32'h3ab83698),
	.w2(32'hbbfd459a),
	.w3(32'hbb5757c5),
	.w4(32'h3bcd12b8),
	.w5(32'h3aa055d9),
	.w6(32'hbab89e04),
	.w7(32'h3bdfa2e9),
	.w8(32'hbac75601),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ee2dc),
	.w1(32'hbbb0be1a),
	.w2(32'hbc0edc34),
	.w3(32'h3b6c8e69),
	.w4(32'hbb53e896),
	.w5(32'hbbd48737),
	.w6(32'h3b675a1e),
	.w7(32'hbb0b6a3c),
	.w8(32'h391ff115),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc274c68),
	.w1(32'h397b31d1),
	.w2(32'hbb3c6283),
	.w3(32'hbbc69840),
	.w4(32'h3a324833),
	.w5(32'hbaa55e27),
	.w6(32'hbb8545aa),
	.w7(32'hbad9eabd),
	.w8(32'hb90a8f68),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845293),
	.w1(32'hbb012961),
	.w2(32'h3b13223d),
	.w3(32'hbae5006b),
	.w4(32'hbbd72f4f),
	.w5(32'hbb1784dc),
	.w6(32'hbae1f48b),
	.w7(32'hbb6409d3),
	.w8(32'hba3ad9b1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bff4),
	.w1(32'hbb72a66d),
	.w2(32'hbbd41496),
	.w3(32'hbb1705ad),
	.w4(32'hbbef6117),
	.w5(32'hbc36b0ab),
	.w6(32'hba67a585),
	.w7(32'hbbd93c61),
	.w8(32'hbbeed5a1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f99c9),
	.w1(32'hba7181c6),
	.w2(32'h3a146945),
	.w3(32'hbbea9709),
	.w4(32'hbb9a6e68),
	.w5(32'h3b31d81b),
	.w6(32'hbb0aa0c4),
	.w7(32'hbbe752e8),
	.w8(32'hbb613803),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc8f8b),
	.w1(32'hbb0e745c),
	.w2(32'hbbc4ba42),
	.w3(32'h3902b456),
	.w4(32'hba1e6dcc),
	.w5(32'h3add689c),
	.w6(32'hbae31702),
	.w7(32'hbb4702bb),
	.w8(32'h3ae371a4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849871),
	.w1(32'hbc47b7c2),
	.w2(32'hbc150629),
	.w3(32'hbadf5d49),
	.w4(32'hbbbf2baf),
	.w5(32'hbc0dd0ae),
	.w6(32'h3a1cc73d),
	.w7(32'hbc0b63d4),
	.w8(32'hbc1987dc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35e4c),
	.w1(32'h39718e64),
	.w2(32'h3988174d),
	.w3(32'hbc2405c3),
	.w4(32'h3bd6adc9),
	.w5(32'h3afd8a22),
	.w6(32'hbc3353a6),
	.w7(32'h3bd87781),
	.w8(32'h3b6c3258),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f0179),
	.w1(32'hbabe6e57),
	.w2(32'hbbb81acf),
	.w3(32'h3b397256),
	.w4(32'h3a92b024),
	.w5(32'hbb1f0275),
	.w6(32'h3b51b52f),
	.w7(32'h3a8e5171),
	.w8(32'hba94f09a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd9aa0),
	.w1(32'hbad72328),
	.w2(32'hbb765964),
	.w3(32'hbb8edc4a),
	.w4(32'hbb145302),
	.w5(32'hba739de8),
	.w6(32'hbb841386),
	.w7(32'h3a829921),
	.w8(32'h3b924ec0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0796e2),
	.w1(32'h39a2a9e7),
	.w2(32'h3aef73cf),
	.w3(32'hba3f9303),
	.w4(32'h39fb46b9),
	.w5(32'h3afce500),
	.w6(32'h3a53305f),
	.w7(32'hbab9adc9),
	.w8(32'h3a86bf58),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1824a4),
	.w1(32'hbba98302),
	.w2(32'hbc13227e),
	.w3(32'h3b9fc42c),
	.w4(32'hba11ae41),
	.w5(32'h36e76d9e),
	.w6(32'h3b3a14e9),
	.w7(32'hbbc99951),
	.w8(32'hba966a4a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb681),
	.w1(32'hbb45313c),
	.w2(32'hbb8387bb),
	.w3(32'hbb7637a7),
	.w4(32'hbaeaaec9),
	.w5(32'hbc0b80ad),
	.w6(32'hbb4649e6),
	.w7(32'hb984492e),
	.w8(32'hb983d570),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b536),
	.w1(32'h3b040d8e),
	.w2(32'h3988fdcb),
	.w3(32'hbc4d4fa3),
	.w4(32'hba8b26b0),
	.w5(32'hbac839f1),
	.w6(32'hbb82f745),
	.w7(32'hb9ae9c7f),
	.w8(32'hbb99df10),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b2716),
	.w1(32'h3adb0107),
	.w2(32'h3afae66b),
	.w3(32'hbb00239d),
	.w4(32'h3b5d4ae1),
	.w5(32'h3b0697df),
	.w6(32'hbb8cbb83),
	.w7(32'h3b35dbed),
	.w8(32'hbb12de3b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a5e9),
	.w1(32'h3bef6e8e),
	.w2(32'h3b98861d),
	.w3(32'h3b189c54),
	.w4(32'h3c4159c0),
	.w5(32'h3bf7071f),
	.w6(32'hbb659eee),
	.w7(32'h3be7d631),
	.w8(32'h3b2225ed),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be44288),
	.w1(32'h3c1f05f5),
	.w2(32'h3c302a81),
	.w3(32'h3c4ba65d),
	.w4(32'h3c84cbff),
	.w5(32'h3c9b0e82),
	.w6(32'h3b997895),
	.w7(32'hbba70ab4),
	.w8(32'hb98f4f09),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c499203),
	.w1(32'hbb8bc599),
	.w2(32'hbc104cc0),
	.w3(32'h3c8ef6db),
	.w4(32'h3b56681c),
	.w5(32'hb9f74832),
	.w6(32'h3b3a852f),
	.w7(32'h3c451231),
	.w8(32'h3bfefaec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1dffe),
	.w1(32'h3b1164f1),
	.w2(32'h3ad478d5),
	.w3(32'h3b923642),
	.w4(32'h3aec49fd),
	.w5(32'h3b76f03d),
	.w6(32'h3c269d87),
	.w7(32'h3b5b1658),
	.w8(32'hbad6eef8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4bd6),
	.w1(32'h3bbb11ee),
	.w2(32'h3b582bd1),
	.w3(32'h3bbb1e8b),
	.w4(32'h39a3a6b1),
	.w5(32'h3b4a0030),
	.w6(32'h3b7d21c9),
	.w7(32'h3a8c172d),
	.w8(32'hba933567),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06c3e5),
	.w1(32'h39009840),
	.w2(32'hba6edb30),
	.w3(32'hbac2859e),
	.w4(32'h3b4b7235),
	.w5(32'h3b25bf15),
	.w6(32'hb8b8dc48),
	.w7(32'h3b470cea),
	.w8(32'h3b91c50b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb9f4),
	.w1(32'h3bc68ecb),
	.w2(32'h3c2ee103),
	.w3(32'hbaa52130),
	.w4(32'hb6d4c15a),
	.w5(32'h3c0930b2),
	.w6(32'h3b0598e7),
	.w7(32'hbb3e7c72),
	.w8(32'h3bbee268),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4fbaa),
	.w1(32'h3c6771c4),
	.w2(32'h3bc781aa),
	.w3(32'h3a884783),
	.w4(32'h3c36df3e),
	.w5(32'h3b17f518),
	.w6(32'h3ba7b433),
	.w7(32'h3cba91b2),
	.w8(32'h3bf65c30),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65f9ce),
	.w1(32'hbb3c20b9),
	.w2(32'hbbf3c7b7),
	.w3(32'h3af45d51),
	.w4(32'h3af9aae4),
	.w5(32'h3ae2994b),
	.w6(32'h3c114646),
	.w7(32'hbabdf44a),
	.w8(32'hbb4bef3b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f461),
	.w1(32'hb9700ecd),
	.w2(32'hba8aa350),
	.w3(32'hbb0dcbef),
	.w4(32'h3a61b6f7),
	.w5(32'h3af95273),
	.w6(32'hbb884548),
	.w7(32'hbb84cdb3),
	.w8(32'hbb83c637),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f626c9),
	.w1(32'hb954c146),
	.w2(32'hbb87a8f4),
	.w3(32'hbb115e36),
	.w4(32'h3bc64cae),
	.w5(32'h3b422466),
	.w6(32'hbbb56e5d),
	.w7(32'h3bf80dc1),
	.w8(32'h3bf1d852),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82fc54),
	.w1(32'hbbc177db),
	.w2(32'hbab73053),
	.w3(32'hbb5874dc),
	.w4(32'h3b476983),
	.w5(32'hba3100ad),
	.w6(32'h3b8a9f35),
	.w7(32'h3bb51b2e),
	.w8(32'h3bb683a0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad57bee),
	.w1(32'hbb17be06),
	.w2(32'hbb1372d4),
	.w3(32'h3b466ee4),
	.w4(32'h3ba6fddc),
	.w5(32'h3be3483d),
	.w6(32'h3b5d5e05),
	.w7(32'h3c207461),
	.w8(32'h3bcad8c6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6911e),
	.w1(32'h39318475),
	.w2(32'h3a82326e),
	.w3(32'h3b48aa77),
	.w4(32'h3b93aa07),
	.w5(32'h3b30eb7c),
	.w6(32'h3ba1caef),
	.w7(32'h3abc0d40),
	.w8(32'h3bad8fd4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d485),
	.w1(32'hbb38e48e),
	.w2(32'hbb8bb54f),
	.w3(32'hba16f531),
	.w4(32'hbb4f5e63),
	.w5(32'hbbb079db),
	.w6(32'hbb5aa9f3),
	.w7(32'hbacfee27),
	.w8(32'hbbdac833),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab68637),
	.w1(32'hba0749dc),
	.w2(32'hbb9470b1),
	.w3(32'hbb8f43e9),
	.w4(32'h3b27eefa),
	.w5(32'hbb367f15),
	.w6(32'hbbed7c4c),
	.w7(32'hb996dd58),
	.w8(32'hbad2d17a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba741e9),
	.w1(32'hba82d011),
	.w2(32'h3af626ab),
	.w3(32'hbaa507f0),
	.w4(32'hbafe8a03),
	.w5(32'hbb4895c7),
	.w6(32'hba8c309c),
	.w7(32'h3a86a4ce),
	.w8(32'h3b6fe90f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c6a4c),
	.w1(32'h3c10959e),
	.w2(32'h3bb5623e),
	.w3(32'h3b0d2044),
	.w4(32'h3bb73e24),
	.w5(32'h3b7b473c),
	.w6(32'h3b8d37fd),
	.w7(32'hba6c5337),
	.w8(32'hbb8cd4c9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16eba7),
	.w1(32'h3b9c5464),
	.w2(32'h3b809a24),
	.w3(32'hba1323db),
	.w4(32'h3b0b1227),
	.w5(32'hbbe4d0a9),
	.w6(32'hbc0f4c02),
	.w7(32'hbaadc052),
	.w8(32'hbb821ab0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c82552),
	.w1(32'h3a9d1001),
	.w2(32'hb9c0c7cf),
	.w3(32'hbb9499c0),
	.w4(32'h3b03ea6e),
	.w5(32'h3b9b417c),
	.w6(32'h390bd5b2),
	.w7(32'hba38a64f),
	.w8(32'h3b84a1b0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac68965),
	.w1(32'h3b61aa9a),
	.w2(32'h39c8f128),
	.w3(32'h3b7207ba),
	.w4(32'h3b9a49cf),
	.w5(32'h3bb68356),
	.w6(32'h3b858f79),
	.w7(32'h3bebeba1),
	.w8(32'h3bc77f2e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad20f83),
	.w1(32'hba3ae353),
	.w2(32'hb9176503),
	.w3(32'h3baa664b),
	.w4(32'h3a925034),
	.w5(32'hbad2f75a),
	.w6(32'hbb24233d),
	.w7(32'h3a04d517),
	.w8(32'hbb43a577),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d22d),
	.w1(32'hba91f1b5),
	.w2(32'hbb375d6b),
	.w3(32'hba8f61f5),
	.w4(32'hba61536a),
	.w5(32'hbaf6f026),
	.w6(32'hbb0bbcc8),
	.w7(32'hba0475ad),
	.w8(32'h3ab69ba5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac936af),
	.w1(32'hbaa8d628),
	.w2(32'hb8a56897),
	.w3(32'hbace46bb),
	.w4(32'h3a760451),
	.w5(32'h3a9d1b74),
	.w6(32'hb9a51e34),
	.w7(32'h3a876499),
	.w8(32'h3b5bf5bb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacaca8),
	.w1(32'hba06dffb),
	.w2(32'hbb144da9),
	.w3(32'hba8d1414),
	.w4(32'hbac97947),
	.w5(32'hbb95dd86),
	.w6(32'hba748986),
	.w7(32'h399fd286),
	.w8(32'hb77baf9c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8ed8),
	.w1(32'h3c69754b),
	.w2(32'h3c5762da),
	.w3(32'hbb1fb792),
	.w4(32'h3c531361),
	.w5(32'h3ca5eb52),
	.w6(32'h3a034aec),
	.w7(32'h3c05f615),
	.w8(32'h3c8c1535),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8863),
	.w1(32'h3b8fba31),
	.w2(32'h3ba57fa5),
	.w3(32'h3c7503fd),
	.w4(32'h3b55335a),
	.w5(32'h3b7c35d4),
	.w6(32'h3c70bf35),
	.w7(32'h3b27c537),
	.w8(32'h3b9576e2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87453f),
	.w1(32'h3b5fa3e0),
	.w2(32'h3bc3e0bb),
	.w3(32'h3b2bc120),
	.w4(32'h3b8b5e55),
	.w5(32'h3be5dcf4),
	.w6(32'h3bad0efe),
	.w7(32'h3b367fdf),
	.w8(32'hbb569f95),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09097),
	.w1(32'h3bc9f2fb),
	.w2(32'h3b5a5e7d),
	.w3(32'h3b88e4a3),
	.w4(32'hba157076),
	.w5(32'h3aa3c8d3),
	.w6(32'h3aa982ba),
	.w7(32'h3b54b568),
	.w8(32'hbab445b3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb625f3),
	.w1(32'hbb52245f),
	.w2(32'hba959515),
	.w3(32'hbc09ebdd),
	.w4(32'h3b06efca),
	.w5(32'hbb19c398),
	.w6(32'hba8a34a2),
	.w7(32'h3b44d98b),
	.w8(32'h3ab0ad69),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dc652),
	.w1(32'hbb6344e4),
	.w2(32'hbbe7f1b1),
	.w3(32'h3973fd90),
	.w4(32'hbc37f31e),
	.w5(32'hbb80d0f2),
	.w6(32'h3ade61cf),
	.w7(32'hbbf745fe),
	.w8(32'hbb9ff3b6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c77b1),
	.w1(32'h3c82da8a),
	.w2(32'h3c3a58e2),
	.w3(32'hbbd0a842),
	.w4(32'h3c460d9f),
	.w5(32'h3c1bc3df),
	.w6(32'hbb9239e4),
	.w7(32'h3c2e0269),
	.w8(32'h3beb8bd9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4edca),
	.w1(32'h3ad91c6d),
	.w2(32'hbb261b83),
	.w3(32'h3c02971a),
	.w4(32'h3a82a39b),
	.w5(32'hbb845db0),
	.w6(32'h3b76c2dd),
	.w7(32'h38159d11),
	.w8(32'hbad1d562),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b5d3),
	.w1(32'h3b2ee861),
	.w2(32'h3b2f17f2),
	.w3(32'hb67ddc52),
	.w4(32'h3b0176d4),
	.w5(32'h3a821872),
	.w6(32'hbac3e7c8),
	.w7(32'hbaa4c17a),
	.w8(32'h3aadeb64),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa130),
	.w1(32'h3af2259a),
	.w2(32'hbaa16102),
	.w3(32'h3b2803c3),
	.w4(32'h3ba6a354),
	.w5(32'h3c3906f1),
	.w6(32'h3a2fa68f),
	.w7(32'h3c8b711c),
	.w8(32'h3c9b4381),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd543),
	.w1(32'hbb8250f6),
	.w2(32'hbbc513b7),
	.w3(32'h3b6e4c25),
	.w4(32'hbb89862b),
	.w5(32'hbbb1ac11),
	.w6(32'h3c9db78c),
	.w7(32'h3af467e5),
	.w8(32'hbb866a62),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7c948),
	.w1(32'h3b9ffba5),
	.w2(32'h3bbe1f68),
	.w3(32'hbbc77499),
	.w4(32'h3b51f3b3),
	.w5(32'h3c092012),
	.w6(32'hbbafadb2),
	.w7(32'h3b641576),
	.w8(32'h3c8c9057),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb311852),
	.w1(32'hb996afbd),
	.w2(32'hbb129819),
	.w3(32'hb997d1ad),
	.w4(32'hba0099cb),
	.w5(32'hb98c22b4),
	.w6(32'h3c34f75c),
	.w7(32'hba1d0336),
	.w8(32'hbb12bd02),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e86b1c),
	.w1(32'hba3718ec),
	.w2(32'hbb3aef3b),
	.w3(32'hbb6a0b12),
	.w4(32'h3aeacd38),
	.w5(32'h3abdb66a),
	.w6(32'hbbc21aee),
	.w7(32'h3b20b87c),
	.w8(32'h3b0796ae),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9cd81),
	.w1(32'hbb7f39fa),
	.w2(32'hb9d05a21),
	.w3(32'h3bf7b735),
	.w4(32'h399c0a28),
	.w5(32'hbaed976b),
	.w6(32'h3bdcbb8b),
	.w7(32'hbbcf3f5b),
	.w8(32'hbc00ff05),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396fdc84),
	.w1(32'hbb3e357f),
	.w2(32'h39957934),
	.w3(32'hba8e32ff),
	.w4(32'h37b4c36a),
	.w5(32'hbb3d2593),
	.w6(32'hbb8a8edd),
	.w7(32'hbb992999),
	.w8(32'hbb265139),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22375b),
	.w1(32'h3b03eb67),
	.w2(32'hbbac47ef),
	.w3(32'h3a8aefc5),
	.w4(32'h3bfb325c),
	.w5(32'hbbb98185),
	.w6(32'h396605e6),
	.w7(32'h3c05261e),
	.w8(32'hbb08c92d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4347ad),
	.w1(32'h3b435f41),
	.w2(32'h3b5c4120),
	.w3(32'hbb9e6798),
	.w4(32'h3ba425d0),
	.w5(32'h3b807834),
	.w6(32'hbc012a79),
	.w7(32'h39aff890),
	.w8(32'h3ab3f020),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0adb93),
	.w1(32'h3b1c3173),
	.w2(32'h3bc89717),
	.w3(32'h3bfff88d),
	.w4(32'h3a91f3f5),
	.w5(32'h3b9d88d5),
	.w6(32'h3bd030de),
	.w7(32'hbb935874),
	.w8(32'h3b17804f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfa658),
	.w1(32'hba1e9747),
	.w2(32'hbac027bd),
	.w3(32'h3af20478),
	.w4(32'hb9191f40),
	.w5(32'h3940e264),
	.w6(32'hba67d006),
	.w7(32'h3b587f7f),
	.w8(32'h398dec95),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac0d46),
	.w1(32'h3bd5bf49),
	.w2(32'h3b90318e),
	.w3(32'hbb4e8027),
	.w4(32'h3bce7a60),
	.w5(32'hb92c8a08),
	.w6(32'hbbac3a31),
	.w7(32'h3b76c3e3),
	.w8(32'hbb825fef),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38edb80c),
	.w1(32'h3b721b93),
	.w2(32'h3a5fddd0),
	.w3(32'h3b4ac433),
	.w4(32'h3bf2f015),
	.w5(32'h3bb27a4d),
	.w6(32'hbb2a2f7f),
	.w7(32'h3bc81b63),
	.w8(32'h3bc38f7c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b929983),
	.w1(32'hbb9feeb1),
	.w2(32'hbbb6453f),
	.w3(32'h3c05889b),
	.w4(32'hbb00275d),
	.w5(32'hbb930983),
	.w6(32'h3c1efcf3),
	.w7(32'hbb0803ba),
	.w8(32'hbb119bad),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81bbc4),
	.w1(32'h3bb5f918),
	.w2(32'h3c003168),
	.w3(32'h3b66aab4),
	.w4(32'h3b67438f),
	.w5(32'h3c153ee3),
	.w6(32'h3bb6860e),
	.w7(32'hba5f2769),
	.w8(32'h3c0cb652),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e7c4),
	.w1(32'hbc11d280),
	.w2(32'hbc1463c0),
	.w3(32'h3bc0a4af),
	.w4(32'hbc5d10f2),
	.w5(32'hbc70713d),
	.w6(32'h3bbc1376),
	.w7(32'hbc02b4b6),
	.w8(32'hbc039405),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc458b3f),
	.w1(32'hbb417933),
	.w2(32'hbb59ff13),
	.w3(32'hbc10a618),
	.w4(32'hbb419d39),
	.w5(32'hbaec9343),
	.w6(32'hbbeebc46),
	.w7(32'hbb20f6df),
	.w8(32'hbb66301d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b28a),
	.w1(32'h3a95cd46),
	.w2(32'h3add33f1),
	.w3(32'hbaea0333),
	.w4(32'h3b48dcf2),
	.w5(32'hba700feb),
	.w6(32'hbb816bbb),
	.w7(32'h3bed6b58),
	.w8(32'hbae1615f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a617fa4),
	.w1(32'hbbc6e045),
	.w2(32'hbb9f3197),
	.w3(32'hbb1a4e64),
	.w4(32'h3a771be1),
	.w5(32'h3ba17f0e),
	.w6(32'hbaa10a10),
	.w7(32'h3b6c3347),
	.w8(32'h3c141df4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca082a),
	.w1(32'hbad0ad78),
	.w2(32'hbb1e2176),
	.w3(32'h3b9bad2d),
	.w4(32'h3b48b07d),
	.w5(32'hba8967bb),
	.w6(32'h3c33fdac),
	.w7(32'hbb0ce505),
	.w8(32'h393cb740),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec01d3),
	.w1(32'h3b076714),
	.w2(32'h3b00e22f),
	.w3(32'hba4952ad),
	.w4(32'h3b27fd41),
	.w5(32'h3bb18329),
	.w6(32'h3af55021),
	.w7(32'hba9b117e),
	.w8(32'hbb1756de),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e6bd),
	.w1(32'hbc001acc),
	.w2(32'hbb9950b3),
	.w3(32'h3c38d069),
	.w4(32'hbbe1fb89),
	.w5(32'hbb080e8c),
	.w6(32'h390c062c),
	.w7(32'hbbd48bce),
	.w8(32'hbb5b98df),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a66f2),
	.w1(32'h3af027db),
	.w2(32'h3c09de05),
	.w3(32'hba967511),
	.w4(32'h3b0ab2e0),
	.w5(32'h3c13d7c2),
	.w6(32'hbb80d442),
	.w7(32'h3985629c),
	.w8(32'h3c85e6bc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee6f8),
	.w1(32'hbadc97d6),
	.w2(32'hba9afbab),
	.w3(32'h3bb1420e),
	.w4(32'hbb4da691),
	.w5(32'h3990980a),
	.w6(32'h3c4519e7),
	.w7(32'h3a148591),
	.w8(32'h3b000999),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57bf48),
	.w1(32'h3b8f184b),
	.w2(32'h3bbd0be2),
	.w3(32'h3b087d5a),
	.w4(32'h3b93a8a2),
	.w5(32'h3ba89735),
	.w6(32'h3b29e0ef),
	.w7(32'h3b273d0c),
	.w8(32'h3ab599ad),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2513d),
	.w1(32'h3b404f47),
	.w2(32'h3a465624),
	.w3(32'h3b4f3f9b),
	.w4(32'hb9543d74),
	.w5(32'hbb232e81),
	.w6(32'h3a929ddc),
	.w7(32'h3a2e2cbb),
	.w8(32'hba763b68),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39626edd),
	.w1(32'h3a1fd869),
	.w2(32'hba23094e),
	.w3(32'hbb1fc3ff),
	.w4(32'h3b242442),
	.w5(32'hbb27d8aa),
	.w6(32'hbb96954d),
	.w7(32'h39121548),
	.w8(32'h3a9097ac),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4401e0),
	.w1(32'hbb9943a8),
	.w2(32'hba2913aa),
	.w3(32'hbae961a1),
	.w4(32'hb9e023ff),
	.w5(32'h3b9f267c),
	.w6(32'hbaf7931e),
	.w7(32'hbb50b6ef),
	.w8(32'h3b937838),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ce57),
	.w1(32'hbba11ec6),
	.w2(32'hbb75feec),
	.w3(32'h3a8b4574),
	.w4(32'hbb1d46ce),
	.w5(32'hbb255281),
	.w6(32'hbbaf93a2),
	.w7(32'hbb9172f0),
	.w8(32'hbb156fe4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395620c2),
	.w1(32'hbc1221e6),
	.w2(32'hbc132d5e),
	.w3(32'h3b837133),
	.w4(32'h397b32d7),
	.w5(32'hb8ed9590),
	.w6(32'h3b548182),
	.w7(32'hbc024f3e),
	.w8(32'hbb06a5ca),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35c91a),
	.w1(32'hbb796126),
	.w2(32'h3ae8e17a),
	.w3(32'hbcb9d1ee),
	.w4(32'h3c0cea7c),
	.w5(32'h3bdaf926),
	.w6(32'hbc91a33f),
	.w7(32'h3b97aa19),
	.w8(32'hbbdb11fa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcfdb1),
	.w1(32'h3b6e6612),
	.w2(32'h3bef54d2),
	.w3(32'hbc084b5a),
	.w4(32'h3b61a833),
	.w5(32'hbc0295a8),
	.w6(32'hbb8fb762),
	.w7(32'hba142fb7),
	.w8(32'h3c303937),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bb0df),
	.w1(32'h3a8c7935),
	.w2(32'h3aa557c2),
	.w3(32'hbb670f7e),
	.w4(32'hba8dde2c),
	.w5(32'hbc16eb0c),
	.w6(32'hbb2aaf82),
	.w7(32'h3bb4cda7),
	.w8(32'h3be2f98e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d00c),
	.w1(32'h3b07c0e0),
	.w2(32'h3b74b398),
	.w3(32'h3acb0ec6),
	.w4(32'h3abe0890),
	.w5(32'h3b92a47b),
	.w6(32'hbb03c8af),
	.w7(32'h3b4bc0f6),
	.w8(32'hbb2f1df0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a071e92),
	.w1(32'h3bee50a7),
	.w2(32'h3c3245c4),
	.w3(32'h3b31c1cc),
	.w4(32'hbc7e60dd),
	.w5(32'hbb0a8f52),
	.w6(32'h3a7335a5),
	.w7(32'h3b079da1),
	.w8(32'h3b013043),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137239),
	.w1(32'hbbb80b06),
	.w2(32'hba674d26),
	.w3(32'h3b93c54d),
	.w4(32'hbaa3c3b9),
	.w5(32'hbb29665b),
	.w6(32'h3ac9d4f3),
	.w7(32'hbbd1578a),
	.w8(32'hbb87f816),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba57cab),
	.w1(32'h3c039ac0),
	.w2(32'h3b6f4bcb),
	.w3(32'hba5afa40),
	.w4(32'h3b500a06),
	.w5(32'h3c6d541e),
	.w6(32'h38b08942),
	.w7(32'h3b81480d),
	.w8(32'h3b84ad4e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a48c),
	.w1(32'hbc19eea6),
	.w2(32'hbc15a12e),
	.w3(32'h3b8203a0),
	.w4(32'hbbc08665),
	.w5(32'hbc035d20),
	.w6(32'h3ab4d252),
	.w7(32'hbb1db264),
	.w8(32'h3b11c0d2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5fb5a),
	.w1(32'h39327551),
	.w2(32'hba5e4dff),
	.w3(32'hbc7241d8),
	.w4(32'h3b230ec3),
	.w5(32'hbb348c36),
	.w6(32'hbbf175eb),
	.w7(32'h3b33c72a),
	.w8(32'h3a522c97),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5c7a5),
	.w1(32'hbc6bcbc0),
	.w2(32'hbc62050f),
	.w3(32'h3a1168ec),
	.w4(32'hbc4a5076),
	.w5(32'h3a957aa4),
	.w6(32'h3b1502c9),
	.w7(32'hbba0b42f),
	.w8(32'hbb822de8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847955),
	.w1(32'h3c52a8cb),
	.w2(32'h3c89489e),
	.w3(32'hbc25b558),
	.w4(32'h3c7fd8d9),
	.w5(32'hbb3fa452),
	.w6(32'hbbef4928),
	.w7(32'h3c694239),
	.w8(32'h3c911e69),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a3384),
	.w1(32'hbacb1531),
	.w2(32'hbb64e6b9),
	.w3(32'h3c8e8ce1),
	.w4(32'h3c0b8f41),
	.w5(32'h3c1940d5),
	.w6(32'h3c18dad6),
	.w7(32'h3b775650),
	.w8(32'h3ab5f814),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0815a6),
	.w1(32'hbbaf50ce),
	.w2(32'hbb0e0a45),
	.w3(32'hbcb79f10),
	.w4(32'h3b606f92),
	.w5(32'hb9cca8a3),
	.w6(32'hbc1cda34),
	.w7(32'hbaf377dd),
	.w8(32'h3b0266b2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c548c),
	.w1(32'hba185076),
	.w2(32'hbc528dac),
	.w3(32'hb99980f5),
	.w4(32'hbc76eeb3),
	.w5(32'h3b1e3046),
	.w6(32'h3b378dfd),
	.w7(32'hbc06a3e9),
	.w8(32'hbbd2435c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d2b5),
	.w1(32'hbc20b325),
	.w2(32'hbc18a4a5),
	.w3(32'hbbb81129),
	.w4(32'hbbddb838),
	.w5(32'hbadd4c00),
	.w6(32'hbb9edc23),
	.w7(32'hbc0d0310),
	.w8(32'hba8c9c96),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818c7a),
	.w1(32'hbc27a8c8),
	.w2(32'hbc24c122),
	.w3(32'hbadb3f53),
	.w4(32'hbb00857f),
	.w5(32'hbbcfd4f6),
	.w6(32'h3a338998),
	.w7(32'hbc467fd2),
	.w8(32'hbbf1e050),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09769b),
	.w1(32'hbbdaa5fc),
	.w2(32'hbbbca7ea),
	.w3(32'hbbd0471b),
	.w4(32'hbc81eb67),
	.w5(32'h3b158c35),
	.w6(32'hbbecbfc6),
	.w7(32'hbbd9d78d),
	.w8(32'hbc187c1a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc470fc7),
	.w1(32'h3ae1e0b0),
	.w2(32'h3ae91108),
	.w3(32'hbb97cbc8),
	.w4(32'hbbcf68f9),
	.w5(32'h3ba15481),
	.w6(32'hbc7413cf),
	.w7(32'hbc0fbdeb),
	.w8(32'hbac370a7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e9c05),
	.w1(32'hbb192d90),
	.w2(32'h3a2229de),
	.w3(32'h3b15f2eb),
	.w4(32'hb989d6f4),
	.w5(32'h3c712761),
	.w6(32'hb605f750),
	.w7(32'h3bfb19c0),
	.w8(32'h3bbd23b8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c465),
	.w1(32'h3be329bf),
	.w2(32'hbb4aa78b),
	.w3(32'h3c13a0c9),
	.w4(32'h3c1d687c),
	.w5(32'hbc4da58d),
	.w6(32'h3a970415),
	.w7(32'h3b8ed1ab),
	.w8(32'h3b953c08),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53478e),
	.w1(32'hb953079c),
	.w2(32'hbc044fe0),
	.w3(32'hbbf8acd2),
	.w4(32'hbbfd9b58),
	.w5(32'h3bae0b40),
	.w6(32'hbb9443c3),
	.w7(32'hbc214063),
	.w8(32'hbb729db3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45694b),
	.w1(32'h3a8dd37b),
	.w2(32'h3bb7c55b),
	.w3(32'hbb5095bd),
	.w4(32'h3bb8b24f),
	.w5(32'hba4acc1f),
	.w6(32'hbbdbf8fc),
	.w7(32'h3c12b48c),
	.w8(32'hbb247d63),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3be575),
	.w1(32'h3b59b25b),
	.w2(32'h3b037e4e),
	.w3(32'h3c2203f4),
	.w4(32'h3b7a10e6),
	.w5(32'hbb9acdc8),
	.w6(32'h3ba64a41),
	.w7(32'h3b508aa8),
	.w8(32'hbaee79ee),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf16c00),
	.w1(32'hba6c3448),
	.w2(32'hba9abac5),
	.w3(32'h3ba1bb7e),
	.w4(32'hbb2cdb64),
	.w5(32'h3b646ac8),
	.w6(32'h3c00363e),
	.w7(32'hbb458452),
	.w8(32'hbb2566fe),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dcb66),
	.w1(32'h3a82be6a),
	.w2(32'h3b92b803),
	.w3(32'h3b95f9dd),
	.w4(32'hbbbcd42f),
	.w5(32'h3c116b95),
	.w6(32'h3b179cd0),
	.w7(32'hbb5bc1c8),
	.w8(32'hbc2832c0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34239b),
	.w1(32'hb627ad53),
	.w2(32'hbc19020a),
	.w3(32'h3a56dd17),
	.w4(32'hbc08b767),
	.w5(32'h3b42089a),
	.w6(32'hbab7d942),
	.w7(32'hbbb82f29),
	.w8(32'hbb33d402),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc839735),
	.w1(32'hbb3b85c0),
	.w2(32'hbc390817),
	.w3(32'h3ad970ae),
	.w4(32'h3af801aa),
	.w5(32'h3c4e18d0),
	.w6(32'hbc293a2f),
	.w7(32'hbbef1298),
	.w8(32'hbb92c821),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a11dc),
	.w1(32'h3b484ed1),
	.w2(32'hb914e67d),
	.w3(32'hbbeba99c),
	.w4(32'hbc37e636),
	.w5(32'h3b94a56e),
	.w6(32'hbb3410de),
	.w7(32'hbbc271be),
	.w8(32'h3b8ba48a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b733),
	.w1(32'h3c100313),
	.w2(32'h3c1bed8d),
	.w3(32'hbb23fd67),
	.w4(32'h3bc83528),
	.w5(32'h3bbc5eeb),
	.w6(32'hbadb5404),
	.w7(32'h3bf09c31),
	.w8(32'h3b9e2cb6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d7b24),
	.w1(32'h3b74e832),
	.w2(32'hbb8c3d5c),
	.w3(32'h3c0ccbe0),
	.w4(32'hbb1dc13c),
	.w5(32'hbc170c53),
	.w6(32'h3b1b522c),
	.w7(32'hbbd765a7),
	.w8(32'h3b66a6d6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1343cc),
	.w1(32'hba23e6f3),
	.w2(32'hbaa53b95),
	.w3(32'hb9b66ee7),
	.w4(32'hbb03c748),
	.w5(32'h3b9ec744),
	.w6(32'h3c03bfc2),
	.w7(32'h3b83252c),
	.w8(32'hb9fe1c0e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5b6f),
	.w1(32'hbb88b549),
	.w2(32'hbc110e01),
	.w3(32'h3a380c6b),
	.w4(32'hbb1da205),
	.w5(32'hba88d180),
	.w6(32'h3c2de609),
	.w7(32'hbbfbd169),
	.w8(32'hbbaf881d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c0f8d),
	.w1(32'h3b5ef7c5),
	.w2(32'h3b243578),
	.w3(32'hbc0dc2b8),
	.w4(32'hbb737f6d),
	.w5(32'hbbb49325),
	.w6(32'hbc1f6b45),
	.w7(32'hbb8fead9),
	.w8(32'h3b4900ed),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb673e6a),
	.w1(32'hbbffbecf),
	.w2(32'hbbe9d03d),
	.w3(32'hba84d598),
	.w4(32'h3af30ff3),
	.w5(32'hbbc4887d),
	.w6(32'hbb63b655),
	.w7(32'hbc738190),
	.w8(32'hbb4d4806),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaafc41),
	.w1(32'h3b12fb8a),
	.w2(32'hb9d0408a),
	.w3(32'hbc879985),
	.w4(32'h3afc6e3d),
	.w5(32'hbb25f96c),
	.w6(32'hbbeb9424),
	.w7(32'h3c2774b4),
	.w8(32'h3b269a30),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85fbb4),
	.w1(32'hbb160707),
	.w2(32'hbb586d17),
	.w3(32'hbbbdce80),
	.w4(32'hbb28241f),
	.w5(32'h3c35a9fa),
	.w6(32'h3bcb1d0c),
	.w7(32'h3af03f8c),
	.w8(32'h3ad0f617),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f169),
	.w1(32'h3b1b0928),
	.w2(32'hbb4e8dbe),
	.w3(32'hbbff2976),
	.w4(32'h3ca9cc54),
	.w5(32'h38ac9e2e),
	.w6(32'h3bc508b3),
	.w7(32'h3ba77b67),
	.w8(32'h3aa4d308),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d7c71),
	.w1(32'hbc0b3cff),
	.w2(32'hbba9c916),
	.w3(32'hbc90fbeb),
	.w4(32'hbbb1e635),
	.w5(32'hbc0fe045),
	.w6(32'hbc128cb0),
	.w7(32'h3a0b0c33),
	.w8(32'h3ab812f7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaee312),
	.w1(32'hbb8c8af6),
	.w2(32'hbae2595c),
	.w3(32'h3c0574df),
	.w4(32'h384a21d9),
	.w5(32'h39cb9c0e),
	.w6(32'hbbc78464),
	.w7(32'hbbc7d6f1),
	.w8(32'hbb8d16dc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7c213),
	.w1(32'hbb1a1769),
	.w2(32'hbc378635),
	.w3(32'hbb6284dc),
	.w4(32'hbbc13c64),
	.w5(32'h3b17b6bc),
	.w6(32'h3a791aab),
	.w7(32'h3b7ed38b),
	.w8(32'hbc13ca38),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89eb8),
	.w1(32'hbbc69dcf),
	.w2(32'h3c221631),
	.w3(32'hbac19dd5),
	.w4(32'h3ba06a00),
	.w5(32'hbbf450a9),
	.w6(32'hbc2d7cbd),
	.w7(32'hbb857747),
	.w8(32'hbb79705e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a71bc3),
	.w1(32'hbae965c7),
	.w2(32'hbba7fe08),
	.w3(32'hbab1786c),
	.w4(32'h3c764aa7),
	.w5(32'hbc016aaf),
	.w6(32'h3c0b1db9),
	.w7(32'h3c422f6e),
	.w8(32'h3b82553c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba814393),
	.w1(32'h3bf997bf),
	.w2(32'h3c0cfcdb),
	.w3(32'hbc6025c4),
	.w4(32'hbb8e07d5),
	.w5(32'h3c2ad71c),
	.w6(32'hbb853c0e),
	.w7(32'h3b7d2684),
	.w8(32'hbb65256b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5228b3),
	.w1(32'hbc11d76c),
	.w2(32'hbbc62bba),
	.w3(32'h3a3be001),
	.w4(32'h3c22578a),
	.w5(32'hb9ebbcce),
	.w6(32'h3adbbf06),
	.w7(32'h3b4f6cf9),
	.w8(32'hb9ace390),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4821e),
	.w1(32'h3b037b52),
	.w2(32'hbb3335ae),
	.w3(32'h392db8b9),
	.w4(32'hbc0f6ef3),
	.w5(32'h3c8c3492),
	.w6(32'h3b1ab426),
	.w7(32'h3b70ed8c),
	.w8(32'hbbef4d8a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4949d0),
	.w1(32'hbc0cb1d1),
	.w2(32'h3b4ca887),
	.w3(32'h3c227dcf),
	.w4(32'h3be68d97),
	.w5(32'h3bc97e35),
	.w6(32'h3c646f89),
	.w7(32'hba4665c0),
	.w8(32'hbbab1be3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc1a44),
	.w1(32'hbb79eeb8),
	.w2(32'hbc16a809),
	.w3(32'hba905c59),
	.w4(32'hbb60371a),
	.w5(32'h3c6c341f),
	.w6(32'h3b70fee5),
	.w7(32'h3bb5292c),
	.w8(32'hbbf0cb05),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b462147),
	.w1(32'hbbcebb1e),
	.w2(32'hbbb1e486),
	.w3(32'hbad0e237),
	.w4(32'hbbf01a84),
	.w5(32'h3afdf5e0),
	.w6(32'hbaeee671),
	.w7(32'hbbee6729),
	.w8(32'hbbf793c6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92667f),
	.w1(32'h3adb9348),
	.w2(32'h3b22a03d),
	.w3(32'h3a814a5d),
	.w4(32'hbb1880b9),
	.w5(32'hbc595732),
	.w6(32'h387c9aae),
	.w7(32'hbb433693),
	.w8(32'hbb408ed3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a4d0d),
	.w1(32'hbba69ca1),
	.w2(32'hbc24aefd),
	.w3(32'hb98c685f),
	.w4(32'hbc395030),
	.w5(32'hbc1c569e),
	.w6(32'hbb61a90d),
	.w7(32'hbb532eed),
	.w8(32'hbbc51373),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc414e8b),
	.w1(32'hbba9d74f),
	.w2(32'hbb750887),
	.w3(32'hbb6f5966),
	.w4(32'hbbc8f527),
	.w5(32'h3c88795c),
	.w6(32'hbc27ffde),
	.w7(32'hbb93a8e0),
	.w8(32'hbc206eba),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47f816),
	.w1(32'h3b637896),
	.w2(32'hbb8d2372),
	.w3(32'hba19cd6a),
	.w4(32'h3c1594d5),
	.w5(32'hbbb636e7),
	.w6(32'hbb8af211),
	.w7(32'hbb899c06),
	.w8(32'h3c81f130),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca57c),
	.w1(32'hbb1b6af0),
	.w2(32'hb90a1090),
	.w3(32'h3bebb2bb),
	.w4(32'h3a94eda5),
	.w5(32'h3c383d33),
	.w6(32'hbb61e0d6),
	.w7(32'h3a7979d6),
	.w8(32'hbbf68ca5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb262e2f),
	.w1(32'h3c8d448d),
	.w2(32'hbb0a7a79),
	.w3(32'hbbdb80f5),
	.w4(32'h3cd7e1fd),
	.w5(32'hbbd31737),
	.w6(32'h3b59f05e),
	.w7(32'h3c9dd27e),
	.w8(32'h3baf3a13),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937ede),
	.w1(32'hbb835ff1),
	.w2(32'hba0578fe),
	.w3(32'hbc7b95ca),
	.w4(32'h3bcf2c21),
	.w5(32'hbc161a5b),
	.w6(32'hbc19cc8a),
	.w7(32'hbbcafc0e),
	.w8(32'h3bbf04e6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa558f5),
	.w1(32'hbb1f0805),
	.w2(32'hbb073375),
	.w3(32'hbbe7af2d),
	.w4(32'h3bdfeadb),
	.w5(32'h3a135809),
	.w6(32'hbc07ab95),
	.w7(32'h3bff13b1),
	.w8(32'hbadeb958),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c639),
	.w1(32'hbbd97523),
	.w2(32'hbbe0276d),
	.w3(32'h3a8fad21),
	.w4(32'hbc64cedc),
	.w5(32'h3bab1cd1),
	.w6(32'h3bfc124f),
	.w7(32'hbb980a54),
	.w8(32'hbc0134cb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc051ea2),
	.w1(32'h3b2392d4),
	.w2(32'h39a60af1),
	.w3(32'hbbb24969),
	.w4(32'h3aa06637),
	.w5(32'h3b5df5f4),
	.w6(32'hbaa3b28d),
	.w7(32'h3c0751e9),
	.w8(32'h3b2edb73),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule