module layer_8_featuremap_5(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ee060),
	.w1(32'hba40b2ed),
	.w2(32'h3bbbba31),
	.w3(32'hbc472a05),
	.w4(32'hbaac587d),
	.w5(32'h3bbb205a),
	.w6(32'hbb5a7b9f),
	.w7(32'hbb013131),
	.w8(32'h3bb2fd45),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaa14a),
	.w1(32'h3a49656f),
	.w2(32'hbb453693),
	.w3(32'hbaab6913),
	.w4(32'hba3b465d),
	.w5(32'hbb9968a7),
	.w6(32'hbaa01a0a),
	.w7(32'h3b342e13),
	.w8(32'h39bd00c6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e23ec),
	.w1(32'h3b8ef13a),
	.w2(32'hba885f53),
	.w3(32'hbba90bfd),
	.w4(32'h3b3c3572),
	.w5(32'hbae21527),
	.w6(32'hbaf269cb),
	.w7(32'h3b31a4fd),
	.w8(32'hbb0fa679),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26386d),
	.w1(32'hbaf5c967),
	.w2(32'hbc07ccd6),
	.w3(32'hbb792166),
	.w4(32'hbb5d8178),
	.w5(32'hbc084be8),
	.w6(32'hbb274b12),
	.w7(32'h3b34e45b),
	.w8(32'hbb93bbf3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1406d4),
	.w1(32'hb8aefb07),
	.w2(32'h3aaab153),
	.w3(32'hbc5c6b96),
	.w4(32'h3a96871f),
	.w5(32'h3b620f96),
	.w6(32'hbc1cde26),
	.w7(32'hba16c963),
	.w8(32'h3ae21684),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa3f82),
	.w1(32'h3b25981d),
	.w2(32'h3b71ea31),
	.w3(32'h3b22bcfe),
	.w4(32'h3aef8f32),
	.w5(32'h3a92e6d2),
	.w6(32'h3a95b4b4),
	.w7(32'h3bab4624),
	.w8(32'h3af929c4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb15f0),
	.w1(32'hbad47fae),
	.w2(32'h3b6f4c65),
	.w3(32'h3aacd29b),
	.w4(32'h3af923fb),
	.w5(32'h3c25a264),
	.w6(32'h3af49456),
	.w7(32'hbbdbfa29),
	.w8(32'hba8efa34),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bc37f),
	.w1(32'hbb9a66ab),
	.w2(32'hbb9eaad2),
	.w3(32'h3a932197),
	.w4(32'hbaadeb36),
	.w5(32'hbbe02ee5),
	.w6(32'hbbe26dbc),
	.w7(32'hba86ede7),
	.w8(32'hbb95fec6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc246),
	.w1(32'hbb5c01a3),
	.w2(32'hbc1bb1a6),
	.w3(32'hbb4303da),
	.w4(32'hbc15681d),
	.w5(32'hbc9706af),
	.w6(32'hbb2026bb),
	.w7(32'hbbec055f),
	.w8(32'hbc721d7e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2aeb6),
	.w1(32'hb920dcf1),
	.w2(32'hbae388ec),
	.w3(32'hbc5abb99),
	.w4(32'hbb157edd),
	.w5(32'hbb510c49),
	.w6(32'hbc206d25),
	.w7(32'h3b214469),
	.w8(32'h3b27415b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bd1c),
	.w1(32'h3bc06088),
	.w2(32'h3b855bd2),
	.w3(32'h3ac092da),
	.w4(32'h3bc14740),
	.w5(32'h3bb63aee),
	.w6(32'h3bbb8b4d),
	.w7(32'h3b25c447),
	.w8(32'h3b9f4284),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d93a7),
	.w1(32'h3b6ff59e),
	.w2(32'h3bb2570d),
	.w3(32'h3b3b4dbd),
	.w4(32'h3c0a4613),
	.w5(32'h3b848d81),
	.w6(32'h3b2222d6),
	.w7(32'h3b928c96),
	.w8(32'h3bbe4038),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badda1b),
	.w1(32'h3b14f5c1),
	.w2(32'h3ba23dc3),
	.w3(32'h3ba95363),
	.w4(32'hbb19c5f0),
	.w5(32'h3b380f38),
	.w6(32'h3baca303),
	.w7(32'hbb274fad),
	.w8(32'hbb3c05f9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d650),
	.w1(32'h3c69a489),
	.w2(32'h3c3771f6),
	.w3(32'hbad44521),
	.w4(32'h3c952a8e),
	.w5(32'h3c8dbaf9),
	.w6(32'hbba083ae),
	.w7(32'h3c38fcd9),
	.w8(32'h3c322f2e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd9f7),
	.w1(32'hbc61f907),
	.w2(32'hbc769e84),
	.w3(32'h3c1edded),
	.w4(32'hbc9ae7a7),
	.w5(32'hbcb29700),
	.w6(32'h3bd8e1eb),
	.w7(32'hbc8dfc66),
	.w8(32'hbc905fe7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c3985),
	.w1(32'hba44879d),
	.w2(32'hbaccf27b),
	.w3(32'hbc8a9813),
	.w4(32'h3a2865a9),
	.w5(32'hba5c7b19),
	.w6(32'hbc7f8c26),
	.w7(32'hbaccd380),
	.w8(32'hbac4d891),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1d380),
	.w1(32'h3bf502aa),
	.w2(32'h3c05962e),
	.w3(32'h3938d37e),
	.w4(32'h3ab9af1a),
	.w5(32'hbb5f0ed8),
	.w6(32'hb81abfd9),
	.w7(32'hbb59c586),
	.w8(32'hbbba505c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae575),
	.w1(32'hbb76f2f0),
	.w2(32'hbb2c2395),
	.w3(32'hbba62694),
	.w4(32'hbab8e6dc),
	.w5(32'h3a8e607c),
	.w6(32'hbba34d98),
	.w7(32'hbb86b2c3),
	.w8(32'hbb877773),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e9b14),
	.w1(32'hbb2fba75),
	.w2(32'hbb36eeb8),
	.w3(32'hbb069dad),
	.w4(32'hbaa28e83),
	.w5(32'hbaaca0e7),
	.w6(32'hbbb3a698),
	.w7(32'hbb44b904),
	.w8(32'hba92c15d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6aeb0),
	.w1(32'hbb11e800),
	.w2(32'hbbeef140),
	.w3(32'hbc1b158f),
	.w4(32'hbbfcd86a),
	.w5(32'hbc802637),
	.w6(32'hbba59a5c),
	.w7(32'hbb4a2407),
	.w8(32'hbc210210),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5a07a),
	.w1(32'hbbc57b8c),
	.w2(32'h39a7b0f4),
	.w3(32'hbbd37c08),
	.w4(32'h3bb4e74e),
	.w5(32'h3c86c53f),
	.w6(32'hbb2bdbf4),
	.w7(32'h3b309d78),
	.w8(32'h3c4a0567),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cf31),
	.w1(32'hbb007f43),
	.w2(32'hbb95ceab),
	.w3(32'h3c0b07a1),
	.w4(32'h3aedf750),
	.w5(32'h3ad2d6b2),
	.w6(32'h3b9b758d),
	.w7(32'h3b443de2),
	.w8(32'h3a163fe0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a523a),
	.w1(32'h3ac1ab97),
	.w2(32'h3b79ce2c),
	.w3(32'h3b853391),
	.w4(32'hbbb4b113),
	.w5(32'hbb9a12d2),
	.w6(32'h3b219880),
	.w7(32'hbb22ebe8),
	.w8(32'hbc02af19),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914d05e),
	.w1(32'h3b1440f9),
	.w2(32'h3c58157a),
	.w3(32'hbba49e85),
	.w4(32'h3c675215),
	.w5(32'h3cf7d0f7),
	.w6(32'hbb439790),
	.w7(32'h3c052813),
	.w8(32'h3cbd7008),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be50727),
	.w1(32'h3bdff1eb),
	.w2(32'h3ac5651a),
	.w3(32'h3cb6a7ed),
	.w4(32'h3b9ccca5),
	.w5(32'h3b54afad),
	.w6(32'h3c9117f0),
	.w7(32'h3a3f681e),
	.w8(32'hbb133775),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bea2a),
	.w1(32'hba8ca5b1),
	.w2(32'h3aaa5152),
	.w3(32'h3b8c04c6),
	.w4(32'hba6b7d4f),
	.w5(32'h3875881f),
	.w6(32'h3b4de65b),
	.w7(32'h3b1e7bb0),
	.w8(32'h3b3ca785),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c616d),
	.w1(32'hbbd56e7e),
	.w2(32'hb9e0aee9),
	.w3(32'h3a9b2ce6),
	.w4(32'hbb55a504),
	.w5(32'h3bdedb8e),
	.w6(32'h3a63ce8f),
	.w7(32'hbb52a782),
	.w8(32'h3be07410),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4abf9),
	.w1(32'h3aa5c112),
	.w2(32'h3a36f4d3),
	.w3(32'hbb510e88),
	.w4(32'hbb9d70c1),
	.w5(32'hbb13f4d0),
	.w6(32'hbb8cdacb),
	.w7(32'h3a5b54e9),
	.w8(32'h3a144b62),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421b6e),
	.w1(32'hbc3a6efb),
	.w2(32'hbc5a1680),
	.w3(32'hbbdf4cc9),
	.w4(32'hbc4dd15b),
	.w5(32'hbc92a4af),
	.w6(32'hbb684e97),
	.w7(32'hbc4be372),
	.w8(32'hbc6192a0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc899403),
	.w1(32'hbb61d32a),
	.w2(32'hbb860c08),
	.w3(32'hbc8c9c2b),
	.w4(32'hbb7b9284),
	.w5(32'hbbadb3f5),
	.w6(32'hbc7781e4),
	.w7(32'hbb819aae),
	.w8(32'hbb988c59),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fb29),
	.w1(32'hba3e98bc),
	.w2(32'hbb902695),
	.w3(32'hbb123a74),
	.w4(32'hba4ebeb5),
	.w5(32'hbc041022),
	.w6(32'hbb5d761f),
	.w7(32'hbad027d3),
	.w8(32'hbba35a4c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad3afa),
	.w1(32'h3c273630),
	.w2(32'h3c95a983),
	.w3(32'hbb65edd8),
	.w4(32'h3c837c67),
	.w5(32'h3cc812a4),
	.w6(32'hba3f850b),
	.w7(32'h3c37cd72),
	.w8(32'h3ca30083),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6340c3),
	.w1(32'hbb27195d),
	.w2(32'hbb88c8ee),
	.w3(32'h3ca03df0),
	.w4(32'hbad9b253),
	.w5(32'hbb2f3493),
	.w6(32'h3c683b0c),
	.w7(32'hbbfdcf58),
	.w8(32'hbc15c3e5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53252),
	.w1(32'h3ab7883c),
	.w2(32'hba44c113),
	.w3(32'hbbc9b8c6),
	.w4(32'hbb33cb23),
	.w5(32'hbab1ecb3),
	.w6(32'hbc3437b3),
	.w7(32'h398773d0),
	.w8(32'hbb703ed1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa5c3),
	.w1(32'hbbd0d8cd),
	.w2(32'hbc021f6c),
	.w3(32'hbbd85c24),
	.w4(32'hbbda243e),
	.w5(32'hbc058a03),
	.w6(32'hbbbf9b20),
	.w7(32'hbb9b2f7e),
	.w8(32'hbba19311),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6fd3),
	.w1(32'hbc300b7f),
	.w2(32'hbc3c579a),
	.w3(32'hbbbaa5c2),
	.w4(32'hbc32fbda),
	.w5(32'hbc2678e7),
	.w6(32'hbb760574),
	.w7(32'hbc2fa008),
	.w8(32'hbc2e922c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588925),
	.w1(32'hb93b53d2),
	.w2(32'hbc199205),
	.w3(32'hbc39f1e9),
	.w4(32'hb9a7dc16),
	.w5(32'hbc154632),
	.w6(32'hbc225df9),
	.w7(32'hbb2de812),
	.w8(32'hbbdcb82c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6d6c0),
	.w1(32'hba7ad0ef),
	.w2(32'h38e1e44d),
	.w3(32'hbc169b06),
	.w4(32'h3ac8fb53),
	.w5(32'h39769fe5),
	.w6(32'hbb9ff190),
	.w7(32'hbb86b38a),
	.w8(32'hbae2b1ee),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44a8c0),
	.w1(32'h3be0915b),
	.w2(32'h3c1868e3),
	.w3(32'h3b961dcd),
	.w4(32'h3bc48b66),
	.w5(32'h3b927a85),
	.w6(32'hba299b97),
	.w7(32'h3bad3c7b),
	.w8(32'h3b99b792),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf710),
	.w1(32'h3b897968),
	.w2(32'h3b6c960f),
	.w3(32'h3c117b7a),
	.w4(32'h3b8c82c7),
	.w5(32'h3a417f1a),
	.w6(32'h3bcbfe98),
	.w7(32'h3adc8b90),
	.w8(32'h3aa6b562),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f4464),
	.w1(32'h3a008506),
	.w2(32'h3ba11545),
	.w3(32'h3a412d5b),
	.w4(32'h3b8072e4),
	.w5(32'h3c72e669),
	.w6(32'h39d60c75),
	.w7(32'hba716b72),
	.w8(32'h39fa8722),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b016),
	.w1(32'h3bf2d5ca),
	.w2(32'h3bc93200),
	.w3(32'h3bed6d9a),
	.w4(32'h3c24782e),
	.w5(32'h3c23218e),
	.w6(32'hbaa6bb2c),
	.w7(32'h3c26b2f3),
	.w8(32'h3c51787d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11afb7),
	.w1(32'hbcb3a141),
	.w2(32'hbce31d40),
	.w3(32'h3c479467),
	.w4(32'hbcdbabd2),
	.w5(32'hbd0e7cca),
	.w6(32'h3c6c8e97),
	.w7(32'hbcc973e2),
	.w8(32'hbd00c9e3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccce90),
	.w1(32'h3be4548a),
	.w2(32'h3c02452f),
	.w3(32'hbd011c90),
	.w4(32'h3bd9d604),
	.w5(32'h3bc22dcb),
	.w6(32'hbce94b33),
	.w7(32'h3ba76265),
	.w8(32'h3bbc124f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f2637),
	.w1(32'h3b2c07a1),
	.w2(32'h3b076c39),
	.w3(32'h3bfb9c52),
	.w4(32'hbb1dd608),
	.w5(32'hbbb72953),
	.w6(32'h3bcc6529),
	.w7(32'hbb2a6fca),
	.w8(32'h3bb4b00b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e219a),
	.w1(32'h39ec6203),
	.w2(32'h3b2fbfd1),
	.w3(32'hbb942f00),
	.w4(32'h3b9ef661),
	.w5(32'h3c2dd406),
	.w6(32'h3a9cd0e0),
	.w7(32'hbabe014b),
	.w8(32'h3baed0c8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29d96),
	.w1(32'hbacce943),
	.w2(32'h394c678f),
	.w3(32'h3c012af5),
	.w4(32'hbb311b05),
	.w5(32'hbb9c1f8a),
	.w6(32'h3bdf1294),
	.w7(32'hbb7d36c6),
	.w8(32'hbb932cab),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad087fe),
	.w1(32'h3b506329),
	.w2(32'h39bda0ce),
	.w3(32'h3b24fc25),
	.w4(32'h3be60ff7),
	.w5(32'h3bd30df2),
	.w6(32'h3b02dce8),
	.w7(32'h3c037b31),
	.w8(32'h3b3ab8c4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fe2c8),
	.w1(32'hbbafb54a),
	.w2(32'hbbcb9ef8),
	.w3(32'h3bc5e6e9),
	.w4(32'hbb9c6e81),
	.w5(32'hbbab8f36),
	.w6(32'h3c08ae66),
	.w7(32'hbb999e9b),
	.w8(32'hbbb994d3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2eeeb),
	.w1(32'h3a90bed6),
	.w2(32'h3aa3cc11),
	.w3(32'hbb7e8824),
	.w4(32'hbb4b4b89),
	.w5(32'hbc1945f8),
	.w6(32'hbb8d4b97),
	.w7(32'hbc06a349),
	.w8(32'hbbf32772),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a314),
	.w1(32'h3aa1395f),
	.w2(32'h3be87106),
	.w3(32'hbbf8cfc0),
	.w4(32'h3c23c655),
	.w5(32'h3c986017),
	.w6(32'hbc0c6a75),
	.w7(32'h3c0ce582),
	.w8(32'h3c9414dd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa94c8),
	.w1(32'hbc152b0e),
	.w2(32'hbc14bbfc),
	.w3(32'h3c87706c),
	.w4(32'hbc03e518),
	.w5(32'hbbf8e86a),
	.w6(32'h3c434c3a),
	.w7(32'hbbf14338),
	.w8(32'hbbb93e5e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaf627),
	.w1(32'h3afe109e),
	.w2(32'h3b112c0a),
	.w3(32'hbbcc6ffe),
	.w4(32'h3b85be5c),
	.w5(32'h3b5cd147),
	.w6(32'hbb9029c3),
	.w7(32'hba6459e6),
	.w8(32'h3bbcb055),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d05cb),
	.w1(32'hbc1a3703),
	.w2(32'hbba7c313),
	.w3(32'h3b147301),
	.w4(32'hbbc65798),
	.w5(32'hbbf992d9),
	.w6(32'h3b5df278),
	.w7(32'hbb8a126e),
	.w8(32'hbb836918),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db6c3),
	.w1(32'hba873f06),
	.w2(32'h3ab4ae43),
	.w3(32'hba390b39),
	.w4(32'hbb6d36be),
	.w5(32'h3a372931),
	.w6(32'hbb1796f4),
	.w7(32'hbb7e914c),
	.w8(32'h38d86bfe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32d58c),
	.w1(32'hbbfb4cac),
	.w2(32'hbbd54cc3),
	.w3(32'h3b986969),
	.w4(32'hbbb1f1d8),
	.w5(32'hbb4eafc0),
	.w6(32'h3c125247),
	.w7(32'hbb9c533d),
	.w8(32'hbb1322f2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74420),
	.w1(32'hbc13fe23),
	.w2(32'hbbd16677),
	.w3(32'hbb3845e3),
	.w4(32'hbbcb76a5),
	.w5(32'hbaa633f8),
	.w6(32'hbb32e065),
	.w7(32'hbbbf6aee),
	.w8(32'h3ac4c9c8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd67476),
	.w1(32'h3b707686),
	.w2(32'hba54df63),
	.w3(32'hbb55c99a),
	.w4(32'hbaf97975),
	.w5(32'hba0f44d5),
	.w6(32'hba7b1965),
	.w7(32'hbb7bf38a),
	.w8(32'hbb9d53ef),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89a979),
	.w1(32'hbba6c32f),
	.w2(32'hbc0e32f1),
	.w3(32'hba8dd986),
	.w4(32'hbc202f4f),
	.w5(32'hbc65b9d9),
	.w6(32'hbb5fe65f),
	.w7(32'hbbdce5ad),
	.w8(32'hbc32e842),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd15aa9),
	.w1(32'h3c94653a),
	.w2(32'h3c4c75e1),
	.w3(32'hbc2dadad),
	.w4(32'h3bed8361),
	.w5(32'h3c04768c),
	.w6(32'hbc0563f0),
	.w7(32'h3bed2794),
	.w8(32'h3bd57ff4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2a567),
	.w1(32'hbaa8683c),
	.w2(32'h3a9864a9),
	.w3(32'h3c057092),
	.w4(32'h3972403e),
	.w5(32'h3a65336a),
	.w6(32'h3c5fff54),
	.w7(32'h3a4e5007),
	.w8(32'h3b370225),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ee4c9),
	.w1(32'h3bc7f5df),
	.w2(32'h3b05d032),
	.w3(32'h3b99a794),
	.w4(32'h3b7e191e),
	.w5(32'h3a1af0b7),
	.w6(32'h3bdd5cc6),
	.w7(32'h3c2082bb),
	.w8(32'h3ad75a68),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76322),
	.w1(32'h3ba82339),
	.w2(32'hbbbc5001),
	.w3(32'h3ba4488f),
	.w4(32'hbc2a1403),
	.w5(32'hbcdd2ed9),
	.w6(32'h3c1c8e8b),
	.w7(32'hbbbe0d13),
	.w8(32'hbcb0e225),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af644ce),
	.w1(32'hbbcd4a2b),
	.w2(32'hbc16cccb),
	.w3(32'hbc881846),
	.w4(32'hbc23c261),
	.w5(32'hbc06a54e),
	.w6(32'hbc4c33f9),
	.w7(32'hba8ac26a),
	.w8(32'hbacdfe2f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b3e1),
	.w1(32'hbc1355ca),
	.w2(32'hbc15ae8e),
	.w3(32'hbb86048d),
	.w4(32'hbbce10a2),
	.w5(32'hbbe65321),
	.w6(32'hbb56a9bf),
	.w7(32'hbbf07341),
	.w8(32'hbc12c72e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dbb5a),
	.w1(32'hbc20222f),
	.w2(32'hbc5d862f),
	.w3(32'hbc1be3b4),
	.w4(32'hbc2f5d9e),
	.w5(32'hbc7e372f),
	.w6(32'hbc43261a),
	.w7(32'hbc06246e),
	.w8(32'hbc23432e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54bd5f),
	.w1(32'hbb85298a),
	.w2(32'hbca80821),
	.w3(32'hbc551489),
	.w4(32'hbca024da),
	.w5(32'hbd299c6b),
	.w6(32'hbc0dbed4),
	.w7(32'hbc656195),
	.w8(32'hbd12f37d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71f34),
	.w1(32'hbd09d45b),
	.w2(32'hbd7a537e),
	.w3(32'hbcdeb0e4),
	.w4(32'hbd8c359b),
	.w5(32'hbdd9dee9),
	.w6(32'hbcb7089d),
	.w7(32'hbd4500ea),
	.w8(32'hbda730ef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e2c98),
	.w1(32'h3b39ac46),
	.w2(32'h3a033512),
	.w3(32'hbda08b08),
	.w4(32'h3968a2e4),
	.w5(32'hbabe3923),
	.w6(32'hbd6f1305),
	.w7(32'hba69d70f),
	.w8(32'hbbce4c3c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3118b5),
	.w1(32'hbc6ba90e),
	.w2(32'hbc043ddd),
	.w3(32'hbb87ffb1),
	.w4(32'hbbe2e29a),
	.w5(32'hbc8c82bf),
	.w6(32'hbbfdaf02),
	.w7(32'hbb81a8f4),
	.w8(32'hbb10ea4e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9de60),
	.w1(32'h3b672e81),
	.w2(32'h3aa377a9),
	.w3(32'hbcba2b8e),
	.w4(32'hbb5bfb8f),
	.w5(32'h3b006ccf),
	.w6(32'hba8fdd72),
	.w7(32'hbbe00e51),
	.w8(32'hbbbc7682),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23cc02),
	.w1(32'hbbbb3ca2),
	.w2(32'hbc7fcaaf),
	.w3(32'h3b3eea76),
	.w4(32'hbbd53041),
	.w5(32'hbb3865d7),
	.w6(32'hbb6e3976),
	.w7(32'hbad6cc23),
	.w8(32'hbbf87555),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeec69),
	.w1(32'hbb36ea9f),
	.w2(32'hbba6c755),
	.w3(32'hbbad0e72),
	.w4(32'h3aacd4d8),
	.w5(32'hbafb26f8),
	.w6(32'hbb862e48),
	.w7(32'h3b7df440),
	.w8(32'h3b01f382),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947ff8),
	.w1(32'hbb32f75b),
	.w2(32'hbc83f743),
	.w3(32'hb99ec3ed),
	.w4(32'hbad72c37),
	.w5(32'hbbdc367b),
	.w6(32'h3a772984),
	.w7(32'h3b5c03a3),
	.w8(32'h3bed590d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca558f3),
	.w1(32'hbb772344),
	.w2(32'hbb554222),
	.w3(32'hbb5a6b99),
	.w4(32'hbc10cc15),
	.w5(32'hbc0435c0),
	.w6(32'h3c6957a0),
	.w7(32'h3a2fcec7),
	.w8(32'h3b3f6875),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa1d1a),
	.w1(32'h3c6141de),
	.w2(32'h3a5791d5),
	.w3(32'hbbec3b7c),
	.w4(32'h3c173d83),
	.w5(32'h3b461ad5),
	.w6(32'hbb76bd1d),
	.w7(32'h3b6e6c32),
	.w8(32'h3c6b4e20),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c1417),
	.w1(32'h3b3d813e),
	.w2(32'hbc3602c4),
	.w3(32'h3c3562ab),
	.w4(32'h3a9ad880),
	.w5(32'h3bbfc201),
	.w6(32'h3b9bbd8a),
	.w7(32'hbabdb7cc),
	.w8(32'hb9e13cea),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce972f2),
	.w1(32'h3b97ff75),
	.w2(32'h3bb6acd9),
	.w3(32'h3ce80d46),
	.w4(32'h3b34961b),
	.w5(32'h3ae4d9f8),
	.w6(32'h3b957683),
	.w7(32'hbabb609b),
	.w8(32'h39474466),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd489a3),
	.w1(32'h39105c1f),
	.w2(32'h3a47f2e4),
	.w3(32'hbba3071c),
	.w4(32'hba948bd8),
	.w5(32'h3b50013d),
	.w6(32'hba53a224),
	.w7(32'h3b3eebca),
	.w8(32'h39def127),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122bcb),
	.w1(32'hbb137ab4),
	.w2(32'hb8bf8901),
	.w3(32'h3ba5611d),
	.w4(32'hbc448bcb),
	.w5(32'hbc392392),
	.w6(32'hbb0a6092),
	.w7(32'h3c0b8d65),
	.w8(32'h3ab016fe),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7113),
	.w1(32'h3c94afe6),
	.w2(32'hbc19fce3),
	.w3(32'hbc351931),
	.w4(32'hbbba0643),
	.w5(32'h3c6a44a1),
	.w6(32'h3911564d),
	.w7(32'h3c2b2c4a),
	.w8(32'h3c0a088f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b0cbf),
	.w1(32'h3acc7d0a),
	.w2(32'h3a57c5b2),
	.w3(32'h3cb11c9e),
	.w4(32'h3a5bfc45),
	.w5(32'h3af78915),
	.w6(32'hba06fee5),
	.w7(32'h3b43c053),
	.w8(32'h3a90f61f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fdb4e),
	.w1(32'h3d8025cb),
	.w2(32'h3cb7debb),
	.w3(32'hbae3b6d3),
	.w4(32'hbd88a9fc),
	.w5(32'hbd4c024e),
	.w6(32'hb975a430),
	.w7(32'h3cbff002),
	.w8(32'h3c8bfaa9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc06352),
	.w1(32'hba683313),
	.w2(32'hbbb0d003),
	.w3(32'h3cc48709),
	.w4(32'hbb4f7b95),
	.w5(32'h3acd4753),
	.w6(32'hbc1414b3),
	.w7(32'h3b10f231),
	.w8(32'h3aa6c0b2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922653),
	.w1(32'hbbc37c68),
	.w2(32'h3a589421),
	.w3(32'h3b7317ab),
	.w4(32'h3a2e80f2),
	.w5(32'hbb675c2b),
	.w6(32'hbaef1d9c),
	.w7(32'hbac065d9),
	.w8(32'h3a903ddd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e96fe),
	.w1(32'h3bbade01),
	.w2(32'h3c34e04f),
	.w3(32'hbbf37646),
	.w4(32'h3be1641e),
	.w5(32'h3c7ccb3f),
	.w6(32'h3b22f73c),
	.w7(32'h3b9803d8),
	.w8(32'h3c041c20),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1324b),
	.w1(32'h3c5c2087),
	.w2(32'h3d455d29),
	.w3(32'h3c8d08b2),
	.w4(32'hbc30fadd),
	.w5(32'hbdcece3d),
	.w6(32'hbc69dd0d),
	.w7(32'hbd0b5229),
	.w8(32'h3c3f073f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53c14a),
	.w1(32'h3a881996),
	.w2(32'h3b51668b),
	.w3(32'hbd488257),
	.w4(32'hbac6f20e),
	.w5(32'h3aa90fcc),
	.w6(32'h3cf41f2d),
	.w7(32'hbb690d90),
	.w8(32'hbafd26ec),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02ec48),
	.w1(32'hbb91b6c4),
	.w2(32'h3bba71a9),
	.w3(32'h3ad30c3f),
	.w4(32'hbb7ce75d),
	.w5(32'hbba0577a),
	.w6(32'hba98d8e7),
	.w7(32'hbb892e19),
	.w8(32'hba9300ff),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd02b),
	.w1(32'hbc1f23d0),
	.w2(32'hba8cb83e),
	.w3(32'hbb82d8ae),
	.w4(32'h3a457dc3),
	.w5(32'hbb194689),
	.w6(32'h3a55e38f),
	.w7(32'hbb80b85a),
	.w8(32'h3961d65a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d4fc),
	.w1(32'hbb432e5a),
	.w2(32'h3b6c2271),
	.w3(32'h3b847102),
	.w4(32'hb9d950b9),
	.w5(32'h390bd390),
	.w6(32'h3a1a8a2c),
	.w7(32'h3bf2f961),
	.w8(32'h3c1cdd38),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f13c1),
	.w1(32'h3d0d9752),
	.w2(32'hbbe2603e),
	.w3(32'hbba2139c),
	.w4(32'hbd4d0047),
	.w5(32'h3c834a1f),
	.w6(32'h3b94129e),
	.w7(32'h3c9f83e8),
	.w8(32'h3d23eae8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4de1f),
	.w1(32'h3a84450b),
	.w2(32'h3b2d80c4),
	.w3(32'h3d835b63),
	.w4(32'hbb02e4eb),
	.w5(32'hbb0b04bd),
	.w6(32'hbc12913e),
	.w7(32'hbbf61d0e),
	.w8(32'hbba67274),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053f56),
	.w1(32'hbaa30ac7),
	.w2(32'hbab67774),
	.w3(32'hbb1c0e26),
	.w4(32'hba2f035c),
	.w5(32'h3b1b653a),
	.w6(32'hbb7fd195),
	.w7(32'hbacae752),
	.w8(32'hbaece506),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a411307),
	.w1(32'hbb051312),
	.w2(32'hbcb4989f),
	.w3(32'hbb04cddf),
	.w4(32'hbc31020a),
	.w5(32'hbc1c5cbe),
	.w6(32'hbab8a39a),
	.w7(32'hbba8a6a2),
	.w8(32'hbc1786fc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89136e),
	.w1(32'hba976ac4),
	.w2(32'h3b144f6f),
	.w3(32'hbc83ad73),
	.w4(32'h3c0e9172),
	.w5(32'h3bcc138f),
	.w6(32'hbabfc35e),
	.w7(32'h3b7ebafe),
	.w8(32'h3b74f927),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0683f),
	.w1(32'h3b6f7f9f),
	.w2(32'h387a49a8),
	.w3(32'hbaacc9ee),
	.w4(32'h3a040cea),
	.w5(32'h3b0b4c28),
	.w6(32'h3becd5ee),
	.w7(32'h3a632e31),
	.w8(32'hb96d7fba),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac266a0),
	.w1(32'h3bfc411d),
	.w2(32'h3b50a29c),
	.w3(32'h3a842c59),
	.w4(32'h3bab8d79),
	.w5(32'hbbbf23bd),
	.w6(32'hbaedfac2),
	.w7(32'hbbb8882e),
	.w8(32'hbafaba8b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be15224),
	.w1(32'hb9fd5437),
	.w2(32'hbb014a28),
	.w3(32'hba06eaed),
	.w4(32'hbb016b81),
	.w5(32'hbad157d4),
	.w6(32'h3c52a253),
	.w7(32'hbabf125c),
	.w8(32'hbb2f4ce6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8b375),
	.w1(32'h3b8fb3e7),
	.w2(32'h3bb7eeab),
	.w3(32'hba99077c),
	.w4(32'h3ad95ff3),
	.w5(32'h3ad46cf3),
	.w6(32'hbab4a206),
	.w7(32'h3af4c79d),
	.w8(32'h3a844fd4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19e369),
	.w1(32'h3aa1ab7e),
	.w2(32'h3b811ad8),
	.w3(32'h39eb1fbe),
	.w4(32'h3babf6d0),
	.w5(32'h3cad665e),
	.w6(32'h3b69fd25),
	.w7(32'h3bab01b2),
	.w8(32'h3ad5e2c1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c4d4),
	.w1(32'hbd093644),
	.w2(32'hbcd190c1),
	.w3(32'h3c9bc1de),
	.w4(32'h3c55d415),
	.w5(32'h3c8fde7a),
	.w6(32'hbc0c454c),
	.w7(32'hbc6120d6),
	.w8(32'hbc85ae12),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4f281),
	.w1(32'h3999c639),
	.w2(32'hbc147f54),
	.w3(32'hbc9a70aa),
	.w4(32'h3c4da574),
	.w5(32'h3cf131b1),
	.w6(32'hb8f75643),
	.w7(32'h3c56e303),
	.w8(32'h3c303513),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee5a54),
	.w1(32'hbc3ae2c2),
	.w2(32'hbc45c90b),
	.w3(32'h3c19b6ca),
	.w4(32'hbbed1682),
	.w5(32'hbc25aa27),
	.w6(32'h3bc3cfed),
	.w7(32'hbb9659ef),
	.w8(32'hbbce3aee),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58c998),
	.w1(32'h3b3a6f6c),
	.w2(32'hbbf50e7f),
	.w3(32'hbbe49840),
	.w4(32'h3bf402dc),
	.w5(32'h3be97b56),
	.w6(32'h3a00f46b),
	.w7(32'h3b7fed45),
	.w8(32'h3b737808),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcafee2),
	.w1(32'h3ba3df14),
	.w2(32'h3af28b74),
	.w3(32'h3b20c2cb),
	.w4(32'h381ad475),
	.w5(32'h3905acbb),
	.w6(32'h3bd08bb3),
	.w7(32'h3ad1a555),
	.w8(32'h3ae85721),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8af051),
	.w1(32'h3b84e590),
	.w2(32'h3acd4ec8),
	.w3(32'hba3e550e),
	.w4(32'h3b0cc40b),
	.w5(32'h39c45ad0),
	.w6(32'h39c91e95),
	.w7(32'hba7d8e2f),
	.w8(32'hbaa96b55),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff4a4),
	.w1(32'hbb48c131),
	.w2(32'h3d020cf1),
	.w3(32'h3a9294c3),
	.w4(32'h3d3fb3f8),
	.w5(32'h3cf0f775),
	.w6(32'hba88df31),
	.w7(32'hbb6051cd),
	.w8(32'hbbd9ebac),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7e59a),
	.w1(32'hbb75b906),
	.w2(32'hbc74224d),
	.w3(32'hba487ed5),
	.w4(32'h3bb63f4f),
	.w5(32'h3c333632),
	.w6(32'h3d029619),
	.w7(32'hbb2ad232),
	.w8(32'hbc43376e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b2d2),
	.w1(32'hbbbc2ad9),
	.w2(32'h3bd8f1ac),
	.w3(32'hbba51256),
	.w4(32'h3ba5261a),
	.w5(32'h3bed78cc),
	.w6(32'h3b99dee3),
	.w7(32'h3be3a4d5),
	.w8(32'hbb79a20c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c392ec6),
	.w1(32'hbca15caa),
	.w2(32'hbb876d9c),
	.w3(32'hbbbffbf5),
	.w4(32'hbb824375),
	.w5(32'hbb6769df),
	.w6(32'h3bcc8cd0),
	.w7(32'hbbac7140),
	.w8(32'h3b3d872d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b566fb9),
	.w1(32'h3bd916ee),
	.w2(32'hbbefac0b),
	.w3(32'hbc94254b),
	.w4(32'hbca8b184),
	.w5(32'hbbdd7806),
	.w6(32'h3c43f4e6),
	.w7(32'hbaf4d2fc),
	.w8(32'hbb98aade),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83f61),
	.w1(32'h3b0ce7a7),
	.w2(32'hb9e2d03f),
	.w3(32'hbba3b0c1),
	.w4(32'hbbe26461),
	.w5(32'hbae61d56),
	.w6(32'hbc6c2faf),
	.w7(32'hbae61845),
	.w8(32'hbb1b03b4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55a54d),
	.w1(32'hbbe18f0c),
	.w2(32'hbae10be8),
	.w3(32'h3a37493b),
	.w4(32'hba482234),
	.w5(32'h3b8c2f4b),
	.w6(32'hbb4b6320),
	.w7(32'hbb4d99e3),
	.w8(32'h3aefb0c9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ca2f),
	.w1(32'h3b719800),
	.w2(32'hbb230350),
	.w3(32'hbb8fb446),
	.w4(32'hbbfac2e1),
	.w5(32'hbae9a53b),
	.w6(32'h3aa722d1),
	.w7(32'h3bb1b0d7),
	.w8(32'hbad5e1d6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0436a8),
	.w1(32'h3b662206),
	.w2(32'h3a91db40),
	.w3(32'h3ba5c0fa),
	.w4(32'h3a9643e4),
	.w5(32'h3acfa8b0),
	.w6(32'hbb018816),
	.w7(32'h3b23d79a),
	.w8(32'h3a0b121d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3f0a0),
	.w1(32'h3c4b3d48),
	.w2(32'h3ba771ff),
	.w3(32'h3b5dc3d2),
	.w4(32'hbc695ba2),
	.w5(32'hbc47fb0d),
	.w6(32'hba177a21),
	.w7(32'hbb6e4026),
	.w8(32'h34222e40),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f5f3d),
	.w1(32'h3c24ed64),
	.w2(32'h3d538e2e),
	.w3(32'h3a0e72ae),
	.w4(32'hbc61049c),
	.w5(32'hbd834d2e),
	.w6(32'h39ae0820),
	.w7(32'h3b3a708d),
	.w8(32'h3c89c138),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa42bf),
	.w1(32'h3cba1ef8),
	.w2(32'h3c9b7bcc),
	.w3(32'hbd47db30),
	.w4(32'hbbd46c7b),
	.w5(32'hbc48800d),
	.w6(32'h3cae1a40),
	.w7(32'h3c037230),
	.w8(32'h3c4c7349),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf3ac1),
	.w1(32'h3a68c16a),
	.w2(32'h397e0882),
	.w3(32'hbc15fb89),
	.w4(32'hba45a0c4),
	.w5(32'h3a526ce3),
	.w6(32'h3b62ec4b),
	.w7(32'h39843a54),
	.w8(32'hba48302b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906cae6),
	.w1(32'h3b0b564d),
	.w2(32'h3be12b18),
	.w3(32'hbb022c97),
	.w4(32'hbb4f9e2f),
	.w5(32'hbb07a201),
	.w6(32'hbac743d3),
	.w7(32'h3b011673),
	.w8(32'hbb314340),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980b97f),
	.w1(32'hbb5d45f9),
	.w2(32'hbb7ac92a),
	.w3(32'h3ad82c01),
	.w4(32'hbc234a3c),
	.w5(32'h3ad2f8d8),
	.w6(32'hbb73746a),
	.w7(32'hbb5ee725),
	.w8(32'hb93ba27f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7810d),
	.w1(32'hbadc4d2a),
	.w2(32'h3a668272),
	.w3(32'h3a99bc9e),
	.w4(32'h3b1e0723),
	.w5(32'h3b0cd4e7),
	.w6(32'hbb10f634),
	.w7(32'h3a090643),
	.w8(32'hbb062cb0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d73ae),
	.w1(32'hbbcd21bc),
	.w2(32'hbc880f62),
	.w3(32'hba22dba2),
	.w4(32'hbce90e43),
	.w5(32'hbc9074ca),
	.w6(32'hbb61bd75),
	.w7(32'hbc1ba6c4),
	.w8(32'hbcc33a31),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc529e8),
	.w1(32'hbb9055cd),
	.w2(32'hbbad81f3),
	.w3(32'hbca01c06),
	.w4(32'hb9809ff3),
	.w5(32'hbacdd98d),
	.w6(32'hbc015016),
	.w7(32'h39940c4a),
	.w8(32'h3b8a3df7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7dc50),
	.w1(32'hb954af19),
	.w2(32'hbc130ef9),
	.w3(32'hbc523664),
	.w4(32'h3bc4ef99),
	.w5(32'h3b9c18fa),
	.w6(32'h3c1c10ca),
	.w7(32'h3b4fa798),
	.w8(32'hbb205d97),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7881e),
	.w1(32'hbac00fc2),
	.w2(32'h3a7ba558),
	.w3(32'h3b426a79),
	.w4(32'h3b2c1e71),
	.w5(32'hba975821),
	.w6(32'hba03f75b),
	.w7(32'h3b7893c6),
	.w8(32'h3b2855df),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9785d),
	.w1(32'hbca86673),
	.w2(32'hbd51e680),
	.w3(32'hbb0d7275),
	.w4(32'hbbb40264),
	.w5(32'h3d6bb771),
	.w6(32'h3b165a80),
	.w7(32'h3c6ecd6a),
	.w8(32'hbc89d178),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule