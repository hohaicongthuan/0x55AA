module layer_10_featuremap_384(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10c393),
	.w1(32'hbb243d63),
	.w2(32'h39cc29c3),
	.w3(32'hb97561be),
	.w4(32'hbb93efca),
	.w5(32'h3ab4a223),
	.w6(32'hbbaf8afa),
	.w7(32'hbb49e483),
	.w8(32'h3a8e8e34),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2adbf5),
	.w1(32'hbb288b1f),
	.w2(32'h3b424fe7),
	.w3(32'h3ad12bc7),
	.w4(32'hbb953a79),
	.w5(32'hba4914ce),
	.w6(32'h3b086562),
	.w7(32'hbba734c0),
	.w8(32'hbacad065),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1860a),
	.w1(32'h3bcd4081),
	.w2(32'h3c331c93),
	.w3(32'h3b1f0e38),
	.w4(32'h3c010a17),
	.w5(32'h3c8dc1a6),
	.w6(32'hb9d797a1),
	.w7(32'h3ad5689c),
	.w8(32'h3c8760f2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6442),
	.w1(32'h3ac17892),
	.w2(32'h3a9f60cb),
	.w3(32'h3b8f9c3b),
	.w4(32'hbabe6e4f),
	.w5(32'hbb758599),
	.w6(32'h3c056116),
	.w7(32'hba91fd8a),
	.w8(32'hb9c668d6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea6446),
	.w1(32'hbadc9af7),
	.w2(32'hbab99e02),
	.w3(32'hbc1dcc92),
	.w4(32'hba269b8d),
	.w5(32'hbae42a44),
	.w6(32'hbbd698e5),
	.w7(32'hba367163),
	.w8(32'hbb405c8e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2049),
	.w1(32'hbb45dc81),
	.w2(32'hbb928534),
	.w3(32'hbb13d076),
	.w4(32'hbb6c2d4c),
	.w5(32'hbba18b0f),
	.w6(32'hbaa2d466),
	.w7(32'hbb3b3e6e),
	.w8(32'hb987ad3e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7c954),
	.w1(32'hbc3fc53d),
	.w2(32'hbc2825ae),
	.w3(32'h3849161f),
	.w4(32'hbc3d54df),
	.w5(32'hbc16646c),
	.w6(32'hba1b66d2),
	.w7(32'hbc13f905),
	.w8(32'hbc01ec99),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd4da4),
	.w1(32'h3ac51d7f),
	.w2(32'h3bb8acc7),
	.w3(32'hbc054743),
	.w4(32'hbb0d15c9),
	.w5(32'hbaebab01),
	.w6(32'hbbaf11cc),
	.w7(32'hbb5214a3),
	.w8(32'hbb6d853a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0b04),
	.w1(32'h3c831bc0),
	.w2(32'h3b6db2ec),
	.w3(32'h399f403a),
	.w4(32'h3c3b7fe5),
	.w5(32'h3b93b0e7),
	.w6(32'h3b0e652e),
	.w7(32'h3c2ac0c2),
	.w8(32'hb9f5519b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bfdf2),
	.w1(32'hbb417cf7),
	.w2(32'hbbf4f3b6),
	.w3(32'h3ba5281f),
	.w4(32'hbaa0da89),
	.w5(32'hbba8c79e),
	.w6(32'h3c0752b5),
	.w7(32'hbb28fe8e),
	.w8(32'hbb925bad),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dc940),
	.w1(32'hbc0023be),
	.w2(32'h3b396ac1),
	.w3(32'hbc146e18),
	.w4(32'hbb6a3eba),
	.w5(32'h3b99179e),
	.w6(32'hbbee5148),
	.w7(32'h396ec3d6),
	.w8(32'h39dcd198),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fbfe0),
	.w1(32'hbbd0653e),
	.w2(32'hbb1b15d9),
	.w3(32'h3b53d374),
	.w4(32'hbbfad667),
	.w5(32'hbb99b91f),
	.w6(32'hbb6aa563),
	.w7(32'hbbb837b1),
	.w8(32'hbba10759),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8317),
	.w1(32'hbb67f517),
	.w2(32'h3b94538d),
	.w3(32'h3b4d3894),
	.w4(32'hbb6bb60a),
	.w5(32'h3b89d64a),
	.w6(32'h3a50cbb3),
	.w7(32'hbb042cb4),
	.w8(32'h3ba37b2d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2423d),
	.w1(32'h3a8960ce),
	.w2(32'hbafea8a1),
	.w3(32'h3c30eee7),
	.w4(32'h3ad150ce),
	.w5(32'hbaf0e796),
	.w6(32'h3b9fa8f5),
	.w7(32'h3b581525),
	.w8(32'h3b3e22e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffe1f2),
	.w1(32'hbb6fadbf),
	.w2(32'hbb59612b),
	.w3(32'h3b720b3e),
	.w4(32'hbbe3a411),
	.w5(32'hbac05fe3),
	.w6(32'h3a673664),
	.w7(32'hbbd45623),
	.w8(32'hbbbaffe7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc117c53),
	.w1(32'hbba97e9f),
	.w2(32'hba3e8fcc),
	.w3(32'hbc189b76),
	.w4(32'hbbbbac79),
	.w5(32'hb901898f),
	.w6(32'hbc387ca2),
	.w7(32'hbbaeea08),
	.w8(32'hbb891c71),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa763c7),
	.w1(32'hbb0ee93e),
	.w2(32'hbb1ccfa0),
	.w3(32'hbb26ddb6),
	.w4(32'h39a315fb),
	.w5(32'h38d3b58a),
	.w6(32'hbb36d3b3),
	.w7(32'h3aec1178),
	.w8(32'h3b139214),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fc885),
	.w1(32'hb9973f69),
	.w2(32'h3bbae6b0),
	.w3(32'hbaea3086),
	.w4(32'hba740de4),
	.w5(32'h3c009a79),
	.w6(32'h3aed06d8),
	.w7(32'h3a860d4c),
	.w8(32'h3bc028bb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6cc5),
	.w1(32'h3b229ca1),
	.w2(32'hba75600e),
	.w3(32'h3beb0fa0),
	.w4(32'h3aeba281),
	.w5(32'h3b03a665),
	.w6(32'h3be858a1),
	.w7(32'h3a5fe09c),
	.w8(32'h39e31fb0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49df59),
	.w1(32'hbb816486),
	.w2(32'h3acd6b2a),
	.w3(32'h3b01bf4a),
	.w4(32'hbaf74d45),
	.w5(32'h3a1e6748),
	.w6(32'h3b639de2),
	.w7(32'hbb3b7e91),
	.w8(32'hbb9b7ba1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab42ba6),
	.w1(32'hbbeaf11a),
	.w2(32'hbba026de),
	.w3(32'h3ae9a840),
	.w4(32'hbbce80cc),
	.w5(32'hbbcf4c38),
	.w6(32'hba2a46b4),
	.w7(32'hbbb85db1),
	.w8(32'hbbac0a23),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c4a7),
	.w1(32'hbac82615),
	.w2(32'h3b17e228),
	.w3(32'hbb99d985),
	.w4(32'hbb8c2518),
	.w5(32'hbb156f39),
	.w6(32'hbb659fc6),
	.w7(32'hbb6ec872),
	.w8(32'hbaac0412),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecff64),
	.w1(32'h3ac16720),
	.w2(32'h3b01cfb7),
	.w3(32'h3a361950),
	.w4(32'h3755301a),
	.w5(32'hba86363d),
	.w6(32'h3b257ebd),
	.w7(32'hbb385304),
	.w8(32'hba89eccb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae371d9),
	.w1(32'h3b016ca8),
	.w2(32'hbb4af9af),
	.w3(32'h3b08753f),
	.w4(32'h3bc27aea),
	.w5(32'h3ac2b902),
	.w6(32'hbb25129d),
	.w7(32'h3b7fa985),
	.w8(32'h3b1a694f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47ffe0),
	.w1(32'hba82eaf6),
	.w2(32'h3b94d63a),
	.w3(32'hbc15613f),
	.w4(32'hbb30bc73),
	.w5(32'h3b791be4),
	.w6(32'hbc103c8a),
	.w7(32'hbb8bc474),
	.w8(32'hbac0a9be),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be70e),
	.w1(32'hb9d845e5),
	.w2(32'hbb7350cb),
	.w3(32'hbb0b53c9),
	.w4(32'h3b545490),
	.w5(32'hba903b37),
	.w6(32'hbba7c43d),
	.w7(32'h3b6aea67),
	.w8(32'hb9e5a684),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61ae75),
	.w1(32'hbb0d9719),
	.w2(32'hbb7a5459),
	.w3(32'h3ac292d6),
	.w4(32'hb90a07ea),
	.w5(32'hbbb3357b),
	.w6(32'h3ac66472),
	.w7(32'hbad34f07),
	.w8(32'hbb7325e0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03536),
	.w1(32'hbbab75e8),
	.w2(32'hbab8d552),
	.w3(32'hbb90013a),
	.w4(32'hbb3f68b0),
	.w5(32'h3ba3abd5),
	.w6(32'hbaa356e4),
	.w7(32'hba65ef30),
	.w8(32'h3a221991),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44dc88),
	.w1(32'h39829554),
	.w2(32'h39f9afd8),
	.w3(32'h3b1daea0),
	.w4(32'h3b4e9521),
	.w5(32'hb95bac39),
	.w6(32'h3b33457c),
	.w7(32'hb9bcc015),
	.w8(32'hbaf3e671),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba766245),
	.w1(32'h3a1a4ad1),
	.w2(32'h39e070dd),
	.w3(32'hbb16481e),
	.w4(32'hb98c12f2),
	.w5(32'hbb200346),
	.w6(32'hbbadfbe9),
	.w7(32'hbb17f767),
	.w8(32'hba95f733),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2adcf4),
	.w1(32'hba78b304),
	.w2(32'hbb0c92cf),
	.w3(32'hba697062),
	.w4(32'h3a979a6b),
	.w5(32'h3b0f694b),
	.w6(32'hbb005c8d),
	.w7(32'hbb2254fb),
	.w8(32'hbaae712e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a500),
	.w1(32'h3c1056f5),
	.w2(32'h3c6f2c8d),
	.w3(32'h3aa2b02d),
	.w4(32'h3a82515b),
	.w5(32'h3c21e79c),
	.w6(32'h3aeabc37),
	.w7(32'hba81c210),
	.w8(32'h3bd43a82),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900a21),
	.w1(32'hbb934b03),
	.w2(32'hbb12fbfe),
	.w3(32'hb96272c3),
	.w4(32'hbb3614dd),
	.w5(32'hba7a6bab),
	.w6(32'hba0248a1),
	.w7(32'hbac83077),
	.w8(32'hb9d48f8d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe21021),
	.w1(32'h389eddca),
	.w2(32'hbb863e35),
	.w3(32'hbbc7935e),
	.w4(32'h3a90ffec),
	.w5(32'hba3ed2c0),
	.w6(32'hbab93801),
	.w7(32'hba2b7746),
	.w8(32'hbb44dc72),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9543a8),
	.w1(32'hbbe0a134),
	.w2(32'h3ba88f14),
	.w3(32'hbb52d5f8),
	.w4(32'h38ecb145),
	.w5(32'h3bace705),
	.w6(32'hbb99fa67),
	.w7(32'h3c11502c),
	.w8(32'h3c38054e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ead1c),
	.w1(32'hbb9bb42e),
	.w2(32'hbc0286f8),
	.w3(32'h3c56e4c5),
	.w4(32'hbbcc20d3),
	.w5(32'hbc184f3d),
	.w6(32'h3c155dbc),
	.w7(32'hbb62819c),
	.w8(32'hbb99b35e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bd64c),
	.w1(32'hbc66292b),
	.w2(32'hbbcb4ccf),
	.w3(32'hbb830a7e),
	.w4(32'hbc4c6d89),
	.w5(32'hbbb81306),
	.w6(32'hba7d46b6),
	.w7(32'hbc61e14e),
	.w8(32'hbc2792b4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9add131),
	.w1(32'hbc0b6f8e),
	.w2(32'hbb186c05),
	.w3(32'hbba8d9cc),
	.w4(32'hbc42eddd),
	.w5(32'hbbcad448),
	.w6(32'hbbbee3a6),
	.w7(32'hbc38e944),
	.w8(32'hbbf1ea26),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd002fa),
	.w1(32'hbb505b2c),
	.w2(32'hbb9e8ec6),
	.w3(32'hbbc7642e),
	.w4(32'hbb1448d2),
	.w5(32'hbb391332),
	.w6(32'hbb81825e),
	.w7(32'hbb534f88),
	.w8(32'hbb4efd90),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6101),
	.w1(32'hbb86d03f),
	.w2(32'hbb2f41cc),
	.w3(32'hba7e3b69),
	.w4(32'hbbae5ab0),
	.w5(32'hbbaabbad),
	.w6(32'hb952d9dc),
	.w7(32'hbb2c68a5),
	.w8(32'h3a500924),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39416166),
	.w1(32'h3bc09b42),
	.w2(32'h3b034e23),
	.w3(32'hbbaaa63b),
	.w4(32'h3b6be1fe),
	.w5(32'hbba69a42),
	.w6(32'hbab4cead),
	.w7(32'h3c4e5780),
	.w8(32'h3c33fb14),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bdb36),
	.w1(32'hbaa70ca2),
	.w2(32'h3bdc912a),
	.w3(32'h3c946f24),
	.w4(32'hbb0b1cb2),
	.w5(32'h3bf431b3),
	.w6(32'h3c400350),
	.w7(32'hba53534a),
	.w8(32'h3ae903b1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857568),
	.w1(32'h397e2709),
	.w2(32'h3b83818f),
	.w3(32'h39897269),
	.w4(32'hbb6726f7),
	.w5(32'h3b414512),
	.w6(32'hbc07ba27),
	.w7(32'hbb23bbd3),
	.w8(32'h3a77d426),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523a77),
	.w1(32'hbb12ad70),
	.w2(32'hba4eda88),
	.w3(32'hbb9247c8),
	.w4(32'hbb4e8b77),
	.w5(32'hbb7248d9),
	.w6(32'hbb838ed6),
	.w7(32'hbafbacc4),
	.w8(32'hbaa782c7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf47302),
	.w1(32'h39f6a8e6),
	.w2(32'hb97aeaf3),
	.w3(32'hbbe62db9),
	.w4(32'h3ae18663),
	.w5(32'h3ad142cc),
	.w6(32'hbbafa564),
	.w7(32'h3a1d1cdf),
	.w8(32'h3918546b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d411f),
	.w1(32'hbbc01eb3),
	.w2(32'hbba62d7f),
	.w3(32'hbafeee34),
	.w4(32'hbbe8ad79),
	.w5(32'hbb344dc9),
	.w6(32'hba7d1e38),
	.w7(32'hbb4173b8),
	.w8(32'hbb8ae221),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc93645),
	.w1(32'hbb776459),
	.w2(32'hbc059a60),
	.w3(32'hbc062147),
	.w4(32'hba7c561f),
	.w5(32'hbb2363da),
	.w6(32'hbb9c901a),
	.w7(32'hbb2fac71),
	.w8(32'hbb2cd2f4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f1f07),
	.w1(32'hbb386e9b),
	.w2(32'hbb57815b),
	.w3(32'h38aa7d1a),
	.w4(32'hba309d05),
	.w5(32'hba0dc3b3),
	.w6(32'hbba4be00),
	.w7(32'h3af2a876),
	.w8(32'hba2296f2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ac35),
	.w1(32'h3a33e2ce),
	.w2(32'hbbc1da9a),
	.w3(32'hbb1d6f44),
	.w4(32'h3b5706de),
	.w5(32'hbbe7a3aa),
	.w6(32'hbb5f7cbf),
	.w7(32'h3ba0ae43),
	.w8(32'hbb8d4f2d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb50a4),
	.w1(32'h3b90accb),
	.w2(32'h3bb47b26),
	.w3(32'hba2c007d),
	.w4(32'h3b61ff57),
	.w5(32'h398d5fdb),
	.w6(32'h3b8b0987),
	.w7(32'h39ff9dc8),
	.w8(32'h3bc3dd32),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b017522),
	.w1(32'h3b3656ef),
	.w2(32'hbbd3fa56),
	.w3(32'h3b401a06),
	.w4(32'h3ba3e645),
	.w5(32'hbab73f1b),
	.w6(32'h3bbc0997),
	.w7(32'h3b816fcd),
	.w8(32'hbb05036b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c29e),
	.w1(32'hbb81cd36),
	.w2(32'h3aba144f),
	.w3(32'hb9d7abca),
	.w4(32'hbbc78bd4),
	.w5(32'h3ae6fa51),
	.w6(32'hbab19484),
	.w7(32'hbb98b81b),
	.w8(32'hbac7ebe0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87435),
	.w1(32'h3ad18e19),
	.w2(32'hbae75da4),
	.w3(32'hbad88177),
	.w4(32'h3a95435d),
	.w5(32'hbba9cd6d),
	.w6(32'hbaefae94),
	.w7(32'h3b8ca814),
	.w8(32'hbacc81f9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd265),
	.w1(32'hbb653a21),
	.w2(32'hba10821b),
	.w3(32'hbb6fe574),
	.w4(32'hbb5e8786),
	.w5(32'hbb8080c3),
	.w6(32'hbaab8dd9),
	.w7(32'h3b213f31),
	.w8(32'hbb745cfb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e31a5),
	.w1(32'hbb0b02d0),
	.w2(32'hbbb18935),
	.w3(32'hbbd22139),
	.w4(32'hbba0df85),
	.w5(32'hbbca96dc),
	.w6(32'hbbe5ae39),
	.w7(32'hbb4db68e),
	.w8(32'hbaffcb87),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6191c),
	.w1(32'hbb76a215),
	.w2(32'h3b139d0c),
	.w3(32'hbc133f57),
	.w4(32'hbbb19203),
	.w5(32'h3b5f209d),
	.w6(32'hbb68b523),
	.w7(32'hbb8e5b40),
	.w8(32'h3b1ab76d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd6c3),
	.w1(32'hbabc1f50),
	.w2(32'h395d2bc3),
	.w3(32'h3be2ab1c),
	.w4(32'h3aa2fd54),
	.w5(32'h3b0818f9),
	.w6(32'h3c09aa39),
	.w7(32'hbaa8262c),
	.w8(32'hba9c6997),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad336f0),
	.w1(32'hbaea656b),
	.w2(32'hbb5fcbe8),
	.w3(32'hba97288f),
	.w4(32'hbbb349d7),
	.w5(32'h3b514e1a),
	.w6(32'hbb15c46b),
	.w7(32'hbbe711c0),
	.w8(32'hbb2735f8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292c23),
	.w1(32'hbb07bff4),
	.w2(32'hbb91eaed),
	.w3(32'hbb13731a),
	.w4(32'hbb7a9f33),
	.w5(32'hbb9c0669),
	.w6(32'hbb0c248d),
	.w7(32'hbb6ac477),
	.w8(32'hbba9f31d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17ba4f),
	.w1(32'hba9a68b4),
	.w2(32'hbaa1e670),
	.w3(32'hb91e52ee),
	.w4(32'hbb9a1222),
	.w5(32'hbbabb515),
	.w6(32'hbb20043d),
	.w7(32'hbbe92b4d),
	.w8(32'hbb9bdeea),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a822ba4),
	.w1(32'h3ae40eaa),
	.w2(32'hbb4bf3be),
	.w3(32'hbb3bde9c),
	.w4(32'h3b844952),
	.w5(32'h3b7f78f9),
	.w6(32'hbb4c1c11),
	.w7(32'h3b1f7985),
	.w8(32'h3ab5c8fe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b343f1),
	.w1(32'hbb154aa9),
	.w2(32'h3a85cae9),
	.w3(32'h3af32e88),
	.w4(32'hbb678f06),
	.w5(32'h3a8b9118),
	.w6(32'hba729fef),
	.w7(32'hbb4b9d8e),
	.w8(32'hbb828222),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eafd0),
	.w1(32'h3c525fde),
	.w2(32'h3c9a862c),
	.w3(32'hbb099c17),
	.w4(32'h3c1badbd),
	.w5(32'h3ca16b03),
	.w6(32'hbba2cde1),
	.w7(32'h3c165fce),
	.w8(32'h3c8ec028),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c028034),
	.w1(32'hbac72b3a),
	.w2(32'hbb0a001f),
	.w3(32'h3bcba9df),
	.w4(32'h3a04f00f),
	.w5(32'hba96c58f),
	.w6(32'h3b12bce4),
	.w7(32'hb9b83d98),
	.w8(32'hbb43330a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb6807),
	.w1(32'h3c0afba1),
	.w2(32'h3bc2853a),
	.w3(32'h3b839e7b),
	.w4(32'h3c266bd6),
	.w5(32'h3ba4629c),
	.w6(32'h3b47cd48),
	.w7(32'h3c1d7fdd),
	.w8(32'h3b98c574),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afae1b6),
	.w1(32'hba83816d),
	.w2(32'hbb727c73),
	.w3(32'hbac0a399),
	.w4(32'h3a15091f),
	.w5(32'hbb847bc3),
	.w6(32'h39ff8924),
	.w7(32'hbad29b9f),
	.w8(32'hbbc02349),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ac27),
	.w1(32'hbbcbe49e),
	.w2(32'hbb9e0d31),
	.w3(32'hbba3a2f0),
	.w4(32'hbc4b368e),
	.w5(32'hbbf36f0c),
	.w6(32'hbb972826),
	.w7(32'hbc4228be),
	.w8(32'hbc232b39),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890717e),
	.w1(32'h3c09cd01),
	.w2(32'hb88eb50c),
	.w3(32'h3aec68a1),
	.w4(32'h3bab0d26),
	.w5(32'h3bd8d13e),
	.w6(32'hbb41040a),
	.w7(32'h3a621fd7),
	.w8(32'h39982ebb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1120fa),
	.w1(32'hbb947b5c),
	.w2(32'hbb9b2e94),
	.w3(32'h3c06f189),
	.w4(32'hbbc66784),
	.w5(32'hbb8eca5f),
	.w6(32'h3bd9a4e8),
	.w7(32'hbb666690),
	.w8(32'hbb82665e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c01292),
	.w1(32'hba05cb16),
	.w2(32'hbb9b365f),
	.w3(32'hbb194b0f),
	.w4(32'hbb3d536c),
	.w5(32'hbb406298),
	.w6(32'hbb160581),
	.w7(32'hbb676209),
	.w8(32'hbb779c15),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16ffb),
	.w1(32'hbb3452b0),
	.w2(32'hbba29d34),
	.w3(32'hbb8643bc),
	.w4(32'hbae82d4c),
	.w5(32'hbb09cf77),
	.w6(32'hbb631d7e),
	.w7(32'hba807430),
	.w8(32'h3b112d6a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a8b48),
	.w1(32'h3aa6c9ed),
	.w2(32'h39a7eca8),
	.w3(32'h390a8645),
	.w4(32'hbbfd1106),
	.w5(32'hbc1da063),
	.w6(32'h3b4317b3),
	.w7(32'hbbeb1c2a),
	.w8(32'hbc0180b4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb153d76),
	.w1(32'h3a5cf9d2),
	.w2(32'hba8d66cd),
	.w3(32'hbb463edf),
	.w4(32'h3aceade6),
	.w5(32'hbbd30a1f),
	.w6(32'hbb9a2208),
	.w7(32'h398e6fca),
	.w8(32'hbbb16909),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd93ee),
	.w1(32'hbb1a0e0b),
	.w2(32'hb9639e66),
	.w3(32'h3b629fb7),
	.w4(32'hbb4c614f),
	.w5(32'hbc029d06),
	.w6(32'hbb9abef5),
	.w7(32'h3b73c3c5),
	.w8(32'h3b7fd92d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88b539),
	.w1(32'h3a5acb1c),
	.w2(32'hbb016a4b),
	.w3(32'hbb01261e),
	.w4(32'hb9d30604),
	.w5(32'h398531a4),
	.w6(32'h39bd4ed7),
	.w7(32'hbabb4f56),
	.w8(32'hbb84a92f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d405),
	.w1(32'hbb83196d),
	.w2(32'hbb9477fe),
	.w3(32'h3b75b938),
	.w4(32'h3a8b5d32),
	.w5(32'hbbcee587),
	.w6(32'hbb79a393),
	.w7(32'hbb6440d4),
	.w8(32'h3b00cb13),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86c930),
	.w1(32'hb9b17ded),
	.w2(32'h3b6c0e37),
	.w3(32'hbb6208a2),
	.w4(32'h39b18b64),
	.w5(32'h3b3cbbc8),
	.w6(32'hbb9bcff2),
	.w7(32'h3b1261b5),
	.w8(32'h3b7ba5a7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bba2d),
	.w1(32'h3c4d8302),
	.w2(32'h3c24e9bc),
	.w3(32'hbb908dbe),
	.w4(32'h3b83d4a3),
	.w5(32'h3b5cbf81),
	.w6(32'h3b8f0ce5),
	.w7(32'hbaa0787c),
	.w8(32'hbbe1a039),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf868f),
	.w1(32'h3aba6046),
	.w2(32'hba03687c),
	.w3(32'h3bcad78e),
	.w4(32'hba0eb6c1),
	.w5(32'h3b8648fe),
	.w6(32'hbb9d5fb7),
	.w7(32'h3b80f08f),
	.w8(32'h3a3c69c3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a86da),
	.w1(32'h3a5bc371),
	.w2(32'h3b1f5a70),
	.w3(32'h3b9b3b78),
	.w4(32'h3a3e8366),
	.w5(32'hba255081),
	.w6(32'hbba98f73),
	.w7(32'hbb5d0ba1),
	.w8(32'hba24152b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a600206),
	.w1(32'h3be3bc72),
	.w2(32'h3c116709),
	.w3(32'hbb815c45),
	.w4(32'hbaf44080),
	.w5(32'hbb1231a6),
	.w6(32'h3b250c7a),
	.w7(32'hba1903db),
	.w8(32'hba0c5a5b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8654),
	.w1(32'h3ab1ce7d),
	.w2(32'hbaab80b9),
	.w3(32'hba9c6b4b),
	.w4(32'hbb511a6f),
	.w5(32'hbb8fa796),
	.w6(32'hbb964d46),
	.w7(32'hbb5fda90),
	.w8(32'hbb73ed08),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26661d),
	.w1(32'h3bae935d),
	.w2(32'h3b752bfc),
	.w3(32'hbb9d725c),
	.w4(32'hbabbb9f8),
	.w5(32'hba746046),
	.w6(32'hbb599e9e),
	.w7(32'hbafb60a1),
	.w8(32'hbb8f8904),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba19c74),
	.w1(32'hbb6ba410),
	.w2(32'hbbb2821f),
	.w3(32'hba9824d8),
	.w4(32'hbbf390ab),
	.w5(32'hbc232fbe),
	.w6(32'hbab0c17b),
	.w7(32'hbae22601),
	.w8(32'hbbc37936),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099d0b),
	.w1(32'h3ae1caa2),
	.w2(32'h3b076448),
	.w3(32'hbbc8feb6),
	.w4(32'hbb7bc466),
	.w5(32'hbb0800b0),
	.w6(32'hbc211c66),
	.w7(32'hbbe65dd8),
	.w8(32'hbb9f655d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7030d7),
	.w1(32'hbb4bab05),
	.w2(32'hbb771d4c),
	.w3(32'h3b845ec2),
	.w4(32'hbb5a8fbe),
	.w5(32'hbbef2843),
	.w6(32'hbb2e67db),
	.w7(32'h3b9a23d0),
	.w8(32'hba9fbb07),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaece55),
	.w1(32'h3aa50e7b),
	.w2(32'hb902a564),
	.w3(32'hbbde8194),
	.w4(32'hbb83b439),
	.w5(32'hbb81d106),
	.w6(32'hbaf966a4),
	.w7(32'h3af7f1ad),
	.w8(32'hba816464),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccddea),
	.w1(32'h3a3bc7ac),
	.w2(32'h3ba401aa),
	.w3(32'hbb8befed),
	.w4(32'hbb10f0c0),
	.w5(32'h3bb32c02),
	.w6(32'hbbbd5aef),
	.w7(32'h3b072820),
	.w8(32'hbb8bf0d7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d5e7),
	.w1(32'hbb0834e7),
	.w2(32'hbbac7ef5),
	.w3(32'hba9a2a4d),
	.w4(32'hbbb4c532),
	.w5(32'hbb170641),
	.w6(32'h3761f6b4),
	.w7(32'h3acf9e4f),
	.w8(32'h3a65ca62),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238007),
	.w1(32'hba9965f4),
	.w2(32'h3aba1bd4),
	.w3(32'hbbaa9d81),
	.w4(32'hbb65bda8),
	.w5(32'h39d4fcda),
	.w6(32'hbbc1b1a2),
	.w7(32'hba258ccf),
	.w8(32'hba1c3c89),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9943be9),
	.w1(32'h398a1612),
	.w2(32'hbb8084eb),
	.w3(32'h3b429789),
	.w4(32'h3a55d6d8),
	.w5(32'hbb7f6d35),
	.w6(32'h3ac2c856),
	.w7(32'hbb15bda9),
	.w8(32'hba2f0ca6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08c8c),
	.w1(32'hbb60d0e3),
	.w2(32'hbb1dd27e),
	.w3(32'hbba6c939),
	.w4(32'hbbe83b21),
	.w5(32'hbba2fb15),
	.w6(32'hbb859658),
	.w7(32'hba6505d5),
	.w8(32'hbb283936),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb396b6a),
	.w1(32'hba883372),
	.w2(32'hbac1b249),
	.w3(32'hbbd29388),
	.w4(32'hbb619da9),
	.w5(32'h3b5a43dd),
	.w6(32'h3adf5222),
	.w7(32'hbc044994),
	.w8(32'hbb998ab0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a72a34),
	.w1(32'hbbedc2ef),
	.w2(32'hbc0838a1),
	.w3(32'hbb110e7c),
	.w4(32'h3bfb548f),
	.w5(32'h3bd8e501),
	.w6(32'hbbbdb22f),
	.w7(32'h3c0d7045),
	.w8(32'h3c4250be),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf792bc),
	.w1(32'hbb71a9bc),
	.w2(32'hbbe7d911),
	.w3(32'h3a96eb9e),
	.w4(32'hbc53ba1d),
	.w5(32'hbc4d644f),
	.w6(32'h3bd8a490),
	.w7(32'hbb830dbf),
	.w8(32'hbba30de6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036587),
	.w1(32'hbb195805),
	.w2(32'h3bccb172),
	.w3(32'hbc395fc8),
	.w4(32'hbb2c2138),
	.w5(32'hbbd086ce),
	.w6(32'hbc28d0b7),
	.w7(32'h39e5a7ae),
	.w8(32'hbb6c569d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6bbe7),
	.w1(32'hbb82b5bc),
	.w2(32'hbb42b8fb),
	.w3(32'hbbca9fe8),
	.w4(32'hbbf03a55),
	.w5(32'hbc31447b),
	.w6(32'h3b174880),
	.w7(32'h3abd6c0c),
	.w8(32'hbaca656a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c72e9),
	.w1(32'hbc08a40c),
	.w2(32'hbb42b167),
	.w3(32'hbbf9b1b4),
	.w4(32'hba7b2051),
	.w5(32'hbb2d9d59),
	.w6(32'hbb1a4e40),
	.w7(32'hbbc0e708),
	.w8(32'hbb690434),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab86433),
	.w1(32'h3b42ad90),
	.w2(32'h3bfc3bb4),
	.w3(32'hba7d257a),
	.w4(32'h3c1d9d53),
	.w5(32'h3c773542),
	.w6(32'hba8f7253),
	.w7(32'h3ae7042d),
	.w8(32'h3becf8fe),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec20ec),
	.w1(32'hbbcbeb2a),
	.w2(32'hbbc301e8),
	.w3(32'h3b956ae4),
	.w4(32'hbc46be07),
	.w5(32'hbc4f4f37),
	.w6(32'h3adbabf1),
	.w7(32'hbbd31e54),
	.w8(32'hbb95faab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506781),
	.w1(32'hbb6013b9),
	.w2(32'hbb4a38e7),
	.w3(32'hbc276aa2),
	.w4(32'hba5eb5cb),
	.w5(32'hbb1c1a50),
	.w6(32'hbbaa5ee8),
	.w7(32'h3c1ccf48),
	.w8(32'h3c671677),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2874a),
	.w1(32'h39f27056),
	.w2(32'hba8b31ba),
	.w3(32'hbb18298d),
	.w4(32'hbb87b0e3),
	.w5(32'hbb460bd8),
	.w6(32'h3a8dd2d6),
	.w7(32'hbb9142f6),
	.w8(32'hbbadeed2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fc8d),
	.w1(32'h3ba2e884),
	.w2(32'h3c122b0c),
	.w3(32'hba87374a),
	.w4(32'h3b37b85e),
	.w5(32'h3bbce749),
	.w6(32'h3b02b874),
	.w7(32'h3b0673bf),
	.w8(32'hbbaee996),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fe2ea),
	.w1(32'h3c4b0bc4),
	.w2(32'h3becbe02),
	.w3(32'h3b8ad21c),
	.w4(32'hbb86f0cc),
	.w5(32'hbb5c0dd7),
	.w6(32'h3b9d56e6),
	.w7(32'h3bad725f),
	.w8(32'h3a60e567),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebf810),
	.w1(32'hbb6b3506),
	.w2(32'hbafec08c),
	.w3(32'h3bb02daa),
	.w4(32'hbb9dfba3),
	.w5(32'hbb37b704),
	.w6(32'hbb4a8c4a),
	.w7(32'hbb1d47b9),
	.w8(32'h3b84fc40),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba439d64),
	.w1(32'hbb202ddb),
	.w2(32'hbb46f69c),
	.w3(32'h3b463600),
	.w4(32'hbadf1222),
	.w5(32'hba8a870a),
	.w6(32'h3a1990f4),
	.w7(32'hba6d4c21),
	.w8(32'hbab0f866),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5662b0),
	.w1(32'hbb751ef2),
	.w2(32'hbade674b),
	.w3(32'hbbb5ded9),
	.w4(32'hbc244611),
	.w5(32'hbc0c6fcd),
	.w6(32'hbb65bd7b),
	.w7(32'hbb9077e3),
	.w8(32'h398e4baf),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348a96),
	.w1(32'h38bc60f9),
	.w2(32'hbaed43c5),
	.w3(32'hbba4f4af),
	.w4(32'hbb61d910),
	.w5(32'hbb426ce7),
	.w6(32'h3b8beacd),
	.w7(32'hbb7d701d),
	.w8(32'hbb27d0c6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578edc),
	.w1(32'hb9e40234),
	.w2(32'h3a36a30d),
	.w3(32'hbb7a31a1),
	.w4(32'h3ad20937),
	.w5(32'hbafb01ca),
	.w6(32'hbbc68e12),
	.w7(32'hba523901),
	.w8(32'h3b971362),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b2c9d),
	.w1(32'h3b5e482d),
	.w2(32'hba22c11a),
	.w3(32'hba9dbc68),
	.w4(32'h3c10594b),
	.w5(32'h3b6c328f),
	.w6(32'h3b8814d8),
	.w7(32'hba1d3598),
	.w8(32'h3c0761cc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b937),
	.w1(32'hbba3cc4e),
	.w2(32'hba41948d),
	.w3(32'h3b24e6d5),
	.w4(32'hbbd8ff48),
	.w5(32'hbbb516b7),
	.w6(32'h3c273f41),
	.w7(32'h39b3eecb),
	.w8(32'h3a8c1da1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367654),
	.w1(32'h39fe5b53),
	.w2(32'h3b0dd663),
	.w3(32'hbbcc67d7),
	.w4(32'hbb709055),
	.w5(32'hbc00e862),
	.w6(32'hbb8087a5),
	.w7(32'hbb1d181e),
	.w8(32'hbbb56e7c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c55f82),
	.w1(32'hba3bb714),
	.w2(32'h3ba600eb),
	.w3(32'hbba08d22),
	.w4(32'hbb808934),
	.w5(32'hbaa43baf),
	.w6(32'hbb3bced9),
	.w7(32'hbb8b93ce),
	.w8(32'hbbce9019),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba16e3b),
	.w1(32'h3b6b8344),
	.w2(32'h3c152495),
	.w3(32'hbb1bb882),
	.w4(32'hbbbaa0ab),
	.w5(32'hbc65e12d),
	.w6(32'hbb0d96c2),
	.w7(32'h3be7ddcc),
	.w8(32'h3c958831),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b875515),
	.w1(32'hbbc229c5),
	.w2(32'hbb7b7354),
	.w3(32'h3be25f23),
	.w4(32'hbbb5c046),
	.w5(32'hbb927bae),
	.w6(32'h3bf2dcd6),
	.w7(32'hbaa89930),
	.w8(32'hbad30a79),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b979),
	.w1(32'h3bad5349),
	.w2(32'h3b4cfe02),
	.w3(32'hbb48ec00),
	.w4(32'h39a4e085),
	.w5(32'hbb322cd7),
	.w6(32'hbb505c9c),
	.w7(32'h3b85f453),
	.w8(32'hbac3f8b8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1add2e),
	.w1(32'hba8438e4),
	.w2(32'hb9cef0b0),
	.w3(32'hba743743),
	.w4(32'hbbafdc38),
	.w5(32'hbb74ad8f),
	.w6(32'hbb2de27b),
	.w7(32'hbbb67627),
	.w8(32'h3b453c11),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdf421),
	.w1(32'hbc2a9969),
	.w2(32'hbc4bb643),
	.w3(32'hbbdeb64c),
	.w4(32'hb9071747),
	.w5(32'h3a492ba4),
	.w6(32'h3a313b14),
	.w7(32'hba3e74bd),
	.w8(32'h3adf4f46),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23630d),
	.w1(32'hba949a07),
	.w2(32'h3a88f898),
	.w3(32'hbb6fc0b2),
	.w4(32'h38e1dbdc),
	.w5(32'h3bb137d1),
	.w6(32'hbb989eea),
	.w7(32'h3990638b),
	.w8(32'hbbaa7304),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115003),
	.w1(32'h3b82df43),
	.w2(32'h3baa8b27),
	.w3(32'h3b7415f8),
	.w4(32'h3a7f3918),
	.w5(32'hbbbb2ef9),
	.w6(32'hba8b0b56),
	.w7(32'h3a02631e),
	.w8(32'h3bdcfdac),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085c0e),
	.w1(32'h3ac47251),
	.w2(32'h3b92b7dd),
	.w3(32'hbb3f9d24),
	.w4(32'h3b5cf315),
	.w5(32'h3b13ef18),
	.w6(32'h3c80ec84),
	.w7(32'h3b8ced1b),
	.w8(32'h3b452e0d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be81029),
	.w1(32'hbb0e25a5),
	.w2(32'h3a96627b),
	.w3(32'hbaf1cd2c),
	.w4(32'hb9b85962),
	.w5(32'hb93d5578),
	.w6(32'h3b3144c3),
	.w7(32'hbbc66611),
	.w8(32'h39673161),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b116c),
	.w1(32'hba2f8d50),
	.w2(32'hbafe6b7e),
	.w3(32'hbb828856),
	.w4(32'hbba7260f),
	.w5(32'hbbc9752d),
	.w6(32'hbacecb0e),
	.w7(32'hbb82dedc),
	.w8(32'hbbe18d36),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92802e),
	.w1(32'h3b01a9e8),
	.w2(32'h3ae6becb),
	.w3(32'hbc1a3c90),
	.w4(32'hbb6906b4),
	.w5(32'hbb7996ae),
	.w6(32'hba173184),
	.w7(32'h3a0cb7bc),
	.w8(32'hba410e61),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39183e52),
	.w1(32'h3b0c48dd),
	.w2(32'h3a8f10c1),
	.w3(32'hbbd6ef6e),
	.w4(32'hbb839651),
	.w5(32'hbba38e5f),
	.w6(32'h3a33ca33),
	.w7(32'hbbb85313),
	.w8(32'h3ae32f12),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba5da0),
	.w1(32'hba8c22e4),
	.w2(32'hba3390b7),
	.w3(32'hbbb1a954),
	.w4(32'hba2a745c),
	.w5(32'hba6e4752),
	.w6(32'hbacffa29),
	.w7(32'h3b038adb),
	.w8(32'h3bf83db8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19dc98),
	.w1(32'hbb83d91b),
	.w2(32'hbb0b78b4),
	.w3(32'h3bcbd193),
	.w4(32'hbc10359b),
	.w5(32'hbb94231d),
	.w6(32'hbb5c7d84),
	.w7(32'hb8841f0c),
	.w8(32'h3b47668e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ffba0),
	.w1(32'hbb1b39ac),
	.w2(32'hbb1d77e5),
	.w3(32'hbbccfb2c),
	.w4(32'h3b080689),
	.w5(32'h380ab7f2),
	.w6(32'hbb47c875),
	.w7(32'h3b27e44b),
	.w8(32'hbb98ac9a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f3416),
	.w1(32'h3b7b5a5c),
	.w2(32'h3b5b901a),
	.w3(32'h3ab3e93d),
	.w4(32'h3b42cbc3),
	.w5(32'hba67e321),
	.w6(32'hbb9adeea),
	.w7(32'h3b3d912e),
	.w8(32'h3ace8cde),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c834f),
	.w1(32'h3a25a6fc),
	.w2(32'h3b0fd2cd),
	.w3(32'h3a95e9aa),
	.w4(32'hbaf3731d),
	.w5(32'hbb57e9db),
	.w6(32'hba628d2b),
	.w7(32'h391c199e),
	.w8(32'hbab4fc14),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872b3f),
	.w1(32'hbbd95a51),
	.w2(32'hbbdbb3fd),
	.w3(32'hb9c93984),
	.w4(32'h3bda802a),
	.w5(32'hbc134a40),
	.w6(32'hbb39a69c),
	.w7(32'h3bf066a3),
	.w8(32'h3c9cf0a0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbc86e),
	.w1(32'h3a13504d),
	.w2(32'hbb569270),
	.w3(32'hbbb6f7b0),
	.w4(32'hbadcaacc),
	.w5(32'hbc131a56),
	.w6(32'h3c3eced2),
	.w7(32'hba96f8c8),
	.w8(32'h39723541),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fadb5),
	.w1(32'h3adb3e26),
	.w2(32'hb9ea2980),
	.w3(32'hbb86e780),
	.w4(32'hbabd57e6),
	.w5(32'hbb343ed6),
	.w6(32'hbb9d381a),
	.w7(32'hbb884b0b),
	.w8(32'hba5655b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5fd70),
	.w1(32'h3b039620),
	.w2(32'hbae88b35),
	.w3(32'h39b60276),
	.w4(32'hbb60e241),
	.w5(32'h3aae63a5),
	.w6(32'h3b1bd7b3),
	.w7(32'hbb77b5d8),
	.w8(32'hbb1f86de),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ebc5a),
	.w1(32'hbb14b867),
	.w2(32'h3aead472),
	.w3(32'hbad783c7),
	.w4(32'hb9c73458),
	.w5(32'hba9d05c2),
	.w6(32'hbaa859ec),
	.w7(32'hbb5243b1),
	.w8(32'hbbd03f19),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533ec0),
	.w1(32'hbc2d1165),
	.w2(32'hbc4d892e),
	.w3(32'h3b8d833f),
	.w4(32'h3b99af03),
	.w5(32'h3b409dc7),
	.w6(32'hbb416419),
	.w7(32'h3b423bf5),
	.w8(32'h3bc2e675),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ec50),
	.w1(32'hbad47984),
	.w2(32'hbad2d420),
	.w3(32'hbb8b24dc),
	.w4(32'hbbc7ee0e),
	.w5(32'hbc6c6d11),
	.w6(32'h3aa12b88),
	.w7(32'hbb591b77),
	.w8(32'h3a1741b3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0dd1),
	.w1(32'hbadb07c7),
	.w2(32'hbb4aca85),
	.w3(32'hbb2fbbcf),
	.w4(32'hb900e16f),
	.w5(32'hbaceef9e),
	.w6(32'hbc10b7a5),
	.w7(32'hbaa7a663),
	.w8(32'h3b860ff0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba161f8e),
	.w1(32'h3aba15fd),
	.w2(32'hb9c7d024),
	.w3(32'hba96b636),
	.w4(32'h3b10613e),
	.w5(32'hb9fd3cb9),
	.w6(32'h388804a7),
	.w7(32'hbc12608e),
	.w8(32'hbc06b904),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c7413),
	.w1(32'h3b8c26ca),
	.w2(32'h3b993dd3),
	.w3(32'h3b05c40a),
	.w4(32'h3acab22a),
	.w5(32'h3b431785),
	.w6(32'hbbaf96c6),
	.w7(32'h3af38d01),
	.w8(32'h3b09cbc4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd14434),
	.w1(32'h39e82191),
	.w2(32'h3ba78c6e),
	.w3(32'hbb266301),
	.w4(32'hbc144743),
	.w5(32'hbb3a679c),
	.w6(32'h3ba69e78),
	.w7(32'h3bc7b555),
	.w8(32'h3c0c321a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c2826),
	.w1(32'h3b54b056),
	.w2(32'hbac2e260),
	.w3(32'hb7f52d2a),
	.w4(32'hbabdce3c),
	.w5(32'h3b321112),
	.w6(32'hbbad2f6a),
	.w7(32'hba8dce96),
	.w8(32'hbb9dc6b8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92391e),
	.w1(32'hbb743f11),
	.w2(32'hbbcc0de1),
	.w3(32'h3a638f8e),
	.w4(32'hbb308d6c),
	.w5(32'hbc1fc46d),
	.w6(32'hbb4947f5),
	.w7(32'hbaa68787),
	.w8(32'hbb400045),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37abf7),
	.w1(32'hbb530bf8),
	.w2(32'hbb29da8f),
	.w3(32'hbbba19b6),
	.w4(32'hbc03613c),
	.w5(32'hbc006778),
	.w6(32'h3b92f26b),
	.w7(32'hbb3aea40),
	.w8(32'hbb4e11ce),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c8624),
	.w1(32'h3b7b4ece),
	.w2(32'h3b8a15a1),
	.w3(32'hbc0d24a0),
	.w4(32'h38ccf5c8),
	.w5(32'hbb46f7c5),
	.w6(32'hb894e129),
	.w7(32'hbad19a26),
	.w8(32'hbad8e39d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94eda9),
	.w1(32'h3b1e0240),
	.w2(32'h3af82ecd),
	.w3(32'hb9d60828),
	.w4(32'h3ab08210),
	.w5(32'hba503733),
	.w6(32'hbab8787c),
	.w7(32'h390ff76e),
	.w8(32'hbae0b28c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d221),
	.w1(32'h3b2bd0b2),
	.w2(32'h3b709cd8),
	.w3(32'hb9e36a0a),
	.w4(32'hbbb1e913),
	.w5(32'hbc04dbe3),
	.w6(32'hba988dfb),
	.w7(32'hb88b9a00),
	.w8(32'h3a9cb591),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab35a13),
	.w1(32'h3b8cb54f),
	.w2(32'hbbb97cc3),
	.w3(32'hbbafa09e),
	.w4(32'hbba49b87),
	.w5(32'hbc3e9d7d),
	.w6(32'hbb0e0655),
	.w7(32'hb9a5c27c),
	.w8(32'hbc024612),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8d796),
	.w1(32'hbb5dc440),
	.w2(32'hbb5e4b3c),
	.w3(32'hbbde1b97),
	.w4(32'hbbf34586),
	.w5(32'hbb6c62f6),
	.w6(32'hbbca0466),
	.w7(32'hb9e9ebaa),
	.w8(32'h3ba1f4dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc0b1),
	.w1(32'hbab3e8f5),
	.w2(32'hbb83af04),
	.w3(32'hbbeca276),
	.w4(32'hbad10feb),
	.w5(32'hbaa57920),
	.w6(32'h3b291c17),
	.w7(32'hbb18fc01),
	.w8(32'hbae7e8b7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38922399),
	.w1(32'hb95a29ff),
	.w2(32'hbbb4ada0),
	.w3(32'hba8fb652),
	.w4(32'hbb7d9230),
	.w5(32'hbb509488),
	.w6(32'hbb732dd5),
	.w7(32'hbb6c9921),
	.w8(32'hbac0e2cc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb36b),
	.w1(32'h3becf043),
	.w2(32'h3b99f81e),
	.w3(32'hbb8addd3),
	.w4(32'hbb21f7bc),
	.w5(32'hbba5a0f3),
	.w6(32'hbbed1728),
	.w7(32'h3b12210b),
	.w8(32'h3add1165),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb020c7),
	.w1(32'hbb1278d7),
	.w2(32'hbb23d145),
	.w3(32'hbbad0062),
	.w4(32'hbbe13e04),
	.w5(32'hbbd45ed6),
	.w6(32'h3b1bf029),
	.w7(32'h3b3bde17),
	.w8(32'h3bee05f9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fb6cd),
	.w1(32'h3a9116fb),
	.w2(32'hba40fef2),
	.w3(32'hbb9cadd8),
	.w4(32'hbb235483),
	.w5(32'h3a383e2a),
	.w6(32'h3bd8155a),
	.w7(32'h3a5003d2),
	.w8(32'h3b8bb9e8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b27c8),
	.w1(32'hbb6ef7f7),
	.w2(32'hba27b1b9),
	.w3(32'hbb20f200),
	.w4(32'hbaf10318),
	.w5(32'hbb49aac4),
	.w6(32'h3b549925),
	.w7(32'hbacab6c5),
	.w8(32'hbb42b736),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cf2ba),
	.w1(32'h396fe7bd),
	.w2(32'h3accad59),
	.w3(32'hbb8500c1),
	.w4(32'h3a20e319),
	.w5(32'hb6f92ef0),
	.w6(32'hbb62fc10),
	.w7(32'hbada5fef),
	.w8(32'h3adf679b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a6865),
	.w1(32'hbb624c93),
	.w2(32'hbb306c1a),
	.w3(32'hbb84147a),
	.w4(32'hbb8cccbd),
	.w5(32'hbb9f9dcd),
	.w6(32'h3aa1b570),
	.w7(32'hbb866aef),
	.w8(32'hbb2f3fd3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68fcb3),
	.w1(32'h3b24e0fc),
	.w2(32'h3b503fcb),
	.w3(32'hbac1f06c),
	.w4(32'hba9a384d),
	.w5(32'h3bf07cbc),
	.w6(32'hbaa09a7b),
	.w7(32'hb94ff7ba),
	.w8(32'hb97c8c07),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6171a1),
	.w1(32'hba6d6312),
	.w2(32'hbb5a9325),
	.w3(32'h3b2b7e02),
	.w4(32'h3aefc630),
	.w5(32'h3a5104d6),
	.w6(32'hb9380350),
	.w7(32'hbae4689c),
	.w8(32'hbb3d1e3e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd7708),
	.w1(32'hb8474ee1),
	.w2(32'hba8ea401),
	.w3(32'h3bcda38f),
	.w4(32'h3a3e0e60),
	.w5(32'hbc1ad876),
	.w6(32'hb8e61eb7),
	.w7(32'hbb2d2e97),
	.w8(32'h3a75444e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd8cca),
	.w1(32'hbbba8f26),
	.w2(32'hbb69b579),
	.w3(32'hbb9f22ea),
	.w4(32'hbb51462f),
	.w5(32'hbb8ce5e4),
	.w6(32'h3bec22f4),
	.w7(32'hbb1c956f),
	.w8(32'hbacf6671),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd5ab4),
	.w1(32'h3b9ffadb),
	.w2(32'h3bcdd16d),
	.w3(32'hbbc0403a),
	.w4(32'hbb4f2306),
	.w5(32'hbb9a336a),
	.w6(32'hbb813971),
	.w7(32'hbbab1169),
	.w8(32'hbbbd8f66),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8fe7),
	.w1(32'h3c4ea65e),
	.w2(32'h3b9fbf7b),
	.w3(32'hbb51ce0f),
	.w4(32'h3bd5275b),
	.w5(32'h3c5a47b3),
	.w6(32'hbba3fb16),
	.w7(32'hbbf9c947),
	.w8(32'hbc50a7b5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3451),
	.w1(32'h3a8d59bf),
	.w2(32'h3b1fbce4),
	.w3(32'h3b4723e1),
	.w4(32'hbb5332fe),
	.w5(32'hbb857614),
	.w6(32'hbc0fb8b3),
	.w7(32'hbb1a8e36),
	.w8(32'hbb794e6e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83b31a),
	.w1(32'hbbb56944),
	.w2(32'hbb19aa65),
	.w3(32'hbb6fd10d),
	.w4(32'h39a0f52c),
	.w5(32'hb80cabe4),
	.w6(32'hbb82e514),
	.w7(32'hbbb4f6f0),
	.w8(32'hbbe560dc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17a19),
	.w1(32'hba82a724),
	.w2(32'hbb9e3af4),
	.w3(32'hb997976a),
	.w4(32'hbb1a98c4),
	.w5(32'hbc11ef76),
	.w6(32'hbb1c78fd),
	.w7(32'hbb872342),
	.w8(32'hbbb9541a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce7312),
	.w1(32'hba781498),
	.w2(32'h3aa751f1),
	.w3(32'hb9946b4b),
	.w4(32'hbba147c7),
	.w5(32'hbba1a714),
	.w6(32'hbb184b7c),
	.w7(32'hbbf2a266),
	.w8(32'h3a1789b1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab6938),
	.w1(32'h3b0834ea),
	.w2(32'h3a63971f),
	.w3(32'hbc01d192),
	.w4(32'hbb3c9b43),
	.w5(32'hbb2dc651),
	.w6(32'h3aaae532),
	.w7(32'hb8909002),
	.w8(32'hbb0b0bc9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d7624),
	.w1(32'hbb78726c),
	.w2(32'hbc0c951e),
	.w3(32'hba1662c0),
	.w4(32'hba6e8d37),
	.w5(32'h3c0bf25f),
	.w6(32'hbb787c72),
	.w7(32'hbb646615),
	.w8(32'hbc1acbae),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb304a00),
	.w1(32'hbb34ec40),
	.w2(32'hbb8d267b),
	.w3(32'h3b2128df),
	.w4(32'hbad911fc),
	.w5(32'hbb5d8eaa),
	.w6(32'h39869584),
	.w7(32'hbb6d7b28),
	.w8(32'hbb68ab23),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ffd97),
	.w1(32'hbb2ce918),
	.w2(32'hba3e8729),
	.w3(32'hb98ae92b),
	.w4(32'hbbb510fc),
	.w5(32'hbc04ee5a),
	.w6(32'h3c073c2d),
	.w7(32'h390e1a42),
	.w8(32'hbb25fcd2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81cb17),
	.w1(32'h3a38878c),
	.w2(32'h37117a18),
	.w3(32'hba988b99),
	.w4(32'hbb10f449),
	.w5(32'hbb24307b),
	.w6(32'hbbdda4dc),
	.w7(32'hba1ed2f0),
	.w8(32'h3aac6a4c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0b339),
	.w1(32'h3abe6c6f),
	.w2(32'h3a790eb5),
	.w3(32'hbb04afec),
	.w4(32'hbaa3bf45),
	.w5(32'hbba11d21),
	.w6(32'h381943ec),
	.w7(32'h3917e80a),
	.w8(32'h39c1b62e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6e5f),
	.w1(32'hbb694776),
	.w2(32'hbba0e252),
	.w3(32'h3b6ba89a),
	.w4(32'hbb92a862),
	.w5(32'hbbc36bde),
	.w6(32'h3b683489),
	.w7(32'hbb1415b3),
	.w8(32'hbb52f33f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6f0b6),
	.w1(32'h398bc574),
	.w2(32'h3af156f4),
	.w3(32'hbb70ef6a),
	.w4(32'hba534a2f),
	.w5(32'h3a923cd8),
	.w6(32'h39f6955c),
	.w7(32'h3bb1242f),
	.w8(32'h3c00cd8e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949402),
	.w1(32'hbb79a4da),
	.w2(32'hbb53fac9),
	.w3(32'h3b5979e5),
	.w4(32'hbb629a03),
	.w5(32'hbbe881dc),
	.w6(32'h3b792b74),
	.w7(32'hbb986391),
	.w8(32'hbbbb94c6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965f953),
	.w1(32'hba5f2940),
	.w2(32'hbbc6522d),
	.w3(32'hbb7f500a),
	.w4(32'hbb7140ad),
	.w5(32'h3b17d160),
	.w6(32'hbac377a1),
	.w7(32'hbae3ba16),
	.w8(32'h3a14cb21),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0952d9),
	.w1(32'hbbc2d283),
	.w2(32'hba1dab23),
	.w3(32'hbba5b360),
	.w4(32'hbb1b03f5),
	.w5(32'h3bc45fc7),
	.w6(32'hbc05d51b),
	.w7(32'hbb4bc663),
	.w8(32'h3bd326a0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeed6ae),
	.w1(32'hbb906013),
	.w2(32'hbb32095e),
	.w3(32'hbb9af069),
	.w4(32'hbbcd8f42),
	.w5(32'hbad0f764),
	.w6(32'h3c1a7d34),
	.w7(32'hbba5ebd0),
	.w8(32'h3b98bfc0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9f995),
	.w1(32'hbbaa81da),
	.w2(32'hbbe6db0d),
	.w3(32'hbb6e75c0),
	.w4(32'hbb614040),
	.w5(32'hbbd71524),
	.w6(32'hba1443eb),
	.w7(32'hbb2bd2bd),
	.w8(32'hbba1e19f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab1526),
	.w1(32'h3b5a71d7),
	.w2(32'h3b04a1b3),
	.w3(32'hbbc5e15b),
	.w4(32'hba14d88a),
	.w5(32'h3bd94ea0),
	.w6(32'hba8bbfb4),
	.w7(32'hbb26896e),
	.w8(32'hbbc2a605),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28d256),
	.w1(32'h3b8e8ea0),
	.w2(32'hba5e6857),
	.w3(32'h3a873a58),
	.w4(32'hbaeeb2f1),
	.w5(32'h3b0195f9),
	.w6(32'hbb3f762a),
	.w7(32'hbb9b5c27),
	.w8(32'hbc323f63),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f3186),
	.w1(32'hba2287ab),
	.w2(32'hbb4be95f),
	.w3(32'h3a60ddb6),
	.w4(32'hbbb4a078),
	.w5(32'hbbc62bf2),
	.w6(32'hbbeda156),
	.w7(32'hbb971ba3),
	.w8(32'hbbd01f02),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc80d5),
	.w1(32'h3baf2928),
	.w2(32'h3b78d265),
	.w3(32'hbb147682),
	.w4(32'hbb818298),
	.w5(32'hbb8fa001),
	.w6(32'hbbbfc22c),
	.w7(32'h3ad0eb83),
	.w8(32'hbb98338c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb9fb),
	.w1(32'hba1874db),
	.w2(32'h3a77d9d8),
	.w3(32'h3b58ec9c),
	.w4(32'hbbe9d8af),
	.w5(32'hbb9db264),
	.w6(32'hbbb0da08),
	.w7(32'h3aac16f6),
	.w8(32'h3a497466),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdd322),
	.w1(32'hbb9d0a96),
	.w2(32'hbb658a37),
	.w3(32'h3adbbbed),
	.w4(32'hbaea30e1),
	.w5(32'hbbad9bbf),
	.w6(32'hb7d711a5),
	.w7(32'hbaa6bd86),
	.w8(32'hbbe4a36d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744757),
	.w1(32'hb942cdad),
	.w2(32'hbb1986ff),
	.w3(32'hbbc7a2d9),
	.w4(32'hba89307a),
	.w5(32'hbb644576),
	.w6(32'hbb5c8a56),
	.w7(32'hbb18a8e8),
	.w8(32'hbb672446),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48849b),
	.w1(32'hba28b6a4),
	.w2(32'h3ac2f754),
	.w3(32'hba49ce6e),
	.w4(32'hbb968a8a),
	.w5(32'hbb820e62),
	.w6(32'hbb3d31d5),
	.w7(32'hbb664713),
	.w8(32'hbb85efbd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f3b2),
	.w1(32'hba879665),
	.w2(32'hbaa9d301),
	.w3(32'hbb9da5eb),
	.w4(32'hbbd39334),
	.w5(32'hbb4391b4),
	.w6(32'hbba22041),
	.w7(32'h3b8c9237),
	.w8(32'h3bb947a2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fe2f9),
	.w1(32'hbb825b32),
	.w2(32'hba2a6ec7),
	.w3(32'hbb9ab4e3),
	.w4(32'hba259cce),
	.w5(32'hbbacd3dd),
	.w6(32'h3ab97719),
	.w7(32'hbbaaef8c),
	.w8(32'hb9a2b8a7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e94c9),
	.w1(32'hb7d147d7),
	.w2(32'hbb8077c2),
	.w3(32'hbb2e0ee8),
	.w4(32'hbb98e999),
	.w5(32'hbc568636),
	.w6(32'h3b44ea5f),
	.w7(32'h3a4722d1),
	.w8(32'hbb56e47a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4a59b),
	.w1(32'h3a971b8f),
	.w2(32'h3a4f09b6),
	.w3(32'hbbc0dfd3),
	.w4(32'h3a7fdaf1),
	.w5(32'h3b3d64f1),
	.w6(32'h399811a4),
	.w7(32'h3a0316f7),
	.w8(32'h3b48b282),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c548),
	.w1(32'h3c14146e),
	.w2(32'h3bfc5ebf),
	.w3(32'h39963fa5),
	.w4(32'hbae943ed),
	.w5(32'hbaff8e44),
	.w6(32'h3aa10046),
	.w7(32'h3b1199eb),
	.w8(32'h3b122d7a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd071cf),
	.w1(32'hb7cf0038),
	.w2(32'h3a8ab97c),
	.w3(32'h3ac4e13c),
	.w4(32'hbb5e13a4),
	.w5(32'hbb22f72f),
	.w6(32'hbb22b642),
	.w7(32'hbba58bee),
	.w8(32'hbb701a41),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aad6f),
	.w1(32'h3b1209d4),
	.w2(32'hb91e8c6f),
	.w3(32'hbbb89545),
	.w4(32'h3aadfc79),
	.w5(32'h3b0824f1),
	.w6(32'h3b0d8a4d),
	.w7(32'h3c17b9a6),
	.w8(32'h3c494b3e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc516e),
	.w1(32'h3af611e6),
	.w2(32'h3b88359d),
	.w3(32'h39c1eb64),
	.w4(32'h3aa2ee08),
	.w5(32'h3bee4713),
	.w6(32'h3b356e6f),
	.w7(32'h3b46d1d1),
	.w8(32'h3bf12429),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9ccb),
	.w1(32'hbc0f80e2),
	.w2(32'hbbcd1540),
	.w3(32'h3b845e5d),
	.w4(32'hbb96946d),
	.w5(32'hbc123b42),
	.w6(32'h3b3cd305),
	.w7(32'hbbd57061),
	.w8(32'hbba3ac2f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c084b),
	.w1(32'hba1d0cbe),
	.w2(32'h392a9c7d),
	.w3(32'hbb94f74d),
	.w4(32'hb8cce63e),
	.w5(32'h39fdc9f2),
	.w6(32'hbaf33aea),
	.w7(32'h3a00a8c3),
	.w8(32'h38924bb0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943b70f),
	.w1(32'hba2b51a9),
	.w2(32'hba1ca0a7),
	.w3(32'h39e71ae5),
	.w4(32'hba3238c9),
	.w5(32'hb9c5b497),
	.w6(32'h3a05a8ea),
	.w7(32'hba31d653),
	.w8(32'hba9d2858),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9766036),
	.w1(32'hb9d93b71),
	.w2(32'hb9c6d21a),
	.w3(32'hba398a5a),
	.w4(32'hbaafe7e3),
	.w5(32'hba8819a6),
	.w6(32'hba319ad0),
	.w7(32'h388e2ac5),
	.w8(32'h389eaa64),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a96e22),
	.w1(32'h3a8ddf3a),
	.w2(32'h3a9af2e7),
	.w3(32'hb96ae041),
	.w4(32'h3ae40d98),
	.w5(32'h3ab99e67),
	.w6(32'h3984c290),
	.w7(32'h3b011159),
	.w8(32'h3accc721),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a284a2e),
	.w1(32'h3a6cfb29),
	.w2(32'h3a022531),
	.w3(32'h3a46c59f),
	.w4(32'h398143f4),
	.w5(32'h38f3ddca),
	.w6(32'h3abfab68),
	.w7(32'h388231af),
	.w8(32'h36c00185),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38870037),
	.w1(32'hb88bee17),
	.w2(32'hb87f0380),
	.w3(32'hb82f9790),
	.w4(32'hba301f34),
	.w5(32'h38998f3e),
	.w6(32'hb91d82d7),
	.w7(32'hb90a8744),
	.w8(32'h399001a2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dab11f),
	.w1(32'h3a450d87),
	.w2(32'h3a8e1344),
	.w3(32'hb963e326),
	.w4(32'h38a307ff),
	.w5(32'h3a65e13c),
	.w6(32'h37687566),
	.w7(32'h3898fa91),
	.w8(32'h39940203),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7664f4),
	.w1(32'h3aef82d8),
	.w2(32'h3ab8d26a),
	.w3(32'h39c0e7af),
	.w4(32'h3b2a13f5),
	.w5(32'h3b08bc3c),
	.w6(32'h3a108fbd),
	.w7(32'h3aec472b),
	.w8(32'h3b00aad4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93a45d),
	.w1(32'h3a19db99),
	.w2(32'h39f3f0a8),
	.w3(32'h3ab3ae57),
	.w4(32'hba232961),
	.w5(32'h387531bf),
	.w6(32'h3a7c4d81),
	.w7(32'h39b14735),
	.w8(32'h38aa36fc),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2f251),
	.w1(32'hb9d431aa),
	.w2(32'hb9d9b7ff),
	.w3(32'h39e74091),
	.w4(32'h380805ff),
	.w5(32'h37b49f86),
	.w6(32'h39819b41),
	.w7(32'hb8f6cf40),
	.w8(32'h3a2faaba),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a153fc),
	.w1(32'h3a325cf7),
	.w2(32'hb99cba2f),
	.w3(32'h3a8530e2),
	.w4(32'h395be164),
	.w5(32'h35c25e03),
	.w6(32'h3a820983),
	.w7(32'h39b93c2d),
	.w8(32'hb97059ff),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a0baf),
	.w1(32'h3af68787),
	.w2(32'h3aed5fa9),
	.w3(32'hb9360fe0),
	.w4(32'h3b263711),
	.w5(32'h3ae34bca),
	.w6(32'h3891f550),
	.w7(32'h3ae0d7f9),
	.w8(32'h3b0f9725),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a883e01),
	.w1(32'hb8b53286),
	.w2(32'h39020ffe),
	.w3(32'h3b17e604),
	.w4(32'hb9985d47),
	.w5(32'h38d88b41),
	.w6(32'h3afd0674),
	.w7(32'hb97ae726),
	.w8(32'hb98fe9df),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf831f),
	.w1(32'h385686c4),
	.w2(32'h39aee404),
	.w3(32'h397301cb),
	.w4(32'hb803c30c),
	.w5(32'h398af59a),
	.w6(32'hb9ac8e42),
	.w7(32'h3a0e84a5),
	.w8(32'h3a370cfe),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917d3ee),
	.w1(32'h39b64bc3),
	.w2(32'h3ac69e9d),
	.w3(32'h382b3741),
	.w4(32'hb79b658c),
	.w5(32'h3aad6451),
	.w6(32'h3a42f5e5),
	.w7(32'hb9109ae2),
	.w8(32'h399eebfb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa22eb6),
	.w1(32'hb9dcb366),
	.w2(32'hb9b1c70c),
	.w3(32'h3ab5b8c0),
	.w4(32'hba066813),
	.w5(32'hba1c2575),
	.w6(32'h3a7ce823),
	.w7(32'h3a531553),
	.w8(32'hba08d8db),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be1099),
	.w1(32'hb9c9f830),
	.w2(32'hb97559ef),
	.w3(32'hb9d5ee31),
	.w4(32'hba6fe2aa),
	.w5(32'hba02ce30),
	.w6(32'h38ef9c87),
	.w7(32'hba85c89e),
	.w8(32'hba4aff2b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f988e5),
	.w1(32'hba0b407c),
	.w2(32'hba588db6),
	.w3(32'hb9f7ee9e),
	.w4(32'hbaa12fd8),
	.w5(32'hba070080),
	.w6(32'h38f9c00a),
	.w7(32'hb98b09f8),
	.w8(32'hba91009a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968e71),
	.w1(32'h38fca04c),
	.w2(32'hb92a47f2),
	.w3(32'hb9bfdb4f),
	.w4(32'hba74c9c2),
	.w5(32'hb8abd59b),
	.w6(32'hba98faa5),
	.w7(32'hb9d97679),
	.w8(32'hba229dab),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a48ba8),
	.w1(32'h39007bf8),
	.w2(32'h39a8df2d),
	.w3(32'hba748a0e),
	.w4(32'h3a75c4b7),
	.w5(32'h3adac7ce),
	.w6(32'hbabd2241),
	.w7(32'h39321da1),
	.w8(32'h3ab4d0b3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a009dad),
	.w1(32'hb8ec3082),
	.w2(32'hb95b8316),
	.w3(32'h3a50a17d),
	.w4(32'hb890017c),
	.w5(32'h38b0ad2c),
	.w6(32'h39ae303a),
	.w7(32'hba8772de),
	.w8(32'hb9888469),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39072e39),
	.w1(32'hba954269),
	.w2(32'hba349b4e),
	.w3(32'hba5a0334),
	.w4(32'hba77a4e3),
	.w5(32'hba76270d),
	.w6(32'hba6d15a1),
	.w7(32'hba56cdc9),
	.w8(32'hbad7d006),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2bbf8),
	.w1(32'hba805294),
	.w2(32'hba477b27),
	.w3(32'hba9c739d),
	.w4(32'hbaa70dab),
	.w5(32'hb9ddeee2),
	.w6(32'hba9616fb),
	.w7(32'hba7e4f19),
	.w8(32'hba814220),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98bd53),
	.w1(32'h37dd9002),
	.w2(32'h391b54f2),
	.w3(32'hba972b21),
	.w4(32'hb998acf9),
	.w5(32'h37434b21),
	.w6(32'hb9c524bc),
	.w7(32'h3a004711),
	.w8(32'h3a2338cf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8b276),
	.w1(32'h39cffef9),
	.w2(32'h3a0eceea),
	.w3(32'h3849f7a8),
	.w4(32'h39c28728),
	.w5(32'h3985eaf1),
	.w6(32'h3a97e45d),
	.w7(32'hba443b93),
	.w8(32'hb9cca74b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa398a8),
	.w1(32'hb965afc0),
	.w2(32'h39e8dc80),
	.w3(32'h3a653dd9),
	.w4(32'hba3f8e6d),
	.w5(32'h3920873d),
	.w6(32'h3968ce60),
	.w7(32'hba26887e),
	.w8(32'hba0097f3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3a003),
	.w1(32'h3a40fbd5),
	.w2(32'h3933991b),
	.w3(32'hba310fca),
	.w4(32'h3a101005),
	.w5(32'h3a37532a),
	.w6(32'hb990d3a1),
	.w7(32'h39676934),
	.w8(32'hba3cbe1b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d80f7f),
	.w1(32'hba8223dd),
	.w2(32'hba8d85a6),
	.w3(32'hba61af09),
	.w4(32'hba863839),
	.w5(32'hba761f76),
	.w6(32'hb91ebdd8),
	.w7(32'hba7257b0),
	.w8(32'hba2fdcb3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccee4a),
	.w1(32'hb993431d),
	.w2(32'h3a090c6a),
	.w3(32'hba268370),
	.w4(32'h37ee634f),
	.w5(32'h39ad4ced),
	.w6(32'hb897d3bc),
	.w7(32'hba21f17d),
	.w8(32'hb9d41436),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99f45f),
	.w1(32'hbaa0941a),
	.w2(32'hba326c2e),
	.w3(32'h3a57e68c),
	.w4(32'hba5e300b),
	.w5(32'hb9bfe1df),
	.w6(32'h39b9c593),
	.w7(32'hbaaab919),
	.w8(32'hbafeb45d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba806050),
	.w1(32'hba74f687),
	.w2(32'hba2a8e68),
	.w3(32'hbaaf93e8),
	.w4(32'hba77a16d),
	.w5(32'hb9cca10d),
	.w6(32'hbb0c0d28),
	.w7(32'hb9ebcfaa),
	.w8(32'hba24c59c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b1df4),
	.w1(32'h384c03fe),
	.w2(32'h392a6967),
	.w3(32'hba828b70),
	.w4(32'hba23b9eb),
	.w5(32'h38cc764f),
	.w6(32'hba39c2e0),
	.w7(32'hb9f20e36),
	.w8(32'hba2c632f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc8b96),
	.w1(32'hb9ab8432),
	.w2(32'h392758a2),
	.w3(32'hb94e27ec),
	.w4(32'hba72dc27),
	.w5(32'hb9345477),
	.w6(32'hba8f39fc),
	.w7(32'hba70bd8e),
	.w8(32'hba752691),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcac32),
	.w1(32'h3a22a6b2),
	.w2(32'hb8a060f8),
	.w3(32'hb97ce286),
	.w4(32'hb9786ea3),
	.w5(32'h38887bb5),
	.w6(32'h396ca69d),
	.w7(32'hb9ad268b),
	.w8(32'hba55205f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0af84),
	.w1(32'hb9c78165),
	.w2(32'hbab3b7c5),
	.w3(32'hbb05adb9),
	.w4(32'hb9fa6886),
	.w5(32'hbaa52d5e),
	.w6(32'hba95476f),
	.w7(32'hb9b043f7),
	.w8(32'hbac55c04),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c33d8),
	.w1(32'hb93e1d8d),
	.w2(32'hb927ad9e),
	.w3(32'hba42f35f),
	.w4(32'hba92a742),
	.w5(32'hba139500),
	.w6(32'hba2dba36),
	.w7(32'hb83ac815),
	.w8(32'h396413c6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a24089),
	.w1(32'hb992da76),
	.w2(32'h37f1a3fd),
	.w3(32'hba899330),
	.w4(32'hb8bc1e0b),
	.w5(32'hb9055db4),
	.w6(32'hb9b112aa),
	.w7(32'h39952f5b),
	.w8(32'h3921acb8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec9341),
	.w1(32'h3a5bf3e5),
	.w2(32'h39e5c95c),
	.w3(32'h38a73d8f),
	.w4(32'h3a8ea303),
	.w5(32'h3a284dd7),
	.w6(32'h3a55a735),
	.w7(32'h3a1f3638),
	.w8(32'h3a2ca4b2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f480eb),
	.w1(32'hba936eb1),
	.w2(32'hba3be799),
	.w3(32'h3a594745),
	.w4(32'hba5ad93f),
	.w5(32'hba710276),
	.w6(32'h399c937a),
	.w7(32'hb937463b),
	.w8(32'hb9effe6e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e68b),
	.w1(32'hba5af3aa),
	.w2(32'hba1254fd),
	.w3(32'hba17e41a),
	.w4(32'hbaaa3f88),
	.w5(32'hba87c2b0),
	.w6(32'hb95f7d22),
	.w7(32'hba6fd463),
	.w8(32'hba5fad6c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9852526),
	.w1(32'hb9ce4770),
	.w2(32'h39781d94),
	.w3(32'hbaae5cc7),
	.w4(32'hbabc50be),
	.w5(32'hb92761d4),
	.w6(32'hba945bb0),
	.w7(32'h39ea1320),
	.w8(32'hba14eeaa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8496510),
	.w1(32'hba628e9d),
	.w2(32'hb8b2dc90),
	.w3(32'hba4f1c10),
	.w4(32'h390c155d),
	.w5(32'hb8b6f15f),
	.w6(32'h389fd087),
	.w7(32'hb93011e6),
	.w8(32'hb9e63791),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f84471),
	.w1(32'hb9db4461),
	.w2(32'h3a3823de),
	.w3(32'h3a1c0947),
	.w4(32'hb996a690),
	.w5(32'h3a3b04fb),
	.w6(32'hb9a98ace),
	.w7(32'hba193e5c),
	.w8(32'hb9668936),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ae5c),
	.w1(32'h3a278a68),
	.w2(32'h392c475f),
	.w3(32'h38a93abf),
	.w4(32'h3a712a9a),
	.w5(32'h39cbe358),
	.w6(32'h3923a68e),
	.w7(32'h3a458bf2),
	.w8(32'h398acc86),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c8412),
	.w1(32'hb9b1c686),
	.w2(32'hbacf3d3c),
	.w3(32'hba0b46e9),
	.w4(32'hb9824cf5),
	.w5(32'hba2d9518),
	.w6(32'hb5f22e14),
	.w7(32'hbac2a912),
	.w8(32'h3a542f66),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba186b63),
	.w1(32'hb907ea36),
	.w2(32'hb9becc46),
	.w3(32'h38acae6a),
	.w4(32'hb6f1bb4e),
	.w5(32'hb9c23bdf),
	.w6(32'h3a34dd76),
	.w7(32'hb920ae26),
	.w8(32'hba4293b8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98805d5),
	.w1(32'h3984103e),
	.w2(32'h396a7f53),
	.w3(32'h39a6f2ce),
	.w4(32'h39ce2c2a),
	.w5(32'h3a575434),
	.w6(32'h39ae4989),
	.w7(32'h3a0ccce9),
	.w8(32'h3a171f94),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a560bf2),
	.w1(32'hb95afa93),
	.w2(32'h3a3f9229),
	.w3(32'h3a37b1a5),
	.w4(32'hb997eb99),
	.w5(32'h3a5f3738),
	.w6(32'h3aa4fc98),
	.w7(32'h3a21f4f3),
	.w8(32'hb78e5bec),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39719d0b),
	.w1(32'h3a0bb81c),
	.w2(32'h395dde73),
	.w3(32'h39b664ce),
	.w4(32'h39e01655),
	.w5(32'h398da0ec),
	.w6(32'h3a357e4b),
	.w7(32'hb9ac1ab6),
	.w8(32'h39ca952a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e99c0),
	.w1(32'h3757cb09),
	.w2(32'hb99ed590),
	.w3(32'h3a8c8b42),
	.w4(32'hba43aa4a),
	.w5(32'hba3f8ae0),
	.w6(32'h3a2e6aa5),
	.w7(32'hb9301f36),
	.w8(32'h38a193c3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bac19),
	.w1(32'hba3df3bb),
	.w2(32'hbabadf97),
	.w3(32'hba148ee5),
	.w4(32'hbac3ebcf),
	.w5(32'hbab7b331),
	.w6(32'hb9a9b5fd),
	.w7(32'hbadaefec),
	.w8(32'hbb024e04),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeef61d),
	.w1(32'h3ab47bbf),
	.w2(32'h3ab82256),
	.w3(32'hbab05cd7),
	.w4(32'h3b02aaa1),
	.w5(32'h3aee6b5e),
	.w6(32'hbac2ff6a),
	.w7(32'h3ac001b7),
	.w8(32'h3ad327f1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5444f3),
	.w1(32'hb945ff73),
	.w2(32'h39953c2e),
	.w3(32'h3ad2d7eb),
	.w4(32'hb94cf6a2),
	.w5(32'h38d70d78),
	.w6(32'h3a5b720f),
	.w7(32'hb9d9a5a0),
	.w8(32'h39d4b35b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9a0ae),
	.w1(32'hb997a31b),
	.w2(32'h38f38abe),
	.w3(32'hb99ae4a3),
	.w4(32'hb9679a8e),
	.w5(32'h3a0253f3),
	.w6(32'hb9c5a2cc),
	.w7(32'hb9faf054),
	.w8(32'hba0ad8dc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa9510),
	.w1(32'hbaa1b28b),
	.w2(32'hba58d36f),
	.w3(32'hba344096),
	.w4(32'hba86f431),
	.w5(32'hba255756),
	.w6(32'hba0f5681),
	.w7(32'hba621cb8),
	.w8(32'hba429756),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d79a2a),
	.w1(32'hb9a06da7),
	.w2(32'h398cbc8f),
	.w3(32'hba507c69),
	.w4(32'hbaa49c86),
	.w5(32'h392b4d55),
	.w6(32'hba324126),
	.w7(32'hb93a58d0),
	.w8(32'hb9ae800c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc8fe9),
	.w1(32'h352e3709),
	.w2(32'hb9f39fc7),
	.w3(32'hb9d7a1d2),
	.w4(32'hba2f5491),
	.w5(32'hba91431c),
	.w6(32'hb975d287),
	.w7(32'hb9bbd93f),
	.w8(32'hb97fb166),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391723ad),
	.w1(32'hba8a79fa),
	.w2(32'hba51d414),
	.w3(32'hba627c78),
	.w4(32'hbac326f9),
	.w5(32'hb9f99eac),
	.w6(32'hb9335fd9),
	.w7(32'hba5e51b7),
	.w8(32'hbaa90d3d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba136048),
	.w1(32'h39a4fc8a),
	.w2(32'h3985c834),
	.w3(32'hbac7d70b),
	.w4(32'h399793db),
	.w5(32'h39b7c7d1),
	.w6(32'hba9e1021),
	.w7(32'h36273966),
	.w8(32'h3a279761),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule