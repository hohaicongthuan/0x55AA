module layer_10_featuremap_39(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83c2e5),
	.w1(32'hbc0a2452),
	.w2(32'hbadfa007),
	.w3(32'hbc84b8ef),
	.w4(32'hbc132430),
	.w5(32'hbb56aaa2),
	.w6(32'hbc6ef4df),
	.w7(32'hba402649),
	.w8(32'hbbf90396),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5caaa),
	.w1(32'h3bcccdf6),
	.w2(32'hb9963966),
	.w3(32'hbc17c9e4),
	.w4(32'h3b5496fe),
	.w5(32'h389092f8),
	.w6(32'hbc405f9f),
	.w7(32'hbb8c4c15),
	.w8(32'h3c051f78),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd590c),
	.w1(32'hbcbb17e6),
	.w2(32'hbc1ed29f),
	.w3(32'hbc492f88),
	.w4(32'hbc866318),
	.w5(32'hbc16f1ce),
	.w6(32'hbcfb772c),
	.w7(32'hbbd6a253),
	.w8(32'hbc747b21),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb73d),
	.w1(32'hbaec3250),
	.w2(32'h3b46d49b),
	.w3(32'hbc0f02c8),
	.w4(32'hbc72e873),
	.w5(32'h3ad3b633),
	.w6(32'hbabcd38e),
	.w7(32'hbc0be249),
	.w8(32'h3a5006ca),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9852a4),
	.w1(32'h3c523e7e),
	.w2(32'hbb58db82),
	.w3(32'hbb2992f1),
	.w4(32'h3a0238df),
	.w5(32'hb9e87237),
	.w6(32'h3bc488d8),
	.w7(32'h3ab30850),
	.w8(32'h3ca52b51),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d005bf1),
	.w1(32'h3b89aecd),
	.w2(32'h3bd04a03),
	.w3(32'h3d8bb49b),
	.w4(32'h3b958493),
	.w5(32'h3be61440),
	.w6(32'h3d77f296),
	.w7(32'hbbb79b6b),
	.w8(32'h3b503d57),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c2698),
	.w1(32'hbacda4c7),
	.w2(32'hba305d62),
	.w3(32'h3b78c153),
	.w4(32'hbbc34441),
	.w5(32'hba61e7f9),
	.w6(32'hba800b6d),
	.w7(32'hbc2cd43f),
	.w8(32'hbb2b0958),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec2ddb),
	.w1(32'h3b151579),
	.w2(32'h3b8868fe),
	.w3(32'hbc1a9e3e),
	.w4(32'h3995c582),
	.w5(32'h3b8bc763),
	.w6(32'hbb0c6dad),
	.w7(32'h3a032e55),
	.w8(32'h3be1d7bc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa566e6),
	.w1(32'hbbb3599b),
	.w2(32'hbb97559a),
	.w3(32'h3a2f771f),
	.w4(32'hbbaa53bb),
	.w5(32'hbb61dd72),
	.w6(32'hbaa72030),
	.w7(32'hbad1fec9),
	.w8(32'hbb400491),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16b285),
	.w1(32'hbbc9757d),
	.w2(32'h3a55fd21),
	.w3(32'hbc0ef7e6),
	.w4(32'hbb309179),
	.w5(32'h3b73d34a),
	.w6(32'h3a20ecd8),
	.w7(32'h3b683d96),
	.w8(32'h3b8382cb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39449757),
	.w1(32'hbb8fe73d),
	.w2(32'hbbd7cd5b),
	.w3(32'h3a4f2270),
	.w4(32'hbb67a5b2),
	.w5(32'hbc7af81b),
	.w6(32'h3a3b2ec4),
	.w7(32'hba180fce),
	.w8(32'hbc17b723),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82767e),
	.w1(32'hba85948e),
	.w2(32'hbb9db2a4),
	.w3(32'hbb97a129),
	.w4(32'hbbb35f64),
	.w5(32'hbba1e10a),
	.w6(32'h3c342b06),
	.w7(32'hbb68bdab),
	.w8(32'hbb92c619),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976e05),
	.w1(32'hbb2f4ccc),
	.w2(32'hbb550b9a),
	.w3(32'hbb27cbca),
	.w4(32'hbac16179),
	.w5(32'hb97c14c0),
	.w6(32'hbb0d0b92),
	.w7(32'hba58b32b),
	.w8(32'h39554e75),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15cfba),
	.w1(32'h3a212619),
	.w2(32'h3b92dd09),
	.w3(32'hbbbe778f),
	.w4(32'h3b7b81a5),
	.w5(32'h3b727328),
	.w6(32'hbbe565bd),
	.w7(32'hb6be4833),
	.w8(32'h3b8c34a8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4ed15),
	.w1(32'hbbb2497c),
	.w2(32'h3a985138),
	.w3(32'h3b20bd76),
	.w4(32'hbc495914),
	.w5(32'h3922001f),
	.w6(32'hbbc866e2),
	.w7(32'hbba9df67),
	.w8(32'h3bf82518),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31444e),
	.w1(32'hbb4f8b43),
	.w2(32'h3b2005c8),
	.w3(32'h3b375565),
	.w4(32'hbbfbbf05),
	.w5(32'h3badcfb2),
	.w6(32'h3b14c393),
	.w7(32'hbbba5bbb),
	.w8(32'h3bb147da),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cb7a5),
	.w1(32'hbba035dd),
	.w2(32'hbbb82fc6),
	.w3(32'h3a06b56c),
	.w4(32'hbb25e791),
	.w5(32'hbb972674),
	.w6(32'hba6dbf88),
	.w7(32'hbaa48ba6),
	.w8(32'hb5cbc1bf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29969),
	.w1(32'hbba1504d),
	.w2(32'h3b8c617b),
	.w3(32'hbbf24115),
	.w4(32'hbb6ea76b),
	.w5(32'h3bce94b6),
	.w6(32'h38f07d66),
	.w7(32'h3bb0b9a3),
	.w8(32'h3a72b43e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dbecc),
	.w1(32'hbba6ce0d),
	.w2(32'hbbd15d6f),
	.w3(32'hbaa46dfe),
	.w4(32'hbbde017b),
	.w5(32'hbbcb53b8),
	.w6(32'hbba90bfe),
	.w7(32'hbb48aac2),
	.w8(32'hbaf3d04b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037344),
	.w1(32'h39c6035a),
	.w2(32'hbb3c7465),
	.w3(32'h3b020f76),
	.w4(32'hbc9a7251),
	.w5(32'hbc00b0f7),
	.w6(32'hbb9e428a),
	.w7(32'hbba08e44),
	.w8(32'hbc4933fc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15cf16),
	.w1(32'h3b19f561),
	.w2(32'h3c12c84c),
	.w3(32'h3b58f802),
	.w4(32'h3b194f96),
	.w5(32'h3c0ec631),
	.w6(32'h3bdf2f47),
	.w7(32'hb8e04d64),
	.w8(32'h3bf3450d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d287a),
	.w1(32'h3bc48a8f),
	.w2(32'hb9c8fd68),
	.w3(32'h3c611003),
	.w4(32'hbc253948),
	.w5(32'h3b31c1bb),
	.w6(32'h3bd166ee),
	.w7(32'hbb2f2aae),
	.w8(32'h3bdcb62e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf414b),
	.w1(32'hbbe45b40),
	.w2(32'h3b3f4220),
	.w3(32'h3c22d7e9),
	.w4(32'hbc5f16ec),
	.w5(32'h3b668b79),
	.w6(32'hbb0d7c40),
	.w7(32'hbc172d28),
	.w8(32'h3b8226f9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d36fc),
	.w1(32'h3979e4e8),
	.w2(32'h3b6b6719),
	.w3(32'h3b1ef616),
	.w4(32'hbaaf3da9),
	.w5(32'h3a50267e),
	.w6(32'h3b2479e0),
	.w7(32'hba55b837),
	.w8(32'h3b1413c4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd985b5),
	.w1(32'hbb5a07ac),
	.w2(32'hbb512154),
	.w3(32'hbb8ccc35),
	.w4(32'h3ac6fe45),
	.w5(32'h3b23ef6a),
	.w6(32'hbbee8e8c),
	.w7(32'hba576443),
	.w8(32'h3c5943ae),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8d49a),
	.w1(32'hbb8234f5),
	.w2(32'h3a91b90c),
	.w3(32'h3cb92ed8),
	.w4(32'hbbc7a3ce),
	.w5(32'h3b945ade),
	.w6(32'h3c87b98f),
	.w7(32'hba09972e),
	.w8(32'h3a65fbdd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aced8dc),
	.w1(32'hbbdc9930),
	.w2(32'h39530997),
	.w3(32'hbc9226e3),
	.w4(32'hbbf15a3d),
	.w5(32'hba5cee07),
	.w6(32'hbc67deac),
	.w7(32'hbc912e27),
	.w8(32'h39b968cd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eaff8),
	.w1(32'h3a87de27),
	.w2(32'hbbb3d130),
	.w3(32'h3c87c95f),
	.w4(32'h3b461ff0),
	.w5(32'hbbeb83d4),
	.w6(32'hb8c9fe2c),
	.w7(32'hb984fa90),
	.w8(32'hbc5e0d01),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe66db6),
	.w1(32'hbc6e76cc),
	.w2(32'hbbd229d5),
	.w3(32'h3bc6d47b),
	.w4(32'hbc0a0b00),
	.w5(32'hbbbb73a0),
	.w6(32'hbbce764e),
	.w7(32'hbc3e6379),
	.w8(32'hbb26c6e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26649a),
	.w1(32'hbb66b839),
	.w2(32'h3bf43e37),
	.w3(32'hbbd8d29a),
	.w4(32'hbb484bab),
	.w5(32'h3b26d75e),
	.w6(32'hbb878669),
	.w7(32'hba17120d),
	.w8(32'h3b45c77e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4eb3),
	.w1(32'h3b396c7b),
	.w2(32'h3b026112),
	.w3(32'h3bbc3143),
	.w4(32'h3be1b03e),
	.w5(32'hbbb9c404),
	.w6(32'h3bb7c925),
	.w7(32'h3b9ce921),
	.w8(32'hbb162e08),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7ea41),
	.w1(32'hbaf6f499),
	.w2(32'hba15c483),
	.w3(32'hbc2f35af),
	.w4(32'h39734de3),
	.w5(32'h390bfdea),
	.w6(32'hbb61bf09),
	.w7(32'h3b77d35a),
	.w8(32'hbb0da88a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084329),
	.w1(32'hbae7747d),
	.w2(32'h3c12725e),
	.w3(32'hbbaf23dd),
	.w4(32'hbaa9f4d6),
	.w5(32'h3b35d100),
	.w6(32'hbbfae958),
	.w7(32'hbb209fb5),
	.w8(32'h3b8b6daf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a46e),
	.w1(32'h3b42a0e7),
	.w2(32'hbb6b47f9),
	.w3(32'h3ac87392),
	.w4(32'h3b28ed7a),
	.w5(32'hbb2ad504),
	.w6(32'h3b7a7307),
	.w7(32'h3b8ec19b),
	.w8(32'hbba4e6f5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcff853),
	.w1(32'hbc01c0cd),
	.w2(32'hba8ac761),
	.w3(32'hbbe9900e),
	.w4(32'hbb743d52),
	.w5(32'h3a7adc97),
	.w6(32'hbab57a22),
	.w7(32'hbb589a52),
	.w8(32'h3a6e9dee),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bcaed),
	.w1(32'h3a4e55f0),
	.w2(32'h3a8be952),
	.w3(32'h3b3b34f5),
	.w4(32'h3b7f6b59),
	.w5(32'hbba5a653),
	.w6(32'h3b616729),
	.w7(32'h3b96a6f7),
	.w8(32'hbc2bb38b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4e7b5),
	.w1(32'hbab040b6),
	.w2(32'h3b52daef),
	.w3(32'h38d496f3),
	.w4(32'hb9dfcdc6),
	.w5(32'hbc1c9c78),
	.w6(32'hba99d699),
	.w7(32'h3ab8b797),
	.w8(32'hbc0baae9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e886),
	.w1(32'hbbfe0f77),
	.w2(32'hbade6855),
	.w3(32'hb99c0572),
	.w4(32'h3a7af84b),
	.w5(32'hbc33a095),
	.w6(32'h3b6a11be),
	.w7(32'h3b72bc75),
	.w8(32'h3b18e744),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c3d5d),
	.w1(32'hbba8089a),
	.w2(32'hb9e49848),
	.w3(32'hbbfc3095),
	.w4(32'hbbe85ce9),
	.w5(32'hbc445d40),
	.w6(32'h3b2dd42a),
	.w7(32'h3ad753ce),
	.w8(32'hbc3c0cf6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb470a),
	.w1(32'hba9e5b3f),
	.w2(32'hba9bb867),
	.w3(32'h38d008de),
	.w4(32'h3b8318b0),
	.w5(32'h3b44fa15),
	.w6(32'hbb8dc260),
	.w7(32'hbadc602b),
	.w8(32'h3af32cc0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd390),
	.w1(32'hbb662aa7),
	.w2(32'hbb055e97),
	.w3(32'h3c5688cf),
	.w4(32'h3c8158e6),
	.w5(32'h3b2ed805),
	.w6(32'h3c709ad5),
	.w7(32'h3c92d130),
	.w8(32'h3a5c5a48),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f9ca8),
	.w1(32'hbaf41800),
	.w2(32'hbbf05577),
	.w3(32'h3b40f7bd),
	.w4(32'h3bce0ae9),
	.w5(32'hbc0af50e),
	.w6(32'h3b6d5472),
	.w7(32'h3b81e786),
	.w8(32'hbc12cbe6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79cd1f),
	.w1(32'hbc04a073),
	.w2(32'h3b13a5bf),
	.w3(32'hbc683aeb),
	.w4(32'hbbe05daa),
	.w5(32'h3a1bd773),
	.w6(32'hbc68b597),
	.w7(32'hbbc8dbb1),
	.w8(32'h38dbc60b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d550),
	.w1(32'h3ae742fa),
	.w2(32'hbb8f76a8),
	.w3(32'h3c221406),
	.w4(32'h3c037e1f),
	.w5(32'hbc5c9021),
	.w6(32'h3c130513),
	.w7(32'h3c1372b6),
	.w8(32'hbbdffa5f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ca01f),
	.w1(32'hbbfe3254),
	.w2(32'hbc18a9fd),
	.w3(32'hbbd72a53),
	.w4(32'hbbed9981),
	.w5(32'hbc13d15d),
	.w6(32'hba09271c),
	.w7(32'hbad80d80),
	.w8(32'hbbc02734),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc207631),
	.w1(32'hbc04f734),
	.w2(32'hbc0cc9b3),
	.w3(32'hbbb42182),
	.w4(32'hbbfb6a93),
	.w5(32'hbc800584),
	.w6(32'hbbfcb909),
	.w7(32'hbbf58c74),
	.w8(32'hbc4565fa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb492403),
	.w1(32'hbb9535a9),
	.w2(32'h3bda3985),
	.w3(32'hbc0a129b),
	.w4(32'hbb112665),
	.w5(32'h399d0b55),
	.w6(32'hbb1f1854),
	.w7(32'hbaba08bb),
	.w8(32'h3b019c9b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19878b),
	.w1(32'hbb5b4fc0),
	.w2(32'hbb51d8a3),
	.w3(32'hbbcf2227),
	.w4(32'hbaa6eacf),
	.w5(32'hbab024b7),
	.w6(32'hbb70d683),
	.w7(32'h3b0aab5c),
	.w8(32'hbacf2154),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba871d06),
	.w1(32'hba2a876a),
	.w2(32'hbbf33cb6),
	.w3(32'h3b0265af),
	.w4(32'h3b862cbe),
	.w5(32'hbb69ffaa),
	.w6(32'h3b5cd65c),
	.w7(32'h3bcc177a),
	.w8(32'hbb66a92d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a7f19),
	.w1(32'h3a743055),
	.w2(32'hbbdc4e1d),
	.w3(32'h3b144fb1),
	.w4(32'h3b51cf38),
	.w5(32'hbc638eaa),
	.w6(32'hbb282311),
	.w7(32'hbb32d3d5),
	.w8(32'hbc11d45d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80eeed),
	.w1(32'hbc2ef302),
	.w2(32'hbc13e99d),
	.w3(32'hbc6ae5a8),
	.w4(32'hbc605ebe),
	.w5(32'hbc250ae2),
	.w6(32'hbc7ef9a1),
	.w7(32'hbc15d74c),
	.w8(32'hbbe1e05b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15216),
	.w1(32'hbb0fea57),
	.w2(32'hbbc045c9),
	.w3(32'h3b5a22ce),
	.w4(32'hbb3e524b),
	.w5(32'hbc55308a),
	.w6(32'h3b1ca9a8),
	.w7(32'h3b51e9e8),
	.w8(32'hbbf0df45),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4484a1),
	.w1(32'hbbf6f18d),
	.w2(32'h3badf03e),
	.w3(32'hbc22112e),
	.w4(32'hbc258ef7),
	.w5(32'h3bf989bb),
	.w6(32'hbc4cc5fc),
	.w7(32'hbb3d5c66),
	.w8(32'hb943a34f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39e79),
	.w1(32'hbb4392c0),
	.w2(32'hbc17748f),
	.w3(32'h3ba508cc),
	.w4(32'h3b57b854),
	.w5(32'hbc474b20),
	.w6(32'hbaf59da3),
	.w7(32'hbbec78df),
	.w8(32'hbb2812f3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26b9f1),
	.w1(32'hbba631bb),
	.w2(32'h3a8f63e7),
	.w3(32'hbbfdd813),
	.w4(32'hbc0a5e28),
	.w5(32'hbc184bcd),
	.w6(32'hbb68a045),
	.w7(32'hba753012),
	.w8(32'hba3eee9c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8410d6),
	.w1(32'hbb939b68),
	.w2(32'hbad6ca7f),
	.w3(32'hbc16aa91),
	.w4(32'hbb6f8f67),
	.w5(32'h3929d4af),
	.w6(32'h3c0a43f1),
	.w7(32'h3b87f150),
	.w8(32'hbbc1bb3e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eb9ef),
	.w1(32'hbb1507db),
	.w2(32'h3b9c9395),
	.w3(32'hbb88e3d6),
	.w4(32'hb9a08add),
	.w5(32'hbbd805ee),
	.w6(32'hbbed3dc1),
	.w7(32'hbbc68d7b),
	.w8(32'hbb1cd0c9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf23c8),
	.w1(32'hba1e3125),
	.w2(32'hb9e73271),
	.w3(32'hbb2ae85e),
	.w4(32'h3b46a150),
	.w5(32'hbbd2cdd8),
	.w6(32'h3932c1cc),
	.w7(32'h3bf50e3b),
	.w8(32'hb9d68ef2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32733b),
	.w1(32'hbc103c49),
	.w2(32'h3b6f78c5),
	.w3(32'h3bd1f1b1),
	.w4(32'h3c306ca1),
	.w5(32'hbb798380),
	.w6(32'h3c7e4e20),
	.w7(32'h3d1235df),
	.w8(32'hb7274238),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ec25),
	.w1(32'h3af1de5c),
	.w2(32'h3b44fe67),
	.w3(32'hbb623ffe),
	.w4(32'hbabe8638),
	.w5(32'hbc443ddd),
	.w6(32'h3a024ec2),
	.w7(32'h3ae92bb3),
	.w8(32'hbc222d0e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfabc60),
	.w1(32'hbc29a504),
	.w2(32'h3b3927bc),
	.w3(32'hbb514a86),
	.w4(32'hbbb10bdf),
	.w5(32'hbb04dacb),
	.w6(32'hbaabee25),
	.w7(32'hbb9b36e1),
	.w8(32'hb83dcdb0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7bb9),
	.w1(32'h39b4634a),
	.w2(32'hbb121f9c),
	.w3(32'h3ba2b1e1),
	.w4(32'h3bcbbe01),
	.w5(32'hbb0ce49b),
	.w6(32'h3c280ea3),
	.w7(32'h3ba0405e),
	.w8(32'h3a874019),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa01e27),
	.w1(32'hb9928c9f),
	.w2(32'hbaa3e15c),
	.w3(32'hbb2b8412),
	.w4(32'hbae693b8),
	.w5(32'hbc387638),
	.w6(32'hbaa2e5b7),
	.w7(32'hba4fe99a),
	.w8(32'h3a05e6bd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00a775),
	.w1(32'hbb7a1895),
	.w2(32'hbb895511),
	.w3(32'hbb962bb6),
	.w4(32'h3b5ffd11),
	.w5(32'hbc350a82),
	.w6(32'hbb16552d),
	.w7(32'h3a945628),
	.w8(32'hbb938719),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b222),
	.w1(32'hbba09641),
	.w2(32'hbab40d0f),
	.w3(32'hbbbc2f2f),
	.w4(32'h3ae82b5a),
	.w5(32'hbb00c148),
	.w6(32'hbb957cd7),
	.w7(32'h391e0868),
	.w8(32'hb8c0a284),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebc5b7),
	.w1(32'hbb884aad),
	.w2(32'h3bafe780),
	.w3(32'hbb010fbf),
	.w4(32'hbae3ac41),
	.w5(32'hbbb8ab29),
	.w6(32'h3b285769),
	.w7(32'h39c06d42),
	.w8(32'hbbbcf37f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb479b90),
	.w1(32'hbbd6c8fd),
	.w2(32'hbc0f2fee),
	.w3(32'h3b34f35c),
	.w4(32'hbbaccce9),
	.w5(32'hbc6f51bf),
	.w6(32'h3a5613a1),
	.w7(32'hbbd9ca4e),
	.w8(32'hbc4b9b89),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18e634),
	.w1(32'hbb292597),
	.w2(32'hbb6844d4),
	.w3(32'hbbe3d803),
	.w4(32'hbbd14041),
	.w5(32'hbbbbe431),
	.w6(32'hbbe42653),
	.w7(32'hbb419ef0),
	.w8(32'hbb691f94),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38e126),
	.w1(32'hbae4756b),
	.w2(32'hbb143956),
	.w3(32'hba6f16d7),
	.w4(32'hbb9d91b9),
	.w5(32'h3ae8afe3),
	.w6(32'hbb1ac2f3),
	.w7(32'hbba022d4),
	.w8(32'h3b2857ab),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c095a),
	.w1(32'hbb84fe33),
	.w2(32'hb9a5eba4),
	.w3(32'h3be2c0f1),
	.w4(32'h3af93f1a),
	.w5(32'hbc5799ca),
	.w6(32'h3c123c34),
	.w7(32'h39cdac94),
	.w8(32'hbc192451),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975f6e8),
	.w1(32'hbc34b941),
	.w2(32'h3b735092),
	.w3(32'h3b9fd121),
	.w4(32'hbbb13bbb),
	.w5(32'hb9e84390),
	.w6(32'h3c2af560),
	.w7(32'hbb538371),
	.w8(32'hbacb5a93),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc3707),
	.w1(32'hbacbe4e6),
	.w2(32'hbc132308),
	.w3(32'hb9c3ea2e),
	.w4(32'h37d2a219),
	.w5(32'hbc545ce2),
	.w6(32'hb9c6e781),
	.w7(32'hbb11e4d7),
	.w8(32'hbc274172),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f50c),
	.w1(32'hbb9f5c86),
	.w2(32'hba2ef760),
	.w3(32'hbbdae6c3),
	.w4(32'hbba6c7bc),
	.w5(32'hbba8106d),
	.w6(32'hbb8ee2b2),
	.w7(32'hbab6915f),
	.w8(32'hbae0af15),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01d8eb),
	.w1(32'hbb769474),
	.w2(32'hbc0f707d),
	.w3(32'h38b5949a),
	.w4(32'h3b3460b0),
	.w5(32'hba96af52),
	.w6(32'h3aff61f9),
	.w7(32'h3b3459a5),
	.w8(32'hbb7e3a67),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecd1d7),
	.w1(32'hbbcd5b71),
	.w2(32'hbbc3ef53),
	.w3(32'h3c1448a9),
	.w4(32'h3bf3becf),
	.w5(32'hbc139bbf),
	.w6(32'h3bb1ab19),
	.w7(32'h3b07a61b),
	.w8(32'hbc1bf673),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdfb49),
	.w1(32'hbc0388a4),
	.w2(32'hbb92f7d5),
	.w3(32'hbaacd7f4),
	.w4(32'hbb3942a1),
	.w5(32'hbbe35151),
	.w6(32'hbb378e7f),
	.w7(32'hbb9e9bd8),
	.w8(32'hbc1af421),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd432),
	.w1(32'hbbe70baf),
	.w2(32'hbbfe1e07),
	.w3(32'hbbdb9c2f),
	.w4(32'hba77ab06),
	.w5(32'hbc01e21f),
	.w6(32'hbc42ad1a),
	.w7(32'hbbf5cb3c),
	.w8(32'hbc26dd3f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc865f1e),
	.w1(32'hbbd9e1b7),
	.w2(32'h3b95a7ec),
	.w3(32'hbbc91e41),
	.w4(32'hbadd5a46),
	.w5(32'hbaa5e078),
	.w6(32'hbc46e3ec),
	.w7(32'hbbb600ad),
	.w8(32'h3b1f4919),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb50d),
	.w1(32'h3b3caf87),
	.w2(32'h3a2bd178),
	.w3(32'hbc050da9),
	.w4(32'h3a5a1898),
	.w5(32'h3bd3d19a),
	.w6(32'hbb842dd0),
	.w7(32'h3b58ab9c),
	.w8(32'h3aaa6945),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01733e),
	.w1(32'h3a4d76f1),
	.w2(32'h3a0fb742),
	.w3(32'h3d3ce709),
	.w4(32'h3c204d63),
	.w5(32'hbb2e12bc),
	.w6(32'h3c18e304),
	.w7(32'hba87a5bf),
	.w8(32'hba98ec59),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44dc8a),
	.w1(32'hb7009975),
	.w2(32'h3c0abb37),
	.w3(32'h3b32039a),
	.w4(32'h382d85ce),
	.w5(32'hb8d3d644),
	.w6(32'h3be90503),
	.w7(32'h3af3bf42),
	.w8(32'h3ab6d848),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b03ba),
	.w1(32'h3b6d3932),
	.w2(32'hb95f2d03),
	.w3(32'h3c6d7c53),
	.w4(32'h3c11d327),
	.w5(32'hba64ad24),
	.w6(32'h3c32b5f0),
	.w7(32'h3ab77089),
	.w8(32'h3ba094ca),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56d759),
	.w1(32'h3b5413f5),
	.w2(32'hbbb2bbc7),
	.w3(32'h3be8db62),
	.w4(32'h3a3f4e78),
	.w5(32'hbc15bbc8),
	.w6(32'h3c119bcf),
	.w7(32'h3b989424),
	.w8(32'hbba4d229),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44443),
	.w1(32'hbc2178d7),
	.w2(32'hbb487af6),
	.w3(32'hbc036d8e),
	.w4(32'hbc129b4c),
	.w5(32'hbc0c28dd),
	.w6(32'hbbc8af7b),
	.w7(32'hbb9fdf76),
	.w8(32'hbc02073a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7947b),
	.w1(32'hbbcf1ed4),
	.w2(32'hbc0ceeaa),
	.w3(32'hbbee8a83),
	.w4(32'hbbcf1057),
	.w5(32'hbc3efa37),
	.w6(32'hbbff337e),
	.w7(32'hbbfd3652),
	.w8(32'hbabd3371),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b9bd1),
	.w1(32'hba8b6598),
	.w2(32'h3b20e729),
	.w3(32'hbc55a952),
	.w4(32'hba833fca),
	.w5(32'h3a2f93e2),
	.w6(32'hbbb98a3d),
	.w7(32'h3b33fd2e),
	.w8(32'h3b29c228),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea313b),
	.w1(32'h3b8c29a9),
	.w2(32'hbb4a3981),
	.w3(32'hba89813c),
	.w4(32'h3c1ba6c2),
	.w5(32'hbada830d),
	.w6(32'h3bbf966c),
	.w7(32'h3c79dbcc),
	.w8(32'hba2ab66d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1313f0),
	.w1(32'hbac50453),
	.w2(32'hbc055610),
	.w3(32'hba5b8684),
	.w4(32'h3997652c),
	.w5(32'hbc30e41c),
	.w6(32'hb9a7d226),
	.w7(32'h3ab0336e),
	.w8(32'hbc009177),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18f47c),
	.w1(32'hbbf769ec),
	.w2(32'h3a907fa5),
	.w3(32'hbc0b8be0),
	.w4(32'hbc45b43a),
	.w5(32'hbb7a709b),
	.w6(32'hbc1b3d8b),
	.w7(32'hbc15f1cb),
	.w8(32'hbbdd0bb9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac84780),
	.w1(32'hbbc04b1c),
	.w2(32'h3c1bfb35),
	.w3(32'h36cce145),
	.w4(32'hbbc5f107),
	.w5(32'hbc5b9251),
	.w6(32'hba17ff3e),
	.w7(32'hbb89396b),
	.w8(32'h3b8bd51d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39324598),
	.w1(32'hbb1d3877),
	.w2(32'h3b34effb),
	.w3(32'hbc011d06),
	.w4(32'hbc0c433b),
	.w5(32'hbca252b8),
	.w6(32'h3c02f3d2),
	.w7(32'h3bbe5c90),
	.w8(32'hbc4c0e48),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc993238),
	.w1(32'hbc72994c),
	.w2(32'hba163f57),
	.w3(32'hbc88b1b7),
	.w4(32'hbc6965b1),
	.w5(32'h3c1583f0),
	.w6(32'hbc459b44),
	.w7(32'hbc24062a),
	.w8(32'h3bd41755),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7a3e0),
	.w1(32'h3a8edd61),
	.w2(32'h3b99b963),
	.w3(32'h3c87211a),
	.w4(32'h3c65a9b3),
	.w5(32'h3aa2c604),
	.w6(32'h3c4db4d7),
	.w7(32'h3c16fea3),
	.w8(32'h398b4d81),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3c836),
	.w1(32'hba8cee01),
	.w2(32'hbb2e789b),
	.w3(32'h3bbb0d6a),
	.w4(32'h3b157822),
	.w5(32'hbb72b213),
	.w6(32'h3b53e627),
	.w7(32'h3a72e996),
	.w8(32'hbafcc266),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891e23),
	.w1(32'hbb8d08cd),
	.w2(32'hbb1ae67d),
	.w3(32'h3aede718),
	.w4(32'hbb92e27d),
	.w5(32'h3b2fdc8c),
	.w6(32'hbb3736ab),
	.w7(32'hbbae1cf7),
	.w8(32'hba25316f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe71498),
	.w1(32'hbaa3b9cc),
	.w2(32'hbb664b5b),
	.w3(32'h38bc9265),
	.w4(32'h3b82b63e),
	.w5(32'h3b1b3f59),
	.w6(32'hbaf899ff),
	.w7(32'hb9a6ff12),
	.w8(32'hbafe7765),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3a1a),
	.w1(32'hba94ce8a),
	.w2(32'hbbd796b1),
	.w3(32'h3c3ccd2d),
	.w4(32'h3c4eb2fb),
	.w5(32'hbc762282),
	.w6(32'h3a23e9ad),
	.w7(32'h3ab642c9),
	.w8(32'hbc17d5ff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43bc28),
	.w1(32'hbbd7fdfa),
	.w2(32'h3b4c6c0c),
	.w3(32'hbca3eadc),
	.w4(32'hbc418568),
	.w5(32'h3b565921),
	.w6(32'hbc2e5844),
	.w7(32'hbc3c1908),
	.w8(32'hba16373f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d82cf),
	.w1(32'h3b444b04),
	.w2(32'h3bb5d568),
	.w3(32'hb8a0fc50),
	.w4(32'h3b213c32),
	.w5(32'h3b8ca224),
	.w6(32'hbb13ddd2),
	.w7(32'h3a28acdf),
	.w8(32'hba9c6862),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6f7c5),
	.w1(32'h3b8bf017),
	.w2(32'hbbf9b133),
	.w3(32'hbc15b54d),
	.w4(32'h3c622671),
	.w5(32'hbb3439b9),
	.w6(32'hbc4ab08e),
	.w7(32'h3c3d865b),
	.w8(32'hbc285441),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc687fc8),
	.w1(32'hbc127b9f),
	.w2(32'hbbda5716),
	.w3(32'h3ae1d114),
	.w4(32'h3bd41dc1),
	.w5(32'hbbadd1ab),
	.w6(32'hbc1c5480),
	.w7(32'hbb8f09e1),
	.w8(32'hbc5962c9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8259a7),
	.w1(32'hbc3978c9),
	.w2(32'h3afb4b3d),
	.w3(32'hbbe84fd4),
	.w4(32'hbb07f6e7),
	.w5(32'h3af539c9),
	.w6(32'hbc640e18),
	.w7(32'hbbc6f2f5),
	.w8(32'h3b46078c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592276),
	.w1(32'h3aabb9cb),
	.w2(32'h38a18951),
	.w3(32'h3b6e27ec),
	.w4(32'hba78f3cd),
	.w5(32'hb906faf0),
	.w6(32'h3bb62a29),
	.w7(32'h3818ed61),
	.w8(32'h3add5c1e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cf513),
	.w1(32'h3bd07330),
	.w2(32'hba97382e),
	.w3(32'hbb8fddcb),
	.w4(32'h3b0dff07),
	.w5(32'hbbba8628),
	.w6(32'hbb7d6ebc),
	.w7(32'h3bab6e38),
	.w8(32'hba50cc1b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3baf2e),
	.w1(32'hbb97619c),
	.w2(32'h3b1509bf),
	.w3(32'hbbc92ebb),
	.w4(32'hbc1a9c38),
	.w5(32'hbae079f0),
	.w6(32'hbb7c242a),
	.w7(32'hbb824233),
	.w8(32'h389cfca0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b570ad3),
	.w1(32'h3b36074e),
	.w2(32'hbb38a34f),
	.w3(32'hbb1b323e),
	.w4(32'hbae7e4ac),
	.w5(32'hbb4bae70),
	.w6(32'hbb1ceb10),
	.w7(32'hba4fc288),
	.w8(32'hbafa8aa9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a0ad0),
	.w1(32'h3b9257ac),
	.w2(32'hbb4c563f),
	.w3(32'hb9163df5),
	.w4(32'h3bbec39c),
	.w5(32'hba048f88),
	.w6(32'hb9bf7790),
	.w7(32'h3bdbf803),
	.w8(32'hbb945cc0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc41068),
	.w1(32'h3b598c0a),
	.w2(32'hbbc97ae2),
	.w3(32'hbbdb8714),
	.w4(32'h3c084280),
	.w5(32'hbc5b30ea),
	.w6(32'hbb79b4a8),
	.w7(32'h3bbbb0a8),
	.w8(32'hbc07f6ae),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc846fe),
	.w1(32'hb9e5877e),
	.w2(32'h3b50b4e7),
	.w3(32'hbc213797),
	.w4(32'hbbe7cfd8),
	.w5(32'h3c03efc5),
	.w6(32'hbb88e5bc),
	.w7(32'hbb1e45e3),
	.w8(32'hbba408fd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fafe9),
	.w1(32'hba109ef5),
	.w2(32'hbba0cca4),
	.w3(32'h3bec6086),
	.w4(32'h3c7b1dc3),
	.w5(32'hbc5eea8e),
	.w6(32'hbbb3b8d2),
	.w7(32'hba86467c),
	.w8(32'hbc064b2c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f22be),
	.w1(32'hbb8768a6),
	.w2(32'h3b0ed592),
	.w3(32'hbc8e1f6e),
	.w4(32'hbc25f60d),
	.w5(32'h3a0f9137),
	.w6(32'hbc57218c),
	.w7(32'hbc17f7be),
	.w8(32'h398b8457),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d2221),
	.w1(32'h3a2d801b),
	.w2(32'h3b8557c4),
	.w3(32'hbb3441fd),
	.w4(32'h3b313dbb),
	.w5(32'hbac19710),
	.w6(32'hbb8a7383),
	.w7(32'h3b055932),
	.w8(32'h37aa3751),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedf7bc),
	.w1(32'hba0660ef),
	.w2(32'h3b137453),
	.w3(32'h3a8954e6),
	.w4(32'hb6dc6287),
	.w5(32'hbb83d58b),
	.w6(32'h3b993c4a),
	.w7(32'h3af87d32),
	.w8(32'hb9e86c74),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaddea9),
	.w1(32'hb9836c09),
	.w2(32'hbad7d09e),
	.w3(32'hbb4f148b),
	.w4(32'hb9c6c067),
	.w5(32'hba0fe15a),
	.w6(32'hbaa61ae1),
	.w7(32'h3b01d8f7),
	.w8(32'hbbf3563d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5124),
	.w1(32'hbbb1768d),
	.w2(32'hbb81feb2),
	.w3(32'hbb00ac13),
	.w4(32'h3ab87b1e),
	.w5(32'hba06b897),
	.w6(32'hba47caee),
	.w7(32'hbaba9e1f),
	.w8(32'hba1a774a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff642d),
	.w1(32'hb9d40f2a),
	.w2(32'hba29c252),
	.w3(32'hbb3ed859),
	.w4(32'h3b702c6d),
	.w5(32'hbb5d538a),
	.w6(32'hbaea02aa),
	.w7(32'h3b381ae0),
	.w8(32'hbbd53cab),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc312eee),
	.w1(32'hbc31f803),
	.w2(32'hbb9c2399),
	.w3(32'h3b8c0d55),
	.w4(32'h3bc62561),
	.w5(32'hbb63ca94),
	.w6(32'h3b1d259d),
	.w7(32'h3aa5563e),
	.w8(32'h3bf8a103),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfc481),
	.w1(32'hbbbb7218),
	.w2(32'hbb1afe42),
	.w3(32'h3b8a7151),
	.w4(32'h3b0c76f3),
	.w5(32'hbc1b6014),
	.w6(32'h3c49cf79),
	.w7(32'h3c226347),
	.w8(32'hbb4d1813),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f95e),
	.w1(32'hbabf60cb),
	.w2(32'hbbf764c6),
	.w3(32'hbbc57790),
	.w4(32'hb8416d82),
	.w5(32'h3b9356a3),
	.w6(32'hbbad49ca),
	.w7(32'hba8e1e2f),
	.w8(32'hbc651f5e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31d238),
	.w1(32'hbb898482),
	.w2(32'hbb5bfd27),
	.w3(32'hba08f4eb),
	.w4(32'h3bc41f05),
	.w5(32'hbbb5b33b),
	.w6(32'hbc3be541),
	.w7(32'hbb934510),
	.w8(32'hbb857819),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e1a9),
	.w1(32'hbb9d5ccd),
	.w2(32'h3ad0507b),
	.w3(32'hbadcafbb),
	.w4(32'hbb8cd7f8),
	.w5(32'h3b222445),
	.w6(32'hbb4e048b),
	.w7(32'hbb962d73),
	.w8(32'h3b9b7c8b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432bbf),
	.w1(32'h3ac097b8),
	.w2(32'hbb397e62),
	.w3(32'h3ae0cd9d),
	.w4(32'h3abdbfea),
	.w5(32'hbbb3a750),
	.w6(32'h3ba9e924),
	.w7(32'h3bc4411f),
	.w8(32'hbb8d9386),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb677c83),
	.w1(32'hbb47d731),
	.w2(32'h3be47e6c),
	.w3(32'hbb833e3b),
	.w4(32'hbb2028ea),
	.w5(32'hb888d932),
	.w6(32'hbb66f50f),
	.w7(32'hbad31d99),
	.w8(32'h3af38988),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74dbe),
	.w1(32'hbc043bd1),
	.w2(32'hbb0c2070),
	.w3(32'hb8de06b0),
	.w4(32'h3b0d649e),
	.w5(32'hbb82de2f),
	.w6(32'h3aad7d13),
	.w7(32'hba89b657),
	.w8(32'hbb31d4da),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c9c5),
	.w1(32'hbac3acd4),
	.w2(32'h3b1529af),
	.w3(32'hb793c7e6),
	.w4(32'hbb8d377d),
	.w5(32'hbbfab639),
	.w6(32'hba7e0da8),
	.w7(32'hbb5976ca),
	.w8(32'hbb35e757),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc2f1b),
	.w1(32'h3b337c0f),
	.w2(32'hbbd3c7ad),
	.w3(32'hbb3b09da),
	.w4(32'hbaaac265),
	.w5(32'hbc33bbf4),
	.w6(32'h3aa3c49d),
	.w7(32'hbb0b6a89),
	.w8(32'hbc1d35b7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf13e4c),
	.w1(32'hbb23c624),
	.w2(32'hbbfc6900),
	.w3(32'hbba49475),
	.w4(32'hbbc892ac),
	.w5(32'hbc4f024a),
	.w6(32'hbaf0053f),
	.w7(32'h3ab594b3),
	.w8(32'hbc2885a8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8894e8),
	.w1(32'hbad1cf6c),
	.w2(32'hbbdc1cdd),
	.w3(32'hbb6dee40),
	.w4(32'hbb18c30d),
	.w5(32'hbbab6a02),
	.w6(32'hb95fa8e6),
	.w7(32'h3b2f10c6),
	.w8(32'hbc4b68dc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8cd9),
	.w1(32'h3b890def),
	.w2(32'hbb866745),
	.w3(32'hbaafdd87),
	.w4(32'h3c20ce35),
	.w5(32'hbb049a3f),
	.w6(32'hbb74ce6b),
	.w7(32'hbae74dfe),
	.w8(32'hbaa184e0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0353c2),
	.w1(32'hbb1f5824),
	.w2(32'hbb2edc5d),
	.w3(32'hbba54fe4),
	.w4(32'hbb7fe81c),
	.w5(32'hbbfc2c56),
	.w6(32'hbb6a30d1),
	.w7(32'hbb7d3bfd),
	.w8(32'hbb36e301),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4631be),
	.w1(32'hbc2ce566),
	.w2(32'hbb9e58c4),
	.w3(32'hbbf7be3b),
	.w4(32'hbb3f81a6),
	.w5(32'hbc0e0db9),
	.w6(32'hbb9c1eb4),
	.w7(32'hba0ce28f),
	.w8(32'hbc23de80),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e7f13),
	.w1(32'hbbe0fc85),
	.w2(32'hbc3bdc44),
	.w3(32'hbbdeffdb),
	.w4(32'hbb8f6c55),
	.w5(32'hbc3c1bee),
	.w6(32'hbc1b1eab),
	.w7(32'hbc1e56e7),
	.w8(32'hbb8c08cc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc538a79),
	.w1(32'hbba9561b),
	.w2(32'hbbb3d0d5),
	.w3(32'hbc040b0e),
	.w4(32'hbc03d918),
	.w5(32'hbba4704d),
	.w6(32'hbc0205c3),
	.w7(32'hbbf3828d),
	.w8(32'hbb4eb62a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc148909),
	.w1(32'h3c0324fb),
	.w2(32'hbb4e5e76),
	.w3(32'hbad56926),
	.w4(32'h3c0f2617),
	.w5(32'hbb1d5a66),
	.w6(32'h3b8c6ae1),
	.w7(32'h3c179468),
	.w8(32'hbb655f81),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7e66),
	.w1(32'hbb273625),
	.w2(32'hbbcc1266),
	.w3(32'h3c2e499f),
	.w4(32'h3bf513e5),
	.w5(32'hba6fcb59),
	.w6(32'h3be1960d),
	.w7(32'h3970a664),
	.w8(32'h3ad28b75),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3160f),
	.w1(32'hbb4545f3),
	.w2(32'h3aae2127),
	.w3(32'h3b2827da),
	.w4(32'hbaeec040),
	.w5(32'hba2d9376),
	.w6(32'h3b4540ea),
	.w7(32'h3a0fbfc4),
	.w8(32'h3b72e213),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350fbc84),
	.w1(32'hb96f07ea),
	.w2(32'hbb818b0f),
	.w3(32'hbb819f5d),
	.w4(32'hba78666e),
	.w5(32'hbc288240),
	.w6(32'h3beb9df8),
	.w7(32'h3b4b8740),
	.w8(32'hbc13fff6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2015ce),
	.w1(32'hbc09d5a9),
	.w2(32'hbc03bfda),
	.w3(32'hbbaa13a4),
	.w4(32'hbbb1951f),
	.w5(32'hbc83d97e),
	.w6(32'hbc194c5d),
	.w7(32'hbbc44de1),
	.w8(32'hbc6e35aa),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507823),
	.w1(32'hbc26c84e),
	.w2(32'hb867861e),
	.w3(32'hbc681c83),
	.w4(32'hbc6009b9),
	.w5(32'hbb1d9482),
	.w6(32'hbc6641ae),
	.w7(32'hbc577858),
	.w8(32'hbbb45f71),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad103d),
	.w1(32'hbac1d6b0),
	.w2(32'hbacf8b10),
	.w3(32'hbba81fe8),
	.w4(32'h38460961),
	.w5(32'h3aaf1242),
	.w6(32'hbbdc98c2),
	.w7(32'hbb80ec40),
	.w8(32'hb9e9964f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bcb1a),
	.w1(32'hbb3ec79f),
	.w2(32'hbbf34bbd),
	.w3(32'h3bcc7cf6),
	.w4(32'h3bb67ce5),
	.w5(32'hbc25de23),
	.w6(32'h3b788e39),
	.w7(32'h3b17a27b),
	.w8(32'hbc46705e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5b5d7),
	.w1(32'hbb590ed9),
	.w2(32'hbc3b9824),
	.w3(32'h3ac883d5),
	.w4(32'hbb86189f),
	.w5(32'hbc0f1b0f),
	.w6(32'h3b8a806f),
	.w7(32'hbc035c18),
	.w8(32'h3beebf96),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670adc),
	.w1(32'hbc1596db),
	.w2(32'h3b80ee84),
	.w3(32'hbc32ae7b),
	.w4(32'hbbf5ea51),
	.w5(32'h3b07b736),
	.w6(32'h3a2d84a1),
	.w7(32'h3ba37d6d),
	.w8(32'h3bee9d14),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5dc5b),
	.w1(32'hbbe20e22),
	.w2(32'hbb82236e),
	.w3(32'h3aa1113e),
	.w4(32'hbb37a3c6),
	.w5(32'hbc27f882),
	.w6(32'h3c4da3b1),
	.w7(32'h3aa09a71),
	.w8(32'hbc203f42),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123805),
	.w1(32'hbbe95b6a),
	.w2(32'h3b0f9150),
	.w3(32'hbc0cf696),
	.w4(32'hbc120bb2),
	.w5(32'h3acd9138),
	.w6(32'hbc128c60),
	.w7(32'hbc1afd0c),
	.w8(32'h3984d5fc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965ff3),
	.w1(32'hba9ae0cc),
	.w2(32'h3a92f1bb),
	.w3(32'h3a9e6455),
	.w4(32'h3aff7161),
	.w5(32'h3b86a3b2),
	.w6(32'h3b4856e3),
	.w7(32'h3c126398),
	.w8(32'hbadc2eef),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23fc5b),
	.w1(32'h3b90b453),
	.w2(32'hbb02d9a9),
	.w3(32'h3bf94a0d),
	.w4(32'h3c2a7d37),
	.w5(32'hbaa75fdf),
	.w6(32'h3b0c7af4),
	.w7(32'h3b839d37),
	.w8(32'hbba2ca1b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68fed),
	.w1(32'hbb984c92),
	.w2(32'h3a3ee6f4),
	.w3(32'h39196c32),
	.w4(32'h3b818f4f),
	.w5(32'hba5b98af),
	.w6(32'hbbdd690d),
	.w7(32'hbba2ca79),
	.w8(32'hbb18b041),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f337),
	.w1(32'hba9da641),
	.w2(32'hba9cbd26),
	.w3(32'h3926cfd3),
	.w4(32'hbb183f7f),
	.w5(32'hbc32709b),
	.w6(32'hbb3663e7),
	.w7(32'hb9c854e3),
	.w8(32'hbb9975d3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44055c),
	.w1(32'hbade3642),
	.w2(32'hbaed0c09),
	.w3(32'hbc8895cc),
	.w4(32'hbc0459de),
	.w5(32'h3b7d7df6),
	.w6(32'hbc01514e),
	.w7(32'hbc0ded13),
	.w8(32'hbb9c692e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1623c7),
	.w1(32'hbba4e92a),
	.w2(32'h3bbc84de),
	.w3(32'h3c209c7f),
	.w4(32'h3b3f9e6f),
	.w5(32'h3b82ae05),
	.w6(32'h3b76b0bc),
	.w7(32'hbb98e5ed),
	.w8(32'h3bdd0254),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8771fc),
	.w1(32'h3b35a8c8),
	.w2(32'hbc0e7c46),
	.w3(32'h3c0f4d8a),
	.w4(32'h3c0c8d68),
	.w5(32'hbc167dc1),
	.w6(32'h3c19d57e),
	.w7(32'h3be0dbd0),
	.w8(32'hbc611f65),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2bb5d),
	.w1(32'hbb4f4ac9),
	.w2(32'hbbb1a261),
	.w3(32'h3c2e3c51),
	.w4(32'h3afcc3c8),
	.w5(32'hbbcafd15),
	.w6(32'hb8780745),
	.w7(32'hbbb0107e),
	.w8(32'hbb0564d8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b9a0),
	.w1(32'hbbfb0bb1),
	.w2(32'hbbc23282),
	.w3(32'hbbc8ca62),
	.w4(32'hbbbd8217),
	.w5(32'hbc05efaa),
	.w6(32'hbb9d80f8),
	.w7(32'hbbcf1509),
	.w8(32'hbc28f6e7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4324a5),
	.w1(32'hbb488fe6),
	.w2(32'hba408368),
	.w3(32'hbbecde19),
	.w4(32'hbbe283a0),
	.w5(32'hbac83731),
	.w6(32'hbc6d5eab),
	.w7(32'hbbfa6aa9),
	.w8(32'h3a4478d1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e71125),
	.w1(32'h3a3a8b98),
	.w2(32'h3c07dc9b),
	.w3(32'h3b66e312),
	.w4(32'hb9c4b8ef),
	.w5(32'h3c3feb0e),
	.w6(32'h3afa3008),
	.w7(32'h3a63bd56),
	.w8(32'h3bf559e5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b19d6),
	.w1(32'h39fb758d),
	.w2(32'hbc09ec18),
	.w3(32'h3c2b2c4c),
	.w4(32'h3b2bbc97),
	.w5(32'hbbc9238a),
	.w6(32'h3b690d98),
	.w7(32'hbb96f581),
	.w8(32'h3ab386f6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1cbd),
	.w1(32'hbba6ca2f),
	.w2(32'hbbb9d617),
	.w3(32'hbcdbbeb8),
	.w4(32'hbccbcf32),
	.w5(32'hbbc381f1),
	.w6(32'hbc99b510),
	.w7(32'hbcb5ffb1),
	.w8(32'hba520614),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc095a8),
	.w1(32'hbafbdc4f),
	.w2(32'hbb8a8db7),
	.w3(32'hbb4ee01f),
	.w4(32'h3b0d4cb9),
	.w5(32'hbbb80e42),
	.w6(32'h3b53e3c6),
	.w7(32'h3bbbdfaf),
	.w8(32'hba627bd7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dcdd7),
	.w1(32'h3b7227c3),
	.w2(32'h3b8bd3e2),
	.w3(32'h3bff8c53),
	.w4(32'h3baa4d99),
	.w5(32'hb9c7681b),
	.w6(32'h3c1c77bb),
	.w7(32'h3c3ba58f),
	.w8(32'hbb71af5e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ee9ea),
	.w1(32'hb9bd94d9),
	.w2(32'hbacb2429),
	.w3(32'h3c81c4de),
	.w4(32'h3c5d522a),
	.w5(32'hbb91e3c2),
	.w6(32'h3c1b12bc),
	.w7(32'h3bb6a8c1),
	.w8(32'hbad30bc0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9248a5),
	.w1(32'h3bcbbad9),
	.w2(32'hbbb3c80c),
	.w3(32'hbb3d513e),
	.w4(32'h3a476acc),
	.w5(32'hbc4cc796),
	.w6(32'hb979866d),
	.w7(32'h3afcdebb),
	.w8(32'hbc037d06),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c6020),
	.w1(32'hbb55d1cf),
	.w2(32'h3b01f5ad),
	.w3(32'hbc54004b),
	.w4(32'h3b863bfe),
	.w5(32'hbb01fff7),
	.w6(32'hbc6511e2),
	.w7(32'h3c0ff07f),
	.w8(32'hbb3e0aaf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07a497),
	.w1(32'h3a953e1b),
	.w2(32'h3a33f3a1),
	.w3(32'hba0e56d9),
	.w4(32'hbb8679a4),
	.w5(32'h3b1d9637),
	.w6(32'hbb9179e2),
	.w7(32'hbb8b280d),
	.w8(32'h3beb2303),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d167b),
	.w1(32'hbb9441cf),
	.w2(32'hbb9ca906),
	.w3(32'hbc22a4fc),
	.w4(32'hbc3107a7),
	.w5(32'hbc241274),
	.w6(32'hbc1b6d4d),
	.w7(32'hbc1e3230),
	.w8(32'hbbdfc4c7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c5ce3),
	.w1(32'hbbd9bce0),
	.w2(32'h3acb2534),
	.w3(32'hbc114717),
	.w4(32'hbba590e0),
	.w5(32'hbb338f71),
	.w6(32'hbb975590),
	.w7(32'hbb2fad42),
	.w8(32'hba9c1ba9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf189a7),
	.w1(32'hbb81c2bd),
	.w2(32'h3c2fe2f1),
	.w3(32'hbc8e1585),
	.w4(32'hbc3e52ee),
	.w5(32'h3c8e5ac9),
	.w6(32'hbc169b89),
	.w7(32'hbc3abf72),
	.w8(32'h3bad6805),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1abbd3),
	.w1(32'hbb09b7c2),
	.w2(32'hbaf06869),
	.w3(32'h3cdb865c),
	.w4(32'hba77d671),
	.w5(32'hba6ce00f),
	.w6(32'h3c90a0c2),
	.w7(32'hbb5ce297),
	.w8(32'hbb331c55),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4aa0c),
	.w1(32'h3a877cde),
	.w2(32'hba3aa58f),
	.w3(32'hba3008fa),
	.w4(32'hbc018b7a),
	.w5(32'hbbad9a5c),
	.w6(32'hbb17efed),
	.w7(32'hbbfa70ff),
	.w8(32'hbacfc570),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe78a37),
	.w1(32'hbaf61aa2),
	.w2(32'hba7bae5e),
	.w3(32'h3b1c1321),
	.w4(32'hb9fb619c),
	.w5(32'hbc011c2d),
	.w6(32'h39abf46a),
	.w7(32'h3b08fe1a),
	.w8(32'h3b562a49),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5edaa2),
	.w1(32'hbb3e7821),
	.w2(32'h3a85fdbf),
	.w3(32'h3be34b5f),
	.w4(32'hbbfce091),
	.w5(32'hbb519b67),
	.w6(32'h3bfd4a46),
	.w7(32'hbb63bffb),
	.w8(32'hbb3fd4c0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5757a0),
	.w1(32'hbb835e0a),
	.w2(32'hbb7781ed),
	.w3(32'hbb3f6adb),
	.w4(32'hbaf34945),
	.w5(32'hbbc1105b),
	.w6(32'hbb85f615),
	.w7(32'hbb277cb3),
	.w8(32'hbbd24674),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0ff0a),
	.w1(32'h3b889c50),
	.w2(32'h3adc598f),
	.w3(32'hbd24a300),
	.w4(32'h3c192ab0),
	.w5(32'hbbb0fbeb),
	.w6(32'hbc73a983),
	.w7(32'h3bec9a4a),
	.w8(32'h3b189e25),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a71cc),
	.w1(32'h3bdd50ba),
	.w2(32'h3b3844c1),
	.w3(32'hbb320400),
	.w4(32'h3ba9d0c3),
	.w5(32'hbb7252a8),
	.w6(32'h3ab60918),
	.w7(32'h3c41f8ef),
	.w8(32'hbbb26a59),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954a53),
	.w1(32'hbacd5f90),
	.w2(32'hbb764c0b),
	.w3(32'h3be6fa31),
	.w4(32'h39ec8ff7),
	.w5(32'hbc7c0c90),
	.w6(32'h3bbc5f49),
	.w7(32'hbab407bc),
	.w8(32'hbc7b4235),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f9a35),
	.w1(32'hbb9c6277),
	.w2(32'h3b7f477d),
	.w3(32'hbcc151f9),
	.w4(32'hbc01c621),
	.w5(32'h3a7fb665),
	.w6(32'hbc270de7),
	.w7(32'hbbfd94e2),
	.w8(32'hbb0dd176),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97c7b),
	.w1(32'hba47e81b),
	.w2(32'hbc2f4180),
	.w3(32'h3bc4d321),
	.w4(32'h3aef93d3),
	.w5(32'hbcac32f3),
	.w6(32'hba1f2933),
	.w7(32'hbb0353e6),
	.w8(32'hbb679fe6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf04fe1),
	.w1(32'h3c7082e3),
	.w2(32'hba3d274a),
	.w3(32'h3d9c0103),
	.w4(32'h3d2e98c5),
	.w5(32'hbc24304d),
	.w6(32'h3d79a63f),
	.w7(32'h3d0cd1cb),
	.w8(32'hbc5ac1d6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9bce7),
	.w1(32'hbc3a197e),
	.w2(32'hbb3faab7),
	.w3(32'hbc8416ba),
	.w4(32'hbbfa13e3),
	.w5(32'hbbadb7dc),
	.w6(32'hbc32ff6f),
	.w7(32'hbb962a53),
	.w8(32'h3c14f964),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a9e33),
	.w1(32'hbc1927cd),
	.w2(32'h3bf583eb),
	.w3(32'h3b0f6f74),
	.w4(32'hbc9529f4),
	.w5(32'h3c494d88),
	.w6(32'hba17e3e8),
	.w7(32'hbc8aa3ae),
	.w8(32'hbb2bdc0b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4306d),
	.w1(32'h3b83c1ff),
	.w2(32'h3b4ea806),
	.w3(32'hbabe3ca4),
	.w4(32'h3b9afa9d),
	.w5(32'h3bfae120),
	.w6(32'h3bc28876),
	.w7(32'h3ba646b9),
	.w8(32'h39a16c2e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c342155),
	.w1(32'h3bfb3ca7),
	.w2(32'hbcb54ecb),
	.w3(32'h3c8bddf4),
	.w4(32'h3c425c9d),
	.w5(32'hbb8b2c05),
	.w6(32'h39af0b28),
	.w7(32'hbb324516),
	.w8(32'h3bb6d33c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce7fe29),
	.w1(32'h3bed7cf5),
	.w2(32'h3c062aed),
	.w3(32'h3d64967b),
	.w4(32'h3cea3e79),
	.w5(32'hbb13f2b0),
	.w6(32'h3cc63ccc),
	.w7(32'h3c350cc5),
	.w8(32'hbb85ec8f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49933c),
	.w1(32'h3b845ae0),
	.w2(32'h3b3adf31),
	.w3(32'hbbad0133),
	.w4(32'h3bc29e61),
	.w5(32'hbb215761),
	.w6(32'h38933d6e),
	.w7(32'h3c647577),
	.w8(32'h3aa5df08),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62c3ec),
	.w1(32'h3b9a21bf),
	.w2(32'h3c526aa1),
	.w3(32'h3d2ff72e),
	.w4(32'h3c90f822),
	.w5(32'h3b2cc333),
	.w6(32'h3ccf5824),
	.w7(32'h3c1c6609),
	.w8(32'hbbd4ef77),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b320573),
	.w1(32'hbc3be85f),
	.w2(32'hbb5656f5),
	.w3(32'hbc0bf74c),
	.w4(32'hbbde59d6),
	.w5(32'hbb109ae7),
	.w6(32'hbbca938f),
	.w7(32'h3906d53a),
	.w8(32'hbc0b05b0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ac87),
	.w1(32'h3bac4fe7),
	.w2(32'h3b9e1fb7),
	.w3(32'hbb26bb14),
	.w4(32'h3b7124eb),
	.w5(32'h3b56e3a1),
	.w6(32'hbbf7e4b3),
	.w7(32'hbb0fb4ad),
	.w8(32'hbb61d922),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c344b09),
	.w1(32'h3b880631),
	.w2(32'hbc3e50ee),
	.w3(32'h3c30ce4f),
	.w4(32'h3be97090),
	.w5(32'hbc3b8091),
	.w6(32'h3aafa66a),
	.w7(32'h3a59bf10),
	.w8(32'hbb02b46e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57a61a),
	.w1(32'h3b26aad0),
	.w2(32'hba81e050),
	.w3(32'h3c6f5fad),
	.w4(32'h3cb62959),
	.w5(32'hb91035bd),
	.w6(32'h3c9b0aa7),
	.w7(32'h3c941a1e),
	.w8(32'h3b68e39d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29f94e),
	.w1(32'hbc415b89),
	.w2(32'hbb552bdf),
	.w3(32'hbc341491),
	.w4(32'hbc3f2629),
	.w5(32'hbc0d842f),
	.w6(32'h3b1c8cd8),
	.w7(32'hbc59f64f),
	.w8(32'hbbb324e0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece079),
	.w1(32'h3b8bd528),
	.w2(32'h38859f0b),
	.w3(32'hbc4e3db6),
	.w4(32'hbbdd9515),
	.w5(32'hbc012165),
	.w6(32'hba23574f),
	.w7(32'hbbd62911),
	.w8(32'h3a2532c1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36a412),
	.w1(32'hbbb61b9d),
	.w2(32'hbb7e30ed),
	.w3(32'hbc1537a2),
	.w4(32'hbc16eefe),
	.w5(32'h3a046d25),
	.w6(32'hbb881533),
	.w7(32'hbc03f656),
	.w8(32'hbb4cb416),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34c267),
	.w1(32'h3a1dad13),
	.w2(32'h3a7d2ecd),
	.w3(32'h3be168ca),
	.w4(32'h3b5ec2ba),
	.w5(32'hba364059),
	.w6(32'h3c167ced),
	.w7(32'h3c5b7035),
	.w8(32'hbb4d2d2e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85fbff),
	.w1(32'hba6ad742),
	.w2(32'h3c1f94d2),
	.w3(32'hbb03b5c2),
	.w4(32'hba35ff49),
	.w5(32'h3bf1c9ec),
	.w6(32'hbb8dd89d),
	.w7(32'hbb2c0955),
	.w8(32'h3c4e8e7b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b188537),
	.w1(32'h3ba21664),
	.w2(32'hbb6fa208),
	.w3(32'h3b0c7c73),
	.w4(32'h3ba7d710),
	.w5(32'h3a19c964),
	.w6(32'h3bc49b1f),
	.w7(32'h3be9f344),
	.w8(32'hbb4a591a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d2278),
	.w1(32'hb9c4c8a0),
	.w2(32'h3b48260d),
	.w3(32'h3b725456),
	.w4(32'h3a99041f),
	.w5(32'hbc57b0fb),
	.w6(32'hba834f22),
	.w7(32'hbbd66756),
	.w8(32'hbbde9072),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f4e33),
	.w1(32'hbc48f08a),
	.w2(32'h3b808444),
	.w3(32'hbc72eb2f),
	.w4(32'hbaefb586),
	.w5(32'h3b94c0b3),
	.w6(32'hbc7256fc),
	.w7(32'hbc2a12d3),
	.w8(32'h3b7bf7dc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78a60e),
	.w1(32'h3b11b113),
	.w2(32'h3b9dd9af),
	.w3(32'h3ab3bcd8),
	.w4(32'h3b4c858d),
	.w5(32'h3bdd3c97),
	.w6(32'h3aa2f3df),
	.w7(32'h3b8f81d4),
	.w8(32'h3c3dc4fd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059dbc),
	.w1(32'h3b7940f0),
	.w2(32'h3baee4c9),
	.w3(32'h3b6ac561),
	.w4(32'hbb49e0ab),
	.w5(32'h3b6221a6),
	.w6(32'h3b25d733),
	.w7(32'hba367312),
	.w8(32'h3c059433),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945056),
	.w1(32'h3baf7fc5),
	.w2(32'hbb75bd28),
	.w3(32'hba043644),
	.w4(32'h3b5931b8),
	.w5(32'hbb85dd6b),
	.w6(32'h3bafa48d),
	.w7(32'h3c03f33b),
	.w8(32'hbacf57ec),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bdab5),
	.w1(32'hbc11d7d9),
	.w2(32'h3bde71fe),
	.w3(32'hbc8f87b8),
	.w4(32'hbbb06c33),
	.w5(32'h3ba9266b),
	.w6(32'hbc10d03b),
	.w7(32'h3b0d619e),
	.w8(32'h3b3cb4ef),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6444b4),
	.w1(32'hbc6fd7dd),
	.w2(32'hbba196f6),
	.w3(32'hbbb7a376),
	.w4(32'hbc8c71d7),
	.w5(32'hbc0cdbb1),
	.w6(32'hbb920583),
	.w7(32'hbc808d1e),
	.w8(32'hbb83fec4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e408b),
	.w1(32'hbb305a3f),
	.w2(32'hbc613e30),
	.w3(32'h3b4e1b97),
	.w4(32'h3a244f7e),
	.w5(32'hbc98fe3a),
	.w6(32'h3b61dfea),
	.w7(32'h3a66aaa4),
	.w8(32'hbc89c452),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9f9e2),
	.w1(32'hbbc68726),
	.w2(32'hbbc8692b),
	.w3(32'hbb8f844d),
	.w4(32'hbc04ad7b),
	.w5(32'hb89ed232),
	.w6(32'hbbbbaf77),
	.w7(32'hbbfe3b3e),
	.w8(32'hbb9975cc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982d41),
	.w1(32'h3a7e3b88),
	.w2(32'h39fbc6b9),
	.w3(32'h3b4f51b3),
	.w4(32'h3ba05717),
	.w5(32'hbb58514e),
	.w6(32'h3c30a472),
	.w7(32'h3c37337d),
	.w8(32'hbc1b3290),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d118d),
	.w1(32'h3b71665a),
	.w2(32'hba8a9728),
	.w3(32'hbba74150),
	.w4(32'hbbf02d4f),
	.w5(32'hbc2aded8),
	.w6(32'hbb5dc885),
	.w7(32'hbb063230),
	.w8(32'hbc373492),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e0fca),
	.w1(32'h3bf84394),
	.w2(32'h39d5cd11),
	.w3(32'h3d07a761),
	.w4(32'h3cffb6b4),
	.w5(32'hba584e0c),
	.w6(32'h3ce66940),
	.w7(32'h3c87565b),
	.w8(32'h39ed1161),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9498bd),
	.w1(32'hb96506a1),
	.w2(32'hbaa00b2e),
	.w3(32'h3b0d8db7),
	.w4(32'hbab3fc59),
	.w5(32'h3af457dc),
	.w6(32'hbb477ab8),
	.w7(32'hba0f82ee),
	.w8(32'h3b6f5e98),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1703fd),
	.w1(32'h3b110ff4),
	.w2(32'hbbf7565e),
	.w3(32'h3ad3a3b8),
	.w4(32'hbaf2d5d1),
	.w5(32'hbc37c820),
	.w6(32'h3ba3ca92),
	.w7(32'h3b466fa1),
	.w8(32'hbb34a579),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebbca1),
	.w1(32'hbb91f1e4),
	.w2(32'hbb50ecde),
	.w3(32'hbc2ffab6),
	.w4(32'hbb8fc240),
	.w5(32'h3a8de80f),
	.w6(32'hbaa69aa1),
	.w7(32'hb9d4402b),
	.w8(32'h3c4d0680),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5f2d4),
	.w1(32'h3a9cf7b4),
	.w2(32'hba549dc5),
	.w3(32'h3c0df6f2),
	.w4(32'hbba87e5c),
	.w5(32'hbb59d5bb),
	.w6(32'h3b8b0970),
	.w7(32'hbc7f4bfc),
	.w8(32'hba36ff30),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3699e),
	.w1(32'h3b4237eb),
	.w2(32'h3ab4e1c1),
	.w3(32'h3c21a6bc),
	.w4(32'h3c81db75),
	.w5(32'hbbe97ec6),
	.w6(32'h3cc3d01b),
	.w7(32'h3ca9be34),
	.w8(32'hbbe1855b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c1daa),
	.w1(32'h3bda436a),
	.w2(32'h3baff7db),
	.w3(32'hbbf08a14),
	.w4(32'hbb850da6),
	.w5(32'hbc54f10b),
	.w6(32'h3b9d1fdf),
	.w7(32'hbb818fd6),
	.w8(32'hbaa951fb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aee72),
	.w1(32'hbc045e2a),
	.w2(32'h3be0f8b7),
	.w3(32'h3931e88b),
	.w4(32'hbc40f829),
	.w5(32'h3bfafbbc),
	.w6(32'h3b04413d),
	.w7(32'hbc284c75),
	.w8(32'h3b7fc6cd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499f8b),
	.w1(32'h3b259344),
	.w2(32'hbbf4199e),
	.w3(32'hbb9f9621),
	.w4(32'h3b148d89),
	.w5(32'hbbe5ed04),
	.w6(32'hbb814d27),
	.w7(32'h3b303b27),
	.w8(32'hbb90a616),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb951bff),
	.w1(32'hbbd6530b),
	.w2(32'hbb5d91a3),
	.w3(32'hbbf13e7d),
	.w4(32'hbc0cce6e),
	.w5(32'h3af07187),
	.w6(32'hbb76e438),
	.w7(32'hbb94f77f),
	.w8(32'hbb516448),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092e90),
	.w1(32'h38a7d6d4),
	.w2(32'h3bb3113f),
	.w3(32'h3ad68e13),
	.w4(32'h3b73c89a),
	.w5(32'hbac6233b),
	.w6(32'hba84c4f6),
	.w7(32'hb9ccd650),
	.w8(32'hbb2f2556),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ff7b2),
	.w1(32'hbc37db25),
	.w2(32'hbc16e1ab),
	.w3(32'hbc948a18),
	.w4(32'hbc25dfb5),
	.w5(32'hbc03e54d),
	.w6(32'hbc2d7ea9),
	.w7(32'hbb12dc2b),
	.w8(32'hbbdc5397),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e7d60),
	.w1(32'hbc62d615),
	.w2(32'h3c99b710),
	.w3(32'h3a0a440f),
	.w4(32'h3a201c80),
	.w5(32'h3ccb28f9),
	.w6(32'h3b95cd60),
	.w7(32'h3bd5c893),
	.w8(32'h3c8c03c2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff2246),
	.w1(32'h3ae1ab8c),
	.w2(32'hbc8d9301),
	.w3(32'h3bcdf2f3),
	.w4(32'hba975807),
	.w5(32'hbc9712a9),
	.w6(32'hbad63dda),
	.w7(32'hbb329d18),
	.w8(32'hbc83d09e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85eb36),
	.w1(32'hbc713131),
	.w2(32'hbb7bf167),
	.w3(32'hbc83218b),
	.w4(32'hbc7c6f3d),
	.w5(32'hbb30af58),
	.w6(32'hbc43326a),
	.w7(32'hbc525310),
	.w8(32'hb9b398bd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca960),
	.w1(32'hbbb26e78),
	.w2(32'hbc34b388),
	.w3(32'hbaaf7b05),
	.w4(32'h3ae3d044),
	.w5(32'hbc54d6f3),
	.w6(32'h3b430c6f),
	.w7(32'h3b86e1eb),
	.w8(32'hbc4db234),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb343a07),
	.w1(32'hbba71ff0),
	.w2(32'h3b85c8f5),
	.w3(32'hbc831808),
	.w4(32'hbbaaf60e),
	.w5(32'hbc8051c8),
	.w6(32'hbc0cfe89),
	.w7(32'hbb9328b2),
	.w8(32'hbc583e4c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fd3e1),
	.w1(32'hbc7985c6),
	.w2(32'h3ba01056),
	.w3(32'hbcfb7fc6),
	.w4(32'hbceb4090),
	.w5(32'h3b2e0382),
	.w6(32'hbcd73156),
	.w7(32'hbc98e75e),
	.w8(32'h3c93b032),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d42ad79),
	.w1(32'h3cc8f495),
	.w2(32'hbaf45c76),
	.w3(32'h3d8d6c49),
	.w4(32'h3d0f6f39),
	.w5(32'hba66c202),
	.w6(32'h3d47e7c7),
	.w7(32'h3cdc9087),
	.w8(32'hbb1e24e3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761dbc),
	.w1(32'h3b95ea7e),
	.w2(32'hbb27cf82),
	.w3(32'h3b1f3418),
	.w4(32'h3c48acff),
	.w5(32'hbc5147e2),
	.w6(32'h3b619e57),
	.w7(32'h3a158ad1),
	.w8(32'hbc2a0605),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa39a9),
	.w1(32'hbb35ac12),
	.w2(32'hbb95537d),
	.w3(32'hba091abe),
	.w4(32'h3bb74b58),
	.w5(32'hbc1340d7),
	.w6(32'hbb73a22c),
	.w7(32'hbc2178bf),
	.w8(32'hbc0316bf),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33bc2b),
	.w1(32'h3aac9f59),
	.w2(32'hbb1c6c60),
	.w3(32'hbc1da398),
	.w4(32'h3ba0c9af),
	.w5(32'hbbf39e41),
	.w6(32'hbb959d67),
	.w7(32'h3b82b231),
	.w8(32'hbbe87148),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fa842),
	.w1(32'h3bfad28b),
	.w2(32'hbc64a19c),
	.w3(32'h3af57fbf),
	.w4(32'hbb9a53ec),
	.w5(32'hbc179a9e),
	.w6(32'h3b5b7783),
	.w7(32'hb90b59d4),
	.w8(32'hbc52497a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a2ad),
	.w1(32'hbb6cf206),
	.w2(32'h3c102f1e),
	.w3(32'h3a88d766),
	.w4(32'hbb8f5f9b),
	.w5(32'hba8aaa1e),
	.w6(32'h39dd478b),
	.w7(32'h3b013780),
	.w8(32'hbb8a2e03),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f7c4),
	.w1(32'h3aacb629),
	.w2(32'h3b82bead),
	.w3(32'hbc59edfe),
	.w4(32'hba5a0ade),
	.w5(32'h3bb8a140),
	.w6(32'hbbe6b179),
	.w7(32'hbb8b9bc0),
	.w8(32'h3a73ff48),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c840),
	.w1(32'h3b58c377),
	.w2(32'hbb55f308),
	.w3(32'h3bbdfca6),
	.w4(32'h3b8d6dd9),
	.w5(32'h3a5c6e7a),
	.w6(32'h3a9be426),
	.w7(32'h3bde8dcd),
	.w8(32'h3b511aae),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e960a),
	.w1(32'h3b01a2d5),
	.w2(32'h3bdc0cae),
	.w3(32'h3aaf78be),
	.w4(32'h3b8cebf9),
	.w5(32'h3c0ec602),
	.w6(32'hba8bd9e1),
	.w7(32'h3b880aa2),
	.w8(32'h3a301fd6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b4b0e),
	.w1(32'hbb0144c6),
	.w2(32'h3b4ab24a),
	.w3(32'hbb8ba34b),
	.w4(32'hbb8f1663),
	.w5(32'h3b73d3b5),
	.w6(32'hbbc3f61b),
	.w7(32'hbafb2614),
	.w8(32'h3acf1b29),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9526ae),
	.w1(32'hbad257b2),
	.w2(32'hba6b3acd),
	.w3(32'hba0289e0),
	.w4(32'hbba1fc17),
	.w5(32'hbb61fc28),
	.w6(32'h3aad8822),
	.w7(32'hbb8a0f31),
	.w8(32'hbab0be14),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08b026),
	.w1(32'h3b94970e),
	.w2(32'hbbed4618),
	.w3(32'h3bc8fa25),
	.w4(32'h3b9d9b68),
	.w5(32'hbc0fec6c),
	.w6(32'h3b84c36b),
	.w7(32'h3b5769de),
	.w8(32'hbb9b5605),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23aa59),
	.w1(32'h3bb46116),
	.w2(32'hbb88f7aa),
	.w3(32'hbae99af2),
	.w4(32'hbc84ebb6),
	.w5(32'hbc935f14),
	.w6(32'h3ae6891d),
	.w7(32'hbc6d430e),
	.w8(32'hbb8bcc4f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75afff),
	.w1(32'h3c0d4da9),
	.w2(32'hbb07d13c),
	.w3(32'h3bc5be41),
	.w4(32'h3bfe85c3),
	.w5(32'h39755bb7),
	.w6(32'h3c53004a),
	.w7(32'h3c11e053),
	.w8(32'h3ad20818),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bc2c9),
	.w1(32'h3c0bf0f3),
	.w2(32'hb9b31087),
	.w3(32'h3c3c977d),
	.w4(32'h3b832d87),
	.w5(32'hbc2e5780),
	.w6(32'h3c074957),
	.w7(32'h3b9a7ac5),
	.w8(32'hba86ebfb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841b1b),
	.w1(32'hbab78447),
	.w2(32'h3c22f047),
	.w3(32'hbc11ad47),
	.w4(32'hba4035ae),
	.w5(32'hbbb60136),
	.w6(32'hb9dc43bb),
	.w7(32'hba8d14f0),
	.w8(32'hbc1889df),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc289f0),
	.w1(32'h3c81d7d1),
	.w2(32'hbb7e5a25),
	.w3(32'h3c65853d),
	.w4(32'h3d2d20c8),
	.w5(32'hbc2c0198),
	.w6(32'h3c84b675),
	.w7(32'h3ccc7765),
	.w8(32'hbc3d13d1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc055efd),
	.w1(32'hbbcac0a3),
	.w2(32'h3bcc4c52),
	.w3(32'h3b567a22),
	.w4(32'h3bdf0361),
	.w5(32'hbc0d4869),
	.w6(32'h3c517a1c),
	.w7(32'h3b07c802),
	.w8(32'hbc19e0e9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2fdef),
	.w1(32'h3c2dc7fa),
	.w2(32'hba820149),
	.w3(32'hbc1fc8cc),
	.w4(32'h3cab433b),
	.w5(32'h3a9f7463),
	.w6(32'hbc119cdf),
	.w7(32'h3c61f6a5),
	.w8(32'h3be3b0d3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9f9b0),
	.w1(32'h3bcde077),
	.w2(32'h38b7fa89),
	.w3(32'h3c06fc86),
	.w4(32'h3bb8c225),
	.w5(32'h3baf57fb),
	.w6(32'h3c269cd8),
	.w7(32'h3be90265),
	.w8(32'h3bc227dc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cb6c6),
	.w1(32'hba11a1e3),
	.w2(32'h3b6efc51),
	.w3(32'h3be54944),
	.w4(32'h3b6c8de0),
	.w5(32'hbb2a6cb0),
	.w6(32'h3b531cf2),
	.w7(32'h3b88324e),
	.w8(32'h3b53336c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff01e8),
	.w1(32'h3b845c72),
	.w2(32'hbbab3bbc),
	.w3(32'h3acf77a3),
	.w4(32'hbb17c012),
	.w5(32'h3a32a7a0),
	.w6(32'h3a5c40bb),
	.w7(32'hbb4be99d),
	.w8(32'hb99d11af),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3afb95),
	.w1(32'h3b36fa2a),
	.w2(32'hbb639321),
	.w3(32'hbc286934),
	.w4(32'hbbc813ce),
	.w5(32'hbc0cd0ce),
	.w6(32'hbc48e83b),
	.w7(32'hbba9593a),
	.w8(32'hbb47b826),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb438363),
	.w1(32'h3b32f669),
	.w2(32'hbbea2679),
	.w3(32'hbafce92b),
	.w4(32'hb9d51dd6),
	.w5(32'hbc02cc9c),
	.w6(32'h3beb426a),
	.w7(32'hbb00c87e),
	.w8(32'hbb7facd5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80df15),
	.w1(32'hbb4bed33),
	.w2(32'hbc36f706),
	.w3(32'hbc26f3e3),
	.w4(32'hbbbd1e2c),
	.w5(32'hbc0970f8),
	.w6(32'hbb6811d6),
	.w7(32'hbbe186e0),
	.w8(32'hbc010714),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f30e4),
	.w1(32'hbb0d1304),
	.w2(32'hbb71b887),
	.w3(32'hbb084261),
	.w4(32'hb987bed5),
	.w5(32'hbb969263),
	.w6(32'hbb15ebd1),
	.w7(32'h38bf13dc),
	.w8(32'hbaadb85f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba041311),
	.w1(32'h3a990aa6),
	.w2(32'hbbd8c193),
	.w3(32'hbae85799),
	.w4(32'h3aecdfb9),
	.w5(32'hbbca5a91),
	.w6(32'h3a6fa9e0),
	.w7(32'h3b0e2a2e),
	.w8(32'h3aa167cd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aae83),
	.w1(32'h3c1a44a0),
	.w2(32'h3bc4a78a),
	.w3(32'hbccca81f),
	.w4(32'h3c6d6dd2),
	.w5(32'h3b8ecb5c),
	.w6(32'hbc0f01df),
	.w7(32'h3cbc9de5),
	.w8(32'h3a7594ae),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b590d32),
	.w1(32'hba06aa45),
	.w2(32'h3baf4fa4),
	.w3(32'h3b49df67),
	.w4(32'hba3de2e3),
	.w5(32'h3bb4c53c),
	.w6(32'h3a86ab0b),
	.w7(32'hba8c8e5a),
	.w8(32'h3b8aef46),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd840f),
	.w1(32'h3afe9004),
	.w2(32'h3c1b3313),
	.w3(32'h3ced2fb0),
	.w4(32'h3bacf6b9),
	.w5(32'h3ba5213c),
	.w6(32'h3ccbec79),
	.w7(32'hbb8ae129),
	.w8(32'h3c0af0a8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd6fb8),
	.w1(32'hbb8506ce),
	.w2(32'hbc230aa2),
	.w3(32'hbb820f7b),
	.w4(32'hb9e44602),
	.w5(32'hbbb567f1),
	.w6(32'h3a894f08),
	.w7(32'hbba80d63),
	.w8(32'hbaf86066),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829096),
	.w1(32'h3a80c54d),
	.w2(32'h3b16b535),
	.w3(32'hbba8a205),
	.w4(32'hbaf537d3),
	.w5(32'hbbdf2f0d),
	.w6(32'h3a989258),
	.w7(32'hbbc17d0a),
	.w8(32'h3b85a062),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule