module layer_10_featuremap_183(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77ebd6b),
	.w1(32'hb6e63564),
	.w2(32'h36ec2e62),
	.w3(32'hb7e6c40e),
	.w4(32'h36d84601),
	.w5(32'h3795706b),
	.w6(32'hb7f90ea0),
	.w7(32'h371af6c6),
	.w8(32'h359073ea),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72298b),
	.w1(32'hbad14bbf),
	.w2(32'hbb37a161),
	.w3(32'hb956bca4),
	.w4(32'hbae23863),
	.w5(32'hbaef6f19),
	.w6(32'hbae2eab0),
	.w7(32'hbac04468),
	.w8(32'hbaf77014),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb691b603),
	.w1(32'hb74a077f),
	.w2(32'hb7946087),
	.w3(32'hb61abf5a),
	.w4(32'hb7065e96),
	.w5(32'hb783a4e3),
	.w6(32'hb75ca97c),
	.w7(32'hb76f52c7),
	.w8(32'hb787a7d7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb828bbe6),
	.w1(32'hba1d7707),
	.w2(32'h397f1005),
	.w3(32'hb996a123),
	.w4(32'hba2739c9),
	.w5(32'hb92f7da8),
	.w6(32'hb9501b5b),
	.w7(32'hba24171c),
	.w8(32'hb96fed9d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca658a),
	.w1(32'hb8622119),
	.w2(32'h381982a6),
	.w3(32'hb9132fb6),
	.w4(32'hb89ed7b7),
	.w5(32'hb705010a),
	.w6(32'hb8fdf5f3),
	.w7(32'hb8b8fbdf),
	.w8(32'hb7862179),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fb2da),
	.w1(32'h383f5cf0),
	.w2(32'h379f862c),
	.w3(32'h374c6372),
	.w4(32'h36fe1ac0),
	.w5(32'hb71d0861),
	.w6(32'hb734d6aa),
	.w7(32'hb8244723),
	.w8(32'hb853e9ce),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0695),
	.w1(32'hbac08cef),
	.w2(32'h39ad4fde),
	.w3(32'hbae6e1a4),
	.w4(32'hba1d9ae7),
	.w5(32'h3a8fc35d),
	.w6(32'hbb0ee2a7),
	.w7(32'h38b6f680),
	.w8(32'h3b1752b4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87dc23),
	.w1(32'h3b6202d6),
	.w2(32'h3bc6d1e2),
	.w3(32'h3bcf8bc1),
	.w4(32'h3bcb9be9),
	.w5(32'h3baceddd),
	.w6(32'h3bf8b618),
	.w7(32'h3bd1af39),
	.w8(32'h3b7e3817),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b19191),
	.w1(32'h3a328969),
	.w2(32'h3a5960f3),
	.w3(32'h3a924435),
	.w4(32'h3a8f0970),
	.w5(32'h3a84d558),
	.w6(32'h3a8bcd1d),
	.w7(32'h3a8ae227),
	.w8(32'h3aa6a401),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ac067),
	.w1(32'hbb62dd88),
	.w2(32'hbb2e82f5),
	.w3(32'h3ab65759),
	.w4(32'hbafcf0df),
	.w5(32'hba980c6c),
	.w6(32'h38d4874a),
	.w7(32'hbac71e0e),
	.w8(32'hb9ea4469),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38531aa7),
	.w1(32'hb970b3d2),
	.w2(32'h396c9fbc),
	.w3(32'h398b3da9),
	.w4(32'hb9038c88),
	.w5(32'hb88ef542),
	.w6(32'h38831bb6),
	.w7(32'hb9f77a73),
	.w8(32'hb885149d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b00e),
	.w1(32'hba9adf37),
	.w2(32'h3afa1d34),
	.w3(32'hbb5215e3),
	.w4(32'hbb370be0),
	.w5(32'h3947d16a),
	.w6(32'hbb56f75c),
	.w7(32'hbb540025),
	.w8(32'h3a3b878d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ef4c3),
	.w1(32'hbb36b736),
	.w2(32'hbb2a806f),
	.w3(32'h39d3a3d6),
	.w4(32'hbaa9cc9e),
	.w5(32'hba8a88fd),
	.w6(32'hb8e13533),
	.w7(32'h39294f12),
	.w8(32'h39e0c97f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaedeb3),
	.w1(32'hbabbe669),
	.w2(32'hb904ace9),
	.w3(32'h3a1dd5ca),
	.w4(32'h398f7e85),
	.w5(32'h38084ca2),
	.w6(32'h3a2e000b),
	.w7(32'h3a168952),
	.w8(32'h3a28b463),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ef71e),
	.w1(32'hbac9cccc),
	.w2(32'hbad69d2b),
	.w3(32'hba2234aa),
	.w4(32'hbaed67f0),
	.w5(32'hbaa02261),
	.w6(32'hbacb966a),
	.w7(32'hbae984a8),
	.w8(32'hbb1067fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e988f0),
	.w1(32'hbabb24b0),
	.w2(32'hbaeefbcb),
	.w3(32'h3b001c15),
	.w4(32'h39bafcc1),
	.w5(32'hb96fe242),
	.w6(32'h3b1d8804),
	.w7(32'h3adc47b2),
	.w8(32'h3a7c99af),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be53ca),
	.w1(32'hba81cfee),
	.w2(32'hba38c063),
	.w3(32'hb97cb14e),
	.w4(32'hba97e897),
	.w5(32'hba541b29),
	.w6(32'h39164172),
	.w7(32'hba73ba05),
	.w8(32'hba31e456),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af362b8),
	.w1(32'h3c1bc9a8),
	.w2(32'h3c3ac128),
	.w3(32'h3ba83508),
	.w4(32'h3c128c28),
	.w5(32'h3c1d6e61),
	.w6(32'h3bd73a13),
	.w7(32'h3bc190c3),
	.w8(32'h3bfa15c4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dbd87),
	.w1(32'h3b3b82c3),
	.w2(32'h3b5f1bea),
	.w3(32'h3b309c79),
	.w4(32'h3b7406fa),
	.w5(32'h3b59fd74),
	.w6(32'h3b45593b),
	.w7(32'h3b57504f),
	.w8(32'h3b33a465),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6417f79),
	.w1(32'hb7f5ac8c),
	.w2(32'hb87cc69b),
	.w3(32'hb8002ef5),
	.w4(32'hb80c68ac),
	.w5(32'hb86d1bd1),
	.w6(32'hb7dcbddd),
	.w7(32'hb717820a),
	.w8(32'hb7277b3d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec0f6d),
	.w1(32'h3825c0d2),
	.w2(32'hb843f878),
	.w3(32'hb6fd30a1),
	.w4(32'h38b842e6),
	.w5(32'h36dc91cf),
	.w6(32'h37943b8c),
	.w7(32'h38815a3a),
	.w8(32'hb8320e27),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179add),
	.w1(32'hba50f4a5),
	.w2(32'hba1bbed7),
	.w3(32'hba8ef513),
	.w4(32'hbab6e20a),
	.w5(32'hba70abcd),
	.w6(32'hbabf8de3),
	.w7(32'hbad257f9),
	.w8(32'hba8720c1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8412b3),
	.w1(32'h3c305e35),
	.w2(32'h3c71b890),
	.w3(32'h3c0b8ffe),
	.w4(32'h3c3cf336),
	.w5(32'h3c557a1f),
	.w6(32'h3c316267),
	.w7(32'h3bd4c143),
	.w8(32'h3c37cea9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f43dd),
	.w1(32'hbb48a1b8),
	.w2(32'hbbab6f90),
	.w3(32'hba4c96f1),
	.w4(32'hbb7bebb8),
	.w5(32'hbb8c24ec),
	.w6(32'hbb007308),
	.w7(32'hbb80e665),
	.w8(32'hbb8dddd7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7e397),
	.w1(32'hbae6e5a5),
	.w2(32'hbbc94639),
	.w3(32'hb9c5a39d),
	.w4(32'hbba0917f),
	.w5(32'hbbcf521e),
	.w6(32'hbaab74da),
	.w7(32'hbba366ab),
	.w8(32'hbb9b046f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f5966),
	.w1(32'hba310267),
	.w2(32'hb9d75d0c),
	.w3(32'h38c5fc81),
	.w4(32'hb9833953),
	.w5(32'hb8f9beae),
	.w6(32'h39a014be),
	.w7(32'hb90293c8),
	.w8(32'hb8312082),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8009af8),
	.w1(32'hb677f9e6),
	.w2(32'hb8f09a6a),
	.w3(32'hb89bd26f),
	.w4(32'hb8825311),
	.w5(32'hb90f1d00),
	.w6(32'hb91fc3f3),
	.w7(32'hb90c473f),
	.w8(32'hb9580668),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc22d9),
	.w1(32'hbb244aad),
	.w2(32'hbb369b3e),
	.w3(32'hbb03d79a),
	.w4(32'hbb7ff7fe),
	.w5(32'hbb2bbd40),
	.w6(32'hbb39c636),
	.w7(32'hbb520df9),
	.w8(32'hbae7abea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840862),
	.w1(32'hba35123b),
	.w2(32'hba699e3c),
	.w3(32'hbaf62d2f),
	.w4(32'hbab96243),
	.w5(32'hbad565f2),
	.w6(32'hbb37b966),
	.w7(32'hbb574a2e),
	.w8(32'hbb4fb540),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a82afd),
	.w1(32'hbb9b3d7e),
	.w2(32'hbbcaf0b3),
	.w3(32'hbaad63a2),
	.w4(32'hbb9d612d),
	.w5(32'hbba8302a),
	.w6(32'hbb5a1150),
	.w7(32'hbb953b37),
	.w8(32'hbb81f5c0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b8724c),
	.w1(32'hb89290da),
	.w2(32'hb905851e),
	.w3(32'hb85bd218),
	.w4(32'hb8dd639b),
	.w5(32'hb9097c5d),
	.w6(32'hb8b0932e),
	.w7(32'hb908bd4b),
	.w8(32'hb91d240d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38367dda),
	.w1(32'hb9915aa3),
	.w2(32'hb9bbd9fa),
	.w3(32'hb8304dca),
	.w4(32'hb9e58193),
	.w5(32'hba0e3969),
	.w6(32'hb90240c3),
	.w7(32'hba077a5a),
	.w8(32'hba122201),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38cfc2),
	.w1(32'hbaea3e9d),
	.w2(32'hbb1228bb),
	.w3(32'h3881f2ed),
	.w4(32'hba92bad9),
	.w5(32'hbae1b3a5),
	.w6(32'hb9ce32a4),
	.w7(32'hbae302e3),
	.w8(32'hbb239640),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaab6e5),
	.w1(32'hba394bd6),
	.w2(32'hbabac12e),
	.w3(32'h3a03ec67),
	.w4(32'hb9caa2cd),
	.w5(32'hbaa8c570),
	.w6(32'hb89f1723),
	.w7(32'hb9d81836),
	.w8(32'hba851ede),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d250f2),
	.w1(32'hb8ea9ea9),
	.w2(32'hb9290606),
	.w3(32'hb8a720dc),
	.w4(32'hb88969ea),
	.w5(32'hb8b7a995),
	.w6(32'hb8e0bc74),
	.w7(32'h3987285a),
	.w8(32'h391792c8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba750e4a),
	.w1(32'hba6a34c7),
	.w2(32'h3893332c),
	.w3(32'hb9867a2d),
	.w4(32'hba3dd905),
	.w5(32'h381b1ba5),
	.w6(32'h383b8d48),
	.w7(32'hba234def),
	.w8(32'h39b4c6ad),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cfc97),
	.w1(32'hbb920b6b),
	.w2(32'h3b1920b7),
	.w3(32'hb99ed0f7),
	.w4(32'hbb4c93f7),
	.w5(32'hbb20fa72),
	.w6(32'h38c2d537),
	.w7(32'hbb437f5b),
	.w8(32'h3aab848e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc49f),
	.w1(32'hbb8815ed),
	.w2(32'hbbf50151),
	.w3(32'hbb875a30),
	.w4(32'hbc2e292b),
	.w5(32'hbc00e958),
	.w6(32'hbc1f65ef),
	.w7(32'hbc4c0d01),
	.w8(32'hbc20fffa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83890f),
	.w1(32'hbbbddb21),
	.w2(32'hbbbcb9a8),
	.w3(32'hbbd5b06d),
	.w4(32'hbc1562a6),
	.w5(32'hbbbfa431),
	.w6(32'hbc33e5d8),
	.w7(32'hbc0df253),
	.w8(32'hbbb9aedc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e88a30),
	.w1(32'hba291029),
	.w2(32'hba75d517),
	.w3(32'hba016ee2),
	.w4(32'hbaaabca9),
	.w5(32'hbaa4d118),
	.w6(32'hba871752),
	.w7(32'hbada129e),
	.w8(32'hbaeb2cd9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04e2ea),
	.w1(32'h3a069987),
	.w2(32'h3a3eabc6),
	.w3(32'h3a27343b),
	.w4(32'h3a005d92),
	.w5(32'h3a214e5d),
	.w6(32'h3a23806d),
	.w7(32'h39305f58),
	.w8(32'h39f87c4f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9933e93),
	.w1(32'hb84ebfe3),
	.w2(32'hb8474403),
	.w3(32'hb98f9197),
	.w4(32'hb8703c76),
	.w5(32'hb7a9e439),
	.w6(32'hb967c788),
	.w7(32'h37c8f370),
	.w8(32'h36ffd70f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8adce68),
	.w1(32'hba91edb3),
	.w2(32'hb9a2ade6),
	.w3(32'hb9b24906),
	.w4(32'hba884e0a),
	.w5(32'hb8fdb64c),
	.w6(32'h39b06d41),
	.w7(32'hb8af1ff0),
	.w8(32'h3a4e59ca),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb047c4d),
	.w1(32'hbad57fe2),
	.w2(32'h399354e1),
	.w3(32'h3ad3b806),
	.w4(32'h3b16b8c0),
	.w5(32'h3b01fdca),
	.w6(32'h3ab03182),
	.w7(32'h3a0c0675),
	.w8(32'h3a915395),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab26b08),
	.w1(32'hbb51357f),
	.w2(32'hbb7cf0aa),
	.w3(32'h38ce27dd),
	.w4(32'hbb61c6ae),
	.w5(32'hbb4a129d),
	.w6(32'hbb01edf4),
	.w7(32'hbb87d39b),
	.w8(32'hbb62cbc6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cd61a),
	.w1(32'hbb3d2d49),
	.w2(32'hbb9500bb),
	.w3(32'hb8268593),
	.w4(32'hbb3c6687),
	.w5(32'hbb47a1cb),
	.w6(32'hb9f2df03),
	.w7(32'hbb282eb9),
	.w8(32'hbb4d3aa3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cff53),
	.w1(32'h3acdcfa6),
	.w2(32'h3b39a9e4),
	.w3(32'h3b5c9c5d),
	.w4(32'h3b2ba19f),
	.w5(32'h3b160052),
	.w6(32'h3ba14184),
	.w7(32'h3b15cdf5),
	.w8(32'h3b1696ca),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9848d),
	.w1(32'h3c0d163a),
	.w2(32'h3c6aed62),
	.w3(32'h3bb765c1),
	.w4(32'h3c2bf28b),
	.w5(32'h3c490ec1),
	.w6(32'h3c072309),
	.w7(32'h3c11051d),
	.w8(32'h3c3fc93b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f026f),
	.w1(32'hb9800286),
	.w2(32'h3a75bbd1),
	.w3(32'hb9cad8d0),
	.w4(32'h39b4a917),
	.w5(32'h3a0fc747),
	.w6(32'hb937f3f2),
	.w7(32'h3801ad5e),
	.w8(32'h3a159767),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a060e02),
	.w1(32'h3b065d32),
	.w2(32'h3b2e4595),
	.w3(32'h3a9fc12d),
	.w4(32'h3b1c44f9),
	.w5(32'h3b3ce9af),
	.w6(32'h3b1477aa),
	.w7(32'h3b528814),
	.w8(32'h3b79a4dc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8391a0),
	.w1(32'hb91afe98),
	.w2(32'h39ace8f7),
	.w3(32'hba85b140),
	.w4(32'hb98fcd06),
	.w5(32'hb922ce07),
	.w6(32'hba391176),
	.w7(32'hb91ea250),
	.w8(32'h398fd695),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eea53),
	.w1(32'h3a2b291c),
	.w2(32'hb978a50b),
	.w3(32'h3aa0f0ae),
	.w4(32'hb908ab24),
	.w5(32'h38f9ea5f),
	.w6(32'h3a5a5093),
	.w7(32'hb9bd1eb7),
	.w8(32'h39eef904),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c5b56),
	.w1(32'h3aa257cb),
	.w2(32'h3acbaac7),
	.w3(32'h3a8a4746),
	.w4(32'h3aa87c77),
	.w5(32'h3a994bac),
	.w6(32'h3acb1fb4),
	.w7(32'h3a9527e8),
	.w8(32'h3a8f6db1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a05e5),
	.w1(32'h3bcbaded),
	.w2(32'h3c024c50),
	.w3(32'h3b5d67f4),
	.w4(32'h3bcfe635),
	.w5(32'h3bb1e2cc),
	.w6(32'h3b82ce0d),
	.w7(32'h3ba72614),
	.w8(32'h3b8fa037),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d5170),
	.w1(32'h3ab3cbc6),
	.w2(32'h3ac7356a),
	.w3(32'h38caf070),
	.w4(32'h3a01f999),
	.w5(32'h3a91a955),
	.w6(32'h37eb44f2),
	.w7(32'h38390f3a),
	.w8(32'h3a00c20a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8959ec2),
	.w1(32'hb8d7d3b7),
	.w2(32'hb8a9eaa0),
	.w3(32'hb84323a7),
	.w4(32'hb89b16bb),
	.w5(32'hb888397b),
	.w6(32'h3810a3bd),
	.w7(32'h3650e0b6),
	.w8(32'h37eb1657),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a81085),
	.w1(32'h34f84f34),
	.w2(32'hb7e5d2b3),
	.w3(32'hb6b2505f),
	.w4(32'hb7537740),
	.w5(32'hb7cd044c),
	.w6(32'hb7a0ec08),
	.w7(32'hb7eb69db),
	.w8(32'hb7aaed3e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f6670),
	.w1(32'h37e15ac4),
	.w2(32'hb8d1890c),
	.w3(32'hb925db42),
	.w4(32'hb7958db7),
	.w5(32'hb85c06cc),
	.w6(32'hb95db1a9),
	.w7(32'hb8992c30),
	.w8(32'hb8e4da82),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba241862),
	.w1(32'hba894bc7),
	.w2(32'hba5c1335),
	.w3(32'hba623735),
	.w4(32'hba9be330),
	.w5(32'hba36f264),
	.w6(32'hba24c2e1),
	.w7(32'hba54e34a),
	.w8(32'hb9d4558d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05dfdf),
	.w1(32'hb9cb9b1a),
	.w2(32'hb8e3ca0e),
	.w3(32'hb9b0652e),
	.w4(32'hb9bcc17c),
	.w5(32'h39234527),
	.w6(32'hba364907),
	.w7(32'hb9b355b5),
	.w8(32'hb8aa9a43),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e09970),
	.w1(32'h3b151942),
	.w2(32'h3b6a274b),
	.w3(32'h3ad362b8),
	.w4(32'h3b1d8796),
	.w5(32'h3b460011),
	.w6(32'h3b0a4e48),
	.w7(32'h3b261a3d),
	.w8(32'h3b529555),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080650),
	.w1(32'h3b79dbcc),
	.w2(32'h3b432852),
	.w3(32'h3b9e41eb),
	.w4(32'h3b7e51d1),
	.w5(32'h3b967f6f),
	.w6(32'h3b9c245e),
	.w7(32'h3b5874d9),
	.w8(32'h3b801fc0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d14729),
	.w1(32'h3872a2c0),
	.w2(32'h389a357f),
	.w3(32'h38be188b),
	.w4(32'h37d57ef3),
	.w5(32'hb8943d4c),
	.w6(32'h38a5847f),
	.w7(32'h387be3bc),
	.w8(32'hb8ffa33e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb796613a),
	.w1(32'hb3959b8a),
	.w2(32'hb7aded48),
	.w3(32'hb4e86494),
	.w4(32'h375121b0),
	.w5(32'hb7645486),
	.w6(32'h373d2661),
	.w7(32'h377c3015),
	.w8(32'hb73fcb0b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869bf25),
	.w1(32'hb8eca731),
	.w2(32'hb93fea6d),
	.w3(32'hb842a8f1),
	.w4(32'hb7e3c618),
	.w5(32'hb9265bf5),
	.w6(32'hb8f1cec8),
	.w7(32'hb92a2bac),
	.w8(32'hb9293b6c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7685800),
	.w1(32'hb5e9f7fd),
	.w2(32'hb89e7867),
	.w3(32'hb81ea727),
	.w4(32'hb8081471),
	.w5(32'hb8a2c809),
	.w6(32'hb7efe3ff),
	.w7(32'hb83edb99),
	.w8(32'hb8d60540),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ada32),
	.w1(32'h3abfb121),
	.w2(32'h3a717339),
	.w3(32'hb9fb6cba),
	.w4(32'h3a8941af),
	.w5(32'h3990bf49),
	.w6(32'h3a455b9f),
	.w7(32'h3b061193),
	.w8(32'h3a97dc28),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace0de8),
	.w1(32'hbaebd1b7),
	.w2(32'hbb4ef3d1),
	.w3(32'hba3da132),
	.w4(32'hbb27951b),
	.w5(32'hbaa80d5c),
	.w6(32'hba4d04ca),
	.w7(32'hbb26b3e6),
	.w8(32'hbaee7632),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585253),
	.w1(32'h3bd5981b),
	.w2(32'h3bc6be65),
	.w3(32'h3b3efb69),
	.w4(32'h3b4f4597),
	.w5(32'h3bbe84b4),
	.w6(32'h3bab440a),
	.w7(32'h3b7d813a),
	.w8(32'h3bbbbbc5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b588d36),
	.w1(32'hbb886bb1),
	.w2(32'hbc0ece08),
	.w3(32'hbafdb31c),
	.w4(32'hbc0c6c31),
	.w5(32'hbc2a6b6b),
	.w6(32'hbb5566cb),
	.w7(32'hbbd27a7a),
	.w8(32'hbc0bb5ec),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e0d816),
	.w1(32'h36bbd5f1),
	.w2(32'hb7fd66ea),
	.w3(32'hb69c3706),
	.w4(32'h37d2a49d),
	.w5(32'hb6c12f40),
	.w6(32'h37eadd42),
	.w7(32'h383493a3),
	.w8(32'hb6d6b87d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f63b5a),
	.w1(32'hb71471d9),
	.w2(32'hb8c38157),
	.w3(32'hb73e6491),
	.w4(32'hb60433c5),
	.w5(32'hb8a1454f),
	.w6(32'hb51d2686),
	.w7(32'h3719b098),
	.w8(32'hb88b8eb2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88331bc),
	.w1(32'h365b6b36),
	.w2(32'hb84d5a81),
	.w3(32'hb7913be5),
	.w4(32'h3713dc24),
	.w5(32'hb840ccc9),
	.w6(32'hb7347eaf),
	.w7(32'h38915523),
	.w8(32'h3812041d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3726051a),
	.w1(32'h3a84e110),
	.w2(32'h3af3d082),
	.w3(32'h3996efdd),
	.w4(32'h3a88cd4c),
	.w5(32'h3ad18a53),
	.w6(32'h3aa2e172),
	.w7(32'h3ad79623),
	.w8(32'h3aebaee0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914deb3),
	.w1(32'h384c3bd4),
	.w2(32'h38f4d5d8),
	.w3(32'hb9050d0b),
	.w4(32'h38d7357d),
	.w5(32'h39433468),
	.w6(32'hb8a32d63),
	.w7(32'h392268ca),
	.w8(32'h39106c2b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ef237),
	.w1(32'h3ba6fc31),
	.w2(32'h3bd23fe0),
	.w3(32'h3b1ea6eb),
	.w4(32'h3b99cecd),
	.w5(32'h3b37bf06),
	.w6(32'h3b4cb6c6),
	.w7(32'h3b69bcc1),
	.w8(32'h3b1d5238),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96bda2e),
	.w1(32'h3b910f28),
	.w2(32'h3be9f9a7),
	.w3(32'h3b889266),
	.w4(32'h3c0636a5),
	.w5(32'h3bdece90),
	.w6(32'h3b7a577b),
	.w7(32'h3bedbc73),
	.w8(32'h3bb4a5ab),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bd413),
	.w1(32'hbb65fd07),
	.w2(32'hbb8ec7c9),
	.w3(32'hba2074ef),
	.w4(32'hbb74272c),
	.w5(32'hbb5376ab),
	.w6(32'hbb2e058c),
	.w7(32'hbb614b53),
	.w8(32'hbb58cf6a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b64266),
	.w1(32'h3a965bac),
	.w2(32'h3ab3548c),
	.w3(32'h3acc5152),
	.w4(32'h3ad0031b),
	.w5(32'h3acf6e26),
	.w6(32'h3ad4a50f),
	.w7(32'h3ae67f48),
	.w8(32'h3ad54d38),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b250df),
	.w1(32'h3a1284de),
	.w2(32'hb8ec87b6),
	.w3(32'h3a02d614),
	.w4(32'hb9f55582),
	.w5(32'hba2138ee),
	.w6(32'h3a3f7e7d),
	.w7(32'h3a101cac),
	.w8(32'h3a851bf9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f81d98),
	.w1(32'hba8101a5),
	.w2(32'hbab32285),
	.w3(32'h382b2b69),
	.w4(32'hbacc61c9),
	.w5(32'hba9c2b37),
	.w6(32'hb9b79afc),
	.w7(32'hbad2c96f),
	.w8(32'hbaab7044),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e484b6),
	.w1(32'h3b349165),
	.w2(32'h3b840195),
	.w3(32'h3a8dabfb),
	.w4(32'h3b3a80ca),
	.w5(32'h3b554ad7),
	.w6(32'h3b2a7a67),
	.w7(32'h3b1fb12e),
	.w8(32'h3b499447),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366fdc95),
	.w1(32'h363633dd),
	.w2(32'hb7a19254),
	.w3(32'h3734ad30),
	.w4(32'hb5d2ebb0),
	.w5(32'hb7f76666),
	.w6(32'h3760cd72),
	.w7(32'h35ae1f89),
	.w8(32'hb8173378),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b7f13d),
	.w1(32'hb7910fe2),
	.w2(32'hb7ebd495),
	.w3(32'hb71c2e77),
	.w4(32'hb74dc08c),
	.w5(32'hb7825e6a),
	.w6(32'h34195a22),
	.w7(32'h37172686),
	.w8(32'hb6672861),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7271f73),
	.w1(32'hb96c03cc),
	.w2(32'hb9d3f51e),
	.w3(32'hb929d68b),
	.w4(32'hb9ac8e57),
	.w5(32'hb9cbe32c),
	.w6(32'hb9a2c20d),
	.w7(32'hb9af2af1),
	.w8(32'hb9c88a61),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6cd1e),
	.w1(32'h38b4518b),
	.w2(32'hb9128ba7),
	.w3(32'hb835291a),
	.w4(32'hb804795c),
	.w5(32'hb93af5b1),
	.w6(32'hb898052f),
	.w7(32'hb7f67148),
	.w8(32'hb8f05865),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0490a1),
	.w1(32'hba621170),
	.w2(32'hbb5708e2),
	.w3(32'hb90f8496),
	.w4(32'hbb5550de),
	.w5(32'hbb8183cf),
	.w6(32'hbae30ebb),
	.w7(32'hbb32518b),
	.w8(32'hbb728a13),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f924b),
	.w1(32'hb9594466),
	.w2(32'hb88b0756),
	.w3(32'hb7e177ac),
	.w4(32'hb83ae1bb),
	.w5(32'hb989264a),
	.w6(32'hb9559deb),
	.w7(32'hb9ee3c6d),
	.w8(32'hba09c696),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0248c2),
	.w1(32'h399f9d8b),
	.w2(32'hb965f453),
	.w3(32'h3a2e2b2e),
	.w4(32'hb9cf03c0),
	.w5(32'hba5ca844),
	.w6(32'h391f9c39),
	.w7(32'hba7374d2),
	.w8(32'hbac1d83f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1540fd),
	.w1(32'h3c159625),
	.w2(32'h3c1ad512),
	.w3(32'h3c0be8d8),
	.w4(32'h3c2de98c),
	.w5(32'h3bf465f2),
	.w6(32'h3c24f72e),
	.w7(32'h3c2e7b5e),
	.w8(32'h3bf8dfe1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a369679),
	.w1(32'hbaf531f4),
	.w2(32'hbad56f58),
	.w3(32'hbaedf97d),
	.w4(32'hbb567cc0),
	.w5(32'hbb35bcc0),
	.w6(32'hbb0e0d73),
	.w7(32'hbb4f2276),
	.w8(32'hbb21e48e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e23a8b),
	.w1(32'hbb0a6364),
	.w2(32'hb88fe4b7),
	.w3(32'h398c5f68),
	.w4(32'hb9e6a2da),
	.w5(32'hba36069d),
	.w6(32'h3a9c14a2),
	.w7(32'hbab9e768),
	.w8(32'h3aa57398),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bad60d),
	.w1(32'hbb299b89),
	.w2(32'hbb845ba6),
	.w3(32'hbaf545b0),
	.w4(32'hbb644188),
	.w5(32'hbb6d9f23),
	.w6(32'hbad80fb9),
	.w7(32'hbb8150aa),
	.w8(32'hbb56aebf),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d5678),
	.w1(32'h3abd8944),
	.w2(32'h3b2a3a6d),
	.w3(32'h3b141069),
	.w4(32'h3b266676),
	.w5(32'h3b1dbc20),
	.w6(32'h3af17531),
	.w7(32'h3af20a0b),
	.w8(32'h3b0ec11b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae78b50),
	.w1(32'h3a668989),
	.w2(32'hba30a7b6),
	.w3(32'h3983e077),
	.w4(32'hba5be207),
	.w5(32'hbaa4a29b),
	.w6(32'hb980a3d1),
	.w7(32'hb997a77a),
	.w8(32'h38f864be),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab55969),
	.w1(32'hbb1312e0),
	.w2(32'hbb2a401c),
	.w3(32'hbad526a3),
	.w4(32'hbb839b68),
	.w5(32'hbb651cc4),
	.w6(32'hbb3c4df2),
	.w7(32'hbb91c7a4),
	.w8(32'hbbaa00bc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac29c7d),
	.w1(32'hba2f8c1e),
	.w2(32'hba040c77),
	.w3(32'hba859394),
	.w4(32'hba4462c9),
	.w5(32'hbb08dfc0),
	.w6(32'hba3eaf81),
	.w7(32'hb9cfe582),
	.w8(32'hbae7646c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b58f9),
	.w1(32'h3a4ae464),
	.w2(32'h3b54cdc5),
	.w3(32'h3b05d719),
	.w4(32'h3b632d7b),
	.w5(32'h3b691d71),
	.w6(32'h3b0e73f6),
	.w7(32'h3b7c8367),
	.w8(32'h3b5c6b72),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cd8f1),
	.w1(32'hb9e7c184),
	.w2(32'h39b1917d),
	.w3(32'hb7f64039),
	.w4(32'hba511ba5),
	.w5(32'hb8038c6b),
	.w6(32'h3accc880),
	.w7(32'h3b0e9769),
	.w8(32'h3bab39d2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9ab54),
	.w1(32'h3b94df2f),
	.w2(32'h3c1994a2),
	.w3(32'h3b91471e),
	.w4(32'h3ba6f33d),
	.w5(32'h3b746ade),
	.w6(32'h3bd8f104),
	.w7(32'h3b22c4e4),
	.w8(32'h3b669a05),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae19441),
	.w1(32'hbbd6c07d),
	.w2(32'hbb3fde4b),
	.w3(32'hbb1cd710),
	.w4(32'hbc0c3d5f),
	.w5(32'hbb9f378f),
	.w6(32'hbadbde6d),
	.w7(32'hbb9bb121),
	.w8(32'hba4ad6f9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d9ab4),
	.w1(32'hbb346aea),
	.w2(32'hbbdae1aa),
	.w3(32'hba467aac),
	.w4(32'hbb3576ea),
	.w5(32'hbbb26854),
	.w6(32'hba9f0984),
	.w7(32'hbb1e9783),
	.w8(32'hbb9004a0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1709d3),
	.w1(32'hbac76903),
	.w2(32'h3b9d1dab),
	.w3(32'h380c8382),
	.w4(32'hba676bbe),
	.w5(32'h39acbab9),
	.w6(32'h3a329805),
	.w7(32'hbaaca616),
	.w8(32'h3b6b3340),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852104),
	.w1(32'hbb2afc0c),
	.w2(32'hb9d3a69a),
	.w3(32'hbb708c26),
	.w4(32'hbb28545d),
	.w5(32'hbb2aa5d3),
	.w6(32'hbb615b4b),
	.w7(32'hbb2ddd7c),
	.w8(32'hbb066b1f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f83ff),
	.w1(32'h3c0e9318),
	.w2(32'h3c972397),
	.w3(32'h3bb0c9db),
	.w4(32'h3c077490),
	.w5(32'h3c0cafcd),
	.w6(32'h3ba5cc85),
	.w7(32'h3bc89209),
	.w8(32'h3b9f565c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90003f4),
	.w1(32'hbb5968b1),
	.w2(32'hbb2ce060),
	.w3(32'hbaf10f61),
	.w4(32'hbb483737),
	.w5(32'hba4ca532),
	.w6(32'hbb1af671),
	.w7(32'hbb857d95),
	.w8(32'hbafb09e9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967aac4),
	.w1(32'hb95510c1),
	.w2(32'hb8f70861),
	.w3(32'hb99818a0),
	.w4(32'hb9a4e730),
	.w5(32'hb924971c),
	.w6(32'hb9904a28),
	.w7(32'hb999e255),
	.w8(32'hb956a263),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87b877),
	.w1(32'h394b3b99),
	.w2(32'hb97a3304),
	.w3(32'h395e074b),
	.w4(32'hb9a3faa1),
	.w5(32'hb9bdb6f7),
	.w6(32'h3ad4e238),
	.w7(32'h3a93751e),
	.w8(32'hb5dd3eba),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12fd53),
	.w1(32'hbb93bea8),
	.w2(32'hbb5dd9cb),
	.w3(32'hb9e8a786),
	.w4(32'hba590448),
	.w5(32'hba53c078),
	.w6(32'h38869ba8),
	.w7(32'h39ab8eff),
	.w8(32'h390c9ab6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6edb8e1),
	.w1(32'hba819bb1),
	.w2(32'hbae4cc2f),
	.w3(32'hba5267de),
	.w4(32'hba94efe9),
	.w5(32'hba573b34),
	.w6(32'hbacf4e63),
	.w7(32'hba9f1e93),
	.w8(32'hba54602b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b011952),
	.w1(32'h3a72b85f),
	.w2(32'h3b073932),
	.w3(32'hb858f7d7),
	.w4(32'h38d6afa6),
	.w5(32'h3a9eda1e),
	.w6(32'hba910dd2),
	.w7(32'h3a0144a7),
	.w8(32'h39bde26b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a830af1),
	.w1(32'hbaafefaa),
	.w2(32'hba9c1407),
	.w3(32'h39fbfbc2),
	.w4(32'hbaf01007),
	.w5(32'hbab1a4fe),
	.w6(32'hb930ca81),
	.w7(32'hbaa3f751),
	.w8(32'hb9922ad2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ded20c),
	.w1(32'hbaf619b2),
	.w2(32'hba27bc2f),
	.w3(32'h38feca10),
	.w4(32'hbb1f8a19),
	.w5(32'hba6064de),
	.w6(32'hba833495),
	.w7(32'hbb981b5a),
	.w8(32'hbb29f31a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397af71a),
	.w1(32'h39ca2eaa),
	.w2(32'h3a82ea30),
	.w3(32'h3ac9012a),
	.w4(32'h3aa734d5),
	.w5(32'h3ac387d2),
	.w6(32'h3b1ea0e7),
	.w7(32'h3af28608),
	.w8(32'h3b177219),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4111),
	.w1(32'hba89a6ff),
	.w2(32'hbb207999),
	.w3(32'h38f29ee5),
	.w4(32'hbaaf2ddc),
	.w5(32'hbac45a73),
	.w6(32'hba85352c),
	.w7(32'hbaff50af),
	.w8(32'hbac1bbfa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396126f4),
	.w1(32'hb639d50b),
	.w2(32'h389b3e56),
	.w3(32'h399d686a),
	.w4(32'hb7db02cf),
	.w5(32'h383f1a3a),
	.w6(32'h3901f580),
	.w7(32'h380bfc05),
	.w8(32'h381e6488),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce01e7),
	.w1(32'hb8a85df6),
	.w2(32'h38593eaa),
	.w3(32'h37e82b68),
	.w4(32'hb795a0a4),
	.w5(32'hb839a9f8),
	.w6(32'h3850ede9),
	.w7(32'hb5c1ed4a),
	.w8(32'hb7f97c15),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0c72f),
	.w1(32'hb68a9b90),
	.w2(32'hb7c2f633),
	.w3(32'h375c7bfb),
	.w4(32'h37b41f0f),
	.w5(32'h3777ff6b),
	.w6(32'h365b3e5c),
	.w7(32'hb72066a0),
	.w8(32'hb72b7c51),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b4581),
	.w1(32'h37f8529f),
	.w2(32'h38d34bed),
	.w3(32'h38d6b5d6),
	.w4(32'h38a9d5ea),
	.w5(32'h388f4676),
	.w6(32'h38c02376),
	.w7(32'h38cdf6ec),
	.w8(32'h392e0de1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be78b),
	.w1(32'hbb59ca0b),
	.w2(32'hbba4de13),
	.w3(32'hbb039c8b),
	.w4(32'hbb7efc09),
	.w5(32'hbb8f1b35),
	.w6(32'hbb576d3c),
	.w7(32'hbb901039),
	.w8(32'hbb99b199),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986d4cb),
	.w1(32'hb9658e30),
	.w2(32'h39b2a90b),
	.w3(32'hb942a213),
	.w4(32'hb9e13a66),
	.w5(32'h395ba56f),
	.w6(32'hb9738eb6),
	.w7(32'hb9fa5809),
	.w8(32'h39011599),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b8522),
	.w1(32'h3a805e33),
	.w2(32'h3b11b57a),
	.w3(32'h3a49486a),
	.w4(32'h3a206461),
	.w5(32'h3ab1b452),
	.w6(32'h3b12096c),
	.w7(32'h3aa5afcc),
	.w8(32'h3ad3c01d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a873261),
	.w1(32'hbb324af9),
	.w2(32'hbb6dab65),
	.w3(32'hbabaabea),
	.w4(32'hbb8f99fc),
	.w5(32'hbb65b04e),
	.w6(32'hbb8854cd),
	.w7(32'hbb6e0fbf),
	.w8(32'hbb4910bc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c46d3),
	.w1(32'hb96073e4),
	.w2(32'hb7afc6d6),
	.w3(32'hb94e2ad8),
	.w4(32'hb8db3ec6),
	.w5(32'h38c174c3),
	.w6(32'hb82b84e0),
	.w7(32'h38c66212),
	.w8(32'h389c6b33),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bde4da),
	.w1(32'hb90b2852),
	.w2(32'hb86f56d9),
	.w3(32'h379feefa),
	.w4(32'hb8a7c74c),
	.w5(32'h3839a91e),
	.w6(32'h38c93529),
	.w7(32'hb77a2867),
	.w8(32'h38d8dcdf),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c95b1f),
	.w1(32'hb4ac9a0c),
	.w2(32'hb84be7eb),
	.w3(32'hb581ffaf),
	.w4(32'hb721c202),
	.w5(32'hb7c358ae),
	.w6(32'h389fd684),
	.w7(32'h3741a1d3),
	.w8(32'hb7946699),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8646f3d),
	.w1(32'h3a95706b),
	.w2(32'h3ab77f2f),
	.w3(32'hb9a73f25),
	.w4(32'h3a97a919),
	.w5(32'h3acd4929),
	.w6(32'h3b92a99f),
	.w7(32'h3b533edc),
	.w8(32'h3b87bf9d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b613189),
	.w1(32'hbb02bc5d),
	.w2(32'hbacfd34f),
	.w3(32'h3b93f30f),
	.w4(32'hbb0b99af),
	.w5(32'h39856e20),
	.w6(32'h3a147047),
	.w7(32'hba491c5f),
	.w8(32'h3abc2445),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0f77),
	.w1(32'h3b2aa3f4),
	.w2(32'hbc0160da),
	.w3(32'hb91c1a0f),
	.w4(32'h3beda34c),
	.w5(32'hb90b0bfd),
	.w6(32'hbc1895e3),
	.w7(32'hbc53baf2),
	.w8(32'hbc183d88),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89c00),
	.w1(32'hbb2f7add),
	.w2(32'h3a224736),
	.w3(32'hbb96bcd7),
	.w4(32'hbb0d9cd9),
	.w5(32'h39065470),
	.w6(32'hbb707688),
	.w7(32'hbb0ec314),
	.w8(32'hba94a1f5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48db59),
	.w1(32'h3adbdfed),
	.w2(32'h3b1efb1a),
	.w3(32'hb980e5cf),
	.w4(32'hb99a8797),
	.w5(32'h3a617347),
	.w6(32'h39b2c798),
	.w7(32'h3a329ab9),
	.w8(32'h3ab76d73),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae78634),
	.w1(32'h3b852c07),
	.w2(32'h3bec8879),
	.w3(32'hba632254),
	.w4(32'h3b9f660c),
	.w5(32'h3ba017ee),
	.w6(32'h3b97f887),
	.w7(32'h3c0814b0),
	.w8(32'h3b634782),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050818),
	.w1(32'hbbead806),
	.w2(32'h3b5c2559),
	.w3(32'h3bdc5ba3),
	.w4(32'hbbb8c664),
	.w5(32'h3a5f18fd),
	.w6(32'hbaba50af),
	.w7(32'h3bb2833c),
	.w8(32'hb85c6fcc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77b2d9),
	.w1(32'hbbad94af),
	.w2(32'hbc04cf67),
	.w3(32'h3bb678f9),
	.w4(32'hbbfa798d),
	.w5(32'hbc014978),
	.w6(32'hbb3c71d2),
	.w7(32'hbbabc314),
	.w8(32'hbbbf5b65),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f192b),
	.w1(32'h39cdef20),
	.w2(32'h3bb192a7),
	.w3(32'hbabe9743),
	.w4(32'h3a3beebc),
	.w5(32'h3b8d2955),
	.w6(32'hba6fd3f3),
	.w7(32'h3a04039b),
	.w8(32'h3acb43e8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a1483),
	.w1(32'hbad17bc9),
	.w2(32'hbb99893a),
	.w3(32'hbb0aaf19),
	.w4(32'hbb25614e),
	.w5(32'hbb80ccbb),
	.w6(32'h3acbca9b),
	.w7(32'hbacaa55d),
	.w8(32'hba9c02f5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cd3f5),
	.w1(32'h3b3e7011),
	.w2(32'h3a876115),
	.w3(32'h3a7ee215),
	.w4(32'h3a81b87d),
	.w5(32'hb9f93a22),
	.w6(32'h3b2efff4),
	.w7(32'hb852907e),
	.w8(32'h3b230009),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb21f2),
	.w1(32'hba0c2eb9),
	.w2(32'h3b97fdee),
	.w3(32'h3a99f2ef),
	.w4(32'h3a0c49d1),
	.w5(32'h3b06c5e2),
	.w6(32'hbb917c49),
	.w7(32'hbab50622),
	.w8(32'h3b0fa9a2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b543d77),
	.w1(32'h3b262289),
	.w2(32'h3b61c27f),
	.w3(32'h3af09441),
	.w4(32'h3ad5abcd),
	.w5(32'h3b5e28df),
	.w6(32'h3b3ce3b6),
	.w7(32'h3b33214d),
	.w8(32'h3a112cb6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46bbcf),
	.w1(32'hba88efe9),
	.w2(32'h3b0b10de),
	.w3(32'h3bd30003),
	.w4(32'hbb73ea64),
	.w5(32'hbbb6b1f0),
	.w6(32'h3b9e7647),
	.w7(32'h3c3e0fac),
	.w8(32'h3c09722c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafce003),
	.w1(32'hbab0a061),
	.w2(32'hbabdc0d7),
	.w3(32'hbb0c28e3),
	.w4(32'hba8b02a8),
	.w5(32'hb998ff7d),
	.w6(32'hba127ee3),
	.w7(32'hbae3cc2b),
	.w8(32'h39fdfb42),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986a00),
	.w1(32'hbb83047f),
	.w2(32'hbc60cbf7),
	.w3(32'hb9908f8d),
	.w4(32'hbbae821f),
	.w5(32'hbc4ae0ef),
	.w6(32'hb993c92c),
	.w7(32'hbb9c560a),
	.w8(32'hba0ed22a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24eefd),
	.w1(32'hbb90a88d),
	.w2(32'h3bf99741),
	.w3(32'hbad59925),
	.w4(32'hbbd99643),
	.w5(32'hbacfac68),
	.w6(32'h3a5fa269),
	.w7(32'h3c3dac0f),
	.w8(32'h3b93cffa),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820934),
	.w1(32'hbb13bbf2),
	.w2(32'hbb938438),
	.w3(32'h3ba459e5),
	.w4(32'hbb42d87c),
	.w5(32'hbba3e56f),
	.w6(32'hbad45b63),
	.w7(32'hbb70b2e0),
	.w8(32'hbb6817c5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8add6),
	.w1(32'h3a84b8a7),
	.w2(32'h3b5fbe5c),
	.w3(32'hbb9c8432),
	.w4(32'h392600f2),
	.w5(32'h3b131107),
	.w6(32'hb9dad274),
	.w7(32'h3ab19d14),
	.w8(32'h3a49ec9d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814a8f),
	.w1(32'hba96ca6e),
	.w2(32'h3adb625f),
	.w3(32'h3a723e6b),
	.w4(32'h3a361b27),
	.w5(32'h3b87390d),
	.w6(32'hbb36bda9),
	.w7(32'hb6467f8d),
	.w8(32'h3a86a2fe),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7ec49),
	.w1(32'hbb877bd3),
	.w2(32'hbae85256),
	.w3(32'h3b75c9f3),
	.w4(32'hbb947029),
	.w5(32'hbb372087),
	.w6(32'hbb9dd343),
	.w7(32'hbb96d829),
	.w8(32'hbb977acd),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac928af),
	.w1(32'hba39b0b4),
	.w2(32'hbb86a125),
	.w3(32'hbad301dd),
	.w4(32'hba5c761c),
	.w5(32'hbb4eb5dd),
	.w6(32'h3a19e9bd),
	.w7(32'hba357fbd),
	.w8(32'hba71053f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87950c),
	.w1(32'h3bb8011f),
	.w2(32'h3b80cc73),
	.w3(32'hbabbdbb2),
	.w4(32'h3bbd1386),
	.w5(32'h3b89e24e),
	.w6(32'h3c1811d3),
	.w7(32'h3c0b4ebb),
	.w8(32'h3c374b68),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30393),
	.w1(32'h3ba54f67),
	.w2(32'hba153e49),
	.w3(32'h3c0e2e4d),
	.w4(32'h3bfa6b25),
	.w5(32'h3c3d0437),
	.w6(32'hbb83088f),
	.w7(32'hbc04b2d0),
	.w8(32'hbbde6fb4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a761b),
	.w1(32'hba397f50),
	.w2(32'hbb110ec8),
	.w3(32'h3b6d6be3),
	.w4(32'hba6b9355),
	.w5(32'hba2dd18b),
	.w6(32'hb9b0c02c),
	.w7(32'h3a0632e5),
	.w8(32'h3af17f2c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce6c4),
	.w1(32'h3b552834),
	.w2(32'h3b921e21),
	.w3(32'h3b573c06),
	.w4(32'h3b04804e),
	.w5(32'h3b39d447),
	.w6(32'h3bcebab1),
	.w7(32'h3b51026b),
	.w8(32'h3be1c8eb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0783a4),
	.w1(32'hbbb22830),
	.w2(32'hbbceb920),
	.w3(32'h39af48c3),
	.w4(32'hbc001278),
	.w5(32'hbc07e215),
	.w6(32'hbbde97bb),
	.w7(32'hbbf78b15),
	.w8(32'hbbdaef69),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6cc84),
	.w1(32'h3b6159b4),
	.w2(32'h3b471958),
	.w3(32'hbbc59809),
	.w4(32'h3b2e59d7),
	.w5(32'hb9cff887),
	.w6(32'hb9d8f110),
	.w7(32'h3b13825a),
	.w8(32'h3b84e00a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba324ecf),
	.w1(32'hb9fa180a),
	.w2(32'hbb22b0d6),
	.w3(32'hbb75493e),
	.w4(32'hbb2b41e4),
	.w5(32'hbb686e9f),
	.w6(32'hbacb89a0),
	.w7(32'hbb0dc124),
	.w8(32'hbac1d1ad),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab13e24),
	.w1(32'h3a2ce529),
	.w2(32'h3a50be47),
	.w3(32'h3aedecc1),
	.w4(32'hb8beb83c),
	.w5(32'hba0489d5),
	.w6(32'h3a39af04),
	.w7(32'hba624fd8),
	.w8(32'hba66b07b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1e59),
	.w1(32'h3b93a891),
	.w2(32'h3a0c92d2),
	.w3(32'hbb8db747),
	.w4(32'h3af00993),
	.w5(32'hbb05c00c),
	.w6(32'h3b6b0664),
	.w7(32'hba0a5364),
	.w8(32'hbae12dde),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f7e59),
	.w1(32'hbb99fe93),
	.w2(32'hbb89489a),
	.w3(32'hbacf31af),
	.w4(32'hbb830f3d),
	.w5(32'hbb6b20a8),
	.w6(32'hbb9ce029),
	.w7(32'hbba0077a),
	.w8(32'hbb69e811),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba843b0b),
	.w1(32'h3b846135),
	.w2(32'h3b75c4c3),
	.w3(32'h39af881e),
	.w4(32'h3b86d5b7),
	.w5(32'h3b842276),
	.w6(32'h3bb81485),
	.w7(32'h3b98b448),
	.w8(32'h3bc40245),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f5be),
	.w1(32'hbaf1bb76),
	.w2(32'hbb10f468),
	.w3(32'h3b8e1fd4),
	.w4(32'hbb117490),
	.w5(32'hbb00480e),
	.w6(32'hba94aca1),
	.w7(32'hbad8cbe6),
	.w8(32'hb9feb412),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f861ab),
	.w1(32'h3c084081),
	.w2(32'h3c0e0d14),
	.w3(32'h3965ebe4),
	.w4(32'h3bc966aa),
	.w5(32'h3baf45d3),
	.w6(32'h3b513413),
	.w7(32'h3bee62bb),
	.w8(32'h3c1aaf05),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67132e),
	.w1(32'h3b0f6070),
	.w2(32'h3a5777ea),
	.w3(32'h3b676aa0),
	.w4(32'h3a96dc59),
	.w5(32'hba54c393),
	.w6(32'h3b10d2ef),
	.w7(32'hbb188611),
	.w8(32'hbb587e24),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba123bc4),
	.w1(32'hbb8668aa),
	.w2(32'hbb0d26b9),
	.w3(32'hbb0eb3b1),
	.w4(32'hbb49dbad),
	.w5(32'hba8b00bf),
	.w6(32'hbbb1daa3),
	.w7(32'hbb885e1f),
	.w8(32'hbb598d26),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45578e),
	.w1(32'hbae11cb6),
	.w2(32'hbaedafe3),
	.w3(32'hba54ed22),
	.w4(32'hbb4c698f),
	.w5(32'hbb4c60b8),
	.w6(32'hba0de943),
	.w7(32'hba527727),
	.w8(32'hba3e7117),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb53f),
	.w1(32'hbbd381bf),
	.w2(32'hbb43cad0),
	.w3(32'hbbb623f0),
	.w4(32'hbbce9010),
	.w5(32'hbb8d357e),
	.w6(32'hbc00b63b),
	.w7(32'hbb42a7b0),
	.w8(32'hbb877fda),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb956553),
	.w1(32'hbb0e8db4),
	.w2(32'h393b7018),
	.w3(32'hbb984ffc),
	.w4(32'hbac1337b),
	.w5(32'h3a039319),
	.w6(32'hbb3d5f57),
	.w7(32'hbac076df),
	.w8(32'hba841413),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40e20),
	.w1(32'h38d8bd05),
	.w2(32'hbafd7bb4),
	.w3(32'h3a437a53),
	.w4(32'hba8296bc),
	.w5(32'hbb116dcb),
	.w6(32'h3ac5c0a3),
	.w7(32'hb97dae0a),
	.w8(32'h39d60a52),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912b91a),
	.w1(32'hbbd444a5),
	.w2(32'hbb2614eb),
	.w3(32'hba4772d6),
	.w4(32'hbbe18b18),
	.w5(32'hbb7c0e0d),
	.w6(32'hbbd1bd5b),
	.w7(32'hbbd470c4),
	.w8(32'hbbbb786b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342ae2),
	.w1(32'hbb168e46),
	.w2(32'h3a8e5982),
	.w3(32'hba0dc495),
	.w4(32'h3a9fc058),
	.w5(32'h3b27dc18),
	.w6(32'h3b29cfd2),
	.w7(32'hb93ae7f6),
	.w8(32'h3afbd097),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79fb75),
	.w1(32'hbb3140c3),
	.w2(32'hb9d3f9a4),
	.w3(32'hba90afc7),
	.w4(32'hbb9aee76),
	.w5(32'hbb7bd737),
	.w6(32'hbbd1c639),
	.w7(32'hbb50c1f1),
	.w8(32'hbb6e2337),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35b688),
	.w1(32'hbb9cd44b),
	.w2(32'hbbdde07f),
	.w3(32'hbbafaab9),
	.w4(32'hbbbba2d7),
	.w5(32'hbbd8abcc),
	.w6(32'hbb583349),
	.w7(32'hbbb675ad),
	.w8(32'hbb731638),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cfd77),
	.w1(32'hbba0997a),
	.w2(32'hba847010),
	.w3(32'hbb38e5cf),
	.w4(32'hbafa8c7b),
	.w5(32'h3a1e21e0),
	.w6(32'hbbdbe676),
	.w7(32'hbb95f954),
	.w8(32'hbacfddae),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023e33),
	.w1(32'h3b67b629),
	.w2(32'hb9c17c42),
	.w3(32'h3b5aad1f),
	.w4(32'h3c0db68e),
	.w5(32'h3bf833ea),
	.w6(32'hba8b2212),
	.w7(32'hbb2d082d),
	.w8(32'h3ad063b1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc253c2),
	.w1(32'h3b219aa0),
	.w2(32'h3bb813ab),
	.w3(32'h3bfa1d23),
	.w4(32'h3b83db25),
	.w5(32'h3c004766),
	.w6(32'h3a8475ea),
	.w7(32'h3a951197),
	.w8(32'h3af727c6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e597),
	.w1(32'h3add91bc),
	.w2(32'h3c17730f),
	.w3(32'h3c195400),
	.w4(32'h3b890f56),
	.w5(32'h3ba4bbc4),
	.w6(32'h3bf6d7df),
	.w7(32'h3c721699),
	.w8(32'h3c220f1e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1f980),
	.w1(32'h3b0b734b),
	.w2(32'hb922b91d),
	.w3(32'h3b99a77f),
	.w4(32'h3a865b7d),
	.w5(32'hbae39c30),
	.w6(32'h3abe9498),
	.w7(32'hbadf78bf),
	.w8(32'hbad03412),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379bb567),
	.w1(32'h3a852fa4),
	.w2(32'h3a60f2a6),
	.w3(32'hb8c760c3),
	.w4(32'hb6129d9a),
	.w5(32'hb96f8637),
	.w6(32'hb8cd244e),
	.w7(32'hbafbec97),
	.w8(32'hba02a7c6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73a963),
	.w1(32'h39a7bb52),
	.w2(32'hbb4017dd),
	.w3(32'hba96949e),
	.w4(32'h389e166e),
	.w5(32'hbb183584),
	.w6(32'h3b2f2c39),
	.w7(32'h39edc607),
	.w8(32'h3ab9ebeb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc776f),
	.w1(32'h3b0b0281),
	.w2(32'h3ba97c0f),
	.w3(32'h3a0a52f9),
	.w4(32'h3bac84ee),
	.w5(32'h3bb93be7),
	.w6(32'h3b85d2c9),
	.w7(32'h3c05c4df),
	.w8(32'h3c1da4b0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e7f43),
	.w1(32'h3b918d83),
	.w2(32'hbb6b9add),
	.w3(32'h3c1adbd4),
	.w4(32'h3b84ac64),
	.w5(32'hbbea6cf4),
	.w6(32'hbaa0e152),
	.w7(32'hb9b80e35),
	.w8(32'h3b170a62),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4f013),
	.w1(32'hbc2c8144),
	.w2(32'hbc39b290),
	.w3(32'hbbddba3e),
	.w4(32'hbc2bd36c),
	.w5(32'hbc43c8c1),
	.w6(32'hbc05d247),
	.w7(32'hbc1c8cfc),
	.w8(32'hbc175481),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f5bd),
	.w1(32'hbc171dcd),
	.w2(32'hbbd86c89),
	.w3(32'hbc45dbf2),
	.w4(32'hbc1b385b),
	.w5(32'hbbf5e760),
	.w6(32'hbc10c442),
	.w7(32'hbbea24fa),
	.w8(32'hbc3eb761),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14cc33),
	.w1(32'hbaec5d38),
	.w2(32'hb9b20d09),
	.w3(32'hbc05e086),
	.w4(32'hbb142bfd),
	.w5(32'hbaf2a9ab),
	.w6(32'hbaee39ae),
	.w7(32'hbaf97245),
	.w8(32'hbb0e7a18),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac037),
	.w1(32'h395f525d),
	.w2(32'hba90c5d5),
	.w3(32'hbb77dd37),
	.w4(32'hbae08801),
	.w5(32'hb9a488a7),
	.w6(32'h3a59a662),
	.w7(32'h370b27d4),
	.w8(32'hbaa6bdea),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cf8a0),
	.w1(32'h3b5aa137),
	.w2(32'h3b65ee1a),
	.w3(32'hba3af2fc),
	.w4(32'h3a9c60a7),
	.w5(32'h3a6c8e73),
	.w6(32'h3b937d7d),
	.w7(32'h3ba63123),
	.w8(32'h3bd1e27c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b497),
	.w1(32'hbc1a654d),
	.w2(32'h3b819cf1),
	.w3(32'h3b93a713),
	.w4(32'hbc0cb3d3),
	.w5(32'hb72b7468),
	.w6(32'h3a481925),
	.w7(32'h3c087d79),
	.w8(32'h3b875215),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1255a3),
	.w1(32'hba4245d3),
	.w2(32'hba0e51e2),
	.w3(32'h3c1525b8),
	.w4(32'hba41fe57),
	.w5(32'h3a357606),
	.w6(32'hbb3f5b35),
	.w7(32'hbb5716e4),
	.w8(32'hbafee987),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a66f),
	.w1(32'h3ba832c4),
	.w2(32'h3b628871),
	.w3(32'h39ea2f6a),
	.w4(32'h3b9ede90),
	.w5(32'h3b1c3fa5),
	.w6(32'h3bbf33f7),
	.w7(32'h3bcb0126),
	.w8(32'h3bee8d90),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf5fd),
	.w1(32'hbc04330e),
	.w2(32'hbc0556f7),
	.w3(32'hba68c3dc),
	.w4(32'hbc29e0d8),
	.w5(32'hbc0242c5),
	.w6(32'hbc3f53bb),
	.w7(32'hbc446321),
	.w8(32'hbc1c313a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ca16),
	.w1(32'h3af4e5c1),
	.w2(32'hbb1bd72e),
	.w3(32'hbbdc7e66),
	.w4(32'h3b4c3e0a),
	.w5(32'h3a6f50eb),
	.w6(32'hb93629ac),
	.w7(32'hbb90caf1),
	.w8(32'hbaa664c3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba822b02),
	.w1(32'h3bc8fa35),
	.w2(32'h3bcfcbeb),
	.w3(32'h3966b90c),
	.w4(32'h3bb61cfa),
	.w5(32'h3c054de6),
	.w6(32'hbb084593),
	.w7(32'h3a4af750),
	.w8(32'h3bf543ae),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a49ef),
	.w1(32'hbb1ed56e),
	.w2(32'h3a67c299),
	.w3(32'h3c0edd41),
	.w4(32'hba43eabe),
	.w5(32'h3a8f738c),
	.w6(32'hbb8e4664),
	.w7(32'hbb03d760),
	.w8(32'hb9115816),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf77b2),
	.w1(32'hbad7eb1e),
	.w2(32'h3a3bdf07),
	.w3(32'h39dd9ea1),
	.w4(32'hbb2c594a),
	.w5(32'h396fb0b8),
	.w6(32'hbb20a0ac),
	.w7(32'hbab2308c),
	.w8(32'hb9a1c901),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f9a32),
	.w1(32'hbc30307a),
	.w2(32'hbb08edfd),
	.w3(32'h39596e3c),
	.w4(32'hbbe0bf41),
	.w5(32'hba84a7c8),
	.w6(32'hbbd3ab1b),
	.w7(32'hba32510d),
	.w8(32'hbaa5f82c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea553),
	.w1(32'h3b0c6c62),
	.w2(32'h3b53e704),
	.w3(32'h3a90ecc6),
	.w4(32'h3a141d21),
	.w5(32'h3a3b7314),
	.w6(32'h399f2cd9),
	.w7(32'h3a7542cf),
	.w8(32'h3abfbf3d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b267cf9),
	.w1(32'hbb029ca2),
	.w2(32'hbba5db96),
	.w3(32'h3aa7b9b1),
	.w4(32'hbb034ea5),
	.w5(32'hbba36b15),
	.w6(32'hbad71fee),
	.w7(32'hbb9cd7cf),
	.w8(32'hbbce9de0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0958db),
	.w1(32'hbb2409f5),
	.w2(32'hbb90d417),
	.w3(32'hba1023bd),
	.w4(32'hbb5451e5),
	.w5(32'hbbb2f1c7),
	.w6(32'hb849a91e),
	.w7(32'hbb25c0c9),
	.w8(32'hbae9d8e9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4fe3),
	.w1(32'hbc0dcdb8),
	.w2(32'hb9363ac6),
	.w3(32'hbb0ffce3),
	.w4(32'hbb85c6a4),
	.w5(32'h3a5cc5b4),
	.w6(32'hb9dd481b),
	.w7(32'h3b8b8a17),
	.w8(32'h3bb864d5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a1d7),
	.w1(32'hbb16c0ed),
	.w2(32'hb9a8efa0),
	.w3(32'h3c136a77),
	.w4(32'hbafac04c),
	.w5(32'h36f70bbd),
	.w6(32'hbb9f60ae),
	.w7(32'hbb79270b),
	.w8(32'hbb3c97f8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72f7b1),
	.w1(32'hba49a75c),
	.w2(32'hba4816db),
	.w3(32'h3a556c5d),
	.w4(32'hba83d817),
	.w5(32'hb9c6568e),
	.w6(32'h3b199128),
	.w7(32'h3aa2875f),
	.w8(32'h3b10a6f7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf6c53),
	.w1(32'h3a637072),
	.w2(32'hba1ba4fe),
	.w3(32'h3b33ccb0),
	.w4(32'h3a70d3bf),
	.w5(32'hbab95d0d),
	.w6(32'h3b58147c),
	.w7(32'h392d16b1),
	.w8(32'h3a4cac8e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3ea1b),
	.w1(32'hbab6274c),
	.w2(32'hbb25c6f9),
	.w3(32'hbad77324),
	.w4(32'hbb411a78),
	.w5(32'hbb61f116),
	.w6(32'h393feb4e),
	.w7(32'hb9fa867c),
	.w8(32'h3a0e9d5f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8d016),
	.w1(32'hbbd58b88),
	.w2(32'hbbc9042b),
	.w3(32'hbab28e60),
	.w4(32'hbbde66a8),
	.w5(32'hbbe33f78),
	.w6(32'hbbda3a36),
	.w7(32'hbbf44003),
	.w8(32'hbbf72e9a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7f502),
	.w1(32'h3c2d389b),
	.w2(32'h3bf3a35c),
	.w3(32'hbc05af14),
	.w4(32'h3a88a8be),
	.w5(32'hbc23d3ea),
	.w6(32'h3c072415),
	.w7(32'h3c8e4436),
	.w8(32'h3c577a25),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1495b9),
	.w1(32'hb8b869f0),
	.w2(32'hbb957196),
	.w3(32'hbc0eefe9),
	.w4(32'hba81600b),
	.w5(32'hbb529b78),
	.w6(32'h3b26a8b6),
	.w7(32'hba8bfcfa),
	.w8(32'h3aaeb798),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3522a1),
	.w1(32'hb767a449),
	.w2(32'h393a25cf),
	.w3(32'h3afc1daa),
	.w4(32'hb9937b32),
	.w5(32'h39936f81),
	.w6(32'hbb6ca940),
	.w7(32'hbae5926b),
	.w8(32'h38a46c45),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd0e17),
	.w1(32'hb9c91ae0),
	.w2(32'hba5c0bd3),
	.w3(32'hbb3fe2dc),
	.w4(32'hbb1b03df),
	.w5(32'hbb678d01),
	.w6(32'hbb1fc209),
	.w7(32'hbb0b2a36),
	.w8(32'hbb895c46),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b935),
	.w1(32'h3b8b244d),
	.w2(32'h3b81dbb1),
	.w3(32'h3a2a3f88),
	.w4(32'h3bbf95e5),
	.w5(32'h3ba73546),
	.w6(32'h3c110210),
	.w7(32'h3c01db78),
	.w8(32'h3c11652c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba096f),
	.w1(32'hba84e5b8),
	.w2(32'hbb423499),
	.w3(32'h3be185a5),
	.w4(32'hbab8a28c),
	.w5(32'hbb394d9c),
	.w6(32'h3aa37e95),
	.w7(32'hba8b8a28),
	.w8(32'hbabfd2e4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a222717),
	.w1(32'hbaacc9bf),
	.w2(32'h3ac1e183),
	.w3(32'h3a1e85df),
	.w4(32'hbafbaff6),
	.w5(32'h3a84aa7c),
	.w6(32'hbb0c5210),
	.w7(32'h38e9c49f),
	.w8(32'h3ac8c8c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27cb6f),
	.w1(32'hbae97901),
	.w2(32'hbb1656b6),
	.w3(32'h3ab27b3e),
	.w4(32'hbab9f9c0),
	.w5(32'hbb2b22e6),
	.w6(32'hbb00e626),
	.w7(32'hbb124086),
	.w8(32'hba8b700d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af9fe),
	.w1(32'hbbe00c71),
	.w2(32'hbbabe1af),
	.w3(32'hbb84acb1),
	.w4(32'hbbfcfc67),
	.w5(32'hbb57a72d),
	.w6(32'hbc1a7915),
	.w7(32'hbc1cf0af),
	.w8(32'hbc0d7234),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e45e1),
	.w1(32'h3b5ce087),
	.w2(32'h3b478b05),
	.w3(32'hbb0cc854),
	.w4(32'h3affd9af),
	.w5(32'hb982e095),
	.w6(32'h3c03ed04),
	.w7(32'h3b173e17),
	.w8(32'h3b5cbdc6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1df560),
	.w1(32'h3aeb94c8),
	.w2(32'h39bb6ad0),
	.w3(32'hba47ae16),
	.w4(32'h3a017991),
	.w5(32'h3a65619c),
	.w6(32'h3b26b189),
	.w7(32'h3abdb109),
	.w8(32'h3af92016),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ae77),
	.w1(32'h3ba650ee),
	.w2(32'hb90a9b8f),
	.w3(32'h3b0c13ca),
	.w4(32'h3b9944e8),
	.w5(32'hbb141fea),
	.w6(32'h3b8f29e1),
	.w7(32'h3b9b1cde),
	.w8(32'h3bcb565a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32ee64),
	.w1(32'h3b0aecf0),
	.w2(32'h3a80d112),
	.w3(32'hbb787996),
	.w4(32'h3b1058d5),
	.w5(32'h3abc70a1),
	.w6(32'h3b76062d),
	.w7(32'h3b41f76f),
	.w8(32'h3b91c2aa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d19aa),
	.w1(32'hbb6270c3),
	.w2(32'hbb3105fc),
	.w3(32'h3b75477e),
	.w4(32'hbb7a2954),
	.w5(32'hbb77ab8b),
	.w6(32'hbb37e221),
	.w7(32'hbb608dec),
	.w8(32'hbb8d17e2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92047c),
	.w1(32'hbb0f281c),
	.w2(32'h3ac2306a),
	.w3(32'hbbcbbd03),
	.w4(32'hb827a718),
	.w5(32'h3b15f2a0),
	.w6(32'h3b6dbcea),
	.w7(32'h3af415ce),
	.w8(32'h3bf0fa74),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba324a2),
	.w1(32'h3b831173),
	.w2(32'h3b4edc18),
	.w3(32'h3c071c9e),
	.w4(32'h3b5f18dd),
	.w5(32'h3b079c93),
	.w6(32'h3bd6e448),
	.w7(32'h3b9fa642),
	.w8(32'h3bbfbb53),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914e71a),
	.w1(32'hbab35d22),
	.w2(32'h3bd910c0),
	.w3(32'h3b0de057),
	.w4(32'h3ade7519),
	.w5(32'h3bbbd1e0),
	.w6(32'hb9970200),
	.w7(32'h3afc6da1),
	.w8(32'h3bacfd2b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9603d3),
	.w1(32'hbbf50a4d),
	.w2(32'hbbe77ee2),
	.w3(32'h3b2ed65a),
	.w4(32'hbc1d23f9),
	.w5(32'hbc02752b),
	.w6(32'hbc0e268e),
	.w7(32'hbc2cca92),
	.w8(32'hbc1d8e8a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa80d),
	.w1(32'h3a3d67f8),
	.w2(32'hba989a2f),
	.w3(32'hbbe23005),
	.w4(32'hbabacc39),
	.w5(32'hbae6a19d),
	.w6(32'h3aa08ae5),
	.w7(32'hba5934d7),
	.w8(32'hbb016007),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fcbdb),
	.w1(32'hbb45f8e9),
	.w2(32'hbb0e59c6),
	.w3(32'h3a180a92),
	.w4(32'hbb5d9257),
	.w5(32'hbb260867),
	.w6(32'hbb5cc842),
	.w7(32'hbb489a6d),
	.w8(32'hbb2bae9f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2d80),
	.w1(32'hbbf5140b),
	.w2(32'hbbe9ebe6),
	.w3(32'hbb455762),
	.w4(32'hbc0dfce3),
	.w5(32'hbbcf67f6),
	.w6(32'hbc0adc28),
	.w7(32'hbc21f3fc),
	.w8(32'hbc217780),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb6303),
	.w1(32'hba3caf25),
	.w2(32'hba646eae),
	.w3(32'hbc010c6f),
	.w4(32'h3902f43c),
	.w5(32'h397b5511),
	.w6(32'h3889b8f2),
	.w7(32'hba517be6),
	.w8(32'h3b172e45),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5b62d),
	.w1(32'h3bb9e87b),
	.w2(32'h3ad2754e),
	.w3(32'h3b55ed0c),
	.w4(32'h3bcec24d),
	.w5(32'h3a902892),
	.w6(32'h3b015890),
	.w7(32'h3a94be71),
	.w8(32'h3b15d0e4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c380),
	.w1(32'hbbffca11),
	.w2(32'hbb973608),
	.w3(32'h3b1d9727),
	.w4(32'hbc0834fd),
	.w5(32'hbb9e3e9c),
	.w6(32'hbc0d8cfa),
	.w7(32'hbbeff69a),
	.w8(32'hbbde12e0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb699ad8),
	.w1(32'hbc02d0b3),
	.w2(32'hbbfebc44),
	.w3(32'hbb997496),
	.w4(32'hbbfcd732),
	.w5(32'hbbecb842),
	.w6(32'hbbf3db3b),
	.w7(32'hbc169a97),
	.w8(32'hbbe979b4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb92f),
	.w1(32'hbb12bd11),
	.w2(32'h3c0f9d94),
	.w3(32'hbc1f764a),
	.w4(32'hbb917d50),
	.w5(32'h3b737522),
	.w6(32'h3b87fd0c),
	.w7(32'h3c1c32a2),
	.w8(32'h3a089767),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01232),
	.w1(32'hbbcb658c),
	.w2(32'h3bfbd911),
	.w3(32'h3b9ce9d9),
	.w4(32'hbbe0d7a8),
	.w5(32'h3be28c7f),
	.w6(32'hbc2b63b9),
	.w7(32'h3a793585),
	.w8(32'hba10e467),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3928ea),
	.w1(32'h3b8ed56a),
	.w2(32'h3b41c547),
	.w3(32'h3c3aa097),
	.w4(32'h3bb9d5fb),
	.w5(32'h3b3fa45a),
	.w6(32'h3c46abed),
	.w7(32'h3bac84ae),
	.w8(32'h3c367716),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1f04a),
	.w1(32'hb8857215),
	.w2(32'h39278e09),
	.w3(32'h3b989a91),
	.w4(32'hb8b6c655),
	.w5(32'hb8d1e91c),
	.w6(32'h3b85f1c8),
	.w7(32'h3b7baf95),
	.w8(32'h3b87bc48),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1fa7),
	.w1(32'h3abb2957),
	.w2(32'hbaa919bd),
	.w3(32'h3a8e4101),
	.w4(32'h3a9d236d),
	.w5(32'hba37cccd),
	.w6(32'h3b84f1aa),
	.w7(32'h3ae3d182),
	.w8(32'h3b499ea0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507dc9),
	.w1(32'h3bbf8bb0),
	.w2(32'h3b64cb07),
	.w3(32'h3b41bd08),
	.w4(32'h3b95649b),
	.w5(32'h3aeeda1a),
	.w6(32'h3bba1824),
	.w7(32'h3b97ee81),
	.w8(32'h3bb12a7c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39046f44),
	.w1(32'hba88f645),
	.w2(32'h396a2115),
	.w3(32'hb9dec611),
	.w4(32'hbb1a3749),
	.w5(32'h3a2ce677),
	.w6(32'hbb072aef),
	.w7(32'hbae159ec),
	.w8(32'hba897725),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956df2c),
	.w1(32'h3b924f2b),
	.w2(32'h3b2d1e8a),
	.w3(32'hb9c35085),
	.w4(32'h3b9437ce),
	.w5(32'h3b60f5fa),
	.w6(32'h3bdabb52),
	.w7(32'h3bbb9415),
	.w8(32'h3c079378),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb02c49),
	.w1(32'h3a7af000),
	.w2(32'hbaf10fa1),
	.w3(32'h3bb756da),
	.w4(32'h3a59b268),
	.w5(32'hba90289b),
	.w6(32'h3b7e0741),
	.w7(32'h3ac6b1c3),
	.w8(32'h3b41afb8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2088e4),
	.w1(32'h3bb5fbb9),
	.w2(32'h3bb3ae88),
	.w3(32'h3ad37e51),
	.w4(32'h3c003859),
	.w5(32'h3bff5b07),
	.w6(32'h3b1cb033),
	.w7(32'h3ba60be2),
	.w8(32'h3c2c5a9a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27708a),
	.w1(32'hba1d57da),
	.w2(32'hbbbb4377),
	.w3(32'h3c2dc413),
	.w4(32'hbb2155c1),
	.w5(32'hbbfd3f08),
	.w6(32'h3a1be60c),
	.w7(32'hbb283553),
	.w8(32'hbb3c6ee7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98a99),
	.w1(32'h3c2c5a83),
	.w2(32'hbb6ba5d2),
	.w3(32'hbb9a1376),
	.w4(32'h3c40b760),
	.w5(32'h39c4fd61),
	.w6(32'hba6e2a98),
	.w7(32'hbbc2a5a7),
	.w8(32'hbb860bae),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03312b),
	.w1(32'hbb3dc3de),
	.w2(32'hbba1f2b7),
	.w3(32'hbbf00399),
	.w4(32'hbb466e14),
	.w5(32'hbbbb95eb),
	.w6(32'hbafde20b),
	.w7(32'hbb6aa487),
	.w8(32'hbb6234f5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0227),
	.w1(32'h3b53d3fe),
	.w2(32'h3b7e20d7),
	.w3(32'hbbbeafad),
	.w4(32'h3b45dbb2),
	.w5(32'h3b20ad94),
	.w6(32'h3b807f19),
	.w7(32'h3ba50b01),
	.w8(32'h3b94cd7b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dab64),
	.w1(32'h3bec2f1b),
	.w2(32'h3ad5d85a),
	.w3(32'h3b1a18b2),
	.w4(32'h3bf48d3a),
	.w5(32'h3b4dfe5d),
	.w6(32'h3bfd5013),
	.w7(32'h3b8fe11b),
	.w8(32'h3bd153ad),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8117f8),
	.w1(32'h3afbf646),
	.w2(32'hbb0bb06c),
	.w3(32'h3a87a919),
	.w4(32'h3ae2f20e),
	.w5(32'hba926fb1),
	.w6(32'h3bc43c6d),
	.w7(32'h3b2c291e),
	.w8(32'h3b96d6b5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0f56c),
	.w1(32'h3a4d11c4),
	.w2(32'hba8d9b11),
	.w3(32'h3b31d9b8),
	.w4(32'hb8a62035),
	.w5(32'hba514ee5),
	.w6(32'h3b49c04b),
	.w7(32'h3a8d5a86),
	.w8(32'h3ac9b50b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba5802),
	.w1(32'h3a50f908),
	.w2(32'hbabd276e),
	.w3(32'h3a2bbc88),
	.w4(32'hb996c2a6),
	.w5(32'hba9b5237),
	.w6(32'h3b3cff9f),
	.w7(32'h3a4a7932),
	.w8(32'h3ab86e25),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7c67f),
	.w1(32'h3bb9e50a),
	.w2(32'h3b374629),
	.w3(32'h3b2076d2),
	.w4(32'h3c006e25),
	.w5(32'h3c26a716),
	.w6(32'hbb87b5c9),
	.w7(32'hbbd6c311),
	.w8(32'hbbae0334),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446123),
	.w1(32'hb931f89b),
	.w2(32'h3aec5df9),
	.w3(32'h3b81ca9a),
	.w4(32'h3a699ceb),
	.w5(32'h3b0bd2aa),
	.w6(32'hb96809cf),
	.w7(32'h3b570653),
	.w8(32'h3abc0ddd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3fd7f),
	.w1(32'hbbe66d62),
	.w2(32'hbbbb8c70),
	.w3(32'h394dcf7e),
	.w4(32'hbbfeee94),
	.w5(32'hbbd608b0),
	.w6(32'hbba84597),
	.w7(32'hbb8f77f7),
	.w8(32'hbbb9196f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd6290),
	.w1(32'hbb68528e),
	.w2(32'hbbc10961),
	.w3(32'hbbce6034),
	.w4(32'hbb88dcc5),
	.w5(32'hbbbe66c4),
	.w6(32'hbb5802c5),
	.w7(32'hbbb84e13),
	.w8(32'hbbaac33b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80249),
	.w1(32'h3b025791),
	.w2(32'hba3fa212),
	.w3(32'hbbc54fc1),
	.w4(32'h3ac21e18),
	.w5(32'hb9e7b271),
	.w6(32'h3b4d445d),
	.w7(32'h3ac10fe5),
	.w8(32'h3b0ead94),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df139c),
	.w1(32'h3ab78f05),
	.w2(32'h3b2c93f2),
	.w3(32'h38f89c18),
	.w4(32'h3ae4fb00),
	.w5(32'h3c09a3e5),
	.w6(32'hbc004ff1),
	.w7(32'hbbef1b0e),
	.w8(32'hbc049aff),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800ea1),
	.w1(32'hbc6d9e82),
	.w2(32'hbc62b19a),
	.w3(32'h3b8b21f6),
	.w4(32'hbc6996c0),
	.w5(32'hbc5faa2b),
	.w6(32'hbc4aa77a),
	.w7(32'hbc6affb0),
	.w8(32'hbc588b34),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc559fe9),
	.w1(32'h3ad9086b),
	.w2(32'h3a73df24),
	.w3(32'hbc4ad194),
	.w4(32'h3b056697),
	.w5(32'h3a5dd2e2),
	.w6(32'h3bd681b9),
	.w7(32'h3b692082),
	.w8(32'h3b88a723),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84658d),
	.w1(32'h37ad7cd0),
	.w2(32'h37ca1173),
	.w3(32'hba1c4210),
	.w4(32'h386f8e74),
	.w5(32'h38d0d357),
	.w6(32'hb6d223ea),
	.w7(32'h390f012c),
	.w8(32'h394fd559),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae0902),
	.w1(32'h3a9e946e),
	.w2(32'hba1e1b04),
	.w3(32'h3a81efac),
	.w4(32'hbb06b417),
	.w5(32'hbacbadab),
	.w6(32'h3b4d98b6),
	.w7(32'hbaaea092),
	.w8(32'hbab7f1a1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule