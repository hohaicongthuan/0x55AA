module layer_10_featuremap_204(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5475b1),
	.w1(32'hb91ae0b2),
	.w2(32'hbb2b2891),
	.w3(32'h3a36d590),
	.w4(32'hba3592a9),
	.w5(32'hba78d136),
	.w6(32'h3a7a992b),
	.w7(32'h38508249),
	.w8(32'h3a2a0a08),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab08623),
	.w1(32'hb98f2f0a),
	.w2(32'hbac3256f),
	.w3(32'h39a6c515),
	.w4(32'h3a8e08d6),
	.w5(32'hb9fe0608),
	.w6(32'h3acc3ec2),
	.w7(32'h3a7b3e5c),
	.w8(32'hb7824b78),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71db13),
	.w1(32'h3a3c01d9),
	.w2(32'h3a12e385),
	.w3(32'h3a85f89b),
	.w4(32'h3a1f489c),
	.w5(32'h39140166),
	.w6(32'h3a193956),
	.w7(32'h37d87d21),
	.w8(32'h3982d066),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394306e1),
	.w1(32'hb996a0d6),
	.w2(32'hba575e71),
	.w3(32'h39950bf3),
	.w4(32'hb80e5a46),
	.w5(32'hba0820f0),
	.w6(32'hba312f03),
	.w7(32'hbad9e7ed),
	.w8(32'hba617c41),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba252207),
	.w1(32'hb93b8e19),
	.w2(32'hba8d29a9),
	.w3(32'h39e40b15),
	.w4(32'hb9099975),
	.w5(32'hb9a193c9),
	.w6(32'h3abd833e),
	.w7(32'h3a523288),
	.w8(32'hb9f631ec),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02b856),
	.w1(32'h39cdf1c1),
	.w2(32'hba55091b),
	.w3(32'hb983e0e8),
	.w4(32'h3a6ae594),
	.w5(32'h378c198b),
	.w6(32'h3a37e8ff),
	.w7(32'h3892ba31),
	.w8(32'h39010110),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef42e),
	.w1(32'h3ba1b025),
	.w2(32'h3baef066),
	.w3(32'h3b94ba60),
	.w4(32'h3a4cc433),
	.w5(32'h39188520),
	.w6(32'h3b937f14),
	.w7(32'h3b694edf),
	.w8(32'h39ad84eb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3a70d),
	.w1(32'hbb7f0137),
	.w2(32'hb99eb1ab),
	.w3(32'hbb0c1d65),
	.w4(32'hbc021c6e),
	.w5(32'hbb3a9a50),
	.w6(32'hbacc53a1),
	.w7(32'h3b26ba45),
	.w8(32'hba9c0915),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a851792),
	.w1(32'h39aadef4),
	.w2(32'h3a2dc8ef),
	.w3(32'h3a9c569f),
	.w4(32'h3a09576f),
	.w5(32'h39cfc9c3),
	.w6(32'h3a240c30),
	.w7(32'h3a4d0c7c),
	.w8(32'h3a4a1280),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f13a8),
	.w1(32'h3b1d2ca2),
	.w2(32'hba298078),
	.w3(32'h3af64215),
	.w4(32'h398aaf36),
	.w5(32'hba8161e3),
	.w6(32'h3a49b82c),
	.w7(32'h388d3cf2),
	.w8(32'hba80b3ba),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19a4d8),
	.w1(32'hbb10db4c),
	.w2(32'hbae78a8d),
	.w3(32'hb9bf0bb5),
	.w4(32'hb9ba5f33),
	.w5(32'hba8ebc54),
	.w6(32'hbaa031f9),
	.w7(32'hbb3b5279),
	.w8(32'hbb65a200),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8604c),
	.w1(32'h3bff704f),
	.w2(32'h3bc15dd8),
	.w3(32'h3b857a11),
	.w4(32'h3b1c72a5),
	.w5(32'h3ad3e112),
	.w6(32'hba659fb2),
	.w7(32'hba003b12),
	.w8(32'hba26ff20),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447e45),
	.w1(32'h3b209b3f),
	.w2(32'h3889c21e),
	.w3(32'h3a49ec5f),
	.w4(32'hba1eda8c),
	.w5(32'hba43278c),
	.w6(32'h3a9d9943),
	.w7(32'hb7eafcbb),
	.w8(32'hb9df2464),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4bbf4),
	.w1(32'hba6dce6e),
	.w2(32'hbb3cc05b),
	.w3(32'h3ab675ab),
	.w4(32'hb943f302),
	.w5(32'hbb07cf93),
	.w6(32'h3b152110),
	.w7(32'h39908cda),
	.w8(32'hba87b62f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb2f87),
	.w1(32'hbaf251fc),
	.w2(32'hbb8c0d46),
	.w3(32'h3b14821e),
	.w4(32'hbad10e1c),
	.w5(32'hba6cea03),
	.w6(32'h3a4332b6),
	.w7(32'hb9cfdd02),
	.w8(32'hba28aae0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb42e3),
	.w1(32'h3a8d057c),
	.w2(32'hbb8225a8),
	.w3(32'hba7605c2),
	.w4(32'hbac5887f),
	.w5(32'hbb0c90c1),
	.w6(32'hb9e1c7ba),
	.w7(32'hb9ae7876),
	.w8(32'hba9e202d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a268b),
	.w1(32'h39dba966),
	.w2(32'h39c23a50),
	.w3(32'h3a30c3ac),
	.w4(32'h38efc3ec),
	.w5(32'hb9ba7c4b),
	.w6(32'h3a631c99),
	.w7(32'h3a55c7c1),
	.w8(32'hb6d629c2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9abce9),
	.w1(32'h3b3cfd96),
	.w2(32'h394df3a3),
	.w3(32'hb999fba7),
	.w4(32'hbb5ed88c),
	.w5(32'hbb050348),
	.w6(32'h3aada1c9),
	.w7(32'h39776804),
	.w8(32'hbab2ee5e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170f0b),
	.w1(32'h3b0781c4),
	.w2(32'h3a4a7053),
	.w3(32'h3a29626e),
	.w4(32'hba6614a4),
	.w5(32'hba5559d1),
	.w6(32'h3ab4966e),
	.w7(32'h3a7fea1c),
	.w8(32'h3a17d65b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c79755),
	.w1(32'h391a12af),
	.w2(32'h3a2592ff),
	.w3(32'h39a28355),
	.w4(32'h396f7105),
	.w5(32'h3932f73a),
	.w6(32'h39a32c61),
	.w7(32'h3a013e5a),
	.w8(32'h394f197a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977df58),
	.w1(32'hb94baf7f),
	.w2(32'hba2d0b2b),
	.w3(32'h37ab3a17),
	.w4(32'hb88628e9),
	.w5(32'hba3c8aee),
	.w6(32'hb9bd5085),
	.w7(32'hba40f323),
	.w8(32'hba11b455),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a0d40),
	.w1(32'hba882412),
	.w2(32'h3a540672),
	.w3(32'hba7b771d),
	.w4(32'h39bc648b),
	.w5(32'hba3ff83e),
	.w6(32'h3ac444fb),
	.w7(32'hba901bd8),
	.w8(32'hb9e1a068),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288cc1),
	.w1(32'h3aea342b),
	.w2(32'hbb24f79b),
	.w3(32'h3a01d004),
	.w4(32'h389a854e),
	.w5(32'hb9f3eda2),
	.w6(32'h3aefb091),
	.w7(32'h3aef955e),
	.w8(32'h3b8c5e68),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d59155),
	.w1(32'h3ac14c1c),
	.w2(32'h3a4eda28),
	.w3(32'h39cd9bf2),
	.w4(32'h3aa4d4ed),
	.w5(32'h3a609a26),
	.w6(32'h3b396bb0),
	.w7(32'h3b33ad62),
	.w8(32'h3b2fe873),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161118),
	.w1(32'hbb98d924),
	.w2(32'hbb36fd10),
	.w3(32'hba416752),
	.w4(32'hb9861bfe),
	.w5(32'hba02d361),
	.w6(32'h3afb7b49),
	.w7(32'h3b2ae055),
	.w8(32'h3ac29622),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29a036),
	.w1(32'hb865f401),
	.w2(32'h3ac434ff),
	.w3(32'h3a5c0290),
	.w4(32'hba736fac),
	.w5(32'hba1cc151),
	.w6(32'hb853158b),
	.w7(32'hb9d44422),
	.w8(32'h3938bc66),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d7e2c),
	.w1(32'h3a1ef64f),
	.w2(32'h3a3ff963),
	.w3(32'h39104156),
	.w4(32'h3a146ddf),
	.w5(32'h399c6bc0),
	.w6(32'h3a4d04cd),
	.w7(32'h3a0ac1c8),
	.w8(32'h39e5a00a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9990e8),
	.w1(32'hbb5e8949),
	.w2(32'h3aa0566c),
	.w3(32'h3ad292b1),
	.w4(32'hbaa3241b),
	.w5(32'h3b4f7b2d),
	.w6(32'hb9bd89f8),
	.w7(32'hbb6c39f1),
	.w8(32'hbb08657f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd071),
	.w1(32'hb9f0313c),
	.w2(32'hb861ddb2),
	.w3(32'h3ab2e6fd),
	.w4(32'h390c4f04),
	.w5(32'h3a06829b),
	.w6(32'hb9d7d242),
	.w7(32'hb93a1c71),
	.w8(32'h381a32b5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff3359),
	.w1(32'hbb7b4d1f),
	.w2(32'hbb47d343),
	.w3(32'h3acdcf04),
	.w4(32'hba4b148c),
	.w5(32'hba56cf8a),
	.w6(32'h3afaadfa),
	.w7(32'h3ad57be4),
	.w8(32'h3a9b0390),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9922e65),
	.w1(32'h3a029e56),
	.w2(32'hb8ed275b),
	.w3(32'hba5f21fb),
	.w4(32'h3a462b2a),
	.w5(32'h3955300e),
	.w6(32'h3a16691d),
	.w7(32'h38a9d0d1),
	.w8(32'h375006e9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f45e9),
	.w1(32'h39a09067),
	.w2(32'hb74a37fc),
	.w3(32'hb90f9d3f),
	.w4(32'h398c3119),
	.w5(32'hb925ffb9),
	.w6(32'h39ee6857),
	.w7(32'hb815df33),
	.w8(32'hb8dbb6f4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a593e5c),
	.w1(32'h3a5a13f6),
	.w2(32'h3a5cd377),
	.w3(32'hb78acb9d),
	.w4(32'hb95017f9),
	.w5(32'hba57207b),
	.w6(32'h39ccbf3b),
	.w7(32'h3a80768a),
	.w8(32'hb9a034eb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005675),
	.w1(32'hbb62118d),
	.w2(32'hbb69b520),
	.w3(32'hba6da223),
	.w4(32'hbb175cae),
	.w5(32'hbb65b530),
	.w6(32'hba61fcb3),
	.w7(32'hbab0fb1e),
	.w8(32'h3aa42921),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64e065),
	.w1(32'h3a94dee4),
	.w2(32'hb90a4728),
	.w3(32'h3a04016e),
	.w4(32'hb8fe8399),
	.w5(32'hba5ea787),
	.w6(32'hba081789),
	.w7(32'hbab75c78),
	.w8(32'hbac7e8d1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55c742),
	.w1(32'h3a8ac7b8),
	.w2(32'h3b04d789),
	.w3(32'h3a03871a),
	.w4(32'hb97dfc14),
	.w5(32'hba8f76db),
	.w6(32'h3b034755),
	.w7(32'h3ab714b4),
	.w8(32'h39c61b16),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc303fd8),
	.w1(32'h3b697a57),
	.w2(32'h3b957e90),
	.w3(32'h3b0b63d4),
	.w4(32'h3c160f6a),
	.w5(32'h3b58e163),
	.w6(32'h398c1c34),
	.w7(32'h3bc3a69e),
	.w8(32'h3b808f57),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9894ca),
	.w1(32'hbbb89a0d),
	.w2(32'hbb4bb60a),
	.w3(32'h3b2485fd),
	.w4(32'h3b5f3d90),
	.w5(32'h3b0c8c72),
	.w6(32'h3bd23993),
	.w7(32'h3bd0edee),
	.w8(32'h3b4c7e83),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a380),
	.w1(32'hbb9b6545),
	.w2(32'hbb88565a),
	.w3(32'h3b601632),
	.w4(32'h3b53eaa4),
	.w5(32'h3b131882),
	.w6(32'h3b9ea1af),
	.w7(32'h3b6ef56c),
	.w8(32'h3ab828c5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384e1ed1),
	.w1(32'h39fe9bc6),
	.w2(32'hb905ca72),
	.w3(32'h3a36462d),
	.w4(32'h3aad6b4f),
	.w5(32'h3a537a43),
	.w6(32'h3ae62728),
	.w7(32'h3a6daa0c),
	.w8(32'h3a19b205),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a175179),
	.w1(32'h3a3c8e9d),
	.w2(32'h39f5c82d),
	.w3(32'h3a80180f),
	.w4(32'hb923cfa5),
	.w5(32'hb9e65c61),
	.w6(32'h39c91d7d),
	.w7(32'h39b044e6),
	.w8(32'h3971aa35),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988bc55),
	.w1(32'h38b53b1a),
	.w2(32'hb9814c1f),
	.w3(32'hba68a387),
	.w4(32'h393327a3),
	.w5(32'hb91a7f06),
	.w6(32'hb8c07ce6),
	.w7(32'hba3885ec),
	.w8(32'h380d136a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc89e9),
	.w1(32'hb915a8d7),
	.w2(32'hb9998d03),
	.w3(32'h39cff28f),
	.w4(32'hb991f5eb),
	.w5(32'hb9afcba7),
	.w6(32'hb8bc5e72),
	.w7(32'hb9c5bb7f),
	.w8(32'hba1f398b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27dc42),
	.w1(32'h3a623a3d),
	.w2(32'hbb165add),
	.w3(32'hba2af835),
	.w4(32'hbabad769),
	.w5(32'h3a0e7b25),
	.w6(32'hba4dae5a),
	.w7(32'hbb508d2d),
	.w8(32'h3a788496),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb433650),
	.w1(32'hbac8b4bf),
	.w2(32'h3a9baf84),
	.w3(32'hba482245),
	.w4(32'h3b06079e),
	.w5(32'h3b232c7b),
	.w6(32'h3b111610),
	.w7(32'h3b285b25),
	.w8(32'h3b3cb875),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6c2f5),
	.w1(32'hb9cc8701),
	.w2(32'h3b2e3079),
	.w3(32'hb9b3c3d6),
	.w4(32'h3abe1ab1),
	.w5(32'h3a53d594),
	.w6(32'h3b62f686),
	.w7(32'h3b8aed35),
	.w8(32'h3b8c72b7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925eb87),
	.w1(32'h3a8b561f),
	.w2(32'hba98d86d),
	.w3(32'h39d88c51),
	.w4(32'h3a4a24f3),
	.w5(32'h3a3c1bb3),
	.w6(32'h3aaa9882),
	.w7(32'h3ad194cd),
	.w8(32'h3afca88c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1c3ab),
	.w1(32'h3b8c55c8),
	.w2(32'h3b326df6),
	.w3(32'h3b5f3bed),
	.w4(32'hba56afce),
	.w5(32'hbaec2c20),
	.w6(32'h3a001bf0),
	.w7(32'h392cd85c),
	.w8(32'hba3456bc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a707001),
	.w1(32'hb8f2ecb0),
	.w2(32'h377a1438),
	.w3(32'h3a8787e8),
	.w4(32'hb9367f09),
	.w5(32'hb9910b7a),
	.w6(32'h38d4bb04),
	.w7(32'hb9879463),
	.w8(32'hb9e6fd51),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9d63d),
	.w1(32'h3a6cb86b),
	.w2(32'h39bf6307),
	.w3(32'hb9db18d6),
	.w4(32'h3a9947c6),
	.w5(32'h3a87461f),
	.w6(32'h3ab75a12),
	.w7(32'h3a818c9d),
	.w8(32'h3a8dd8b5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a519eb3),
	.w1(32'h3b0f0d8f),
	.w2(32'h3b030e6b),
	.w3(32'h3a98bb4a),
	.w4(32'h3b18785d),
	.w5(32'h3b1a0c15),
	.w6(32'h3addd207),
	.w7(32'h3b045369),
	.w8(32'h3b249618),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421c8a),
	.w1(32'hb9a18b83),
	.w2(32'hb9c9ed56),
	.w3(32'h3adf6653),
	.w4(32'h3867dce5),
	.w5(32'h3b0fd917),
	.w6(32'hb938d9fa),
	.w7(32'h3a5b4820),
	.w8(32'h3b38ec5a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cba96),
	.w1(32'hb8133b95),
	.w2(32'hbadca8de),
	.w3(32'h3b1a74a9),
	.w4(32'hb9a8c148),
	.w5(32'hba98bb00),
	.w6(32'hb794a62e),
	.w7(32'hba71c381),
	.w8(32'hb99f8b45),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b613c),
	.w1(32'h3b864459),
	.w2(32'h3ac24acc),
	.w3(32'h3adeacb2),
	.w4(32'hba3d7da4),
	.w5(32'hbb0a5328),
	.w6(32'h3a15171f),
	.w7(32'h3948ab7a),
	.w8(32'hbb1cdc82),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182c7a),
	.w1(32'hba6afbac),
	.w2(32'hba3d0c38),
	.w3(32'hbabc33ff),
	.w4(32'hbad30ff9),
	.w5(32'hb9913334),
	.w6(32'hb98785e9),
	.w7(32'hb98893b1),
	.w8(32'h38880d8a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba351211),
	.w1(32'h39260a83),
	.w2(32'h37df98ba),
	.w3(32'hba81b1a3),
	.w4(32'hb90cdf13),
	.w5(32'hba237dc0),
	.w6(32'hb8cd0ae4),
	.w7(32'h390bfe2a),
	.w8(32'hba197e07),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac3770),
	.w1(32'h3acc2485),
	.w2(32'h3a1a34dd),
	.w3(32'hba8b23e9),
	.w4(32'h3ac497a9),
	.w5(32'h3a7cff8e),
	.w6(32'h3aa0cbe2),
	.w7(32'h3a5df146),
	.w8(32'h3a60a7a2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64b1f9),
	.w1(32'h38c69530),
	.w2(32'hbab0ec4f),
	.w3(32'h3a2bc9e1),
	.w4(32'hb917f81b),
	.w5(32'hba26170d),
	.w6(32'h3ab814a8),
	.w7(32'h39c3c224),
	.w8(32'h39021d2f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf23074),
	.w1(32'h3a441fe5),
	.w2(32'h3914812e),
	.w3(32'hb9b702c6),
	.w4(32'h3aad4931),
	.w5(32'h3a50fbfb),
	.w6(32'h3a84909f),
	.w7(32'h3a13cd45),
	.w8(32'h3a135e36),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9faba8),
	.w1(32'h3a960f8b),
	.w2(32'h3a501a5e),
	.w3(32'h3ab61b1d),
	.w4(32'h3a838ff6),
	.w5(32'h3a401d77),
	.w6(32'h3aa0c076),
	.w7(32'h3a59e1c4),
	.w8(32'h3a5f73e9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f4b2),
	.w1(32'h3b1b029c),
	.w2(32'hb98a982d),
	.w3(32'h3a629424),
	.w4(32'hb8b55c6b),
	.w5(32'hba56ab9a),
	.w6(32'h3ae397bf),
	.w7(32'h390d60fd),
	.w8(32'hb861b55d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac14009),
	.w1(32'hbad20801),
	.w2(32'hbabc332b),
	.w3(32'hba63ac51),
	.w4(32'hbb62a5c4),
	.w5(32'h3a86d2a0),
	.w6(32'hb9636022),
	.w7(32'hbb065ae7),
	.w8(32'h38851d1b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c090e1),
	.w1(32'hbaeb0cb6),
	.w2(32'hbac0f814),
	.w3(32'h3a9d3da0),
	.w4(32'hbac12406),
	.w5(32'hbab6b3b1),
	.w6(32'hba3a19a6),
	.w7(32'hbaeec76b),
	.w8(32'hbab0abc3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb82ba),
	.w1(32'hba07a33e),
	.w2(32'hba11894b),
	.w3(32'h397cb597),
	.w4(32'hb80f94f1),
	.w5(32'hb9a020ce),
	.w6(32'hb9f8f0c2),
	.w7(32'hb9e3fafd),
	.w8(32'hb8ffc9ee),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc3337),
	.w1(32'hb93b185d),
	.w2(32'hb9b466b3),
	.w3(32'hb8317252),
	.w4(32'hb89df0ef),
	.w5(32'hb9b9c43e),
	.w6(32'h3992113a),
	.w7(32'h39881f4c),
	.w8(32'h38e8ff29),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cbd07),
	.w1(32'hb6e8ae56),
	.w2(32'h3a5922a3),
	.w3(32'hb89b59b9),
	.w4(32'hba0bf430),
	.w5(32'hba5e1ed3),
	.w6(32'hb9b7a0ab),
	.w7(32'h3963fc40),
	.w8(32'h39eab2a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b792238),
	.w1(32'h3c11eda0),
	.w2(32'h3a3c2e90),
	.w3(32'h3b8fd637),
	.w4(32'h3967fdf6),
	.w5(32'hbb050fd3),
	.w6(32'hbba857f5),
	.w7(32'hbb9457b1),
	.w8(32'hbc2589e3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ddd5c),
	.w1(32'h3a702994),
	.w2(32'hbab43afe),
	.w3(32'hbb98fb00),
	.w4(32'hbbad0f95),
	.w5(32'hbbe94603),
	.w6(32'h3b60d4f4),
	.w7(32'h3b04bd82),
	.w8(32'hb8d159ec),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae66331),
	.w1(32'hb8e59878),
	.w2(32'hbb339d62),
	.w3(32'hbb32412a),
	.w4(32'hbb0cb3cc),
	.w5(32'hb9c4aef4),
	.w6(32'h3a7dac64),
	.w7(32'h39e99cad),
	.w8(32'h3b324e13),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5560),
	.w1(32'hbb774a71),
	.w2(32'hba9ba6c3),
	.w3(32'hb9e5d73c),
	.w4(32'h3a8acf86),
	.w5(32'h3adbe963),
	.w6(32'h3bc6b59e),
	.w7(32'h3bd692fa),
	.w8(32'h3bbbdb1c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addd733),
	.w1(32'h3a42de52),
	.w2(32'h3998d1af),
	.w3(32'h3aebb938),
	.w4(32'h3a590bd6),
	.w5(32'h3a1b7f79),
	.w6(32'h3a6bb6c0),
	.w7(32'h39e6d21d),
	.w8(32'h39d3400e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3d064),
	.w1(32'h3a323542),
	.w2(32'h394d79c2),
	.w3(32'h3a375307),
	.w4(32'h3a6ec94b),
	.w5(32'h3a16f3ba),
	.w6(32'h3a976e47),
	.w7(32'h3a1e0249),
	.w8(32'h3a432887),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d52c6),
	.w1(32'h3a4a1b75),
	.w2(32'h3a19ba18),
	.w3(32'h39eb90e8),
	.w4(32'h3a7fe9bb),
	.w5(32'h3a52c32b),
	.w6(32'h3a73c08d),
	.w7(32'h3a671479),
	.w8(32'h3a624f02),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb44b8),
	.w1(32'h3a77d569),
	.w2(32'h37df0ee0),
	.w3(32'h3a04097a),
	.w4(32'hb874b282),
	.w5(32'hba486349),
	.w6(32'h3a082c01),
	.w7(32'hba22c1e5),
	.w8(32'hba6d99fa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b2d24),
	.w1(32'h3a5f1493),
	.w2(32'h39e52519),
	.w3(32'hb99c94f1),
	.w4(32'h3abe09a5),
	.w5(32'h3abfea22),
	.w6(32'h3aa4c874),
	.w7(32'h3a7f2f55),
	.w8(32'h3a8379fb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f4fec),
	.w1(32'h3b67a745),
	.w2(32'h3b97c6bb),
	.w3(32'h3b51f9c1),
	.w4(32'h3b0da461),
	.w5(32'h3b19dd79),
	.w6(32'h398ab7c8),
	.w7(32'h3a711520),
	.w8(32'h3a8eaf50),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74382d),
	.w1(32'h3b4eb969),
	.w2(32'h3b4526f8),
	.w3(32'h3b09868e),
	.w4(32'hba160931),
	.w5(32'hbae9b7b4),
	.w6(32'h3a2ce393),
	.w7(32'h3aa58126),
	.w8(32'h393f53ec),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc6136),
	.w1(32'hbb0a0dd8),
	.w2(32'hbaaa8667),
	.w3(32'h39e47aea),
	.w4(32'h393f83e2),
	.w5(32'h39488889),
	.w6(32'h3a5e7f22),
	.w7(32'h3aada965),
	.w8(32'h3ac538b4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36c0f2),
	.w1(32'hba8f80c5),
	.w2(32'hbaa7aedb),
	.w3(32'h3873a9e9),
	.w4(32'hbb0f45ab),
	.w5(32'hbaf8e4b9),
	.w6(32'hb8a46f9b),
	.w7(32'hba1e57d0),
	.w8(32'hbae6c961),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908772e),
	.w1(32'h3b9e1c23),
	.w2(32'h3b070f60),
	.w3(32'h3b1534d6),
	.w4(32'h3b12947c),
	.w5(32'h39887219),
	.w6(32'hbade0fa1),
	.w7(32'hbae5d0a1),
	.w8(32'hbb72c048),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b4e5a),
	.w1(32'hbaf81f1b),
	.w2(32'hbaca4313),
	.w3(32'hb9ae57c3),
	.w4(32'h392dcc19),
	.w5(32'h3a388b02),
	.w6(32'hb90ba70d),
	.w7(32'h39ec77f2),
	.w8(32'h3a69a1b9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81bd8f),
	.w1(32'h3b133b5f),
	.w2(32'h3a052cb8),
	.w3(32'h39940116),
	.w4(32'h3a8caf25),
	.w5(32'h39925b40),
	.w6(32'h3ad85780),
	.w7(32'h3a2eee54),
	.w8(32'h3a935706),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49eb82),
	.w1(32'hba999730),
	.w2(32'hba85794f),
	.w3(32'h3aa79286),
	.w4(32'hb9c04d14),
	.w5(32'hb9fda9e1),
	.w6(32'hba89f587),
	.w7(32'hba9cf4d1),
	.w8(32'hba80289b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c9fc9),
	.w1(32'h3a1cc71e),
	.w2(32'h384d9071),
	.w3(32'hba29a99d),
	.w4(32'h3a5400aa),
	.w5(32'h3995fc6f),
	.w6(32'h3a98cc11),
	.w7(32'h3a41555f),
	.w8(32'h3a235d97),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f503a),
	.w1(32'hb9eef938),
	.w2(32'hba40de57),
	.w3(32'h3a4a0fcc),
	.w4(32'h3a0a61ac),
	.w5(32'h39835e41),
	.w6(32'hb9a5e528),
	.w7(32'hba44d489),
	.w8(32'hba250b0e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a9c8b),
	.w1(32'hb9d1877e),
	.w2(32'hba7270f9),
	.w3(32'h3a880d07),
	.w4(32'hb92f48e8),
	.w5(32'hba03b312),
	.w6(32'h39c202d6),
	.w7(32'hb99c5514),
	.w8(32'hb9f006a5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bba2e),
	.w1(32'hbaacf3d9),
	.w2(32'hb9d275d9),
	.w3(32'hba4dc1f6),
	.w4(32'h3b166e91),
	.w5(32'h3a809ea5),
	.w6(32'h3b10fe45),
	.w7(32'h3b07336a),
	.w8(32'h3b2967b8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f9901),
	.w1(32'h39964b20),
	.w2(32'hb715036c),
	.w3(32'h3a28221e),
	.w4(32'h39b42e8e),
	.w5(32'hb90bfbe9),
	.w6(32'h38ae6efd),
	.w7(32'hb94919be),
	.w8(32'hb99af40b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba971cbc),
	.w1(32'hbb091c45),
	.w2(32'hba874cfd),
	.w3(32'hba8599c2),
	.w4(32'hba71bbd6),
	.w5(32'hba6ee7a0),
	.w6(32'h3aa2f850),
	.w7(32'h3a83c322),
	.w8(32'h3a1fd484),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a9ef),
	.w1(32'h3b036a8d),
	.w2(32'h38da08ce),
	.w3(32'h39e819ba),
	.w4(32'hba33c7df),
	.w5(32'hbaf85300),
	.w6(32'h3ace9bd6),
	.w7(32'h3a797564),
	.w8(32'h386766e4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09603a),
	.w1(32'hbafa4fad),
	.w2(32'hbab460cf),
	.w3(32'h3ab5805e),
	.w4(32'h3b0d343b),
	.w5(32'h3ab464c2),
	.w6(32'h3b0e3dde),
	.w7(32'h3ac92670),
	.w8(32'h3a4581a8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43e638),
	.w1(32'h3bbcd910),
	.w2(32'h3abfe675),
	.w3(32'h3b79b34d),
	.w4(32'h3bde1b71),
	.w5(32'h3b05d448),
	.w6(32'h38d802ed),
	.w7(32'h3a661683),
	.w8(32'hbb5bba0f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309572),
	.w1(32'hba904553),
	.w2(32'hba8c7fd3),
	.w3(32'h3a64a7fb),
	.w4(32'h3afdefa4),
	.w5(32'h3ae8fe35),
	.w6(32'h3b885b41),
	.w7(32'h3b5e9ad6),
	.w8(32'h3b59861f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7628),
	.w1(32'hba150b14),
	.w2(32'hbb94c61b),
	.w3(32'h38eb45c7),
	.w4(32'hbb1c734b),
	.w5(32'hbba0dc61),
	.w6(32'hb9849bfd),
	.w7(32'hbaf59ff7),
	.w8(32'hbb95703b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f2ea2),
	.w1(32'h3a3308f3),
	.w2(32'hba937bfa),
	.w3(32'h39f5df09),
	.w4(32'h3b043dc7),
	.w5(32'hb9003148),
	.w6(32'h3aa432a8),
	.w7(32'h377917e0),
	.w8(32'hbac01e91),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8b6c7),
	.w1(32'hb990ed54),
	.w2(32'hbaa75838),
	.w3(32'h3a01bc91),
	.w4(32'h3ac56b53),
	.w5(32'hbaa9bb30),
	.w6(32'h3af6ba34),
	.w7(32'h3a6b8a61),
	.w8(32'hb9d683cc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac401c),
	.w1(32'h3a13b680),
	.w2(32'h39ac4c34),
	.w3(32'hba24c7ec),
	.w4(32'hb988dc5e),
	.w5(32'h39bae919),
	.w6(32'h3a2c42fb),
	.w7(32'hb9cb7806),
	.w8(32'hb9e5abda),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6305),
	.w1(32'h39e0bd8b),
	.w2(32'hba1ee5ba),
	.w3(32'h382b0b96),
	.w4(32'hbb426787),
	.w5(32'hbb0cf207),
	.w6(32'hba247497),
	.w7(32'hba5a3a19),
	.w8(32'h39fc8147),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba155d84),
	.w1(32'h3b834311),
	.w2(32'h3ae5450a),
	.w3(32'h3b70cc74),
	.w4(32'h3baf3373),
	.w5(32'h3b830a6e),
	.w6(32'hbaaabd88),
	.w7(32'hb87fc01c),
	.w8(32'hba1c73a6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4c6bc),
	.w1(32'hbb81a42e),
	.w2(32'hbb79e36a),
	.w3(32'hba7a55ba),
	.w4(32'hb9af2d5f),
	.w5(32'hbc11680a),
	.w6(32'h3b25385b),
	.w7(32'h3abb7c3b),
	.w8(32'h3b0ec7a6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ba26),
	.w1(32'hbba163f3),
	.w2(32'hbb86de01),
	.w3(32'h3a17092c),
	.w4(32'hbab453bd),
	.w5(32'hbb0415cf),
	.w6(32'h3b1330d2),
	.w7(32'hb86b652c),
	.w8(32'hba0baa58),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856b2a),
	.w1(32'hbb0a94c8),
	.w2(32'h3b2c9f35),
	.w3(32'hbaed3cfe),
	.w4(32'h3b13b4bd),
	.w5(32'h3b03a9f1),
	.w6(32'h3b5b1db6),
	.w7(32'h3b8dff59),
	.w8(32'h3b8b2c2b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba970d96),
	.w1(32'h3bb82fc6),
	.w2(32'h3b898bce),
	.w3(32'h3b3378ae),
	.w4(32'h3bcb5692),
	.w5(32'h3aafc61f),
	.w6(32'h39dc8a2a),
	.w7(32'h3b0a7a96),
	.w8(32'h3a60d275),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ddc0e),
	.w1(32'h3aa449b4),
	.w2(32'h39221b64),
	.w3(32'h3ad1a750),
	.w4(32'h3a86816d),
	.w5(32'h3a31e2ce),
	.w6(32'h3aa6ad6e),
	.w7(32'h3a49407a),
	.w8(32'h3a578f0c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4d4a),
	.w1(32'hbbd147a3),
	.w2(32'h3aebedfd),
	.w3(32'hba1c59a2),
	.w4(32'h3ada41e7),
	.w5(32'hbc013a7e),
	.w6(32'h3a9deade),
	.w7(32'h3aaf3800),
	.w8(32'h3b499cf0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2a409),
	.w1(32'h3b430a41),
	.w2(32'h3b31fb15),
	.w3(32'h3b637d7d),
	.w4(32'h3b6791f1),
	.w5(32'h3ac16f7f),
	.w6(32'hb9836ae2),
	.w7(32'h39d3feb5),
	.w8(32'h3ad309ae),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b9b17),
	.w1(32'hb976c988),
	.w2(32'hb98b4b62),
	.w3(32'hb8a00d1b),
	.w4(32'h392bed46),
	.w5(32'hb9bd6601),
	.w6(32'h39a1c5a7),
	.w7(32'hb9d67f58),
	.w8(32'hb9f9dd92),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86367d),
	.w1(32'hbab78432),
	.w2(32'hba98ac0b),
	.w3(32'h390226d6),
	.w4(32'h3a48a077),
	.w5(32'hb929d2ad),
	.w6(32'h3a80c85a),
	.w7(32'h39a5690a),
	.w8(32'hb94e7074),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a562a70),
	.w1(32'h3b16cd3c),
	.w2(32'h3a8304e2),
	.w3(32'hb8fc273f),
	.w4(32'h3a580aa8),
	.w5(32'hb8806cd5),
	.w6(32'h3b0695c9),
	.w7(32'h3aa0dc65),
	.w8(32'h3a400081),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58ecfa),
	.w1(32'h38cec3dc),
	.w2(32'h3a4b756c),
	.w3(32'h3a303ffa),
	.w4(32'h3b3dc39e),
	.w5(32'h3b4ff22b),
	.w6(32'h3b406007),
	.w7(32'h3b44b782),
	.w8(32'h3b61ac47),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4b8cc),
	.w1(32'hbad69992),
	.w2(32'hba3c50ad),
	.w3(32'h3b695d61),
	.w4(32'h3b22c51b),
	.w5(32'h3aeef66d),
	.w6(32'h3add6542),
	.w7(32'h3b1a3069),
	.w8(32'h3aba54ca),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea3815),
	.w1(32'hbb28c44d),
	.w2(32'hbaa51c63),
	.w3(32'h3a04884e),
	.w4(32'hba310e20),
	.w5(32'h39cd1b31),
	.w6(32'h3972ac62),
	.w7(32'h3a9fad6c),
	.w8(32'h395e6c6d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2000f),
	.w1(32'h3b3a0be1),
	.w2(32'h3b8bb668),
	.w3(32'hb8b9cdf9),
	.w4(32'h3a3d1c3d),
	.w5(32'hba4ca0bb),
	.w6(32'h3b89f39c),
	.w7(32'h3b8a8df0),
	.w8(32'h3b14b595),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41d590),
	.w1(32'hba97382e),
	.w2(32'hbbaa0e1d),
	.w3(32'h3a7c429a),
	.w4(32'hbaad45e0),
	.w5(32'hbb2701e9),
	.w6(32'hba3e3a30),
	.w7(32'hbada1c3c),
	.w8(32'hbb059890),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcd18c),
	.w1(32'h3a8cf3ca),
	.w2(32'h3ae582b0),
	.w3(32'h3a609e73),
	.w4(32'h3aff4c8a),
	.w5(32'h3b16c598),
	.w6(32'h3b09c8f9),
	.w7(32'h3b1f7c42),
	.w8(32'h3b228926),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0bc05),
	.w1(32'h3a534400),
	.w2(32'h3a5aa8d2),
	.w3(32'h3ab2b08b),
	.w4(32'h3a9b60ba),
	.w5(32'h3a88c4af),
	.w6(32'h3aaf1782),
	.w7(32'h3a8eba4c),
	.w8(32'h3a993f3a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18d1bc),
	.w1(32'h393a1897),
	.w2(32'hb9545147),
	.w3(32'h3a5243a9),
	.w4(32'h39d08829),
	.w5(32'h3939e79b),
	.w6(32'h3a7272c9),
	.w7(32'h3a4c23e4),
	.w8(32'h397c167d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a84da9),
	.w1(32'h39c0eba2),
	.w2(32'h38dcd05c),
	.w3(32'h3a06c02c),
	.w4(32'h3a0363a9),
	.w5(32'h39a64a77),
	.w6(32'h3a8526f0),
	.w7(32'h3a19b22d),
	.w8(32'h39f227e2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961a853),
	.w1(32'h39d3d05c),
	.w2(32'h39f007f3),
	.w3(32'h39e75cc8),
	.w4(32'h3a1c5fcb),
	.w5(32'h3a2dec99),
	.w6(32'h3a9ca170),
	.w7(32'hb9a78f3c),
	.w8(32'hba183531),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0495c1),
	.w1(32'hba190d52),
	.w2(32'h3ade27e6),
	.w3(32'h39c94b1d),
	.w4(32'h393c5b3d),
	.w5(32'h3ab9e971),
	.w6(32'h3a939031),
	.w7(32'h3b453c79),
	.w8(32'h3b41e9dd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce7ef),
	.w1(32'h3a466464),
	.w2(32'hb9d1ea27),
	.w3(32'h39b96049),
	.w4(32'h3a6bb49c),
	.w5(32'hb897c177),
	.w6(32'h3a18b99d),
	.w7(32'hba23c042),
	.w8(32'hba0ccc9e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f37b2),
	.w1(32'h3af1339e),
	.w2(32'h3a52798d),
	.w3(32'h3a4e0d13),
	.w4(32'hb9605d26),
	.w5(32'hb98636f4),
	.w6(32'hb94bb359),
	.w7(32'hb9bc2613),
	.w8(32'hba3dc1b1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a05c),
	.w1(32'hbb09baee),
	.w2(32'hbb1ae422),
	.w3(32'hbab29bee),
	.w4(32'h3aa0d998),
	.w5(32'hb9bca931),
	.w6(32'h3b76c900),
	.w7(32'h3b418a57),
	.w8(32'h3a88c0a7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a783cb0),
	.w1(32'h39fc7ee5),
	.w2(32'h3af43f32),
	.w3(32'h3a930504),
	.w4(32'h3a5af285),
	.w5(32'hba0c270e),
	.w6(32'h38d81df6),
	.w7(32'hb9de6961),
	.w8(32'hb9a0e911),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4191),
	.w1(32'h39de4724),
	.w2(32'hbaf77c33),
	.w3(32'hba621384),
	.w4(32'h3a8b20c3),
	.w5(32'hb9d99a2e),
	.w6(32'h3a846981),
	.w7(32'hb9c38253),
	.w8(32'hb9622b99),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f8cc),
	.w1(32'h3933df1b),
	.w2(32'hb9c5f4a9),
	.w3(32'hb9f09b79),
	.w4(32'h3a046155),
	.w5(32'hb9489c58),
	.w6(32'h39ae358d),
	.w7(32'hb9b7f331),
	.w8(32'hb9632e79),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdb2e2),
	.w1(32'hbb9451c4),
	.w2(32'h39cc6901),
	.w3(32'hba1e52ff),
	.w4(32'hba8cc3c5),
	.w5(32'hbb2e8196),
	.w6(32'h3b8bdddd),
	.w7(32'h3c025090),
	.w8(32'h3af659a1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd413ec),
	.w1(32'h38c7fe43),
	.w2(32'h3bca645b),
	.w3(32'hbb26d6ca),
	.w4(32'hbb298d04),
	.w5(32'hbb8756a9),
	.w6(32'h3becc878),
	.w7(32'h3c33c838),
	.w8(32'h3aa30dae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb3449),
	.w1(32'h3c31f0e8),
	.w2(32'hbbd5ad80),
	.w3(32'h3b2ab7ef),
	.w4(32'h3c7db55c),
	.w5(32'hbafaec41),
	.w6(32'hbc8397bc),
	.w7(32'hbc8492b7),
	.w8(32'h3b814b19),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6107),
	.w1(32'h3c58e34c),
	.w2(32'h3aab8561),
	.w3(32'hbc21c932),
	.w4(32'h3b80bd9d),
	.w5(32'h3b962359),
	.w6(32'h3b47bb34),
	.w7(32'hbbec9139),
	.w8(32'hbbc8cd75),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb69a6),
	.w1(32'h3b332b21),
	.w2(32'hba591036),
	.w3(32'hb7e0249b),
	.w4(32'hb9f354ea),
	.w5(32'hb8722c2e),
	.w6(32'hbb03da0b),
	.w7(32'hbb6eee35),
	.w8(32'hbb3daf72),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ebd3),
	.w1(32'h3aebbbb7),
	.w2(32'h3c224e72),
	.w3(32'h3a1af2f9),
	.w4(32'hbbc8c263),
	.w5(32'hbc4ed0ba),
	.w6(32'h3bde9c2b),
	.w7(32'hbc2ff8be),
	.w8(32'hbc6de6ea),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe15bab),
	.w1(32'hb950def0),
	.w2(32'h3d141834),
	.w3(32'hbb753997),
	.w4(32'hba864a0f),
	.w5(32'h3ba0b631),
	.w6(32'h3a62dec6),
	.w7(32'h3b67f8e9),
	.w8(32'hbc3bb5bc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b957),
	.w1(32'hb8c0c47d),
	.w2(32'hba931f9f),
	.w3(32'h3b9caf1f),
	.w4(32'h3be6fe32),
	.w5(32'h3b496ae3),
	.w6(32'h3842a9e4),
	.w7(32'hbb4b1877),
	.w8(32'hbc16101d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7e29b),
	.w1(32'h3c493c58),
	.w2(32'h3bacbb17),
	.w3(32'h3b1b94ea),
	.w4(32'hb9d2bc40),
	.w5(32'h3bff5a9d),
	.w6(32'h3b2af08e),
	.w7(32'hbbbf05d7),
	.w8(32'hbbd0efca),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf34997),
	.w1(32'hbbf329ac),
	.w2(32'h3931a1ee),
	.w3(32'h3b5b623f),
	.w4(32'hb9902dee),
	.w5(32'hbb24bc48),
	.w6(32'h3b446513),
	.w7(32'h3bc940d7),
	.w8(32'h3a6a9c56),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad612c),
	.w1(32'h3acfb92e),
	.w2(32'hba963e66),
	.w3(32'hb9c76d5c),
	.w4(32'h3baab343),
	.w5(32'hb998c6b7),
	.w6(32'h3a995670),
	.w7(32'h3b27604d),
	.w8(32'hbb0d68d9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08197e),
	.w1(32'h3c99ac8a),
	.w2(32'h3a31d888),
	.w3(32'hb935149e),
	.w4(32'h3b86d142),
	.w5(32'h3b126674),
	.w6(32'h3b154a0d),
	.w7(32'hbc34e7ad),
	.w8(32'hbbafbd28),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058a6a),
	.w1(32'hbc6c6b85),
	.w2(32'hbc583310),
	.w3(32'h3a8db503),
	.w4(32'hbbf9e280),
	.w5(32'hbc3ba246),
	.w6(32'hbc2b2f2e),
	.w7(32'hbb4a9ddf),
	.w8(32'h3baec95f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc567ced),
	.w1(32'h3c11a589),
	.w2(32'h3c00b8ea),
	.w3(32'hbc06c340),
	.w4(32'h3a372ae6),
	.w5(32'hbbac72f6),
	.w6(32'h3c00c561),
	.w7(32'hba3bdd13),
	.w8(32'hbc51e3bb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ea84),
	.w1(32'hbbaf54dc),
	.w2(32'hbb01ddf7),
	.w3(32'h3b81297f),
	.w4(32'h3ab2e0db),
	.w5(32'h3a8a1831),
	.w6(32'hbadada29),
	.w7(32'h3b73bc06),
	.w8(32'h3adc2cb9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe999f),
	.w1(32'hbc6e2371),
	.w2(32'h3a9e8ecf),
	.w3(32'hba485ab0),
	.w4(32'hbbf5be80),
	.w5(32'hbc36b6d6),
	.w6(32'h3bed962c),
	.w7(32'h3c883918),
	.w8(32'h3bbd418c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e0b0a),
	.w1(32'hbbd3e770),
	.w2(32'h3d2c50ed),
	.w3(32'hbb129549),
	.w4(32'hbc38a836),
	.w5(32'hbbd39f6c),
	.w6(32'h3b56ce04),
	.w7(32'h39d226c6),
	.w8(32'hbcbcacc3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0898b9),
	.w1(32'h3ac44b94),
	.w2(32'hbb267266),
	.w3(32'h3aee3a79),
	.w4(32'h3b6ffe2c),
	.w5(32'h390cbeef),
	.w6(32'hb9dc5beb),
	.w7(32'hbb22bfcd),
	.w8(32'hbb7692e1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eeb6e4),
	.w1(32'h3a9c8db4),
	.w2(32'hba6fd81d),
	.w3(32'hb946a121),
	.w4(32'hbb95b801),
	.w5(32'hbb3710f9),
	.w6(32'hbb8cfb7a),
	.w7(32'hbac08ec7),
	.w8(32'h3b104176),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b78d),
	.w1(32'h3c260ac0),
	.w2(32'h3ae4717a),
	.w3(32'hb9cc8bc1),
	.w4(32'hba26315b),
	.w5(32'h3b3a596a),
	.w6(32'hb8832d04),
	.w7(32'hbc1de39c),
	.w8(32'hbbc8013f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd9f27),
	.w1(32'h3b215a25),
	.w2(32'h3a295efb),
	.w3(32'h3ae561aa),
	.w4(32'h3b48495b),
	.w5(32'h3b27f9d7),
	.w6(32'h3b0adacd),
	.w7(32'hbb9e14cd),
	.w8(32'hbb935e32),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828c37),
	.w1(32'h3aad36ad),
	.w2(32'hbb3c49ad),
	.w3(32'hbb04fe89),
	.w4(32'h3b234405),
	.w5(32'hbb23a014),
	.w6(32'hb97205e8),
	.w7(32'hba8e5a3e),
	.w8(32'hbacddb22),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b6ea7),
	.w1(32'hbc1a1e38),
	.w2(32'hbbb28c66),
	.w3(32'hbb4d036c),
	.w4(32'hbb204659),
	.w5(32'hbb6ca507),
	.w6(32'h3a3f7a82),
	.w7(32'h3bcbc5b0),
	.w8(32'h3c024508),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc47546),
	.w1(32'h3a9f973c),
	.w2(32'hbc3b9f8b),
	.w3(32'hb994c2e2),
	.w4(32'hbaaf8da2),
	.w5(32'h3b765671),
	.w6(32'h3aab334c),
	.w7(32'h3b67d22b),
	.w8(32'hba167b82),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f277),
	.w1(32'h3acee0be),
	.w2(32'hbb1940f5),
	.w3(32'hbbab9087),
	.w4(32'h3b9557cc),
	.w5(32'h3ab5376e),
	.w6(32'h3be247f6),
	.w7(32'h3a80633f),
	.w8(32'h3b17f7d8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27853),
	.w1(32'hbaac46d5),
	.w2(32'hb9c63295),
	.w3(32'h3bcc08e4),
	.w4(32'h3b611bbf),
	.w5(32'hba5c2ee7),
	.w6(32'hb9933db4),
	.w7(32'h3b9d7a08),
	.w8(32'hba863be7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a10b2),
	.w1(32'h3ba43812),
	.w2(32'hbbe37764),
	.w3(32'h3ab26e09),
	.w4(32'h3bc5dd03),
	.w5(32'h3b690275),
	.w6(32'h3baf6f52),
	.w7(32'hbb0ade28),
	.w8(32'hbb482eba),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe133a),
	.w1(32'h3b351765),
	.w2(32'hbb3a022d),
	.w3(32'hbabe829a),
	.w4(32'hbc0ff4a3),
	.w5(32'hbbcc6801),
	.w6(32'hbaac53f1),
	.w7(32'h3a2d41de),
	.w8(32'hbb12dae9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d5187),
	.w1(32'hba864a7b),
	.w2(32'hbb515e11),
	.w3(32'hbace6112),
	.w4(32'h3aa7bc44),
	.w5(32'hbad66d22),
	.w6(32'hb982a6ff),
	.w7(32'h3a71bcfe),
	.w8(32'h3aa7714c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979d4b6),
	.w1(32'h3c4a5c2c),
	.w2(32'h3a84880b),
	.w3(32'hbaf619a1),
	.w4(32'h3b681986),
	.w5(32'hbb2bd841),
	.w6(32'h3b3e5a88),
	.w7(32'hbbcb1886),
	.w8(32'hbb9bc8a4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb297da5),
	.w1(32'h3b9a7f8b),
	.w2(32'hbc0b82f6),
	.w3(32'h3a907289),
	.w4(32'h3ba45e39),
	.w5(32'hbbc83dcd),
	.w6(32'h3c549c3a),
	.w7(32'hbb25fdde),
	.w8(32'h3b0423ac),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3589),
	.w1(32'h3b710b61),
	.w2(32'h3b38d467),
	.w3(32'hbaf1cecb),
	.w4(32'hbb2d0d83),
	.w5(32'h3ab21b24),
	.w6(32'hba97df49),
	.w7(32'h390c499b),
	.w8(32'hbba5a4fa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b546430),
	.w1(32'hbb8e78ca),
	.w2(32'hbb2e34d4),
	.w3(32'h3b4536d5),
	.w4(32'hba052eb5),
	.w5(32'hba8c475f),
	.w6(32'h38413251),
	.w7(32'h3b421112),
	.w8(32'h3bcb6c5c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7386bc),
	.w1(32'hbb32d6a1),
	.w2(32'hbb172c24),
	.w3(32'hba2e7d1f),
	.w4(32'h3a38bf48),
	.w5(32'hba68e35f),
	.w6(32'h374c3e45),
	.w7(32'h3b5d486b),
	.w8(32'h3b31f6da),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7faa00),
	.w1(32'h3c043d52),
	.w2(32'hbc158562),
	.w3(32'h3a4153f1),
	.w4(32'h3b9b04c5),
	.w5(32'hbc08a2a5),
	.w6(32'h3a226d0b),
	.w7(32'hbc138b27),
	.w8(32'hbb8038f7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04a39b),
	.w1(32'h3c17dc49),
	.w2(32'h3c86bbd2),
	.w3(32'hbbbdc3ee),
	.w4(32'h3be4eb2d),
	.w5(32'h3c6f6384),
	.w6(32'h3b72ca49),
	.w7(32'h3c047b41),
	.w8(32'hbbcc2fb7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989406),
	.w1(32'h3c4410e8),
	.w2(32'hbae3e72f),
	.w3(32'hbc03177c),
	.w4(32'h3b31c3bf),
	.w5(32'h3b2495aa),
	.w6(32'h3aa40c20),
	.w7(32'hbc413848),
	.w8(32'hbbd7122c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e5059),
	.w1(32'hb88739f5),
	.w2(32'h3a823871),
	.w3(32'hba543aad),
	.w4(32'h3aad2ca7),
	.w5(32'hba6fa428),
	.w6(32'h3a994e85),
	.w7(32'h3af688a7),
	.w8(32'h3b71c49d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36883),
	.w1(32'h3c73ed9d),
	.w2(32'h3c2f31d6),
	.w3(32'hbaf5f568),
	.w4(32'h3aa70b27),
	.w5(32'h3a53b62c),
	.w6(32'h3bac149e),
	.w7(32'hbb9d7712),
	.w8(32'hbc1da42d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824775),
	.w1(32'h3c081ea2),
	.w2(32'h3ad87f38),
	.w3(32'h3aa1bb3b),
	.w4(32'h3b5fd7bd),
	.w5(32'h3bdccd35),
	.w6(32'h3b009ab9),
	.w7(32'hbbad95d7),
	.w8(32'hbb8f4fdf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b46e7),
	.w1(32'hbb4794ac),
	.w2(32'hba83f2cd),
	.w3(32'h3b433a44),
	.w4(32'h3b1d8d3f),
	.w5(32'hba57eede),
	.w6(32'h3ae9adfb),
	.w7(32'h3b32bb0a),
	.w8(32'h3a5b49ab),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cdeae),
	.w1(32'h3b85b336),
	.w2(32'h3b9a2251),
	.w3(32'h3a8e789a),
	.w4(32'h3ac7f1fa),
	.w5(32'h3b5c2dbd),
	.w6(32'h3b7dc9c7),
	.w7(32'hbb4cc1af),
	.w8(32'hbbb9a465),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c132),
	.w1(32'h3beff9d9),
	.w2(32'h3b90daac),
	.w3(32'hbad163fa),
	.w4(32'h3a8b0658),
	.w5(32'h3adf6d6e),
	.w6(32'h3bc5b71a),
	.w7(32'h3ba91751),
	.w8(32'hba0fff40),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80b30b),
	.w1(32'h3b3ca674),
	.w2(32'h3b0b27fd),
	.w3(32'h3b39610f),
	.w4(32'hbb861f03),
	.w5(32'hbb66109d),
	.w6(32'h3b0ab6da),
	.w7(32'hbb0fd98e),
	.w8(32'hbbbc7014),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ba07),
	.w1(32'hba75ba5e),
	.w2(32'hbb19efcc),
	.w3(32'hbb7505d1),
	.w4(32'h3b47bf21),
	.w5(32'hbae32b5d),
	.w6(32'h3b02bf5c),
	.w7(32'h3b7010cb),
	.w8(32'h3b1ebe6e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a818e8a),
	.w1(32'h3c9ee877),
	.w2(32'h3b8fba3e),
	.w3(32'h38bfc7e0),
	.w4(32'h3bea04cb),
	.w5(32'h3c3f875c),
	.w6(32'h3b96c598),
	.w7(32'hbbf70e28),
	.w8(32'hbaaeb17b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bc33e),
	.w1(32'hbbbbb22f),
	.w2(32'hbc0df83a),
	.w3(32'h3c023545),
	.w4(32'hbb1d3d7e),
	.w5(32'hb9c039b1),
	.w6(32'hbbbf1f6c),
	.w7(32'hbb595cfe),
	.w8(32'h3b6ba7ba),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d50dd),
	.w1(32'hbbb99700),
	.w2(32'hbb92586a),
	.w3(32'hba28a9e5),
	.w4(32'h3b3e6c22),
	.w5(32'h3b8e1115),
	.w6(32'h3a8f160b),
	.w7(32'hbb49a9e2),
	.w8(32'hbbca2b85),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceec6c),
	.w1(32'h3c137f74),
	.w2(32'h3d0d52c9),
	.w3(32'h3a2d83ea),
	.w4(32'hb987d8b5),
	.w5(32'hbb081de3),
	.w6(32'h3c219a5f),
	.w7(32'hbb489662),
	.w8(32'hbc8edf10),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76620a),
	.w1(32'h3ba8d22e),
	.w2(32'hb8bfa0c2),
	.w3(32'h3ad3c195),
	.w4(32'hb97c1439),
	.w5(32'h3b0cf1fa),
	.w6(32'h3be8022d),
	.w7(32'h3ba2eea7),
	.w8(32'h3b36beae),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f8f0),
	.w1(32'h39f15024),
	.w2(32'hbb87b352),
	.w3(32'hbb1747a2),
	.w4(32'h3b1137c8),
	.w5(32'hbb39be40),
	.w6(32'hbaf88789),
	.w7(32'hba17fd50),
	.w8(32'hba59dd94),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fab98),
	.w1(32'hbbcc60d6),
	.w2(32'h3918326a),
	.w3(32'hba176088),
	.w4(32'hba0bc59d),
	.w5(32'hbb5cf1f5),
	.w6(32'h3b53bbaa),
	.w7(32'h3c072ed3),
	.w8(32'h3b73a98e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb511d1),
	.w1(32'hba976d97),
	.w2(32'h39b7ad70),
	.w3(32'h39c3cd4f),
	.w4(32'hbb8ad507),
	.w5(32'hbb647e21),
	.w6(32'h3acbb0e8),
	.w7(32'h3a98fa81),
	.w8(32'hba07a83b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0135b),
	.w1(32'h3c7ca508),
	.w2(32'hbcbd70bf),
	.w3(32'hbb928556),
	.w4(32'h3c4dd60f),
	.w5(32'hbba49b01),
	.w6(32'h39a0f4e3),
	.w7(32'hbc760700),
	.w8(32'hbc1c69bd),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f58f3),
	.w1(32'h3996c092),
	.w2(32'hbc120862),
	.w3(32'hbb6ac24f),
	.w4(32'hbab4dd00),
	.w5(32'hbb340e18),
	.w6(32'hbb29ccf8),
	.w7(32'hbc235ebc),
	.w8(32'hbc2397d2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb65875),
	.w1(32'h3bba26f3),
	.w2(32'h3c961264),
	.w3(32'hbb4960d0),
	.w4(32'h3bd2ef33),
	.w5(32'h3c2f9cad),
	.w6(32'h3bf1d03d),
	.w7(32'h3b95121b),
	.w8(32'hbc2bad58),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819c9f),
	.w1(32'h3b7d923f),
	.w2(32'hbadce6b5),
	.w3(32'h3b495888),
	.w4(32'h3b1635c6),
	.w5(32'hba67ca93),
	.w6(32'hbb9873bc),
	.w7(32'hbbb0a834),
	.w8(32'hbba395e3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb54dd5),
	.w1(32'hbb108d93),
	.w2(32'hbb1c39bc),
	.w3(32'hbb155e7d),
	.w4(32'h3afaee36),
	.w5(32'h39310439),
	.w6(32'h3bb1865d),
	.w7(32'h37f15ef3),
	.w8(32'h3b3c286a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9550ce),
	.w1(32'hbb21fbf0),
	.w2(32'hbbe78aef),
	.w3(32'h3ac05c36),
	.w4(32'h3a4710cc),
	.w5(32'hba9de1b2),
	.w6(32'hba9cfbf7),
	.w7(32'h3b04c973),
	.w8(32'hba207140),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e6aa),
	.w1(32'hbb792ea5),
	.w2(32'h3d070206),
	.w3(32'h3b055a5b),
	.w4(32'hba25a310),
	.w5(32'h3b4ed78b),
	.w6(32'h3c1e70b9),
	.w7(32'h3bdbff6f),
	.w8(32'hbc4c6a62),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06293e),
	.w1(32'h3c4ef531),
	.w2(32'hbb1fd1d6),
	.w3(32'hbb401e90),
	.w4(32'h3b322a02),
	.w5(32'h3b31a310),
	.w6(32'h3aefcab7),
	.w7(32'hbc0faedb),
	.w8(32'hbb6f5205),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af958),
	.w1(32'hb9f70950),
	.w2(32'hbb096d75),
	.w3(32'hba677d2e),
	.w4(32'hb9988288),
	.w5(32'hbb9eedfb),
	.w6(32'h3adafa4a),
	.w7(32'h3b4b99f3),
	.w8(32'h39202bdb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a76fe0),
	.w1(32'h3bc6eefd),
	.w2(32'h3be380b0),
	.w3(32'h3b3d7449),
	.w4(32'h3bac501c),
	.w5(32'h3c102e8e),
	.w6(32'h3afc4305),
	.w7(32'hbb30b7a5),
	.w8(32'hbbd8452a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaba1c8),
	.w1(32'hbb8bbbbc),
	.w2(32'hbb375217),
	.w3(32'h3b14f068),
	.w4(32'h39cb69ab),
	.w5(32'hbb5bed39),
	.w6(32'hbb29109a),
	.w7(32'h3b8dfae0),
	.w8(32'h3bcc0ad1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8cbb3),
	.w1(32'hb98e064c),
	.w2(32'h3b5eb36c),
	.w3(32'hbb0cc2f9),
	.w4(32'hbc04fc09),
	.w5(32'h3a8af6b0),
	.w6(32'hbbebe065),
	.w7(32'hbb89377b),
	.w8(32'hbc1c2b95),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc846203),
	.w1(32'h3c6c142d),
	.w2(32'h3b14ee22),
	.w3(32'hbbf0fd16),
	.w4(32'h3b9e7215),
	.w5(32'h3be6edab),
	.w6(32'h3b1ffa92),
	.w7(32'hbbecfd1a),
	.w8(32'hbb22081f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb326a39),
	.w1(32'h3b5c7da6),
	.w2(32'hb991bfdd),
	.w3(32'h3ba03506),
	.w4(32'h3b23f368),
	.w5(32'hba620c61),
	.w6(32'h3a5b4980),
	.w7(32'hbb34b327),
	.w8(32'hbb87a85e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f7745),
	.w1(32'hba3587d6),
	.w2(32'h3c8ad124),
	.w3(32'h3b611f33),
	.w4(32'h3c030824),
	.w5(32'h3c29b275),
	.w6(32'h3c305e35),
	.w7(32'h3bf6329b),
	.w8(32'hbc07ca5b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a5d8),
	.w1(32'hba87867e),
	.w2(32'h3a4df7da),
	.w3(32'hbb820871),
	.w4(32'hbb597578),
	.w5(32'h36ce872f),
	.w6(32'hbba0ed57),
	.w7(32'hbb5b4b73),
	.w8(32'hbc05743e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb508bc),
	.w1(32'h3adcb7a0),
	.w2(32'hbac02995),
	.w3(32'h3694ca98),
	.w4(32'h3bdca945),
	.w5(32'h3b94285e),
	.w6(32'h3c510869),
	.w7(32'h3bd222a3),
	.w8(32'h3ba745df),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0423a4),
	.w1(32'hbacac362),
	.w2(32'hbafc56d6),
	.w3(32'h3b6a33f0),
	.w4(32'h3b2e8ef9),
	.w5(32'hb9305e19),
	.w6(32'h3aafc769),
	.w7(32'h3aa9615a),
	.w8(32'h3a4876d1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd84c6),
	.w1(32'hbab762ad),
	.w2(32'h3c84ea14),
	.w3(32'h3b23b05e),
	.w4(32'hbbfab7d6),
	.w5(32'h3af635c0),
	.w6(32'h3c50462f),
	.w7(32'h3c6964d3),
	.w8(32'hba23657f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdad5b4),
	.w1(32'h3bd0cbaa),
	.w2(32'h3a57fa6c),
	.w3(32'h3765cbd8),
	.w4(32'h3adbf4ba),
	.w5(32'h3b87a0d9),
	.w6(32'h3a20a1a7),
	.w7(32'hbbfcf729),
	.w8(32'hbb7d5124),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5f84),
	.w1(32'hbbe785c4),
	.w2(32'h3ad42839),
	.w3(32'hb947ff65),
	.w4(32'hbaddd0e8),
	.w5(32'hb988779e),
	.w6(32'hba280d52),
	.w7(32'h3b5eac68),
	.w8(32'hba2b70d7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7940),
	.w1(32'hbbd198a2),
	.w2(32'hbbb407f6),
	.w3(32'hbb1c16a9),
	.w4(32'hb90f85e7),
	.w5(32'hbb915c9b),
	.w6(32'h386f535b),
	.w7(32'h3a624135),
	.w8(32'hb92d3e47),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b2f1a),
	.w1(32'hbb36346a),
	.w2(32'hbb839aaa),
	.w3(32'h3a1fbb6f),
	.w4(32'h3a85c313),
	.w5(32'hba74d029),
	.w6(32'hb941c113),
	.w7(32'h3abaa6f1),
	.w8(32'h3b89fc8c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14b716),
	.w1(32'h3c738045),
	.w2(32'hbb95d3a3),
	.w3(32'hba9d4323),
	.w4(32'h3b685086),
	.w5(32'h3acef377),
	.w6(32'h3b1cbbd2),
	.w7(32'hbc1c3616),
	.w8(32'hbc0115ee),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b89d0),
	.w1(32'h3b455937),
	.w2(32'hbc3002ab),
	.w3(32'hbb290275),
	.w4(32'hbbb32692),
	.w5(32'hbc8af359),
	.w6(32'h3c2af754),
	.w7(32'hbb704a7b),
	.w8(32'hbbc72928),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79f15a),
	.w1(32'hbc2aabf5),
	.w2(32'hb9664e78),
	.w3(32'hbb8d8cf4),
	.w4(32'h38212eb0),
	.w5(32'hbb8381da),
	.w6(32'h3b7a0de4),
	.w7(32'h3c18509e),
	.w8(32'h3ba0c2d7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2ef9f),
	.w1(32'h3ba126dc),
	.w2(32'h3a97c73a),
	.w3(32'hb9590aa8),
	.w4(32'hb9c07404),
	.w5(32'h3b75fc48),
	.w6(32'hbb0373ea),
	.w7(32'hbba07829),
	.w8(32'hbb88ea0f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4f58),
	.w1(32'h39d66f7d),
	.w2(32'hbb23c42c),
	.w3(32'hbaf0085d),
	.w4(32'hbb10039f),
	.w5(32'hbb9c108d),
	.w6(32'hbbc2aa1d),
	.w7(32'hba8ad76e),
	.w8(32'h39cbe2f5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a2094),
	.w1(32'hbbdbdb03),
	.w2(32'hbb608cf1),
	.w3(32'hbadddb14),
	.w4(32'hbb30bc40),
	.w5(32'hbb858b25),
	.w6(32'h3b142030),
	.w7(32'h3ba7cc0c),
	.w8(32'h3bc10f0d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baea6e2),
	.w1(32'h3ae483a6),
	.w2(32'hbb31be01),
	.w3(32'h39157ef8),
	.w4(32'h3bae36df),
	.w5(32'h3b26e1d5),
	.w6(32'h3c41e552),
	.w7(32'h3b86c5ee),
	.w8(32'h3b5d1c8a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa58543),
	.w1(32'h3c19be70),
	.w2(32'h3b733d1d),
	.w3(32'h3ab26edb),
	.w4(32'h3a91f8e5),
	.w5(32'h3bc7bcd0),
	.w6(32'h3b63d5b0),
	.w7(32'hbb7bb81d),
	.w8(32'hbb9fc5b8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc46d9d),
	.w1(32'h3c1244bf),
	.w2(32'h3ae078d0),
	.w3(32'hb9943009),
	.w4(32'h3ac6eba4),
	.w5(32'h3a6ea5ea),
	.w6(32'h3b84dfb7),
	.w7(32'h3988fea0),
	.w8(32'h39ffb6e6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95d8bc),
	.w1(32'h3c39eb24),
	.w2(32'h3b821b16),
	.w3(32'h3a3fba02),
	.w4(32'h3b6f5739),
	.w5(32'h3b8651bc),
	.w6(32'h3b35262a),
	.w7(32'hbb4ab309),
	.w8(32'hbb74c4a1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8799c1),
	.w1(32'hbb9bf10f),
	.w2(32'hbb5fcd99),
	.w3(32'hbad46e0b),
	.w4(32'hbbdb8f16),
	.w5(32'hbb69be44),
	.w6(32'hbb452cd3),
	.w7(32'h3a95fe17),
	.w8(32'h385c9077),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe41293),
	.w1(32'hba2ae61a),
	.w2(32'hbaafeb97),
	.w3(32'hbc066f19),
	.w4(32'hbaa05b4c),
	.w5(32'h3b137a6b),
	.w6(32'h3a578bae),
	.w7(32'h3a3c4d7f),
	.w8(32'hbabb1e81),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e86a21),
	.w1(32'h3c02d93b),
	.w2(32'h3b08fc6f),
	.w3(32'h3bb1ac6d),
	.w4(32'hbae76dee),
	.w5(32'hbb0b1dff),
	.w6(32'hb916776b),
	.w7(32'h3b554c54),
	.w8(32'hbb9e33ce),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338c87),
	.w1(32'hbb863de1),
	.w2(32'hbb8bf7a0),
	.w3(32'hbb8fc027),
	.w4(32'hba97fdfb),
	.w5(32'hbb0701bf),
	.w6(32'hb9803573),
	.w7(32'h3b2bc635),
	.w8(32'h3b9d64ed),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ddd7),
	.w1(32'h3bac10ef),
	.w2(32'hbb86f48a),
	.w3(32'hba19ee09),
	.w4(32'h3ab45145),
	.w5(32'hba853f01),
	.w6(32'hbad09210),
	.w7(32'hbbc1b10f),
	.w8(32'hbbe087b5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9631f0),
	.w1(32'h3a04053f),
	.w2(32'h3b7a7563),
	.w3(32'hbaa4b362),
	.w4(32'h3aaf9c02),
	.w5(32'hbb821a40),
	.w6(32'h3b8ca2df),
	.w7(32'h3c144ed2),
	.w8(32'h3c087bea),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc004),
	.w1(32'hbaa19999),
	.w2(32'hbb7cd00f),
	.w3(32'h37e78581),
	.w4(32'hbb5b1537),
	.w5(32'hbb932821),
	.w6(32'h394cdfaa),
	.w7(32'h3b813e5f),
	.w8(32'h3bdc1cd1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ef96),
	.w1(32'h3b8a693e),
	.w2(32'h3ab2e56e),
	.w3(32'h3a467d2c),
	.w4(32'h3ab24f7a),
	.w5(32'h3b1f6eb1),
	.w6(32'hbafce52f),
	.w7(32'hbb4323de),
	.w8(32'hbb6ba932),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab77ec6),
	.w1(32'h3bc171de),
	.w2(32'hbac6596f),
	.w3(32'h3aebc0bd),
	.w4(32'h3b3f60f2),
	.w5(32'h3b551a0b),
	.w6(32'h3b02d7d3),
	.w7(32'hbb8f929a),
	.w8(32'hbb231dfe),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aa99a),
	.w1(32'h3b14048c),
	.w2(32'hbc15f8fc),
	.w3(32'hbb401067),
	.w4(32'h3c219b9c),
	.w5(32'hbabc65fd),
	.w6(32'h3c883377),
	.w7(32'h3b31d2eb),
	.w8(32'h3b810525),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef63f7),
	.w1(32'h3bb1579d),
	.w2(32'h3b245085),
	.w3(32'h3ad90439),
	.w4(32'h3b335bb5),
	.w5(32'h3b0a3b6d),
	.w6(32'hba6fd84b),
	.w7(32'hbb724af9),
	.w8(32'hbb8a4ce2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbffd66),
	.w1(32'hbb6fd679),
	.w2(32'hbbc74f7b),
	.w3(32'hb97e90d1),
	.w4(32'h3bc5b44f),
	.w5(32'h3bb48d63),
	.w6(32'h39d56c1e),
	.w7(32'h397ff583),
	.w8(32'hbbaf2b71),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc357b3a),
	.w1(32'hbb7adf17),
	.w2(32'hbaf10bc3),
	.w3(32'hbb69c4fb),
	.w4(32'hbb5c9e27),
	.w5(32'hbb89ab8e),
	.w6(32'hbb31173d),
	.w7(32'hba00fab5),
	.w8(32'h3b0b407a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e39e64),
	.w1(32'h3c11f8ce),
	.w2(32'hbad14c2a),
	.w3(32'hbb199784),
	.w4(32'h3c227683),
	.w5(32'hba396d13),
	.w6(32'hb9e42dc3),
	.w7(32'hbaf0aac6),
	.w8(32'hbb8d693e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde51c),
	.w1(32'h3c00c3f3),
	.w2(32'h3ba92868),
	.w3(32'hbb0f270a),
	.w4(32'hbacbc6ac),
	.w5(32'h3a3a73bf),
	.w6(32'h3b4bb3aa),
	.w7(32'hbbe254b4),
	.w8(32'hbc11d38f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c4cc),
	.w1(32'h3c3e825a),
	.w2(32'hba0f28c0),
	.w3(32'hbbbea761),
	.w4(32'h3a7c9514),
	.w5(32'h3ab6b00d),
	.w6(32'h3ba53abd),
	.w7(32'hbb2d987d),
	.w8(32'hbbeba129),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6dcb1),
	.w1(32'hbca30c65),
	.w2(32'h3b3e8768),
	.w3(32'hba7289e2),
	.w4(32'hbb9e50b6),
	.w5(32'hbc6f86fa),
	.w6(32'hbc005835),
	.w7(32'hbc4c603a),
	.w8(32'hbc806f83),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27693d),
	.w1(32'hbbcdaaed),
	.w2(32'h3a0e8f05),
	.w3(32'hbc822a71),
	.w4(32'hb991466c),
	.w5(32'h3c55ae14),
	.w6(32'h3ba97fd7),
	.w7(32'h3c2551b6),
	.w8(32'hbbeee2dd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc556047),
	.w1(32'hbc2657e2),
	.w2(32'h3b5bac6b),
	.w3(32'h3adf8856),
	.w4(32'h39b5e723),
	.w5(32'hbc138a31),
	.w6(32'h3ba24840),
	.w7(32'h3c7d9ef0),
	.w8(32'h3b87a87b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55b609),
	.w1(32'hbb819af1),
	.w2(32'h3a3adbd0),
	.w3(32'h3a2f9822),
	.w4(32'hbb21d583),
	.w5(32'hbb6426a2),
	.w6(32'h3a9101ab),
	.w7(32'h3a6647da),
	.w8(32'hbb8c5968),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1023e7),
	.w1(32'hbbd9c21f),
	.w2(32'hb9e19a9a),
	.w3(32'hbaf2a6e8),
	.w4(32'h39c110ea),
	.w5(32'hbb586410),
	.w6(32'h3b0d53b2),
	.w7(32'h3bb23bbc),
	.w8(32'h3b291ed2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca9569),
	.w1(32'h3b3c7049),
	.w2(32'hbaaa6b3a),
	.w3(32'h3a877994),
	.w4(32'h3b575e60),
	.w5(32'hbae48a5b),
	.w6(32'h398a7fd9),
	.w7(32'h3aada86e),
	.w8(32'h38a44e59),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32610c),
	.w1(32'h3bede832),
	.w2(32'hbb15e4ef),
	.w3(32'hbb2d9ae0),
	.w4(32'h3a54db3f),
	.w5(32'h3ace2c5b),
	.w6(32'hbb4d8079),
	.w7(32'hbbe1445c),
	.w8(32'hbbd24261),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf08ec),
	.w1(32'hbbfc8a4c),
	.w2(32'hbbe075bf),
	.w3(32'hbaba8410),
	.w4(32'hbb0af27a),
	.w5(32'hbb7d35e9),
	.w6(32'hbafe03cc),
	.w7(32'h3b8cddfc),
	.w8(32'h3c1749b5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baba584),
	.w1(32'hbc052910),
	.w2(32'h39a7c9a5),
	.w3(32'hba988ede),
	.w4(32'hba1c673b),
	.w5(32'hbb680a4d),
	.w6(32'h3b2ee2a0),
	.w7(32'h3be8d1c2),
	.w8(32'h3b384fb9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc04bb4),
	.w1(32'h3b907408),
	.w2(32'hbb41c03f),
	.w3(32'hb9f5d009),
	.w4(32'h39fe873a),
	.w5(32'hba9ddf91),
	.w6(32'h3b1e7731),
	.w7(32'hbb435215),
	.w8(32'hbc0739f0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ba8b),
	.w1(32'h3ab91420),
	.w2(32'hbba325e2),
	.w3(32'h3a40be5e),
	.w4(32'h3b9ab2a2),
	.w5(32'hba59c180),
	.w6(32'h3b15788c),
	.w7(32'hba89b6ef),
	.w8(32'hba6b7aa5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac715ba),
	.w1(32'hbafe59b0),
	.w2(32'h3a1c8a13),
	.w3(32'h3bb3ce7e),
	.w4(32'hbb88d977),
	.w5(32'hbbd98a59),
	.w6(32'hbc82036c),
	.w7(32'hbc585a9e),
	.w8(32'h3a9621f4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210a3b),
	.w1(32'h3bc963f6),
	.w2(32'hbb07f8bd),
	.w3(32'hbba016a4),
	.w4(32'h3ba3b3ea),
	.w5(32'h3a51c235),
	.w6(32'h3a01c78a),
	.w7(32'hbb638a71),
	.w8(32'hbbbdea0c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b114005),
	.w1(32'h3c1fcc27),
	.w2(32'hbabe5673),
	.w3(32'h3bb235c0),
	.w4(32'h3b25e254),
	.w5(32'hbb010d08),
	.w6(32'h39e21a50),
	.w7(32'hbbce7f96),
	.w8(32'hbb9f5664),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff62f2),
	.w1(32'hbb83d5ec),
	.w2(32'hbb56d640),
	.w3(32'hbae0e8f4),
	.w4(32'h3b87f5c9),
	.w5(32'hbb04d209),
	.w6(32'hbac4ace0),
	.w7(32'hbae4ad7a),
	.w8(32'h3aa8200c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eccf6),
	.w1(32'hbc35b8be),
	.w2(32'hba723692),
	.w3(32'hba11afd8),
	.w4(32'hba5461af),
	.w5(32'hbbc2a790),
	.w6(32'h3b7e7f85),
	.w7(32'h3c15dde5),
	.w8(32'h3b6c18f4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01632c),
	.w1(32'hbbf1b327),
	.w2(32'hbab13810),
	.w3(32'hb98000f4),
	.w4(32'h3a9cba9e),
	.w5(32'hbab49314),
	.w6(32'hba9fd6f0),
	.w7(32'h3b2ca9e1),
	.w8(32'h3a14f94f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77049),
	.w1(32'hbbca7d09),
	.w2(32'hba814f5b),
	.w3(32'hbaaa85d6),
	.w4(32'h3b055a78),
	.w5(32'hba86f50c),
	.w6(32'hb9daa071),
	.w7(32'h3b173847),
	.w8(32'h3a477685),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5279bd),
	.w1(32'hbc361082),
	.w2(32'hbc4b9e8e),
	.w3(32'hbac275c7),
	.w4(32'h3a663137),
	.w5(32'hbb86b2bd),
	.w6(32'hbc10d5c9),
	.w7(32'hbb24358c),
	.w8(32'h3a9f189b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e51a6),
	.w1(32'h3a00bded),
	.w2(32'h3adaaf04),
	.w3(32'hbc289df5),
	.w4(32'h3bd9057b),
	.w5(32'h3b9250ef),
	.w6(32'h3b3571e4),
	.w7(32'hbc1965a2),
	.w8(32'hbb4e4c21),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1dd22),
	.w1(32'hbba4aa3a),
	.w2(32'h3a6d8b46),
	.w3(32'h3a5638e6),
	.w4(32'hb9dc849d),
	.w5(32'hbb7ce067),
	.w6(32'hbb0051a9),
	.w7(32'hbae8c7de),
	.w8(32'hbb0751d6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc3423),
	.w1(32'hba4ee44d),
	.w2(32'hbba71b58),
	.w3(32'hbb193621),
	.w4(32'h3a345cb1),
	.w5(32'hbb0be5ad),
	.w6(32'hba293007),
	.w7(32'hbb1c647f),
	.w8(32'hbad403a2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6131ae),
	.w1(32'hbbae906c),
	.w2(32'hbb206771),
	.w3(32'hbb796086),
	.w4(32'h3aede6cd),
	.w5(32'hbb1882f0),
	.w6(32'h3943864b),
	.w7(32'h3b763bc7),
	.w8(32'h3ab04128),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f8d52),
	.w1(32'hbb819f4e),
	.w2(32'hbc8908eb),
	.w3(32'hb9f0ad06),
	.w4(32'h3bf56c78),
	.w5(32'hbaed1545),
	.w6(32'hbbd5f258),
	.w7(32'hbc2f4760),
	.w8(32'hbb8e0dbc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9afe2e),
	.w1(32'h3bda0248),
	.w2(32'hb9919d6d),
	.w3(32'hbc173531),
	.w4(32'h3c18461f),
	.w5(32'h3b9a814e),
	.w6(32'h3ad95841),
	.w7(32'hbbabf7a1),
	.w8(32'hbbf5f151),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bf18f),
	.w1(32'hbb95e649),
	.w2(32'hbbd777f5),
	.w3(32'hbb4221e5),
	.w4(32'hbb48fcf9),
	.w5(32'hbb7e7c86),
	.w6(32'hbaa44f69),
	.w7(32'h3a14a339),
	.w8(32'h3b43db90),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b640b1f),
	.w1(32'h38cfeb86),
	.w2(32'h39c28de1),
	.w3(32'hba64998d),
	.w4(32'hb9003774),
	.w5(32'h3a008f16),
	.w6(32'h3820bbb6),
	.w7(32'h391a2abf),
	.w8(32'hba0b5e22),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb03ea),
	.w1(32'hb8bc2235),
	.w2(32'h3b0123c2),
	.w3(32'h39d12be6),
	.w4(32'hb90a6c47),
	.w5(32'hb9ec825f),
	.w6(32'h3b6f5e69),
	.w7(32'h3b6bdac4),
	.w8(32'h3b16932f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule