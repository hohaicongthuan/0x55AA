module layer_10_featuremap_304(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b052b7d),
	.w1(32'hbb61804c),
	.w2(32'h3b4977de),
	.w3(32'hbac817d9),
	.w4(32'h3a6b41ca),
	.w5(32'hbb5f73d8),
	.w6(32'hba2d159e),
	.w7(32'h3b9a9989),
	.w8(32'hba639ca8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6eee4),
	.w1(32'h3b477cf1),
	.w2(32'h3b5d7608),
	.w3(32'hbae71a00),
	.w4(32'h3b51aa8b),
	.w5(32'hbb596465),
	.w6(32'hbbbaf73c),
	.w7(32'hbb75d70a),
	.w8(32'h3bb2a27b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f9595),
	.w1(32'h3ca477bb),
	.w2(32'h3c70d2b7),
	.w3(32'h3b38c1a0),
	.w4(32'h3bec2d88),
	.w5(32'h3b252b37),
	.w6(32'h3cb22ff4),
	.w7(32'h3ca324f1),
	.w8(32'hb9316923),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35b81b),
	.w1(32'h3b8f0cd2),
	.w2(32'h3a94dc1b),
	.w3(32'h398ac1d5),
	.w4(32'h3a7dc144),
	.w5(32'hbb31c966),
	.w6(32'hba0e2db2),
	.w7(32'hb9bdbb5a),
	.w8(32'h399c924b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa95d80),
	.w1(32'hbb6794e1),
	.w2(32'hbab507fb),
	.w3(32'hbbc289a0),
	.w4(32'hbbadaf6b),
	.w5(32'h3ae0a6e4),
	.w6(32'hba076a02),
	.w7(32'h3bd44ce1),
	.w8(32'h3adebad3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54943d),
	.w1(32'h3af78b94),
	.w2(32'h3b71e6c6),
	.w3(32'h3ad0bb2d),
	.w4(32'h3b17f706),
	.w5(32'hba88bf06),
	.w6(32'h3b355761),
	.w7(32'h3be4c5c1),
	.w8(32'hbb0ac507),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bdf5e),
	.w1(32'hbc2218fa),
	.w2(32'hbc206710),
	.w3(32'hbbe4fec8),
	.w4(32'hbc58d3ab),
	.w5(32'h3a4624ab),
	.w6(32'hbbf965bd),
	.w7(32'hbc0e0d98),
	.w8(32'h39057d76),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0c9e1),
	.w1(32'h3c2ff357),
	.w2(32'h3c9c1624),
	.w3(32'hbb9a2fc4),
	.w4(32'h3ca1f83b),
	.w5(32'h3c90ea03),
	.w6(32'h3b8ee810),
	.w7(32'h3b7309dc),
	.w8(32'h3b6f20fd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1757d6),
	.w1(32'hb91046d3),
	.w2(32'h3b274104),
	.w3(32'hbac6c6f0),
	.w4(32'hba1b790e),
	.w5(32'h3b1f48c5),
	.w6(32'hb9ac3886),
	.w7(32'h3b6b33bc),
	.w8(32'h3af9d2e0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94acb6),
	.w1(32'hbacca2fc),
	.w2(32'hb9bcb8c9),
	.w3(32'hbb5734f9),
	.w4(32'hba1169fb),
	.w5(32'h3b26d45e),
	.w6(32'hbb8acf81),
	.w7(32'h3aacf8f6),
	.w8(32'hbb752c9f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980db59),
	.w1(32'h3b823472),
	.w2(32'h3bf4b8ae),
	.w3(32'h3b6b4ef2),
	.w4(32'h3b58b71a),
	.w5(32'h3a0674d6),
	.w6(32'h3a72d505),
	.w7(32'h3b5ade0f),
	.w8(32'hbb4338c5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f05e5),
	.w1(32'hbc482ada),
	.w2(32'hbc77cc50),
	.w3(32'hbb338378),
	.w4(32'hbc79c09b),
	.w5(32'hbc1d929a),
	.w6(32'hbc840125),
	.w7(32'hbc65dfca),
	.w8(32'hbb538954),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098d25),
	.w1(32'h3c276c1d),
	.w2(32'h3b590859),
	.w3(32'hbb675e61),
	.w4(32'hbb601d3b),
	.w5(32'hbbeeb167),
	.w6(32'h3b68c7ea),
	.w7(32'hbb9ef731),
	.w8(32'hbc30d2d6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cdee4),
	.w1(32'hbbc42434),
	.w2(32'hbba3663b),
	.w3(32'hbc4563b0),
	.w4(32'hbb8ff2a5),
	.w5(32'h3b8d64ac),
	.w6(32'hbb7be037),
	.w7(32'hbb2e87d2),
	.w8(32'hba7c247d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0f256),
	.w1(32'hb9ae72de),
	.w2(32'h3acea1f1),
	.w3(32'hbb2b5ced),
	.w4(32'h3ae9eff0),
	.w5(32'h3c0d4185),
	.w6(32'hbb709ed1),
	.w7(32'h3b5f64b3),
	.w8(32'h3ad52d04),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae34086),
	.w1(32'hbc3a9383),
	.w2(32'hba0597bf),
	.w3(32'hbb2170a3),
	.w4(32'h3b2d04cd),
	.w5(32'hb98479ce),
	.w6(32'hbc09930a),
	.w7(32'h3c0d546c),
	.w8(32'h3af14e76),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1338f9),
	.w1(32'hbb59fe04),
	.w2(32'hba62d4aa),
	.w3(32'hbac7d123),
	.w4(32'hbb1c2b10),
	.w5(32'hbb792ebd),
	.w6(32'hbb95250e),
	.w7(32'hb8b2330f),
	.w8(32'hbb4b27f4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb561e41),
	.w1(32'hbac94a7d),
	.w2(32'hba476365),
	.w3(32'hbc1b6b5f),
	.w4(32'h3b7de6ae),
	.w5(32'h3c0aad07),
	.w6(32'hbb2c6f29),
	.w7(32'h3aa1d5fb),
	.w8(32'h3b7eb872),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2f4d),
	.w1(32'hbb1f37fd),
	.w2(32'h3a945658),
	.w3(32'hba99cc54),
	.w4(32'h3b4e51b5),
	.w5(32'hbb932632),
	.w6(32'hbae57a1b),
	.w7(32'h3a9df7a7),
	.w8(32'hbbfb0052),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e58aa),
	.w1(32'h3c7a6b29),
	.w2(32'h3932698c),
	.w3(32'hbaef1d2b),
	.w4(32'hbb80192e),
	.w5(32'h3aab3c97),
	.w6(32'h3b46f24e),
	.w7(32'hbc3ce793),
	.w8(32'hba75f187),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3b96b),
	.w1(32'hbbb4c37d),
	.w2(32'hbb249a6c),
	.w3(32'hbba8a528),
	.w4(32'hbba0a49f),
	.w5(32'hbb1aa398),
	.w6(32'hbc11c2d8),
	.w7(32'hbb3b1bc4),
	.w8(32'hbb51350e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aede7),
	.w1(32'hbb9707ab),
	.w2(32'hbacc95d2),
	.w3(32'hbbf7eda3),
	.w4(32'hbb138936),
	.w5(32'hbb52d950),
	.w6(32'hbbd99df1),
	.w7(32'hbb955a02),
	.w8(32'hbb9a58c6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1276db),
	.w1(32'hbc099bdd),
	.w2(32'hbbf107e1),
	.w3(32'hbc37bd4e),
	.w4(32'hbc2cd45a),
	.w5(32'h3c431c5d),
	.w6(32'hbc233c6b),
	.w7(32'h3b8160b3),
	.w8(32'hbc39e983),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad4c8),
	.w1(32'hbb2eb3bd),
	.w2(32'h3bd3ad5c),
	.w3(32'hbc335749),
	.w4(32'hbbd99136),
	.w5(32'hbb1ec498),
	.w6(32'hbc2702c3),
	.w7(32'hb976a082),
	.w8(32'h3bb81a4b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909140),
	.w1(32'h3b27e0dd),
	.w2(32'h3c845b7b),
	.w3(32'hbc84cf68),
	.w4(32'h3b7d6142),
	.w5(32'h3bc96bd2),
	.w6(32'hbb0c2085),
	.w7(32'h3c93c005),
	.w8(32'hbb97e15b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9697e),
	.w1(32'hbba6b6ef),
	.w2(32'hba43f771),
	.w3(32'h3b5f2d97),
	.w4(32'h3a3f93ea),
	.w5(32'hbb8af093),
	.w6(32'hbba461ae),
	.w7(32'hba9781ac),
	.w8(32'hbb8338a9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31ee02),
	.w1(32'hb78f235d),
	.w2(32'h39fd40b0),
	.w3(32'hb8dc0472),
	.w4(32'h3a9440e7),
	.w5(32'hbb468288),
	.w6(32'hbb0ad4d2),
	.w7(32'h3b30f7fa),
	.w8(32'h3bc5ea63),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912e5cf),
	.w1(32'hbb40ec03),
	.w2(32'hbb6253ae),
	.w3(32'hbbb6b810),
	.w4(32'h3be592e9),
	.w5(32'hbc2f5110),
	.w6(32'hba48dae1),
	.w7(32'h3c842c90),
	.w8(32'hbbe08223),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71f762),
	.w1(32'hbb4b10e5),
	.w2(32'hbae8de7c),
	.w3(32'hbba5177a),
	.w4(32'hbb81f8c0),
	.w5(32'hbc0d8395),
	.w6(32'hbba1ffbe),
	.w7(32'hbba1f5d7),
	.w8(32'hbb5d7ffd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564d65),
	.w1(32'h3be4c6a5),
	.w2(32'h3b874d48),
	.w3(32'hbb96df68),
	.w4(32'h3c19603e),
	.w5(32'h3b92f99b),
	.w6(32'h3a849f01),
	.w7(32'hbb1d69f9),
	.w8(32'h3a6d1fc7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad72e8),
	.w1(32'h3a8830c9),
	.w2(32'h3b251549),
	.w3(32'h3ba7770f),
	.w4(32'h3a351444),
	.w5(32'hbbda0269),
	.w6(32'hba1901fe),
	.w7(32'hbb90b9e2),
	.w8(32'h39519828),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83508d),
	.w1(32'h3b854b7e),
	.w2(32'h3b48c9c5),
	.w3(32'hbbf0ddcc),
	.w4(32'hbbded020),
	.w5(32'hbaa50fb8),
	.w6(32'hbb78ade7),
	.w7(32'h3ae2469d),
	.w8(32'h3ba27101),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaecdd3),
	.w1(32'hba65a1a7),
	.w2(32'hbc217b27),
	.w3(32'h3c809ffe),
	.w4(32'h394459bc),
	.w5(32'hba8f36b1),
	.w6(32'h3b8da2df),
	.w7(32'hbc3d3f75),
	.w8(32'hbb5f8ade),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb794672),
	.w1(32'hbbdcb2a9),
	.w2(32'h3ab40b32),
	.w3(32'hbb6e2701),
	.w4(32'hbb689e35),
	.w5(32'h3b1ec930),
	.w6(32'hbc0c89ea),
	.w7(32'hbae6d522),
	.w8(32'h3a767e8f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d757),
	.w1(32'h3b8ac612),
	.w2(32'h3b746351),
	.w3(32'hbbb63402),
	.w4(32'hbbc38e51),
	.w5(32'hb994e66e),
	.w6(32'hba3cc51c),
	.w7(32'h3b261f32),
	.w8(32'h3b31ec6c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de36e3),
	.w1(32'hbb93766c),
	.w2(32'hbb7cee17),
	.w3(32'hbb5332db),
	.w4(32'hbbdd3fc0),
	.w5(32'h3c163c1d),
	.w6(32'hbb4555cb),
	.w7(32'hbbb15b94),
	.w8(32'hbbb94be4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2126b),
	.w1(32'h3c593337),
	.w2(32'hbc59c3bb),
	.w3(32'h3be93569),
	.w4(32'hbc3a1ae3),
	.w5(32'hbb63bb5b),
	.w6(32'hbc136973),
	.w7(32'hbcb0f024),
	.w8(32'hbc3334ae),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1a52f),
	.w1(32'h3bebfade),
	.w2(32'h3c4c1296),
	.w3(32'hbb3aa383),
	.w4(32'h3bea881b),
	.w5(32'hb9c28ce3),
	.w6(32'hbc17fee6),
	.w7(32'h3ae635cf),
	.w8(32'hbbf5d2a7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc853fad),
	.w1(32'hbb1dae83),
	.w2(32'hbc02f683),
	.w3(32'hbc837b1d),
	.w4(32'hbb1cb1e5),
	.w5(32'hbc1c6879),
	.w6(32'hbc96e85e),
	.w7(32'hbbb73da8),
	.w8(32'hbb1d391e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78189c),
	.w1(32'hbb6cddac),
	.w2(32'hbaf1e9dd),
	.w3(32'hbb8a0507),
	.w4(32'hbb05f2ee),
	.w5(32'h3a32c898),
	.w6(32'hbb86252c),
	.w7(32'hbbdfe615),
	.w8(32'hbab698a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f0b7c),
	.w1(32'hbafc3876),
	.w2(32'h39335719),
	.w3(32'hbaf6e26f),
	.w4(32'hbb291701),
	.w5(32'h3a6a5864),
	.w6(32'hbc02e641),
	.w7(32'h3ab9621b),
	.w8(32'hbb1fa55a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3499c),
	.w1(32'hb9f92b55),
	.w2(32'hb984fbbe),
	.w3(32'hb9802a1b),
	.w4(32'h3963d236),
	.w5(32'h393f4b00),
	.w6(32'hbb56db7e),
	.w7(32'h39be80e2),
	.w8(32'h3b877059),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b798f46),
	.w1(32'hbab1d161),
	.w2(32'h3b512fb2),
	.w3(32'hba9dad02),
	.w4(32'hb91b3bae),
	.w5(32'hbbb65be6),
	.w6(32'h3ad6465f),
	.w7(32'h3b0c084a),
	.w8(32'h3a8a5aea),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86cea9),
	.w1(32'hbb7c7efb),
	.w2(32'h3a61d954),
	.w3(32'hbb13ba96),
	.w4(32'hbb0197f2),
	.w5(32'hbb52b838),
	.w6(32'hbbcdbe4f),
	.w7(32'h3abf836a),
	.w8(32'hbbe93b7f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5389fc),
	.w1(32'h3b7f277c),
	.w2(32'hba15f456),
	.w3(32'h3b59eb80),
	.w4(32'h3ba0cd0f),
	.w5(32'hbaf99eaf),
	.w6(32'hbb5536bb),
	.w7(32'hbb2d31b0),
	.w8(32'hbb6638a1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b16d),
	.w1(32'h3aa0f2cf),
	.w2(32'h3a0a1ad8),
	.w3(32'hbb1b2427),
	.w4(32'h3908de25),
	.w5(32'h3b0fafb3),
	.w6(32'hbc006c98),
	.w7(32'hbc3af644),
	.w8(32'hbc016a31),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66da25),
	.w1(32'h3a8016ed),
	.w2(32'h3a133bf5),
	.w3(32'h3bf4c88d),
	.w4(32'h3bd173ba),
	.w5(32'hb9e64c20),
	.w6(32'hbbaee6ae),
	.w7(32'hbb13eb70),
	.w8(32'hba6b80a6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd2108),
	.w1(32'hbbf4e2b0),
	.w2(32'hbc134968),
	.w3(32'hbc555919),
	.w4(32'hbc4ad926),
	.w5(32'h3b4dcfd0),
	.w6(32'hbc2c5e0f),
	.w7(32'hbc3f45e1),
	.w8(32'hbb5a6499),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aa56f),
	.w1(32'h3bd7517c),
	.w2(32'h3beaf4bc),
	.w3(32'h3af20d0c),
	.w4(32'h3b677f27),
	.w5(32'hbb3a1353),
	.w6(32'h3bec3028),
	.w7(32'h3ba5fc8e),
	.w8(32'hbb545194),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e43c),
	.w1(32'hba9d8ad6),
	.w2(32'h3a8a05af),
	.w3(32'hbb59a80c),
	.w4(32'hbb053bbc),
	.w5(32'hbc139cbb),
	.w6(32'hbb85191d),
	.w7(32'hb9e10dc1),
	.w8(32'h3b8ea92a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcefe06),
	.w1(32'hbbb336ce),
	.w2(32'hbbdc630b),
	.w3(32'hbc1f716b),
	.w4(32'hbc042141),
	.w5(32'hbb500400),
	.w6(32'h3b7e933b),
	.w7(32'hbbbf48d5),
	.w8(32'h3a2aeef9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8704713),
	.w1(32'h3b7e03fb),
	.w2(32'h3b7adaad),
	.w3(32'hbb82784f),
	.w4(32'hba886f94),
	.w5(32'h3c623458),
	.w6(32'hbb6debdc),
	.w7(32'hbb7a5d5e),
	.w8(32'hbb8a4946),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba204c8),
	.w1(32'hbbda50c3),
	.w2(32'h3b8e2281),
	.w3(32'hbb015cd5),
	.w4(32'hbb22c768),
	.w5(32'hbba8904b),
	.w6(32'hbbdeb6d6),
	.w7(32'h3a354e29),
	.w8(32'hbb9b0645),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4874f1),
	.w1(32'hbc6ff869),
	.w2(32'hbc8eb435),
	.w3(32'hbc029836),
	.w4(32'hbc0bcc8f),
	.w5(32'h3b419ad7),
	.w6(32'hbc5f31ea),
	.w7(32'hbc33fcbc),
	.w8(32'hbc37a9fa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375796),
	.w1(32'h3c0eb3d1),
	.w2(32'hbac39efe),
	.w3(32'h3ac7e337),
	.w4(32'hb99265d4),
	.w5(32'h3ac16e03),
	.w6(32'hbb224604),
	.w7(32'hbc6a19a3),
	.w8(32'h3bd8df64),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af37697),
	.w1(32'h3bbc4b00),
	.w2(32'h3c0e2d50),
	.w3(32'hbaec1e32),
	.w4(32'hbb9160d7),
	.w5(32'h3b1316ee),
	.w6(32'h3b512981),
	.w7(32'h3b84204f),
	.w8(32'h3ba1333c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e05c),
	.w1(32'hbb7765e2),
	.w2(32'h393f3ce1),
	.w3(32'hbb547d40),
	.w4(32'hbbb4dd9f),
	.w5(32'hbbe273ed),
	.w6(32'hb9872ad4),
	.w7(32'hba6b518a),
	.w8(32'hbb9aad02),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce818),
	.w1(32'h3a833f73),
	.w2(32'h3a850420),
	.w3(32'hbb197cfe),
	.w4(32'hbb40d9ac),
	.w5(32'hb9ac0673),
	.w6(32'h3b52be25),
	.w7(32'hba1cc47c),
	.w8(32'hbb49ac12),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1095e5),
	.w1(32'hbac2a6cb),
	.w2(32'h3a035ca7),
	.w3(32'hbb30d11a),
	.w4(32'hbb4d1ed7),
	.w5(32'h39a9a115),
	.w6(32'hbbb225d0),
	.w7(32'h39997bd2),
	.w8(32'h38fe9322),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692507),
	.w1(32'h3b44d396),
	.w2(32'h3c0a0eff),
	.w3(32'hbbcd8eb0),
	.w4(32'hb9e30c5e),
	.w5(32'hbba275f7),
	.w6(32'hbb8047ed),
	.w7(32'h3bfaa03f),
	.w8(32'hbbb6ac44),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e1d3c),
	.w1(32'hbab64671),
	.w2(32'hb9470d78),
	.w3(32'hbbb8a9fa),
	.w4(32'hba5ddc2b),
	.w5(32'h3b02c8de),
	.w6(32'hbbba120d),
	.w7(32'hbabdb797),
	.w8(32'hb9254e39),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b2aa),
	.w1(32'hb9d08aea),
	.w2(32'hbb2b77b7),
	.w3(32'h3b53fcd9),
	.w4(32'h3c744995),
	.w5(32'hbb8751e1),
	.w6(32'hbb2f6707),
	.w7(32'h3c3cabac),
	.w8(32'hbb5eab90),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38444e4b),
	.w1(32'h3b8a7654),
	.w2(32'h3b2ba72f),
	.w3(32'hbc2044ac),
	.w4(32'hbc11e9d4),
	.w5(32'hbb137a1e),
	.w6(32'h391545ff),
	.w7(32'h3ac448b4),
	.w8(32'hbaa68d17),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb787ea6),
	.w1(32'hbb6c7df9),
	.w2(32'hbaef673e),
	.w3(32'hbacedc2a),
	.w4(32'hbb70e247),
	.w5(32'hbbf0e122),
	.w6(32'hbb2b70d0),
	.w7(32'hbb451dc0),
	.w8(32'hbb9e92ad),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f76ee),
	.w1(32'h3b9cf940),
	.w2(32'hbb9c8725),
	.w3(32'hbb28acbb),
	.w4(32'hbafd7aac),
	.w5(32'h3c734329),
	.w6(32'hbb18c1d1),
	.w7(32'hbbd6863d),
	.w8(32'hbbfc98ff),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03dad),
	.w1(32'hbb9a5a6f),
	.w2(32'h3b8046c7),
	.w3(32'h3bde8848),
	.w4(32'h3ae8bc1d),
	.w5(32'h3b23e6da),
	.w6(32'hbbfcc7dc),
	.w7(32'hbbbe03ad),
	.w8(32'hbb054d5b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d7325),
	.w1(32'h3b3f64e2),
	.w2(32'hbbf70da0),
	.w3(32'hbbe2ac6e),
	.w4(32'h3c52c8c8),
	.w5(32'h3b510b5f),
	.w6(32'hbc144540),
	.w7(32'h3c5d76b0),
	.w8(32'h3c89ea79),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020dbf),
	.w1(32'h3b19e6e4),
	.w2(32'h3bd7f752),
	.w3(32'hbb82b837),
	.w4(32'h3b80381a),
	.w5(32'h3c0df49d),
	.w6(32'h3c19d2ef),
	.w7(32'hbb35ae53),
	.w8(32'hbc1728dd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb616112),
	.w1(32'h39c08877),
	.w2(32'hbb958b82),
	.w3(32'h3c6f689d),
	.w4(32'h3be03260),
	.w5(32'hb919c361),
	.w6(32'h3c0c328a),
	.w7(32'hbae40dfe),
	.w8(32'hbb91e952),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00c82),
	.w1(32'h39b48cb8),
	.w2(32'h3a4ed7ae),
	.w3(32'hbc2466b8),
	.w4(32'hbb20fad3),
	.w5(32'h3b2fddb4),
	.w6(32'hbcc892ad),
	.w7(32'hbc0674d2),
	.w8(32'hbc64a255),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb012912),
	.w1(32'hbb85354e),
	.w2(32'h3a7217a0),
	.w3(32'h3b00bdc0),
	.w4(32'h3aa39ac6),
	.w5(32'h3be517ff),
	.w6(32'hbb566ebc),
	.w7(32'h3a819657),
	.w8(32'h3b8e9561),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6bcd),
	.w1(32'hbb18e9b9),
	.w2(32'h39a96637),
	.w3(32'hbb2fb4df),
	.w4(32'hbb2bfdea),
	.w5(32'h3bf8f22c),
	.w6(32'hbb69eafe),
	.w7(32'hbb459c2e),
	.w8(32'hbb81ab26),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125823),
	.w1(32'hbb9167c3),
	.w2(32'h3aea5ce8),
	.w3(32'h3bd80ffe),
	.w4(32'hbb0da3bb),
	.w5(32'hbbf7f26d),
	.w6(32'hbc09e4ca),
	.w7(32'hbbbb8c6a),
	.w8(32'hbb4c9b75),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eb4c1),
	.w1(32'h3b7a255d),
	.w2(32'h37b92d25),
	.w3(32'hbbe5f139),
	.w4(32'hbb4e36d6),
	.w5(32'h3b1b649a),
	.w6(32'hbba512aa),
	.w7(32'hbb7c4e20),
	.w8(32'h3b22e720),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aea2a),
	.w1(32'h3a9ae644),
	.w2(32'h3b547501),
	.w3(32'h3acbb5f3),
	.w4(32'hba148aea),
	.w5(32'hbbf942f1),
	.w6(32'h3b044e65),
	.w7(32'h3b6bd3cb),
	.w8(32'h3b2b800a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617eeb),
	.w1(32'h3c12e8f2),
	.w2(32'h3adc4636),
	.w3(32'hbc47a60e),
	.w4(32'hbc154df4),
	.w5(32'h3b433f8a),
	.w6(32'h3a05c9b7),
	.w7(32'hbafe4d23),
	.w8(32'hbbdf22b4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ab2a7),
	.w1(32'hb9b65052),
	.w2(32'h3c2f3796),
	.w3(32'hbbf23eeb),
	.w4(32'hbb727f17),
	.w5(32'h3be45c51),
	.w6(32'hbc0d9661),
	.w7(32'h399d507f),
	.w8(32'h3bacf83a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb972d3c),
	.w1(32'hba8e63a5),
	.w2(32'h3b0226ad),
	.w3(32'hbafa0c6e),
	.w4(32'h385796e0),
	.w5(32'hbaa26707),
	.w6(32'hbbe2424c),
	.w7(32'hbc0500b2),
	.w8(32'hbb927cb5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf52c9d),
	.w1(32'h38340e50),
	.w2(32'hbb45023e),
	.w3(32'hbb5f7791),
	.w4(32'h3ba48f80),
	.w5(32'h3bdb6207),
	.w6(32'hba974372),
	.w7(32'hbb3cada0),
	.w8(32'h3bf6b792),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86feae),
	.w1(32'hba99e13e),
	.w2(32'hbb9f56ce),
	.w3(32'hbb720f19),
	.w4(32'hbb755a3a),
	.w5(32'hbbe90f5d),
	.w6(32'hbabf9766),
	.w7(32'h3bb951d1),
	.w8(32'h3b89edfd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7531cf),
	.w1(32'h3aeaa8f8),
	.w2(32'h3afaa66e),
	.w3(32'hbb7398b9),
	.w4(32'hbae4010e),
	.w5(32'hbb5aae82),
	.w6(32'hbaed6acd),
	.w7(32'hbaff6a0e),
	.w8(32'hbb103299),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c11bc),
	.w1(32'h3a9694e3),
	.w2(32'hb9c4aebe),
	.w3(32'hbbf9d115),
	.w4(32'hbb8c6aa9),
	.w5(32'h3a3e6167),
	.w6(32'hbb0fdcaf),
	.w7(32'hbb23c179),
	.w8(32'h3ba2e658),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19edbc),
	.w1(32'h3c793ca6),
	.w2(32'h3c1f609a),
	.w3(32'h3c40b6e4),
	.w4(32'h3bacbd4f),
	.w5(32'h3baff449),
	.w6(32'h3c9e3252),
	.w7(32'h3b66bbd2),
	.w8(32'h3a2213f3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e06b),
	.w1(32'h3c033e32),
	.w2(32'hba1c6f0c),
	.w3(32'h3b80ed88),
	.w4(32'h3ab78bb0),
	.w5(32'hbb6a126f),
	.w6(32'h3bb611d2),
	.w7(32'h3b15abda),
	.w8(32'h3b5faf90),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98d17b),
	.w1(32'h3c0fffe8),
	.w2(32'h3bc3a65b),
	.w3(32'h3a1197a5),
	.w4(32'h3a737877),
	.w5(32'h3b8a1313),
	.w6(32'h3c3237ad),
	.w7(32'h3ba4da75),
	.w8(32'h3a9a63b5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e956c),
	.w1(32'h3b4732aa),
	.w2(32'h3beb87b6),
	.w3(32'h3a9275d6),
	.w4(32'h3a2e691f),
	.w5(32'hbbf829f5),
	.w6(32'hbb9840aa),
	.w7(32'hbb278d64),
	.w8(32'hbbc5a760),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa75a4),
	.w1(32'h3b27e48e),
	.w2(32'hbad58a33),
	.w3(32'h3b3873e4),
	.w4(32'h3a935b9f),
	.w5(32'hbbcc0ba8),
	.w6(32'hb9805c5f),
	.w7(32'hbc089992),
	.w8(32'hbb430222),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7351b),
	.w1(32'h3bb8525f),
	.w2(32'h3ba059f6),
	.w3(32'hbba5c6f8),
	.w4(32'hbb3c841a),
	.w5(32'hbae18392),
	.w6(32'h3ba57f63),
	.w7(32'hbb121341),
	.w8(32'h3a8f2139),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a0a3),
	.w1(32'h3b3af255),
	.w2(32'h3bbf3517),
	.w3(32'hbb29197c),
	.w4(32'hba17aa63),
	.w5(32'h3b79a6af),
	.w6(32'h3ac24b75),
	.w7(32'h3a9c0f25),
	.w8(32'h3b0f9859),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd6a0),
	.w1(32'h3903badf),
	.w2(32'hbc293422),
	.w3(32'hbb8754ce),
	.w4(32'h3b157e57),
	.w5(32'h3a71fa28),
	.w6(32'h3a8f146c),
	.w7(32'hbb0c5ed3),
	.w8(32'hbbcef902),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229e8e),
	.w1(32'h3b407377),
	.w2(32'hbb8759d4),
	.w3(32'hbb8aecc8),
	.w4(32'hbb928054),
	.w5(32'hbc1cf8b2),
	.w6(32'hbb039a88),
	.w7(32'hbadcc0b4),
	.w8(32'hba44759d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34a72d),
	.w1(32'h3bc87e8d),
	.w2(32'hbc564c2d),
	.w3(32'h39dafd34),
	.w4(32'hbc225c5f),
	.w5(32'hbc4aa406),
	.w6(32'hbbea2207),
	.w7(32'hbbcdbba3),
	.w8(32'h3b5d7f10),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09b71f),
	.w1(32'hbb8c477a),
	.w2(32'hbbefad6e),
	.w3(32'hbc783a25),
	.w4(32'hbc47947e),
	.w5(32'hbbbd26c4),
	.w6(32'hbc3b415d),
	.w7(32'hbb9b79a0),
	.w8(32'h3903a398),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8493c4),
	.w1(32'hbc03b19b),
	.w2(32'hbb35185a),
	.w3(32'hbc19fc5d),
	.w4(32'h3b4f7ce6),
	.w5(32'h3c358ca9),
	.w6(32'h3b32a084),
	.w7(32'h3c50e196),
	.w8(32'h3b7b87f1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44b790),
	.w1(32'hbbc35e1c),
	.w2(32'hb9fb391d),
	.w3(32'h3b3feeeb),
	.w4(32'hb939e9cd),
	.w5(32'hbb0a2965),
	.w6(32'hbbeea275),
	.w7(32'hb8dc4936),
	.w8(32'h3bb77af2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2032ec),
	.w1(32'h3b0e62e8),
	.w2(32'h3bd08dc4),
	.w3(32'hbb17c795),
	.w4(32'h3b35eb93),
	.w5(32'hba863fad),
	.w6(32'hbbe9bbfc),
	.w7(32'hbba2f3b2),
	.w8(32'hbb06ea38),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba1b7),
	.w1(32'h3a33c32a),
	.w2(32'hbb2c9402),
	.w3(32'hbba09e3c),
	.w4(32'hbb40388e),
	.w5(32'hba919f4e),
	.w6(32'hba862ef8),
	.w7(32'hbbc103a9),
	.w8(32'hbb7ec1ca),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bfab2),
	.w1(32'hbc1b6d35),
	.w2(32'hbb476850),
	.w3(32'hbca1468a),
	.w4(32'hbc106d4f),
	.w5(32'h3b39af9a),
	.w6(32'hbc6cc54b),
	.w7(32'hbbc5bf98),
	.w8(32'hbb134eda),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c341c48),
	.w1(32'hba0a9e30),
	.w2(32'hbc6f9919),
	.w3(32'hbaebcd01),
	.w4(32'hbbcb834a),
	.w5(32'hbc5ef587),
	.w6(32'hbc7472c9),
	.w7(32'hbbdb969a),
	.w8(32'hba7f60e8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd08d9),
	.w1(32'h3b7ea8eb),
	.w2(32'h3ae1d931),
	.w3(32'h3c640442),
	.w4(32'hbb9f0893),
	.w5(32'h3c842d54),
	.w6(32'h3c3975ed),
	.w7(32'hb975e0f0),
	.w8(32'hbc4bdd68),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adad4a4),
	.w1(32'h3bb4f2da),
	.w2(32'h3b7a07e4),
	.w3(32'h3c4852d8),
	.w4(32'h3b116f77),
	.w5(32'h3b28490a),
	.w6(32'hbc3e63f0),
	.w7(32'hba8fe485),
	.w8(32'h3aa404b2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64e1d),
	.w1(32'h3bb88a75),
	.w2(32'h3c4a7fd9),
	.w3(32'hbc9ae0a8),
	.w4(32'hbc91215e),
	.w5(32'h3b652c82),
	.w6(32'hbae069dd),
	.w7(32'hbc9b17e1),
	.w8(32'h3c019367),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464f50),
	.w1(32'h3a8bceff),
	.w2(32'hbc8e3634),
	.w3(32'h3c5a688a),
	.w4(32'hbc366b3a),
	.w5(32'hbc0a0760),
	.w6(32'h3a9ff89f),
	.w7(32'hbc5d3b0f),
	.w8(32'hbc37a09a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cd21f),
	.w1(32'hbb8d5ae7),
	.w2(32'hb9fed969),
	.w3(32'hbabe3bd7),
	.w4(32'hbc0d0a4d),
	.w5(32'hb9e1f47c),
	.w6(32'hbbb415b0),
	.w7(32'hbbe505f9),
	.w8(32'h3b85cbc8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccc05e),
	.w1(32'h3c672d37),
	.w2(32'h3b346bff),
	.w3(32'h3cb1a865),
	.w4(32'h3b6e12a3),
	.w5(32'h3be68d53),
	.w6(32'h3b86722f),
	.w7(32'hbbe85f6b),
	.w8(32'hba89d992),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c347),
	.w1(32'hbc53000f),
	.w2(32'h3b0e3160),
	.w3(32'h3c29b827),
	.w4(32'hbb901223),
	.w5(32'hbc8c395d),
	.w6(32'hbb9b682f),
	.w7(32'hbb478f01),
	.w8(32'hba6de706),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85402c),
	.w1(32'h3915c22e),
	.w2(32'hbaadfccb),
	.w3(32'h3aaed0ac),
	.w4(32'h3b5d712d),
	.w5(32'hb9bd79b1),
	.w6(32'h3cf36b4b),
	.w7(32'h3c03b733),
	.w8(32'h3a822574),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b908036),
	.w1(32'hbb6f58d5),
	.w2(32'hbb8191bf),
	.w3(32'h3b8e08a7),
	.w4(32'hbbae2c99),
	.w5(32'h3b940a22),
	.w6(32'h3ab0b372),
	.w7(32'hbc07bc74),
	.w8(32'h3b96d97e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1156b),
	.w1(32'hbbe8a84a),
	.w2(32'hbba12394),
	.w3(32'hbb92f980),
	.w4(32'hbb53f752),
	.w5(32'h3b0b968e),
	.w6(32'hbbdc5390),
	.w7(32'hbbeddc5d),
	.w8(32'hbb68c582),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5eea),
	.w1(32'hbc03a639),
	.w2(32'hbba7c0ec),
	.w3(32'h36ea0f5b),
	.w4(32'h3a466da9),
	.w5(32'hbb544be8),
	.w6(32'hbbc70f9c),
	.w7(32'hbbf9b224),
	.w8(32'hbb82ab0f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2791ce),
	.w1(32'hbaf6fb52),
	.w2(32'hbb2b8b65),
	.w3(32'hbad3ceaa),
	.w4(32'hb9039121),
	.w5(32'hbc357941),
	.w6(32'hbb971237),
	.w7(32'h3b809bf0),
	.w8(32'hbb733900),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01ca25),
	.w1(32'h3b79c904),
	.w2(32'hba79fc91),
	.w3(32'hbbdc3819),
	.w4(32'hbc503f8a),
	.w5(32'hbbc8c0e1),
	.w6(32'hbc5376f7),
	.w7(32'hbc83a98d),
	.w8(32'hbac0fd24),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0d35),
	.w1(32'h3bd38811),
	.w2(32'h3bc5228a),
	.w3(32'hbb8f6cb8),
	.w4(32'h3b60c052),
	.w5(32'h3b1f9d6f),
	.w6(32'h3b73a740),
	.w7(32'h3b21ff9c),
	.w8(32'h3c36db6f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164619),
	.w1(32'h3c08a072),
	.w2(32'h3c54a935),
	.w3(32'hbc2677f4),
	.w4(32'h3b8d3d94),
	.w5(32'h3c3ee297),
	.w6(32'hb988d8dc),
	.w7(32'h3cb5cb41),
	.w8(32'h3c67d816),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02bba1),
	.w1(32'h3ab037e0),
	.w2(32'h3bd70340),
	.w3(32'hb675b946),
	.w4(32'hbc21b829),
	.w5(32'h3c8352fb),
	.w6(32'hbb741d17),
	.w7(32'hbbf22e06),
	.w8(32'hbac4db76),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0e30),
	.w1(32'h3c09bd5d),
	.w2(32'h3c72f108),
	.w3(32'h3b6ce2fa),
	.w4(32'hbc4c8203),
	.w5(32'h39f49d98),
	.w6(32'hbce4d627),
	.w7(32'hbc704a83),
	.w8(32'hbb096a13),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae17157),
	.w1(32'hbb90974c),
	.w2(32'hbab5f05a),
	.w3(32'hbb3d497e),
	.w4(32'hbb6d3057),
	.w5(32'h39cd58d1),
	.w6(32'hbbe11747),
	.w7(32'hbbc2bdd8),
	.w8(32'hbb1d87bc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9858cf6),
	.w1(32'hbaed9f78),
	.w2(32'hbc04c91c),
	.w3(32'hbb056a5d),
	.w4(32'hbbd420d4),
	.w5(32'h39f692a5),
	.w6(32'h3bc393d5),
	.w7(32'hbbea5b24),
	.w8(32'h3c67030b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d40ca),
	.w1(32'hb990cfc3),
	.w2(32'hbb4022ed),
	.w3(32'h3b96cc8d),
	.w4(32'h3aaaccd3),
	.w5(32'hbb2c8c57),
	.w6(32'h3c93fc7c),
	.w7(32'h3c05f419),
	.w8(32'h39960d32),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24a2b3),
	.w1(32'h3c78b882),
	.w2(32'h3b73320c),
	.w3(32'hbb23b268),
	.w4(32'hbb611658),
	.w5(32'hbb65435f),
	.w6(32'h3a66796d),
	.w7(32'hbbd3a064),
	.w8(32'hbc2825df),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb477c50),
	.w1(32'hbbb664b1),
	.w2(32'hbc689c48),
	.w3(32'hbc3f0a07),
	.w4(32'hbb368451),
	.w5(32'hbc11f88a),
	.w6(32'h3c7dd001),
	.w7(32'hbb3e59db),
	.w8(32'hbaf8e9c2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afe03),
	.w1(32'hbc0305f4),
	.w2(32'hbc4482a6),
	.w3(32'hbbed8246),
	.w4(32'hbc0d6c21),
	.w5(32'hbba8fcea),
	.w6(32'hbc482b00),
	.w7(32'hbc09243f),
	.w8(32'h3ba4c26b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f7719),
	.w1(32'hbb21a232),
	.w2(32'hb9c4bb07),
	.w3(32'h38bb0644),
	.w4(32'h3c13325f),
	.w5(32'hbc1e6af9),
	.w6(32'h3c9c7bc5),
	.w7(32'hbb355afc),
	.w8(32'hbb2bf1ba),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19a230),
	.w1(32'hbbd45a3c),
	.w2(32'hbbd670e7),
	.w3(32'hbbfec951),
	.w4(32'hbb7de24c),
	.w5(32'hbae868ba),
	.w6(32'hbaa671a6),
	.w7(32'h38673da7),
	.w8(32'h3ba33a79),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9944d76),
	.w1(32'h3bb1ac3e),
	.w2(32'hbaa192af),
	.w3(32'hbb9de308),
	.w4(32'hbba9f90e),
	.w5(32'h3b843422),
	.w6(32'h3c16833d),
	.w7(32'h3a5db766),
	.w8(32'h3c07a7c2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8465c9),
	.w1(32'hbc00cd8f),
	.w2(32'hbc3dc374),
	.w3(32'h3b53e1e1),
	.w4(32'hbb46aa18),
	.w5(32'hbbabacb4),
	.w6(32'h3c4529b9),
	.w7(32'hbc07ab9a),
	.w8(32'h399c184b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00b0ec),
	.w1(32'hbb3ada78),
	.w2(32'hbb1ad841),
	.w3(32'hbb845d69),
	.w4(32'hbb433329),
	.w5(32'hbb8e5279),
	.w6(32'hbacd38ae),
	.w7(32'hba6f9800),
	.w8(32'h3c14b85e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b622b4),
	.w1(32'h3c08f1d9),
	.w2(32'h3ae80192),
	.w3(32'hbc5f8566),
	.w4(32'hbc65be5c),
	.w5(32'h3bdc0fa3),
	.w6(32'hbbf235f8),
	.w7(32'hbbe69dc2),
	.w8(32'hbc45a3d2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46336e),
	.w1(32'h3a1edf9b),
	.w2(32'hbb6bd432),
	.w3(32'hbbd4a286),
	.w4(32'hbba33be6),
	.w5(32'h3baf6c4a),
	.w6(32'hbbae8fea),
	.w7(32'hbbd0c73b),
	.w8(32'h3aa97f82),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be2e6),
	.w1(32'h3b68923e),
	.w2(32'h3a818577),
	.w3(32'hba9d5763),
	.w4(32'hbbb0358e),
	.w5(32'h3c0748c1),
	.w6(32'hbb956472),
	.w7(32'hbb1ea978),
	.w8(32'hbbe37be0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde5073),
	.w1(32'hbb54c8ba),
	.w2(32'h3c2d0b7a),
	.w3(32'h3bd62afa),
	.w4(32'h3bb42a26),
	.w5(32'hb981d22c),
	.w6(32'hbc4b6530),
	.w7(32'hbc47edb1),
	.w8(32'hbb8a87e1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9376d3),
	.w1(32'hbb7683c6),
	.w2(32'hbaeb9a00),
	.w3(32'hbbb5dfbf),
	.w4(32'hbbab153a),
	.w5(32'hbbec6672),
	.w6(32'hbaf8c108),
	.w7(32'hbb71ae10),
	.w8(32'h3c1129fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba77a7),
	.w1(32'hb9a10977),
	.w2(32'h3af91055),
	.w3(32'hbbf70cb4),
	.w4(32'h3c027824),
	.w5(32'h3b2fd4f2),
	.w6(32'h3c8ffea1),
	.w7(32'h3c031c72),
	.w8(32'h3abd4336),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2b3e),
	.w1(32'hbb9b28db),
	.w2(32'hba8953db),
	.w3(32'h3a542818),
	.w4(32'h3bc4ce2d),
	.w5(32'h3b1b45c0),
	.w6(32'h3af62425),
	.w7(32'h3bb76d98),
	.w8(32'h39a22a5b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc15de),
	.w1(32'hbb55137e),
	.w2(32'hbc012b45),
	.w3(32'hbb759838),
	.w4(32'hbb08f27e),
	.w5(32'hba870462),
	.w6(32'hbb3feaa4),
	.w7(32'hbb580ba5),
	.w8(32'hbc35d72c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa36562),
	.w1(32'hb98ad989),
	.w2(32'h3af8fdd7),
	.w3(32'hbb18603e),
	.w4(32'hbaa1dbde),
	.w5(32'h3a5940f7),
	.w6(32'hbc37ca1e),
	.w7(32'hbc22cc1d),
	.w8(32'h3b810f21),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaddfe),
	.w1(32'h3b250eb5),
	.w2(32'h3ae7021a),
	.w3(32'hbb3b3bac),
	.w4(32'hba98fe55),
	.w5(32'hba7e8e7b),
	.w6(32'hbb186cb4),
	.w7(32'h3b56f5cc),
	.w8(32'h3b1546ea),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0695ef),
	.w1(32'hbc33b0cc),
	.w2(32'hbc30354c),
	.w3(32'hbacbd2c6),
	.w4(32'hbbf8a2a6),
	.w5(32'hb9d4bbe4),
	.w6(32'hbac11665),
	.w7(32'hbb667525),
	.w8(32'hb842ff2b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b358e),
	.w1(32'h3ae368c1),
	.w2(32'h3b934feb),
	.w3(32'h3bfe32f5),
	.w4(32'h3a133f27),
	.w5(32'hbc17b6ba),
	.w6(32'h3ca1c9cf),
	.w7(32'hb91753ee),
	.w8(32'hbc474615),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c625bd4),
	.w1(32'h3c3dc20e),
	.w2(32'h3bbd5a1c),
	.w3(32'hbc7ac392),
	.w4(32'hbb9d46a3),
	.w5(32'h3bac2811),
	.w6(32'h3c976310),
	.w7(32'h3c4d9c2d),
	.w8(32'h3a54785e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b042bc),
	.w1(32'hbb87b741),
	.w2(32'h3b9ed43c),
	.w3(32'h3b98c933),
	.w4(32'hba8c35dc),
	.w5(32'hbc1284b3),
	.w6(32'hbab8aeef),
	.w7(32'hbb447e59),
	.w8(32'hbc52029e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd5e85f),
	.w1(32'h3b904341),
	.w2(32'hbac2fd3d),
	.w3(32'hbc8d1207),
	.w4(32'h3bbb8f0a),
	.w5(32'h3b658c15),
	.w6(32'hbc10f273),
	.w7(32'hbc1508e2),
	.w8(32'h3ae77654),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b393fa),
	.w1(32'hb9964062),
	.w2(32'hb98c3e01),
	.w3(32'h3bd2bd2c),
	.w4(32'h3b27ad0e),
	.w5(32'hbc1387b0),
	.w6(32'hbb4eb8c8),
	.w7(32'h3a14ae35),
	.w8(32'hbba2c1ae),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb768b82),
	.w1(32'h3b87d790),
	.w2(32'h3ab831e2),
	.w3(32'hbb8b43f3),
	.w4(32'h3b01e365),
	.w5(32'hbbcfe21f),
	.w6(32'h3ad74585),
	.w7(32'hba77f216),
	.w8(32'hbb9684ba),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa215c7),
	.w1(32'hbb00593b),
	.w2(32'h3b62a984),
	.w3(32'hbbc92455),
	.w4(32'hbb1de302),
	.w5(32'h3af4ca52),
	.w6(32'hba07f9ba),
	.w7(32'h3b156312),
	.w8(32'h39c184f3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152ff6),
	.w1(32'hbbb077e9),
	.w2(32'hbab1f02f),
	.w3(32'h3bce91db),
	.w4(32'h3b396621),
	.w5(32'hbb3f1277),
	.w6(32'hba145ed9),
	.w7(32'hbab14812),
	.w8(32'h3b4ebf8f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3ecff),
	.w1(32'hbbb97cbb),
	.w2(32'h3a4664ce),
	.w3(32'hb9ae8c48),
	.w4(32'hba54a2df),
	.w5(32'h3c493ad8),
	.w6(32'h3bdff58b),
	.w7(32'hbab4bba2),
	.w8(32'h3aeda169),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074f89),
	.w1(32'h3c2cdec9),
	.w2(32'h3cb0c54b),
	.w3(32'h3c979b3f),
	.w4(32'hbb240c5e),
	.w5(32'hbc01b60c),
	.w6(32'h3c0c0bd6),
	.w7(32'h3a884281),
	.w8(32'hbc059dba),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a4873),
	.w1(32'hbbf0fd25),
	.w2(32'h3aae0e06),
	.w3(32'hb9f07f4f),
	.w4(32'hb9131e40),
	.w5(32'hbaca1b93),
	.w6(32'hba86010e),
	.w7(32'h3821f425),
	.w8(32'hbbb92a49),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd5a72),
	.w1(32'hbae2cd27),
	.w2(32'hbac0f524),
	.w3(32'hbc40f83a),
	.w4(32'hbbd32f42),
	.w5(32'hbc3478ea),
	.w6(32'hbc96a94e),
	.w7(32'hbbf6a306),
	.w8(32'h3bfde2a7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33cf27),
	.w1(32'h3c191be4),
	.w2(32'h3bad75fb),
	.w3(32'h388e9cdd),
	.w4(32'hbbea22f1),
	.w5(32'hbbcd62e5),
	.w6(32'h3c298b2e),
	.w7(32'h3bba95c4),
	.w8(32'h3a2e814c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f046),
	.w1(32'h3b4b3718),
	.w2(32'hbbbc37bb),
	.w3(32'hbbad2312),
	.w4(32'hbc68c4e5),
	.w5(32'h3ccc0ee2),
	.w6(32'hbb270426),
	.w7(32'hbc76e176),
	.w8(32'hbc911cdb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f4000),
	.w1(32'h3cf804b3),
	.w2(32'h3cef0bac),
	.w3(32'h3ca3d461),
	.w4(32'h3cfa721c),
	.w5(32'hbb880dfd),
	.w6(32'hbd26e8c6),
	.w7(32'hbccf1f86),
	.w8(32'hbba7b034),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a818a),
	.w1(32'hbbcc6e43),
	.w2(32'h38b0c3e3),
	.w3(32'h3b3f18ce),
	.w4(32'h3b05eebc),
	.w5(32'h3bf919d0),
	.w6(32'hbaf69ae4),
	.w7(32'h3b6d3522),
	.w8(32'hbade137d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b872c9e),
	.w1(32'hbb14e6eb),
	.w2(32'hb9d11e56),
	.w3(32'h3b8b03a1),
	.w4(32'h3b81c970),
	.w5(32'h37027e7c),
	.w6(32'hbb873d75),
	.w7(32'h39f83ea2),
	.w8(32'h3a2a0457),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ad85),
	.w1(32'hb993d9fc),
	.w2(32'hbb84489f),
	.w3(32'h3b0f499f),
	.w4(32'h3b4e8a34),
	.w5(32'hbc68a37a),
	.w6(32'h39d36247),
	.w7(32'hbb2d2eda),
	.w8(32'hbc87a3fa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc116569),
	.w1(32'hbae75ab4),
	.w2(32'hbc958e91),
	.w3(32'hbc7a34ed),
	.w4(32'h3a0033ad),
	.w5(32'hbc880ebf),
	.w6(32'hbc8a3ed7),
	.w7(32'hbca97904),
	.w8(32'hbbc00e30),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf9fd),
	.w1(32'hbba1749a),
	.w2(32'h3a4bdf10),
	.w3(32'hbc764726),
	.w4(32'hbc0df4f7),
	.w5(32'h3bb48b58),
	.w6(32'hbbd7542a),
	.w7(32'h3aa2eb79),
	.w8(32'h3c328042),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993aac8),
	.w1(32'hbbf7ddd4),
	.w2(32'hbbd025a0),
	.w3(32'h3c07099a),
	.w4(32'h3b9f3ab1),
	.w5(32'hbbd19c79),
	.w6(32'h3c8a166b),
	.w7(32'h3bb708a1),
	.w8(32'h3bec55fc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49450f),
	.w1(32'h3c735e67),
	.w2(32'h3ba28f60),
	.w3(32'hbb8c9e4e),
	.w4(32'hbbe626e3),
	.w5(32'h3bc6ce46),
	.w6(32'h3bdd23d8),
	.w7(32'hbbce54a1),
	.w8(32'h3a93eec9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd6c8),
	.w1(32'h3a74aac1),
	.w2(32'hbb9b8ab9),
	.w3(32'hbc10dfe2),
	.w4(32'hbc0187e4),
	.w5(32'hbbb9e8be),
	.w6(32'hbc64bc5f),
	.w7(32'hbb901d80),
	.w8(32'hbb9574e8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba669e59),
	.w1(32'hba8197f4),
	.w2(32'hbc0fe679),
	.w3(32'hbb0c13b1),
	.w4(32'h3ae26732),
	.w5(32'hbc6ab25f),
	.w6(32'hbbb05c75),
	.w7(32'hbc325dcf),
	.w8(32'hbc80ea90),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5a7e3),
	.w1(32'hbc04aa92),
	.w2(32'hba2fa347),
	.w3(32'hbb9d3f29),
	.w4(32'h3c43bf1c),
	.w5(32'h3c403456),
	.w6(32'hbc9293e0),
	.w7(32'hbc6558a0),
	.w8(32'hbbdff1d6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833cb5),
	.w1(32'h3b2e59a7),
	.w2(32'h3c07ea93),
	.w3(32'h3c4b3f07),
	.w4(32'h39830db4),
	.w5(32'hbc0c3087),
	.w6(32'hbbf8e9e9),
	.w7(32'h39a0c630),
	.w8(32'hbbb4ac50),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06656c),
	.w1(32'h3b6591bc),
	.w2(32'hbb480ab4),
	.w3(32'hbba65289),
	.w4(32'hba9724eb),
	.w5(32'h3b24b422),
	.w6(32'hbc3989ac),
	.w7(32'hbc013170),
	.w8(32'h3b9d6aad),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e2037),
	.w1(32'hbbb7a495),
	.w2(32'hba98448c),
	.w3(32'h3a2fe9c0),
	.w4(32'h3bb602c3),
	.w5(32'hbc47dd35),
	.w6(32'h3a5fee9f),
	.w7(32'h3bb9d28b),
	.w8(32'hbb5300a1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2d92),
	.w1(32'hbac6ef02),
	.w2(32'hbbf9aa1a),
	.w3(32'hbc237972),
	.w4(32'hbc0dc899),
	.w5(32'h39daf3d9),
	.w6(32'h3b192f32),
	.w7(32'hbbfa602a),
	.w8(32'hbc76a8ba),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8252af),
	.w1(32'h3abe0c47),
	.w2(32'hbb795d3d),
	.w3(32'hbaa92870),
	.w4(32'hbb2af802),
	.w5(32'hb9ec08cb),
	.w6(32'hbc421469),
	.w7(32'hbb55150a),
	.w8(32'hbc073ba0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39552),
	.w1(32'h3ca04a84),
	.w2(32'h3bd415cd),
	.w3(32'h3c14d771),
	.w4(32'h3c94af3b),
	.w5(32'h3b2457fa),
	.w6(32'h3c859e91),
	.w7(32'h3c3ebd87),
	.w8(32'hbbb9f37f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af7e5),
	.w1(32'hbb2d8f09),
	.w2(32'h3b0b752a),
	.w3(32'h3aff3b67),
	.w4(32'hbb3aa926),
	.w5(32'h3b730b08),
	.w6(32'hbbb170b4),
	.w7(32'h38c3f3a7),
	.w8(32'h3b956ed8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e5414),
	.w1(32'h3babd431),
	.w2(32'h3c18a051),
	.w3(32'h3b89ef08),
	.w4(32'h3bb94ecc),
	.w5(32'hbb15e72d),
	.w6(32'h39c68cfb),
	.w7(32'h3bb9c642),
	.w8(32'h3b81ce24),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987b44c),
	.w1(32'h3b78ab02),
	.w2(32'hbb58b6ac),
	.w3(32'hbb8dea7f),
	.w4(32'hbb308fc7),
	.w5(32'h3b993991),
	.w6(32'h3c1abe6a),
	.w7(32'hbb55d2e8),
	.w8(32'hbbc0390c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b921),
	.w1(32'h39ebd274),
	.w2(32'hbbd2bf81),
	.w3(32'h3c30d57b),
	.w4(32'h39b966b4),
	.w5(32'hbbc60016),
	.w6(32'hbbacd486),
	.w7(32'hbbd8bec1),
	.w8(32'hbc5d460d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd41d08),
	.w1(32'hbc114e2f),
	.w2(32'hb968028b),
	.w3(32'hbbcdbef4),
	.w4(32'hbb3da1f4),
	.w5(32'h3addca91),
	.w6(32'hbc4de119),
	.w7(32'hbbeec1ef),
	.w8(32'hbbf98859),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4e83),
	.w1(32'hb97f9b63),
	.w2(32'h3a87f831),
	.w3(32'hba3defff),
	.w4(32'hbaae8334),
	.w5(32'hbbaca507),
	.w6(32'hbbaad8ff),
	.w7(32'hbc0241dc),
	.w8(32'h3b3a6c3b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eacee),
	.w1(32'h3c376f73),
	.w2(32'h3c2bfd7d),
	.w3(32'hbc5a118e),
	.w4(32'hbbaa5cd3),
	.w5(32'h3ab6dea2),
	.w6(32'hbadcabea),
	.w7(32'h3b213399),
	.w8(32'h3b29dd8d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1aeac),
	.w1(32'h3bbc22b5),
	.w2(32'h3c0237b2),
	.w3(32'hb9a6bdd3),
	.w4(32'h3ab1a289),
	.w5(32'hbbcc2256),
	.w6(32'hbb6d3737),
	.w7(32'h3c0b3b57),
	.w8(32'hbb66c4fb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a956a92),
	.w1(32'hba6305c9),
	.w2(32'hb98efa00),
	.w3(32'hbc4998bd),
	.w4(32'hbc03d505),
	.w5(32'h3b800ac0),
	.w6(32'hbc42cfa6),
	.w7(32'hbbbb8af1),
	.w8(32'h3b2ad062),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf330f),
	.w1(32'h3bfd11ae),
	.w2(32'h3b3be2ed),
	.w3(32'hbc0e112e),
	.w4(32'hbbbcd7f8),
	.w5(32'hba7a4572),
	.w6(32'h3c7f871b),
	.w7(32'h3bd432ac),
	.w8(32'h3bdf49fd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbf423),
	.w1(32'hbbb720ed),
	.w2(32'h3bf0e530),
	.w3(32'hbb5f4b26),
	.w4(32'hbb01b504),
	.w5(32'hbc5bf911),
	.w6(32'h3c962197),
	.w7(32'h3c40aa15),
	.w8(32'hbbe46003),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f51b),
	.w1(32'h3b3e9e23),
	.w2(32'hbbcef0ba),
	.w3(32'hbbf918b6),
	.w4(32'h3b1ec302),
	.w5(32'hbc53b22e),
	.w6(32'h3cf16f42),
	.w7(32'h3beb8d30),
	.w8(32'hbc3665e4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dbaf1),
	.w1(32'h3b9dd3d3),
	.w2(32'hb9a57950),
	.w3(32'hbc31eecf),
	.w4(32'hbbf38adb),
	.w5(32'h3cb702f4),
	.w6(32'hbbf2ee39),
	.w7(32'h3aecb2c8),
	.w8(32'h3c8ab9b6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc918),
	.w1(32'h3c9712f9),
	.w2(32'h3cbca1d3),
	.w3(32'h3cc049bc),
	.w4(32'h39a127a1),
	.w5(32'hbbd9732f),
	.w6(32'h3ca2f583),
	.w7(32'h3c6fe264),
	.w8(32'hbc68be57),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49ad8d),
	.w1(32'hbbc1b592),
	.w2(32'hbc4793e6),
	.w3(32'h3bb901a0),
	.w4(32'h3c45075e),
	.w5(32'hba898e8b),
	.w6(32'hbc9fb12d),
	.w7(32'hbc59b621),
	.w8(32'hbc187ee9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e7301),
	.w1(32'h3c451701),
	.w2(32'h3b5c2086),
	.w3(32'h3c4783f1),
	.w4(32'h3baf16f3),
	.w5(32'h3a91b887),
	.w6(32'hbc4065ad),
	.w7(32'hbbd47c8b),
	.w8(32'hbc71bbd4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a312539),
	.w1(32'h3bfc2cf4),
	.w2(32'hbb10a469),
	.w3(32'h3c58210f),
	.w4(32'hbc00406c),
	.w5(32'hbc2dfb5f),
	.w6(32'h3be47287),
	.w7(32'hbc19a9c1),
	.w8(32'hbc0fe245),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08729e),
	.w1(32'h3b6fd1ea),
	.w2(32'h3b740b6d),
	.w3(32'hbc40c034),
	.w4(32'hbbb9b49f),
	.w5(32'h3c4f96c1),
	.w6(32'hbbcbb3cf),
	.w7(32'hbaee7166),
	.w8(32'h3b6033f6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dff3d),
	.w1(32'hbbc84e89),
	.w2(32'h3b6e5309),
	.w3(32'hbc63d344),
	.w4(32'h3be33c4b),
	.w5(32'h3ad94506),
	.w6(32'hbc0f4f93),
	.w7(32'hbc02a0a3),
	.w8(32'hbaa6112b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51246e),
	.w1(32'h3aa27bcc),
	.w2(32'hbbd3f91a),
	.w3(32'hbb53adea),
	.w4(32'h3c23a987),
	.w5(32'hbc01a1fe),
	.w6(32'hbbc7db38),
	.w7(32'h3aa1e929),
	.w8(32'hbc458c54),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38259fb4),
	.w1(32'hbb476635),
	.w2(32'hbbda21ce),
	.w3(32'hbb2cc6be),
	.w4(32'hbb58f5b9),
	.w5(32'hbc1866df),
	.w6(32'hbbf6b01b),
	.w7(32'hbb82e8e9),
	.w8(32'h3c1acdbb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec84f0),
	.w1(32'hbc24cbf6),
	.w2(32'hbbe65812),
	.w3(32'hbb8fbba4),
	.w4(32'h3a331529),
	.w5(32'hbc11a4aa),
	.w6(32'h3d11826c),
	.w7(32'h3bbe6ced),
	.w8(32'hbc1cc622),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6181),
	.w1(32'h3c79ec30),
	.w2(32'h3b374d74),
	.w3(32'h3b111421),
	.w4(32'h3b8df502),
	.w5(32'hbc127b5d),
	.w6(32'hbb8aab9a),
	.w7(32'h3aebf1c7),
	.w8(32'hbc125764),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196034),
	.w1(32'hbbb01743),
	.w2(32'hbc3c4003),
	.w3(32'hbadcd76e),
	.w4(32'hbc220ce9),
	.w5(32'h3c4414bd),
	.w6(32'h3b5bf726),
	.w7(32'hbae42225),
	.w8(32'h3cf5e0b0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6c54),
	.w1(32'h3c22336c),
	.w2(32'h3c1cc42d),
	.w3(32'hbab59026),
	.w4(32'h3b783e7f),
	.w5(32'hbb868a2e),
	.w6(32'h3cafbb2f),
	.w7(32'h3cdc986e),
	.w8(32'hbb9ab021),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb027e27),
	.w1(32'hbb453f78),
	.w2(32'h3a228c2b),
	.w3(32'hb931d152),
	.w4(32'hbaee919a),
	.w5(32'h3ba69755),
	.w6(32'hbb8d12eb),
	.w7(32'hbb8234c7),
	.w8(32'h3c106055),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a395e02),
	.w1(32'h3c1422b3),
	.w2(32'h3c9eacc0),
	.w3(32'hb98babe3),
	.w4(32'h3a7b2fb4),
	.w5(32'h3a8201ee),
	.w6(32'hbbeeff53),
	.w7(32'h3aa64390),
	.w8(32'h3ae9c4fc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c23b4),
	.w1(32'h3c691e51),
	.w2(32'h3c199294),
	.w3(32'hbc282680),
	.w4(32'hbc3a925d),
	.w5(32'hbbacf584),
	.w6(32'h3b121dce),
	.w7(32'hbbaae5f3),
	.w8(32'hbb84b359),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9264a),
	.w1(32'hbc716f58),
	.w2(32'hbc09d5a1),
	.w3(32'hbb97bf34),
	.w4(32'hbc46df5a),
	.w5(32'hba9934a8),
	.w6(32'hbd032513),
	.w7(32'hbc57828d),
	.w8(32'hbb609294),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9b6c4),
	.w1(32'h3bbed179),
	.w2(32'h3ba6a27f),
	.w3(32'h3b89d150),
	.w4(32'hba8e6d52),
	.w5(32'hbbca9a55),
	.w6(32'hbbfd21d9),
	.w7(32'h3aac40a2),
	.w8(32'hbc5c52f0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeec396),
	.w1(32'hbaf463f5),
	.w2(32'h3a9dcfac),
	.w3(32'h3a8c378c),
	.w4(32'hb90ed1e5),
	.w5(32'hbbf97e76),
	.w6(32'hbaa01078),
	.w7(32'hbb806149),
	.w8(32'h3b4f35a7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f49ef),
	.w1(32'hb9c8071b),
	.w2(32'h3bb37850),
	.w3(32'hbbba6d2f),
	.w4(32'hbb30ab30),
	.w5(32'hba55dc7e),
	.w6(32'h3be1a403),
	.w7(32'hba253986),
	.w8(32'hb99c1c4a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02ffe8),
	.w1(32'hbaeab572),
	.w2(32'h3b1a10c6),
	.w3(32'h3ad000a9),
	.w4(32'h3b5fc603),
	.w5(32'h3ad15188),
	.w6(32'hbc03c7fd),
	.w7(32'h3b8ba630),
	.w8(32'h3a8c6bec),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937dabb),
	.w1(32'hba05bae7),
	.w2(32'hbae27c4e),
	.w3(32'h3b0979ea),
	.w4(32'h3a887f17),
	.w5(32'hbc31808d),
	.w6(32'hb908593a),
	.w7(32'hbbbe3428),
	.w8(32'hbbcd3a2b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba66b3),
	.w1(32'h3ba2d5ec),
	.w2(32'h3c3efb6a),
	.w3(32'h3a3c80a9),
	.w4(32'h3b3a74b1),
	.w5(32'h3bfd1948),
	.w6(32'h3af465cb),
	.w7(32'h3b5a689b),
	.w8(32'h3cb7d7eb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255e53),
	.w1(32'h3c7f0f3e),
	.w2(32'h3c2c7b0e),
	.w3(32'h3c9733d3),
	.w4(32'h3c7da57a),
	.w5(32'hbc03d84c),
	.w6(32'h3c9da2cc),
	.w7(32'h3cbe3798),
	.w8(32'hbbb114e2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc135aa),
	.w1(32'hbb401f98),
	.w2(32'hba4f48f8),
	.w3(32'h3b193895),
	.w4(32'hbb249f75),
	.w5(32'h3a58c97a),
	.w6(32'h3c1338d9),
	.w7(32'h3a48164d),
	.w8(32'hbb7143e6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2867a),
	.w1(32'h38df664f),
	.w2(32'h3c0e1702),
	.w3(32'h3bb9fc63),
	.w4(32'h3bd40f5e),
	.w5(32'hbb19d4ab),
	.w6(32'hbc633035),
	.w7(32'hba973bd2),
	.w8(32'hbbba3d96),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd90af),
	.w1(32'h3a97bb73),
	.w2(32'hba5601b9),
	.w3(32'hb9283c78),
	.w4(32'hba0812dc),
	.w5(32'h3ab56afc),
	.w6(32'hbb95353a),
	.w7(32'h3afb59e3),
	.w8(32'hbb593cd3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b513b0a),
	.w1(32'hba29a878),
	.w2(32'h3b65d286),
	.w3(32'hbba1dafb),
	.w4(32'hbbf4678e),
	.w5(32'hba8b25eb),
	.w6(32'hbc963870),
	.w7(32'hbc0cbe05),
	.w8(32'hbac20542),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5dbd2),
	.w1(32'h3b21baa8),
	.w2(32'h3bad7b75),
	.w3(32'h3bc17650),
	.w4(32'hba9a7e9e),
	.w5(32'hbbc2b9ad),
	.w6(32'hbb31c182),
	.w7(32'h3ae783c5),
	.w8(32'hba994662),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d057),
	.w1(32'hbc1b30bd),
	.w2(32'hbc06a242),
	.w3(32'h3b1f102e),
	.w4(32'hbbb1fa08),
	.w5(32'hbbd52ea0),
	.w6(32'h3bdcd780),
	.w7(32'hbb876eba),
	.w8(32'h3b855732),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab098ad),
	.w1(32'hbbf06aea),
	.w2(32'hbb444136),
	.w3(32'h38abdc84),
	.w4(32'h3af5f784),
	.w5(32'hbc15a8d1),
	.w6(32'hba470f07),
	.w7(32'hbc3097df),
	.w8(32'hbc074492),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2af57c),
	.w1(32'hbc1c12e3),
	.w2(32'hba849c9b),
	.w3(32'hbc43343f),
	.w4(32'hbc4ee435),
	.w5(32'h3b5d543a),
	.w6(32'h3bbd9de6),
	.w7(32'hbb82633b),
	.w8(32'hb8d15d62),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379eaf90),
	.w1(32'h3bf410d5),
	.w2(32'h3b871d9b),
	.w3(32'h3b9cf48c),
	.w4(32'h3b57dffd),
	.w5(32'h3baf0c10),
	.w6(32'hbaeb85c3),
	.w7(32'hbc10d7d1),
	.w8(32'hbc446090),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc545e7),
	.w1(32'hbb9d1c1d),
	.w2(32'hbaa9be9d),
	.w3(32'hbbd26c1b),
	.w4(32'hbc39802b),
	.w5(32'h3c662ba4),
	.w6(32'hbc9fb6c5),
	.w7(32'h3acf8997),
	.w8(32'h3d19567e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fae22),
	.w1(32'h3af50288),
	.w2(32'h3c03c4eb),
	.w3(32'h3c2676d2),
	.w4(32'h3bd022d4),
	.w5(32'h3b2503f7),
	.w6(32'h3ca45079),
	.w7(32'h3cdf4c58),
	.w8(32'h3a20bb1f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb343a87),
	.w1(32'hbafa75f5),
	.w2(32'h3891b416),
	.w3(32'h3aebad24),
	.w4(32'h3b4f555f),
	.w5(32'hba09e1c8),
	.w6(32'hb9358962),
	.w7(32'h3b0932a9),
	.w8(32'h3b629c8e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc10c1),
	.w1(32'hbb1a1620),
	.w2(32'hbcae08b3),
	.w3(32'h3bd9b3fd),
	.w4(32'hbc6a2d03),
	.w5(32'hba3fff2d),
	.w6(32'h3bca0ff3),
	.w7(32'hbaa4a052),
	.w8(32'hbbde148e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a4c3b),
	.w1(32'h3ae63611),
	.w2(32'hbc04f61c),
	.w3(32'hbc349bb9),
	.w4(32'hbba7deee),
	.w5(32'hbb886540),
	.w6(32'hbc0ca5b4),
	.w7(32'hbbe19e90),
	.w8(32'h3b59b27d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010144),
	.w1(32'h3af1d96d),
	.w2(32'hbbf018da),
	.w3(32'h3a1b4bd3),
	.w4(32'hbc15c85e),
	.w5(32'hbc07eb7e),
	.w6(32'hbbbdfd58),
	.w7(32'hbc320af9),
	.w8(32'hbc51dda9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7716b),
	.w1(32'h3af6482c),
	.w2(32'hbc1d85ea),
	.w3(32'hbc5440e0),
	.w4(32'hbb8e38e5),
	.w5(32'h3bb6d39c),
	.w6(32'hbbcc2904),
	.w7(32'hbabbb64a),
	.w8(32'h3b08c176),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc357c2),
	.w1(32'h3b193b88),
	.w2(32'h3bf7e56b),
	.w3(32'h3bb6458b),
	.w4(32'h3c17fc7d),
	.w5(32'h3a7b1001),
	.w6(32'h3b96b287),
	.w7(32'h3af3f545),
	.w8(32'hbb9202fe),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1198ca),
	.w1(32'hbba0127b),
	.w2(32'hbb9bc80f),
	.w3(32'h3a230de7),
	.w4(32'h3a127ba6),
	.w5(32'hbc1b25e4),
	.w6(32'hbb48eb37),
	.w7(32'hbb7cd82c),
	.w8(32'h3bd10cc0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a94b),
	.w1(32'hbaa00b33),
	.w2(32'h3b196b41),
	.w3(32'hbbff4a74),
	.w4(32'hbb5a545c),
	.w5(32'hbaa433b9),
	.w6(32'h3c76d92f),
	.w7(32'h3b856812),
	.w8(32'hbc21b095),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f5159),
	.w1(32'h3b40b023),
	.w2(32'h3b978058),
	.w3(32'hbafe0016),
	.w4(32'hbb0e8d70),
	.w5(32'h3bfa227c),
	.w6(32'hbc83098c),
	.w7(32'h37ed280e),
	.w8(32'h3c9659f8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e26a4d),
	.w1(32'hbbd8baad),
	.w2(32'hbc6524f1),
	.w3(32'h3d1b28fb),
	.w4(32'h3c77d322),
	.w5(32'hb5546614),
	.w6(32'h3c8afb9a),
	.w7(32'hbbc069fa),
	.w8(32'hb6ed1724),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f5bad),
	.w1(32'hbb58c4cf),
	.w2(32'hbae9a651),
	.w3(32'hbae1a74c),
	.w4(32'hbb3de9b8),
	.w5(32'h3a2797f6),
	.w6(32'hba9c0566),
	.w7(32'hbadb1da3),
	.w8(32'h38adda17),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93c65d),
	.w1(32'hbb2194c7),
	.w2(32'h3aeaa121),
	.w3(32'hbbf35e29),
	.w4(32'hbae01886),
	.w5(32'h3b947965),
	.w6(32'hbaae443a),
	.w7(32'h3a13ecfc),
	.w8(32'hbb235aa2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7203dc0),
	.w1(32'hba192a52),
	.w2(32'h39c07061),
	.w3(32'hba92683f),
	.w4(32'hba95447a),
	.w5(32'h3881397e),
	.w6(32'hbada800d),
	.w7(32'hbb284acb),
	.w8(32'hbb2c0bad),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3844d511),
	.w1(32'h37b40744),
	.w2(32'h37db20d1),
	.w3(32'h38b7e664),
	.w4(32'h38864e98),
	.w5(32'h357749ac),
	.w6(32'hb76b0485),
	.w7(32'hb81eba51),
	.w8(32'hb80da8c6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c18d),
	.w1(32'hbaccc4b5),
	.w2(32'hbbff7445),
	.w3(32'hbbbb9d12),
	.w4(32'hbc073e3a),
	.w5(32'h3b629e8d),
	.w6(32'hbac21b71),
	.w7(32'hbc494a2f),
	.w8(32'hbb85db33),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64b609),
	.w1(32'hbab5f62b),
	.w2(32'hbb36dd39),
	.w3(32'hbb26ae30),
	.w4(32'hbaaaf8fa),
	.w5(32'h3a25f57b),
	.w6(32'hbb1d9a2b),
	.w7(32'hbac1ec95),
	.w8(32'hba01f9c1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391484f6),
	.w1(32'h35425588),
	.w2(32'h379ddf04),
	.w3(32'h3909c0b2),
	.w4(32'h361ebcc3),
	.w5(32'h38e2c51a),
	.w6(32'h38d2dbef),
	.w7(32'h38ddd4be),
	.w8(32'h39457b21),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31a674),
	.w1(32'hba2b1403),
	.w2(32'hbb3fdd43),
	.w3(32'hbb17ec4a),
	.w4(32'hba1b407f),
	.w5(32'h3a37f24e),
	.w6(32'hbab9c3cb),
	.w7(32'h37361b46),
	.w8(32'hba4bba41),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38921125),
	.w1(32'h3811e38d),
	.w2(32'hb93a5b74),
	.w3(32'h37cdef0a),
	.w4(32'hb70f0096),
	.w5(32'hb92823bb),
	.w6(32'hb7e0ae50),
	.w7(32'hb82318ba),
	.w8(32'hb9244e4e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dbbd4),
	.w1(32'hba464f81),
	.w2(32'hba093441),
	.w3(32'hba6d9fa2),
	.w4(32'hba20d172),
	.w5(32'hb96a7c42),
	.w6(32'hb9825d15),
	.w7(32'hb9d040cf),
	.w8(32'hb987d809),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b12bfe),
	.w1(32'h38539aff),
	.w2(32'h383106bd),
	.w3(32'h38112fd1),
	.w4(32'h3802f710),
	.w5(32'hb70b6b6b),
	.w6(32'h37b57135),
	.w7(32'hb7676e0c),
	.w8(32'hb842ece5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bcf634),
	.w1(32'h384d0662),
	.w2(32'h37d455a0),
	.w3(32'hb8717abb),
	.w4(32'h37a8e18a),
	.w5(32'h3895e0c7),
	.w6(32'hb8c252ea),
	.w7(32'hb8bbe5ff),
	.w8(32'hb89bd6b6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4d9af),
	.w1(32'hbb133a2a),
	.w2(32'hbb0c1dac),
	.w3(32'hb99c34a1),
	.w4(32'hbaad8d59),
	.w5(32'hbae794d5),
	.w6(32'hba63af21),
	.w7(32'hbab8b72a),
	.w8(32'hbacd63f8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45b9fa),
	.w1(32'hbb561bc2),
	.w2(32'hbbefb042),
	.w3(32'hbbb970a1),
	.w4(32'hbb734e9c),
	.w5(32'hbb93f63a),
	.w6(32'hbc1eadb8),
	.w7(32'hba92e72a),
	.w8(32'hba159ce4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00f666),
	.w1(32'hbb2ea210),
	.w2(32'hbb30a201),
	.w3(32'hbb1efa71),
	.w4(32'hb9a33d66),
	.w5(32'h3ad9a9ec),
	.w6(32'hbb162fe9),
	.w7(32'hbac844f9),
	.w8(32'hb98cce20),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4eb37),
	.w1(32'hbb389d69),
	.w2(32'hbbccf7e1),
	.w3(32'hbb537b80),
	.w4(32'hbb0b3917),
	.w5(32'hbb64a335),
	.w6(32'hbb9fa9b9),
	.w7(32'hb9d3acd3),
	.w8(32'hbaa66785),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a98cd7),
	.w1(32'hb9a95917),
	.w2(32'hb9502e80),
	.w3(32'hb9511971),
	.w4(32'hb9887cc1),
	.w5(32'hb9528626),
	.w6(32'hb984e5b7),
	.w7(32'hb9662175),
	.w8(32'hb9555591),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba544531),
	.w1(32'hba070fde),
	.w2(32'h3972aa36),
	.w3(32'hb9697e95),
	.w4(32'h396ff4e9),
	.w5(32'h39a6c66a),
	.w6(32'h37977c2c),
	.w7(32'hb988f372),
	.w8(32'hb9433001),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842b774),
	.w1(32'h3888693c),
	.w2(32'h3807b78c),
	.w3(32'h37e4abee),
	.w4(32'h385667f4),
	.w5(32'h3837481c),
	.w6(32'h38397b87),
	.w7(32'h38299445),
	.w8(32'h3809d966),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb727eae9),
	.w1(32'h38148f1d),
	.w2(32'h37e5ce4b),
	.w3(32'hb83dcc1e),
	.w4(32'hb800e82c),
	.w5(32'hb8192ffe),
	.w6(32'hb897994d),
	.w7(32'hb86a44de),
	.w8(32'hb8371710),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd85df),
	.w1(32'hbab83382),
	.w2(32'hbaa6371c),
	.w3(32'hbb8512a9),
	.w4(32'h3bcbb70c),
	.w5(32'h3b8852c9),
	.w6(32'hbb4c5f9f),
	.w7(32'h3b2c150b),
	.w8(32'h3a71ceec),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38270e7a),
	.w1(32'h38470c76),
	.w2(32'h385cacb6),
	.w3(32'hb8aa3692),
	.w4(32'h37c1a4d3),
	.w5(32'h38502137),
	.w6(32'h38da22d7),
	.w7(32'h38eddb27),
	.w8(32'h3993357d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955d582),
	.w1(32'hb9f8bf38),
	.w2(32'hba21e1b9),
	.w3(32'h39127d68),
	.w4(32'hb919cfde),
	.w5(32'hb90812fa),
	.w6(32'h3a609359),
	.w7(32'h3a374db8),
	.w8(32'h3a2576dc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a129c22),
	.w1(32'h3a4add15),
	.w2(32'h3b42714d),
	.w3(32'h3aea1941),
	.w4(32'h3b76486f),
	.w5(32'h3b334441),
	.w6(32'h3a44efa0),
	.w7(32'h3b32f0e4),
	.w8(32'hb9197f75),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81be870),
	.w1(32'hb8158403),
	.w2(32'hb839ed17),
	.w3(32'h3893aa04),
	.w4(32'hb7c9eeea),
	.w5(32'hb8113076),
	.w6(32'h3894715b),
	.w7(32'hb89122db),
	.w8(32'h37a09842),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a64156),
	.w1(32'hbac37c1e),
	.w2(32'hbad4ca19),
	.w3(32'hbb0a434c),
	.w4(32'hbae3bfd4),
	.w5(32'hba6c5b21),
	.w6(32'hbb0f515d),
	.w7(32'hbb10bc80),
	.w8(32'hbaceb4e2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10d9a4),
	.w1(32'h39a30f9c),
	.w2(32'h39f02d76),
	.w3(32'hba1894ac),
	.w4(32'h38c04a84),
	.w5(32'h3a576a58),
	.w6(32'hb9a7cbdd),
	.w7(32'hb81cb149),
	.w8(32'h3a36dcd0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97c37c),
	.w1(32'hba9cf286),
	.w2(32'hbab2a5b1),
	.w3(32'hbb9f28b9),
	.w4(32'h3c6b1cd1),
	.w5(32'h3bbc397b),
	.w6(32'hbb44c3a4),
	.w7(32'h3c81a9d7),
	.w8(32'h3bca02ce),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8862153),
	.w1(32'hb93faf34),
	.w2(32'hb922b675),
	.w3(32'hb7004821),
	.w4(32'hb6562346),
	.w5(32'h35b6a89e),
	.w6(32'hb91c4d3c),
	.w7(32'hb9140f9e),
	.w8(32'hb7673f0c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d68c1),
	.w1(32'h3b2ac44b),
	.w2(32'h3b6f8b53),
	.w3(32'h3b53eb3f),
	.w4(32'h3a0d2071),
	.w5(32'hbadded92),
	.w6(32'h3b154de4),
	.w7(32'hbadd33d1),
	.w8(32'hbbd10703),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule