module layer_10_featuremap_190(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977eeca),
	.w1(32'hba8dd73a),
	.w2(32'hbaa3fcd6),
	.w3(32'hb965299a),
	.w4(32'h3866d1ae),
	.w5(32'hba8dca1d),
	.w6(32'hbaf4554c),
	.w7(32'hbac33567),
	.w8(32'hb91263e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda8fb),
	.w1(32'h386a460c),
	.w2(32'hba267d8f),
	.w3(32'hba9fe4ae),
	.w4(32'h3a79bae0),
	.w5(32'h38a3d98d),
	.w6(32'h38661698),
	.w7(32'h3a985506),
	.w8(32'hb76c2cc0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919617d),
	.w1(32'hb8317089),
	.w2(32'h395610e9),
	.w3(32'hb9226112),
	.w4(32'hb6a3f908),
	.w5(32'h3960cd0c),
	.w6(32'h38ef2f70),
	.w7(32'h3854b3b9),
	.w8(32'hb7da62f5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84e02b1),
	.w1(32'h39e85b01),
	.w2(32'hba32a772),
	.w3(32'hb95c75b8),
	.w4(32'hba251d2a),
	.w5(32'hba41ac5d),
	.w6(32'hb89dfa64),
	.w7(32'hba23d0d1),
	.w8(32'hba1290b4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26c0f8),
	.w1(32'h3926590a),
	.w2(32'h396132a9),
	.w3(32'hba48c9a1),
	.w4(32'hb94a825b),
	.w5(32'hb9311061),
	.w6(32'h37530231),
	.w7(32'h3a3acc80),
	.w8(32'h39f7ca85),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8f1b),
	.w1(32'hb942ef2f),
	.w2(32'hb9737ba7),
	.w3(32'hb73d4639),
	.w4(32'hb98f01ef),
	.w5(32'hb9e352d7),
	.w6(32'hb99f8290),
	.w7(32'hb9e81fe9),
	.w8(32'hb9edf47f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e115b4),
	.w1(32'hbab91447),
	.w2(32'hbb82d1e8),
	.w3(32'hba4588cf),
	.w4(32'hbb06915d),
	.w5(32'hbb6badd2),
	.w6(32'h3a925aca),
	.w7(32'hbaa6d1d3),
	.w8(32'hbb222611),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa951b6),
	.w1(32'hbb5bfddf),
	.w2(32'hbb5d6dc5),
	.w3(32'hbac7155e),
	.w4(32'hbb447c44),
	.w5(32'hbb464fb4),
	.w6(32'hbad28c94),
	.w7(32'hbb07ae4e),
	.w8(32'hbb901d23),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bb7f7),
	.w1(32'hba5769db),
	.w2(32'hbaa43f3d),
	.w3(32'h37c40d3b),
	.w4(32'hbaadcce6),
	.w5(32'hbab27ff2),
	.w6(32'h3900bbe1),
	.w7(32'hba01c02f),
	.w8(32'hba738182),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7d617),
	.w1(32'hb81a3faa),
	.w2(32'hbbb425c9),
	.w3(32'h3b24f239),
	.w4(32'h3b119d07),
	.w5(32'hbb8e7147),
	.w6(32'h3a89b0fc),
	.w7(32'h3a56fcbe),
	.w8(32'hbbaf9c41),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a7c53),
	.w1(32'hb983f317),
	.w2(32'hb9c026fe),
	.w3(32'h3a0b6299),
	.w4(32'h39d3f0e3),
	.w5(32'h3a565022),
	.w6(32'hb9fa093f),
	.w7(32'hba0535b4),
	.w8(32'hb9878001),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19bea5),
	.w1(32'h3b410c54),
	.w2(32'hbb4a7a3a),
	.w3(32'h3a495ad3),
	.w4(32'h378797ae),
	.w5(32'hbb56db7d),
	.w6(32'h39120442),
	.w7(32'hb826423f),
	.w8(32'hbb503cf2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9c68),
	.w1(32'h3a9f86aa),
	.w2(32'hbb912acc),
	.w3(32'h3b4f30dd),
	.w4(32'h3ac863bc),
	.w5(32'hbb8b1b0f),
	.w6(32'h3b49ffd3),
	.w7(32'h3a5c1d1e),
	.w8(32'hbbd607cd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3da7d8),
	.w1(32'hba8381b8),
	.w2(32'hbae91804),
	.w3(32'h3a0a7129),
	.w4(32'hba353d14),
	.w5(32'hba180db7),
	.w6(32'h3ad47b91),
	.w7(32'h398eb5ec),
	.w8(32'hba374d41),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f19ef),
	.w1(32'hba51c41c),
	.w2(32'hbb33cf64),
	.w3(32'h3b2c07fe),
	.w4(32'h3a9f0f07),
	.w5(32'hbac1b9e2),
	.w6(32'hbae12310),
	.w7(32'h382da00b),
	.w8(32'hbb38c331),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab627ab),
	.w1(32'hbb255427),
	.w2(32'hbbbcdeb3),
	.w3(32'hb8915477),
	.w4(32'hbaaa22fc),
	.w5(32'hbb8e6719),
	.w6(32'h3918ee01),
	.w7(32'hbad0220d),
	.w8(32'hbbbd8340),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba651491),
	.w1(32'hba6e6522),
	.w2(32'hb810fcb1),
	.w3(32'hba79b7c2),
	.w4(32'hbaaba10e),
	.w5(32'hb7938936),
	.w6(32'hbaa379f8),
	.w7(32'hba8c8c05),
	.w8(32'hba93f6c5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001996),
	.w1(32'hba506c24),
	.w2(32'hbb9ee57b),
	.w3(32'hb6c16f12),
	.w4(32'hb79a4397),
	.w5(32'hbb6d363e),
	.w6(32'hb9a6346d),
	.w7(32'hbb1552c0),
	.w8(32'hbbb7062c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae96ce8),
	.w1(32'hba217620),
	.w2(32'hbb8404c4),
	.w3(32'h3aa70ba1),
	.w4(32'hba2fb2d1),
	.w5(32'hbb49c3cf),
	.w6(32'h3a0b3577),
	.w7(32'hba07a0ad),
	.w8(32'hbb776fa2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d91caa),
	.w1(32'hb93e5f32),
	.w2(32'hb92c367a),
	.w3(32'hb86bc564),
	.w4(32'hb88e7ef7),
	.w5(32'h384b313b),
	.w6(32'hb8f5b23b),
	.w7(32'hb86a3665),
	.w8(32'hb91a0db3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae95c5),
	.w1(32'hb8a5d885),
	.w2(32'hb9abfb7e),
	.w3(32'hb9577cda),
	.w4(32'h3a070c9c),
	.w5(32'h39f554f6),
	.w6(32'h391693ba),
	.w7(32'hb904c089),
	.w8(32'hb938ca51),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf5eed),
	.w1(32'hba9e82aa),
	.w2(32'hba5bacde),
	.w3(32'h3a832ce0),
	.w4(32'h3a7babff),
	.w5(32'h3a131054),
	.w6(32'hba49c2b1),
	.w7(32'h3a10e14d),
	.w8(32'hb863a801),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba750e93),
	.w1(32'hbb261dfc),
	.w2(32'hbc3fdba9),
	.w3(32'h3ad03850),
	.w4(32'h3abc9301),
	.w5(32'hbc08dc06),
	.w6(32'hba9ec650),
	.w7(32'hb9c018f2),
	.w8(32'hbc34938d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c75b5),
	.w1(32'h3a47a86a),
	.w2(32'hbb70e70f),
	.w3(32'h39fbad49),
	.w4(32'h3b337077),
	.w5(32'hbb3fd9c7),
	.w6(32'h3a02817b),
	.w7(32'h3a2d660f),
	.w8(32'hbba999ad),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f16999),
	.w1(32'h3aa72175),
	.w2(32'hbb248367),
	.w3(32'h3b036da3),
	.w4(32'h3b513d70),
	.w5(32'hba7d5daa),
	.w6(32'hbac6c075),
	.w7(32'hb99fe362),
	.w8(32'hbb7e2d42),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96cff0),
	.w1(32'hba3ce6a3),
	.w2(32'hba209dbd),
	.w3(32'hb9d3a0f4),
	.w4(32'hba96d953),
	.w5(32'hba3ab303),
	.w6(32'hba43c64f),
	.w7(32'hba565d78),
	.w8(32'hbab6bcb2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ac7fb),
	.w1(32'hb93a6056),
	.w2(32'h38222ecf),
	.w3(32'hba256eb3),
	.w4(32'hb84ed218),
	.w5(32'h399d8e5f),
	.w6(32'hb980eb18),
	.w7(32'hb776a5b9),
	.w8(32'h38406de1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7ad37),
	.w1(32'hbaccb857),
	.w2(32'hba302a3f),
	.w3(32'h3acb1416),
	.w4(32'hba4b08ae),
	.w5(32'h3a4dda6c),
	.w6(32'h3913bf9a),
	.w7(32'hbad072f3),
	.w8(32'hba6de868),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd32a5),
	.w1(32'h3b08c6da),
	.w2(32'h3a6730fc),
	.w3(32'h3aca178f),
	.w4(32'h3afb3cac),
	.w5(32'h3ae72b11),
	.w6(32'h36d1d910),
	.w7(32'h38094fea),
	.w8(32'h3a67bd17),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9e963),
	.w1(32'hb98a42a1),
	.w2(32'hbb11236e),
	.w3(32'h3a98a8a0),
	.w4(32'h39b72dc0),
	.w5(32'hbb008cda),
	.w6(32'hba884948),
	.w7(32'hbac719d5),
	.w8(32'hbb8431a5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e51db0),
	.w1(32'hb93d016c),
	.w2(32'hb99fb1d6),
	.w3(32'h37a6ab87),
	.w4(32'h3950f787),
	.w5(32'h3906ea97),
	.w6(32'hb8c1a830),
	.w7(32'hb9630212),
	.w8(32'hb9844da5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cffa23),
	.w1(32'h38363d62),
	.w2(32'h39a9aa4d),
	.w3(32'hb89e5329),
	.w4(32'hb80f6d3a),
	.w5(32'h398c298d),
	.w6(32'hb8c2f1d0),
	.w7(32'hb8bc9267),
	.w8(32'hb85587e8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ed08b),
	.w1(32'hbab3775a),
	.w2(32'hbb2be5eb),
	.w3(32'h3a0c44ca),
	.w4(32'hba4004f9),
	.w5(32'hbb253578),
	.w6(32'hba89cebf),
	.w7(32'hb9e0f822),
	.w8(32'hbb63c8e1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8c92),
	.w1(32'hb996bc85),
	.w2(32'hbab4c2ca),
	.w3(32'hba0de564),
	.w4(32'hb9ad5864),
	.w5(32'hba94def1),
	.w6(32'hbae869be),
	.w7(32'hb9fb1cc0),
	.w8(32'hbb0c3063),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ea929),
	.w1(32'hb89885c2),
	.w2(32'hb92f62eb),
	.w3(32'hba8032ba),
	.w4(32'h39a964e2),
	.w5(32'hb8a76f62),
	.w6(32'h39a7c639),
	.w7(32'h393cdc02),
	.w8(32'h37e09186),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b5181),
	.w1(32'hb9b273df),
	.w2(32'hbaec726b),
	.w3(32'h3a003440),
	.w4(32'hb9b3725a),
	.w5(32'hbaae42c0),
	.w6(32'h3980bf2a),
	.w7(32'hba24fe9d),
	.w8(32'hbade3f16),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61d37a),
	.w1(32'h3bb886b2),
	.w2(32'hbb91312b),
	.w3(32'h3ad44984),
	.w4(32'h3be47e96),
	.w5(32'hbad105dd),
	.w6(32'h3b0558c7),
	.w7(32'h3bdbafa0),
	.w8(32'hbab9875b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb757a),
	.w1(32'h3bcffcd3),
	.w2(32'h3af12a99),
	.w3(32'h3ad1b725),
	.w4(32'h3bdfbdfa),
	.w5(32'h3bb3091b),
	.w6(32'hbb3f0a24),
	.w7(32'h3b596f3d),
	.w8(32'h3b4e5351),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad722eb),
	.w1(32'h3af7af28),
	.w2(32'h3ab62de3),
	.w3(32'h3b5cdfdc),
	.w4(32'h3b8beee7),
	.w5(32'h3b90fdd3),
	.w6(32'hb9804c88),
	.w7(32'h39907554),
	.w8(32'h3abebedb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9726ca),
	.w1(32'hb8dbd6f7),
	.w2(32'h37e85387),
	.w3(32'hba751b44),
	.w4(32'h39de3e09),
	.w5(32'h3a38dd74),
	.w6(32'hbabe23f5),
	.w7(32'hb966fd5b),
	.w8(32'h385dd150),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97638ef),
	.w1(32'hba4c03ef),
	.w2(32'hba7f600d),
	.w3(32'hb97a35e6),
	.w4(32'hb9a7eead),
	.w5(32'hb9f638d1),
	.w6(32'hba25b9d6),
	.w7(32'hba17b0c3),
	.w8(32'hb9956c03),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e83f7),
	.w1(32'h3880be53),
	.w2(32'h38e9459a),
	.w3(32'hb9700514),
	.w4(32'h35bd2f5a),
	.w5(32'h39ef1568),
	.w6(32'hb9b0dd0e),
	.w7(32'hb986eeed),
	.w8(32'hb9120cd5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a928cc2),
	.w1(32'h3b610fd5),
	.w2(32'hb9dcc458),
	.w3(32'h3af51693),
	.w4(32'h3b6db132),
	.w5(32'h39d3c548),
	.w6(32'h3af7aca4),
	.w7(32'h3b804336),
	.w8(32'h3a088629),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29fbe),
	.w1(32'hba895d43),
	.w2(32'hbbcdd886),
	.w3(32'h39c5ead5),
	.w4(32'hb912ad00),
	.w5(32'hbb9343ef),
	.w6(32'h3a8d5285),
	.w7(32'hba13e74b),
	.w8(32'hbb99358c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce982f),
	.w1(32'h3a237fb2),
	.w2(32'hbb2c7d6f),
	.w3(32'h3b207ac6),
	.w4(32'h3b62d792),
	.w5(32'hba99a081),
	.w6(32'h3a1f5492),
	.w7(32'h3b10d116),
	.w8(32'hbb3a2536),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf4572),
	.w1(32'h3a2447a4),
	.w2(32'hbb81714a),
	.w3(32'h3b5edd69),
	.w4(32'h3b8693c9),
	.w5(32'hbb10e216),
	.w6(32'hba33af12),
	.w7(32'h3a58643f),
	.w8(32'hbbb9ed9e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a8924),
	.w1(32'hbb4d130d),
	.w2(32'hbbce06d8),
	.w3(32'hba93a31a),
	.w4(32'hbaa74f18),
	.w5(32'hbb90a6b7),
	.w6(32'hbaf747cb),
	.w7(32'hb9f3e249),
	.w8(32'hbb8219c5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b9a2c),
	.w1(32'hbb09785c),
	.w2(32'hbc1aea70),
	.w3(32'hbab568df),
	.w4(32'hbb49faf5),
	.w5(32'hbbf6e4ef),
	.w6(32'hba009a99),
	.w7(32'hbb20a53f),
	.w8(32'hbbe6740c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39887da9),
	.w1(32'h3a234118),
	.w2(32'h38f7c51f),
	.w3(32'hb7ae5aec),
	.w4(32'h39cc205a),
	.w5(32'h3822a39e),
	.w6(32'h3a1b6f75),
	.w7(32'h3a6719d9),
	.w8(32'h399039aa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9982d8e),
	.w1(32'hb994a2cf),
	.w2(32'hba968087),
	.w3(32'hb8acc3fa),
	.w4(32'hb9961c48),
	.w5(32'hbac54210),
	.w6(32'h3a01a137),
	.w7(32'hb8fcf2e8),
	.w8(32'hba5f519a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45682f),
	.w1(32'h3adcdd76),
	.w2(32'h3a8ce7da),
	.w3(32'h3a53f57f),
	.w4(32'h3ab7aacc),
	.w5(32'h3a7cb98e),
	.w6(32'h3ac1b4da),
	.w7(32'h3a45a675),
	.w8(32'h3a64f604),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a697e05),
	.w1(32'hba171199),
	.w2(32'hbb712640),
	.w3(32'h3b309bab),
	.w4(32'hb90198f4),
	.w5(32'hbb2aba32),
	.w6(32'h39df74a3),
	.w7(32'hb840514e),
	.w8(32'hbb5ae9f9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2ccc3),
	.w1(32'hba5c4439),
	.w2(32'hbb0ca464),
	.w3(32'hba0ff4d7),
	.w4(32'hb9e9686f),
	.w5(32'hbad6ebd8),
	.w6(32'hb9e711a4),
	.w7(32'hba9565bc),
	.w8(32'hbafa9c37),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46c32e),
	.w1(32'hbb3e1b8f),
	.w2(32'hbbe10012),
	.w3(32'hb8929329),
	.w4(32'hbb296b27),
	.w5(32'hbbc40770),
	.w6(32'hba1c8c31),
	.w7(32'hbaa5fe1e),
	.w8(32'hbbcdf6b3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02061a),
	.w1(32'hb9f53450),
	.w2(32'hba1632d3),
	.w3(32'h38af7480),
	.w4(32'hb9ba3418),
	.w5(32'hb9ff74ae),
	.w6(32'h37edc360),
	.w7(32'hb999d504),
	.w8(32'hba55a40a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf405b),
	.w1(32'hba9945d2),
	.w2(32'hbab7cc9d),
	.w3(32'hb913d19c),
	.w4(32'hba078c22),
	.w5(32'hba071e70),
	.w6(32'hb9d16c09),
	.w7(32'hba181c77),
	.w8(32'hba173c58),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab36f7),
	.w1(32'hb90823f1),
	.w2(32'hba33bda9),
	.w3(32'hb985ee50),
	.w4(32'hb8cbe906),
	.w5(32'hb9901d34),
	.w6(32'hb6b6ad16),
	.w7(32'hb9e77117),
	.w8(32'hba26019a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93624f),
	.w1(32'hb9747eec),
	.w2(32'hb9f80d4a),
	.w3(32'hba070101),
	.w4(32'hba3e4374),
	.w5(32'hba10d7a4),
	.w6(32'hba85c67b),
	.w7(32'hb98f4ab9),
	.w8(32'hb9330e5d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39918c7f),
	.w1(32'h3a7c0ace),
	.w2(32'h39d56296),
	.w3(32'hb91a6b73),
	.w4(32'h3a456294),
	.w5(32'h399f36d3),
	.w6(32'h3a1eebeb),
	.w7(32'h3a712e79),
	.w8(32'h3a587a8e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af07eb),
	.w1(32'hb92699ff),
	.w2(32'hb9d829d5),
	.w3(32'hb8a14457),
	.w4(32'h38a2872c),
	.w5(32'hb9ab97b5),
	.w6(32'h3975732f),
	.w7(32'hb7bd2d98),
	.w8(32'hb9b29ea8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39795363),
	.w1(32'h393d337c),
	.w2(32'hbabc8e86),
	.w3(32'h3a7d9bb8),
	.w4(32'h396e285f),
	.w5(32'hba8de8d1),
	.w6(32'h3a461eb8),
	.w7(32'hb8ab645e),
	.w8(32'hbb22fd99),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4398fa),
	.w1(32'hbb27009f),
	.w2(32'hbb28bfb8),
	.w3(32'hbaac36cf),
	.w4(32'hba668d9f),
	.w5(32'hba386b46),
	.w6(32'hba33c3f5),
	.w7(32'hba085607),
	.w8(32'hbaf20973),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9952218),
	.w1(32'hb9e4edde),
	.w2(32'hba6af742),
	.w3(32'hb95af6ad),
	.w4(32'hba074d37),
	.w5(32'hba8a2c13),
	.w6(32'hb99bef96),
	.w7(32'h39057944),
	.w8(32'h39206c71),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9076cd6),
	.w1(32'h398521c4),
	.w2(32'h39274fbb),
	.w3(32'hb92ca37e),
	.w4(32'h39a3cf07),
	.w5(32'h38e5c81e),
	.w6(32'h3a2738f0),
	.w7(32'h39ef473a),
	.w8(32'h3a965ace),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87000f),
	.w1(32'h392ae077),
	.w2(32'h39a95f1e),
	.w3(32'h3a570b89),
	.w4(32'h38d8463f),
	.w5(32'h39b2b935),
	.w6(32'h38d17480),
	.w7(32'h379cdccf),
	.w8(32'h38f6c95d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842888b),
	.w1(32'hba179c8a),
	.w2(32'hba7b5683),
	.w3(32'hb8c34125),
	.w4(32'hb9e8406a),
	.w5(32'hb9c7e9ca),
	.w6(32'hb9f6d9c6),
	.w7(32'hb95a7f58),
	.w8(32'hba02b18d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16590c),
	.w1(32'hbba796dd),
	.w2(32'hbbe921ec),
	.w3(32'hba05f16c),
	.w4(32'hbb58996a),
	.w5(32'hbb94042b),
	.w6(32'hbae0ec87),
	.w7(32'hbb898244),
	.w8(32'hbba913a8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c16d3),
	.w1(32'hb9afa053),
	.w2(32'hbbd1aafe),
	.w3(32'h3b4f48b6),
	.w4(32'h3acae648),
	.w5(32'hbba39f74),
	.w6(32'h37e31eb2),
	.w7(32'hbad8db7c),
	.w8(32'hbbf92737),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390181a2),
	.w1(32'h393460eb),
	.w2(32'hbb773bbe),
	.w3(32'h3ab7ad7f),
	.w4(32'h3aa1a0bb),
	.w5(32'hbb3dc7e5),
	.w6(32'hb96f5557),
	.w7(32'hbab6344e),
	.w8(32'hbb9ed928),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dad18),
	.w1(32'h3b2080da),
	.w2(32'hbb863c26),
	.w3(32'h3b33b4e6),
	.w4(32'h3b8c38e7),
	.w5(32'hbb0319e6),
	.w6(32'hba0f2f34),
	.w7(32'hb879ea5c),
	.w8(32'hbbc7f7be),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32e002),
	.w1(32'h38d29ba9),
	.w2(32'h392a23b6),
	.w3(32'h3aaa0bf1),
	.w4(32'h38d153f4),
	.w5(32'h3918e65d),
	.w6(32'h39a5d583),
	.w7(32'h380b7202),
	.w8(32'h39497cf0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bd8eb),
	.w1(32'hb7be4a10),
	.w2(32'hb8fbac2b),
	.w3(32'h396f392f),
	.w4(32'hb8762ccc),
	.w5(32'h38c104e6),
	.w6(32'h383c5e02),
	.w7(32'hb936b2cf),
	.w8(32'hb943f3c9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930ac1f),
	.w1(32'h387c2311),
	.w2(32'h37c8bef2),
	.w3(32'h38d9b627),
	.w4(32'h38f0db43),
	.w5(32'h385c70c7),
	.w6(32'h393a7a13),
	.w7(32'hb812e825),
	.w8(32'h366a42ac),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a312f),
	.w1(32'hb94f7a3b),
	.w2(32'hba92f2ca),
	.w3(32'h393a51e7),
	.w4(32'h389efdd4),
	.w5(32'h390dc242),
	.w6(32'hb9b3023e),
	.w7(32'hba197829),
	.w8(32'hba8e7fa4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969ebe7),
	.w1(32'hb9a9f29d),
	.w2(32'hb9443a87),
	.w3(32'h39819707),
	.w4(32'hba0a7df6),
	.w5(32'hb9ea018c),
	.w6(32'hb7f1f17e),
	.w7(32'hb91c9667),
	.w8(32'hb99fd9e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba744abd),
	.w1(32'hbaaaf780),
	.w2(32'hbb30b013),
	.w3(32'hbaf37168),
	.w4(32'hbb0e8afb),
	.w5(32'hba08d81b),
	.w6(32'hbaca8008),
	.w7(32'hbaf04e6d),
	.w8(32'hbb5e937a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a336),
	.w1(32'h3a95bb76),
	.w2(32'hbb784038),
	.w3(32'h3b70f4a5),
	.w4(32'h39da8ecc),
	.w5(32'hbb58bcc8),
	.w6(32'h3b2318a4),
	.w7(32'h3af91bb2),
	.w8(32'hbb2794a8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4361),
	.w1(32'h3a1360fe),
	.w2(32'hbb2d07e3),
	.w3(32'hb9d5f5c6),
	.w4(32'h39a3637f),
	.w5(32'hbae9bf81),
	.w6(32'hba8fe6a2),
	.w7(32'hbaa81422),
	.w8(32'hbb813e27),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7601f),
	.w1(32'hb92af638),
	.w2(32'hbabd334d),
	.w3(32'h3a87be09),
	.w4(32'hb981a2ef),
	.w5(32'hbab02a6e),
	.w6(32'h398c60df),
	.w7(32'h3990b2e7),
	.w8(32'hbb052202),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb0cdd),
	.w1(32'h39527aa6),
	.w2(32'hbb3424fe),
	.w3(32'hba4a1d01),
	.w4(32'h3a203ce2),
	.w5(32'hbafab798),
	.w6(32'h3a3ae1bd),
	.w7(32'h36d7c47d),
	.w8(32'hbb130a2d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98eeb3),
	.w1(32'hba6e0ab5),
	.w2(32'hbaeafaca),
	.w3(32'h3a2c2df7),
	.w4(32'hb896d9c5),
	.w5(32'hbaa546cf),
	.w6(32'hb88041c2),
	.w7(32'hba2e5d14),
	.w8(32'hbb07f842),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae746f),
	.w1(32'hba8022c2),
	.w2(32'hbb5d612b),
	.w3(32'hba8c6a1b),
	.w4(32'hba250635),
	.w5(32'hbb06accf),
	.w6(32'hb89a25f5),
	.w7(32'hba8f3e27),
	.w8(32'hbb1ffc50),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913adba),
	.w1(32'hba29cb01),
	.w2(32'hba32151e),
	.w3(32'h3850d2ef),
	.w4(32'hba4bc06a),
	.w5(32'hba09b61c),
	.w6(32'hba083be0),
	.w7(32'hba43ec76),
	.w8(32'hba17b6eb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd129f),
	.w1(32'hb99c5ae6),
	.w2(32'hb8b72ea5),
	.w3(32'hb9af1a9d),
	.w4(32'hb8324761),
	.w5(32'h38a9a683),
	.w6(32'hb93e4bd2),
	.w7(32'hb917ba31),
	.w8(32'hb8922263),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2398a),
	.w1(32'h3aa4ff1b),
	.w2(32'h3ad862a0),
	.w3(32'h3681c7f2),
	.w4(32'h3a1c67e7),
	.w5(32'h3a5e8dbf),
	.w6(32'h393c5ecb),
	.w7(32'h39bc239d),
	.w8(32'h39aa37b9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22838b),
	.w1(32'hb944294a),
	.w2(32'hb9ca3c66),
	.w3(32'h38608514),
	.w4(32'h39c4027f),
	.w5(32'h39e5797e),
	.w6(32'hba0409fb),
	.w7(32'hb9f19742),
	.w8(32'h38a39847),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7d454),
	.w1(32'h3abdcbe9),
	.w2(32'h3a1fbb8a),
	.w3(32'hbad88d76),
	.w4(32'h3a35dea6),
	.w5(32'hb99244bb),
	.w6(32'hbb51a68b),
	.w7(32'hba696370),
	.w8(32'hba5c4699),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bdf61),
	.w1(32'h3a4bd20b),
	.w2(32'hb999eafd),
	.w3(32'h39056142),
	.w4(32'h3a8be78c),
	.w5(32'hb943ba64),
	.w6(32'hba00265e),
	.w7(32'h39a25aeb),
	.w8(32'hb9ed81a8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5959f0),
	.w1(32'hb919a77a),
	.w2(32'hbaf80e8b),
	.w3(32'h3a2f9bdd),
	.w4(32'h3a749776),
	.w5(32'hba9d2b74),
	.w6(32'hba8b9c4c),
	.w7(32'h37a163ae),
	.w8(32'hbb0f04e9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364711),
	.w1(32'hbb4b70eb),
	.w2(32'hbbafb7e3),
	.w3(32'hbb48bf85),
	.w4(32'hbb07504f),
	.w5(32'hbb5850ad),
	.w6(32'hbb388dbe),
	.w7(32'hbabd906a),
	.w8(32'hbb61cb34),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f2429),
	.w1(32'h3abf614e),
	.w2(32'hb976b0d9),
	.w3(32'h3a4e394d),
	.w4(32'h3b10baf6),
	.w5(32'h3aced76a),
	.w6(32'hbaa7044e),
	.w7(32'h3a00dbe0),
	.w8(32'h385e8cac),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09783b),
	.w1(32'h3a1c2707),
	.w2(32'hbbb18ed4),
	.w3(32'h3abfbd75),
	.w4(32'h38b8c788),
	.w5(32'hbba50883),
	.w6(32'h3ab23e0d),
	.w7(32'h381779c9),
	.w8(32'hbb86c14a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c932),
	.w1(32'h3aa49cbd),
	.w2(32'hba641faa),
	.w3(32'h3af08480),
	.w4(32'h3a9e8d32),
	.w5(32'hb987bf7f),
	.w6(32'hbaf1c98e),
	.w7(32'hba41643b),
	.w8(32'hba9ba6d4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ffc76),
	.w1(32'hbb1847fa),
	.w2(32'hbbed3f4e),
	.w3(32'h3a879f07),
	.w4(32'hba34f398),
	.w5(32'hbb900005),
	.w6(32'h3a208eba),
	.w7(32'hba3bf912),
	.w8(32'hbb8845aa),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383bb7b4),
	.w1(32'hba6a9048),
	.w2(32'hbada5899),
	.w3(32'hb983f140),
	.w4(32'hba0c4e9d),
	.w5(32'hbb0e8f70),
	.w6(32'hbab3310c),
	.w7(32'hbaa4b4de),
	.w8(32'hbb315455),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6328b2),
	.w1(32'hba0d5387),
	.w2(32'hbaccfb7e),
	.w3(32'h386f2299),
	.w4(32'h39dfd2df),
	.w5(32'hba3a4d22),
	.w6(32'hbb0d42d2),
	.w7(32'hba695e1d),
	.w8(32'hbb0fc5ff),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87c5cf),
	.w1(32'h3a7e8207),
	.w2(32'h3a1eec73),
	.w3(32'h3a3a043d),
	.w4(32'h3a6e37a5),
	.w5(32'hb95a9e61),
	.w6(32'h3aceb3b8),
	.w7(32'h39b19791),
	.w8(32'hb6a56ed2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7593f2),
	.w1(32'h38acf3a0),
	.w2(32'hbbfb808a),
	.w3(32'h3af2876d),
	.w4(32'h3a28e224),
	.w5(32'hbbff6ffa),
	.w6(32'h3a911be7),
	.w7(32'hba6829dd),
	.w8(32'hbbeeeb90),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72d93f),
	.w1(32'hba85f4e6),
	.w2(32'hbbad44e2),
	.w3(32'h3a0dcdbc),
	.w4(32'hba81bab5),
	.w5(32'hbbad9b51),
	.w6(32'h389d0a91),
	.w7(32'hbb02078f),
	.w8(32'hbb9a3636),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904fe2f),
	.w1(32'h3b79d839),
	.w2(32'hbbbe6f18),
	.w3(32'hbb3a8fcb),
	.w4(32'h3ad81f1a),
	.w5(32'hbb85f198),
	.w6(32'hbb7e3efc),
	.w7(32'hb89fed94),
	.w8(32'hbba10dee),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6a66),
	.w1(32'h3be8fd64),
	.w2(32'h3b0cb97c),
	.w3(32'h3a3b0ef6),
	.w4(32'h3c18ee94),
	.w5(32'h3b7f6081),
	.w6(32'hbb6dd3af),
	.w7(32'h3bd6f11d),
	.w8(32'h3ab31376),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9565f3),
	.w1(32'h3a727f12),
	.w2(32'hbb7f6041),
	.w3(32'h3ac3b1f2),
	.w4(32'h3b2a1d65),
	.w5(32'hbb0f4938),
	.w6(32'hb9c91c62),
	.w7(32'h3903b46d),
	.w8(32'hbbe491c2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972452e),
	.w1(32'h3a6af7ec),
	.w2(32'hbbd833a4),
	.w3(32'h3aad7e18),
	.w4(32'h3b488d30),
	.w5(32'hbb754872),
	.w6(32'h3a292f47),
	.w7(32'h3b775a96),
	.w8(32'hb868864b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c827f),
	.w1(32'h3a40d79f),
	.w2(32'hba230bdc),
	.w3(32'h3af198a2),
	.w4(32'h3aa47124),
	.w5(32'hb9c70fe1),
	.w6(32'h3b1b2fe0),
	.w7(32'h3abb768f),
	.w8(32'h3a8ccccc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2af354),
	.w1(32'h3b0a6e74),
	.w2(32'hbba87caa),
	.w3(32'hbb08a1a2),
	.w4(32'h3ac7bacf),
	.w5(32'hbb1410cd),
	.w6(32'h3966a703),
	.w7(32'h3b047023),
	.w8(32'hbb6d1cf4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05abc8),
	.w1(32'h396e7392),
	.w2(32'hbb53c7b3),
	.w3(32'h3ad15808),
	.w4(32'hb9a49634),
	.w5(32'hbb8bc79e),
	.w6(32'h3b116f26),
	.w7(32'h39d029ab),
	.w8(32'hbb85bd94),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997cbf3),
	.w1(32'hb8d9bf86),
	.w2(32'h394122a2),
	.w3(32'hb96c2727),
	.w4(32'h377543c2),
	.w5(32'h39a3bb5f),
	.w6(32'h398353c1),
	.w7(32'h39b87b56),
	.w8(32'h39ae23d5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989663c),
	.w1(32'hba6433f6),
	.w2(32'hba84e434),
	.w3(32'h372f896a),
	.w4(32'hb95f6fbd),
	.w5(32'hb8e77658),
	.w6(32'hba74de5a),
	.w7(32'hba62e3f5),
	.w8(32'hba83a647),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a812d37),
	.w1(32'h3a13d0b2),
	.w2(32'hbb9681ab),
	.w3(32'h3b36a716),
	.w4(32'h3acc24d5),
	.w5(32'hbb6bc930),
	.w6(32'h3b2b2ebf),
	.w7(32'h3a4441ae),
	.w8(32'hbb95ceb8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fbb16),
	.w1(32'h3af7c5c4),
	.w2(32'hba1e29a3),
	.w3(32'h3b1c064b),
	.w4(32'h3b5ce86e),
	.w5(32'hba31728d),
	.w6(32'h3b1a9c9c),
	.w7(32'h3b180f26),
	.w8(32'hba884668),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39305a67),
	.w1(32'hbada1e3f),
	.w2(32'hbb1482b8),
	.w3(32'h3abb503f),
	.w4(32'hba353be1),
	.w5(32'hbaaf052b),
	.w6(32'hb9b82a2c),
	.w7(32'hba5b0113),
	.w8(32'hbad90e2f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b67aec),
	.w1(32'hb996ee0a),
	.w2(32'hbb6e6df9),
	.w3(32'h3a9b6268),
	.w4(32'h3aa239a4),
	.w5(32'hbb35aa86),
	.w6(32'h3a1fba6b),
	.w7(32'h399edd62),
	.w8(32'hbb03a173),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b50c5),
	.w1(32'h3b0ee706),
	.w2(32'hb7d3b8d8),
	.w3(32'h3ab7a938),
	.w4(32'h3b4679b2),
	.w5(32'h3a8ba5e7),
	.w6(32'hba8a07d9),
	.w7(32'h395e62c1),
	.w8(32'hba7df536),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5499e),
	.w1(32'hbabc69e7),
	.w2(32'hbb1535d2),
	.w3(32'hb9eaa728),
	.w4(32'hba8a1d00),
	.w5(32'hbae65eae),
	.w6(32'h3a8b9771),
	.w7(32'h3925edf8),
	.w8(32'hbae80f0b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954cfe0),
	.w1(32'hba86077d),
	.w2(32'hbb2398a6),
	.w3(32'h39ba6344),
	.w4(32'h3938b536),
	.w5(32'hbb1e0a58),
	.w6(32'hb9c68273),
	.w7(32'hb7339898),
	.w8(32'hbb2d8b0a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968d9a8),
	.w1(32'hb82bd33b),
	.w2(32'hb9aec682),
	.w3(32'hb8542557),
	.w4(32'h39039ff0),
	.w5(32'hb926db72),
	.w6(32'h393e8e46),
	.w7(32'hb7f5f16e),
	.w8(32'h3993c613),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8056487),
	.w1(32'hb8e61fed),
	.w2(32'hb8b831d7),
	.w3(32'h3970f16a),
	.w4(32'hb7ffa100),
	.w5(32'hb6d376ec),
	.w6(32'hb8aad588),
	.w7(32'hb8a2236a),
	.w8(32'hb8799339),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38740a15),
	.w1(32'hb63acd61),
	.w2(32'hb8d9d890),
	.w3(32'h38b8bb9b),
	.w4(32'hb8debc7e),
	.w5(32'hb94c3c1b),
	.w6(32'hb90ad43d),
	.w7(32'hb98f7d4a),
	.w8(32'hb87703ed),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8295710),
	.w1(32'hbae21039),
	.w2(32'hba900a6a),
	.w3(32'hb9b2db6d),
	.w4(32'hb90d8fe0),
	.w5(32'hba07a9bf),
	.w6(32'hbaa56092),
	.w7(32'hba53fb17),
	.w8(32'hba43230a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d4829),
	.w1(32'h3a775f5b),
	.w2(32'hba31adba),
	.w3(32'h3aae3da6),
	.w4(32'h3ae16103),
	.w5(32'hba5248aa),
	.w6(32'hb6fbeb6b),
	.w7(32'h37a350fb),
	.w8(32'hbb543a58),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bd3f7),
	.w1(32'hba6882e0),
	.w2(32'hba6b5ff5),
	.w3(32'h393ecdba),
	.w4(32'hba048eef),
	.w5(32'hba26e14e),
	.w6(32'hba094108),
	.w7(32'hb9a8aceb),
	.w8(32'hb9c72338),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2cb41),
	.w1(32'hba990eb3),
	.w2(32'hbb5c7e6c),
	.w3(32'hbaaec747),
	.w4(32'hbabbf5c0),
	.w5(32'hbb59af30),
	.w6(32'hb9b60439),
	.w7(32'hba9c645d),
	.w8(32'hbb3d1ed3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31f6cd),
	.w1(32'hb9922e8e),
	.w2(32'hbb2020e5),
	.w3(32'h3a0995df),
	.w4(32'h3a6b6941),
	.w5(32'hbad538d3),
	.w6(32'hba24f2ee),
	.w7(32'hb92a37a8),
	.w8(32'hbb56a3fa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aea854),
	.w1(32'hbaa92b6e),
	.w2(32'hba5596a9),
	.w3(32'h38f7c28a),
	.w4(32'hba4f6d94),
	.w5(32'hb9d8aa09),
	.w6(32'hb99871f9),
	.w7(32'hb8f2abf1),
	.w8(32'hb9f8f993),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e269c),
	.w1(32'hb9d891a1),
	.w2(32'hba8e35e0),
	.w3(32'hb95f0840),
	.w4(32'hba288656),
	.w5(32'hbaab7a0a),
	.w6(32'hba37d0aa),
	.w7(32'hba95796f),
	.w8(32'hba890a22),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa53a3),
	.w1(32'hb9d747a5),
	.w2(32'hba065aef),
	.w3(32'hbad7b50b),
	.w4(32'h3909329a),
	.w5(32'h39332112),
	.w6(32'hb952c4cc),
	.w7(32'hb9e600f4),
	.w8(32'hb9bc8f50),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f65869),
	.w1(32'hb8b850c4),
	.w2(32'hba9e1705),
	.w3(32'hba0ce570),
	.w4(32'hb9f2e477),
	.w5(32'hbaa31d31),
	.w6(32'hbaa8073d),
	.w7(32'hba912c76),
	.w8(32'hbaa18dc6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe12e),
	.w1(32'h3a246f46),
	.w2(32'hbb870bed),
	.w3(32'h3b8f0702),
	.w4(32'h3a4d08e4),
	.w5(32'hbb490b38),
	.w6(32'h3a42f5e4),
	.w7(32'hba6e332e),
	.w8(32'hbb82ea55),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a73a04),
	.w1(32'hbb264586),
	.w2(32'hbbabf0ba),
	.w3(32'h3ab2f2bd),
	.w4(32'hbaf9a9ef),
	.w5(32'hbb87f71a),
	.w6(32'h3a1f483a),
	.w7(32'hba61bc2b),
	.w8(32'hbb895bdc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936c800),
	.w1(32'h38fa3198),
	.w2(32'hb97be033),
	.w3(32'h3970fb3f),
	.w4(32'h39a9a43f),
	.w5(32'h38f6f6b2),
	.w6(32'h3a173bfe),
	.w7(32'h39cf1947),
	.w8(32'h3985ae94),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39958e58),
	.w1(32'hb9d451a9),
	.w2(32'hba66f412),
	.w3(32'h38b940d4),
	.w4(32'hb85ad6bf),
	.w5(32'hba1daceb),
	.w6(32'hb9bf3ebc),
	.w7(32'hb9c7dd83),
	.w8(32'hbaa1efef),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7f0e9),
	.w1(32'hb978de47),
	.w2(32'hba1bc5e2),
	.w3(32'hb91a969f),
	.w4(32'h39debd6f),
	.w5(32'h392b36c8),
	.w6(32'hb96708f7),
	.w7(32'h38e0d484),
	.w8(32'h38a8bf1b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02c475),
	.w1(32'h39c47b61),
	.w2(32'hbaa82feb),
	.w3(32'h3a7edb4a),
	.w4(32'h39fa64b6),
	.w5(32'hba80601c),
	.w6(32'h3a429daf),
	.w7(32'h39b212a6),
	.w8(32'hbab42180),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb444d20),
	.w1(32'hbb3ccf53),
	.w2(32'hbb2d43fb),
	.w3(32'hbb240b1a),
	.w4(32'hbaf996db),
	.w5(32'hbac4d779),
	.w6(32'hbafd624d),
	.w7(32'hbadaa5e2),
	.w8(32'hbafa1492),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404001),
	.w1(32'hba889a97),
	.w2(32'hbbb8ef4d),
	.w3(32'h39c2765a),
	.w4(32'hb8fda432),
	.w5(32'hbb9ceb92),
	.w6(32'h398646a0),
	.w7(32'hbb19b1f3),
	.w8(32'hbbb9d695),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f4f57),
	.w1(32'h3a510414),
	.w2(32'hbb021d43),
	.w3(32'h3ad0115f),
	.w4(32'h3b0f790f),
	.w5(32'hba68d91d),
	.w6(32'h39937d5a),
	.w7(32'h3aada9ec),
	.w8(32'hba98c195),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb844d951),
	.w1(32'hba194876),
	.w2(32'hbb7e8bcb),
	.w3(32'h3a28401d),
	.w4(32'hb9c3f072),
	.w5(32'hbb6e9d53),
	.w6(32'hba8a91a6),
	.w7(32'hba18d908),
	.w8(32'hbb23ab98),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96dc88),
	.w1(32'hbac1edd6),
	.w2(32'hbb93e00d),
	.w3(32'hbaca9c95),
	.w4(32'hba7b41a5),
	.w5(32'hbb46d4fd),
	.w6(32'hb9c21fa6),
	.w7(32'hba8791ed),
	.w8(32'hbb542225),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52b52e),
	.w1(32'h3a0a9151),
	.w2(32'hba18bb8a),
	.w3(32'hb9054390),
	.w4(32'h3aa8a89d),
	.w5(32'h3a10fc64),
	.w6(32'hba9bb9c7),
	.w7(32'h39b6dceb),
	.w8(32'hbaade4c6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bd549),
	.w1(32'hbab61ae2),
	.w2(32'hbb98c756),
	.w3(32'h3a55be43),
	.w4(32'hb90da076),
	.w5(32'hbb74179c),
	.w6(32'h3aaa58f5),
	.w7(32'h39cae7e4),
	.w8(32'hbb5f7149),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94848f3),
	.w1(32'h37fef4b6),
	.w2(32'hba24c9e1),
	.w3(32'h393d6b2d),
	.w4(32'h39c90202),
	.w5(32'hba0d23f1),
	.w6(32'h39472465),
	.w7(32'h3921b3ca),
	.w8(32'hba7803e1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4c18b),
	.w1(32'hbb15f9de),
	.w2(32'hbb76e80a),
	.w3(32'h3a530fad),
	.w4(32'hb8ef4fff),
	.w5(32'hbb4646bb),
	.w6(32'hbb0e13cc),
	.w7(32'hbb15b570),
	.w8(32'hbb803cff),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39e0b),
	.w1(32'hba88ddf1),
	.w2(32'hbac3cb5d),
	.w3(32'hbabe62e6),
	.w4(32'hba487acf),
	.w5(32'hb9f67fe5),
	.w6(32'hbb1883c2),
	.w7(32'hba86ee50),
	.w8(32'hba8a6a44),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937d120),
	.w1(32'h38a049b0),
	.w2(32'hb867fb66),
	.w3(32'hb93bb75b),
	.w4(32'h38453572),
	.w5(32'hb89aba22),
	.w6(32'h390c17d4),
	.w7(32'h37ceb6e9),
	.w8(32'h3839228e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378336ac),
	.w1(32'h38bd447d),
	.w2(32'h396d479f),
	.w3(32'h3838558c),
	.w4(32'h39279d95),
	.w5(32'h397d9b16),
	.w6(32'h382e4d2a),
	.w7(32'h38fc9b51),
	.w8(32'h39293e77),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c913c),
	.w1(32'h3a9333b8),
	.w2(32'h39234ae8),
	.w3(32'h38d6ee5e),
	.w4(32'h398d10e6),
	.w5(32'hb99e4446),
	.w6(32'h3984213a),
	.w7(32'h399e18af),
	.w8(32'hba600b1b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fecde),
	.w1(32'hb9d255c4),
	.w2(32'hbb1f1a47),
	.w3(32'hbac2c2dd),
	.w4(32'h3a846ce7),
	.w5(32'hba08dd05),
	.w6(32'hbb3cdecb),
	.w7(32'hba129f83),
	.w8(32'hbaf03e18),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1476d6),
	.w1(32'h3b160be1),
	.w2(32'hbad65458),
	.w3(32'h3b367adf),
	.w4(32'h3acc67f6),
	.w5(32'hba970403),
	.w6(32'h3b0b5c0b),
	.w7(32'h39b6ca7b),
	.w8(32'hbb89666d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c9fcd8),
	.w1(32'hb8111ad8),
	.w2(32'hb950d1ea),
	.w3(32'h378763b4),
	.w4(32'h3787d3c4),
	.w5(32'hb8bcb4c4),
	.w6(32'h387eeec8),
	.w7(32'hb8bf4721),
	.w8(32'hb7fe41b0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9752d9b),
	.w1(32'hba38dd7b),
	.w2(32'hbb9a49cf),
	.w3(32'h3a4b8698),
	.w4(32'h38c32f1f),
	.w5(32'hbb6432ed),
	.w6(32'h39e131cd),
	.w7(32'hba46533a),
	.w8(32'hbbb02e5f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61066b),
	.w1(32'h37418690),
	.w2(32'hbb500d82),
	.w3(32'h3aa789b4),
	.w4(32'h394a247b),
	.w5(32'hbb3aa566),
	.w6(32'hba20152b),
	.w7(32'h37d95f29),
	.w8(32'hbb70e482),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d0111),
	.w1(32'hbaf068aa),
	.w2(32'hbbdf8e37),
	.w3(32'hbb125ad8),
	.w4(32'hbb037e52),
	.w5(32'hbbb5d824),
	.w6(32'h39a8c2a6),
	.w7(32'hba3df5fc),
	.w8(32'hbb9521c6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869600e),
	.w1(32'hba4601be),
	.w2(32'hbaf3640a),
	.w3(32'h3a3d6e36),
	.w4(32'h3a94ed56),
	.w5(32'hba898314),
	.w6(32'hba54adf4),
	.w7(32'hbb0667c8),
	.w8(32'hbb6cedfd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7244e),
	.w1(32'h3a8b62a8),
	.w2(32'h3a3b94a1),
	.w3(32'h37b04cf6),
	.w4(32'h3ac9ce3b),
	.w5(32'h3ac73406),
	.w6(32'h38c74ac1),
	.w7(32'h3a5544c7),
	.w8(32'h3abf31c5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff034c),
	.w1(32'h3aae9e20),
	.w2(32'h3abc53c0),
	.w3(32'h3aba5320),
	.w4(32'h3aaed889),
	.w5(32'h3a973440),
	.w6(32'h3aee6f54),
	.w7(32'h3abfa69a),
	.w8(32'h3a394ce3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada847d),
	.w1(32'h39ac225d),
	.w2(32'hbab9b8a5),
	.w3(32'h398d6a1d),
	.w4(32'h3a90e3b8),
	.w5(32'hba7e1ce0),
	.w6(32'h38784c78),
	.w7(32'h3a914a30),
	.w8(32'hba79680e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d18b4),
	.w1(32'h39c258a1),
	.w2(32'hb9c51266),
	.w3(32'h3a9e52d1),
	.w4(32'h3afa226d),
	.w5(32'h3ae02ef5),
	.w6(32'hbac484cc),
	.w7(32'h38dc7d2a),
	.w8(32'h3ab44779),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5357e),
	.w1(32'h3abb88f0),
	.w2(32'h3a41e937),
	.w3(32'h39c5cd96),
	.w4(32'h3abcf8b3),
	.w5(32'h3a990670),
	.w6(32'hb900cea8),
	.w7(32'h3a7dca88),
	.w8(32'h3a2f2cac),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91837a1),
	.w1(32'hba16f782),
	.w2(32'hba9eecfb),
	.w3(32'hb9a199a4),
	.w4(32'hb9a5e2b7),
	.w5(32'hba45a2da),
	.w6(32'hb9b1d796),
	.w7(32'hba069b85),
	.w8(32'hba3be6e9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e0098),
	.w1(32'hb9026127),
	.w2(32'hb96a2c8d),
	.w3(32'hb6b78c02),
	.w4(32'hb7d80fbc),
	.w5(32'hb8cdf90c),
	.w6(32'hb89b0b8c),
	.w7(32'hb90e5327),
	.w8(32'hb92c4018),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898179e),
	.w1(32'hbaa01622),
	.w2(32'hbb9db521),
	.w3(32'h3aae961c),
	.w4(32'h3992f236),
	.w5(32'hbb71f223),
	.w6(32'hb99d4763),
	.w7(32'hb9b4f88c),
	.w8(32'hbb726205),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1399e),
	.w1(32'h389ed1bf),
	.w2(32'hba4c34bd),
	.w3(32'h38fb2ef2),
	.w4(32'h38478d14),
	.w5(32'hba1fd43d),
	.w6(32'h39a5fda3),
	.w7(32'h39291696),
	.w8(32'hb9b798a6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb5d55),
	.w1(32'h39fa3f85),
	.w2(32'hba75076e),
	.w3(32'h3aa7c9bc),
	.w4(32'h3ab63929),
	.w5(32'hb9b86e32),
	.w6(32'h3a8d2f12),
	.w7(32'h3a7dd16c),
	.w8(32'hbab00200),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9258e3d),
	.w1(32'h392dbe87),
	.w2(32'h39380513),
	.w3(32'hb9ac6800),
	.w4(32'hb9107a3c),
	.w5(32'h390d1ecb),
	.w6(32'hb98201f7),
	.w7(32'h38ee21c1),
	.w8(32'h39ad5bc3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af58e77),
	.w1(32'h39a3a937),
	.w2(32'hbab17e81),
	.w3(32'h3ac4e9ec),
	.w4(32'h399baa96),
	.w5(32'hbb2b0d5e),
	.w6(32'h3a8da9f5),
	.w7(32'hb9cb84bf),
	.w8(32'hbb329068),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0c49e),
	.w1(32'h39d13aa2),
	.w2(32'h3a2166fb),
	.w3(32'h39aa7a5b),
	.w4(32'h3a22e1f8),
	.w5(32'h3a49b2e4),
	.w6(32'h39e67666),
	.w7(32'h39f0c300),
	.w8(32'h3a06da37),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b49147),
	.w1(32'h3880ba4a),
	.w2(32'h3782e16b),
	.w3(32'h39c9e609),
	.w4(32'hb97c947e),
	.w5(32'hb9933962),
	.w6(32'h394c73c7),
	.w7(32'hb9327643),
	.w8(32'hb88532bc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e0f534),
	.w1(32'h39a6d174),
	.w2(32'hbaaa2a54),
	.w3(32'h3ad48a0c),
	.w4(32'h3b36ca83),
	.w5(32'h3a157735),
	.w6(32'h3a934d4a),
	.w7(32'h3b557dc0),
	.w8(32'h3a390c92),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961ebcb),
	.w1(32'hb9b64eec),
	.w2(32'hbbd1158e),
	.w3(32'hb8b3131f),
	.w4(32'h3a58c394),
	.w5(32'hbbaa1b54),
	.w6(32'hba859d0c),
	.w7(32'hba1f6faa),
	.w8(32'hbbc0ad5f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd6a0),
	.w1(32'h3b372ee1),
	.w2(32'h3a8cc809),
	.w3(32'h3a09a5ed),
	.w4(32'h3ad4c646),
	.w5(32'h3a430bda),
	.w6(32'h39adeec4),
	.w7(32'h3a1ee49c),
	.w8(32'h398d5d29),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1defbb),
	.w1(32'h3ab11d72),
	.w2(32'hbab5e77f),
	.w3(32'h3ae87ee5),
	.w4(32'h3b142117),
	.w5(32'hbab2c75a),
	.w6(32'h3aad9acb),
	.w7(32'h3ac69c33),
	.w8(32'hbb4d4317),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21560e),
	.w1(32'h353ae3e8),
	.w2(32'hb99199e6),
	.w3(32'hb703be46),
	.w4(32'hb854b5cd),
	.w5(32'hb81ff81f),
	.w6(32'h3961f4fa),
	.w7(32'h3884362b),
	.w8(32'hb844f460),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40c22d),
	.w1(32'hb8dbafc4),
	.w2(32'hbb489b13),
	.w3(32'h3b6265d1),
	.w4(32'h3a9b42f5),
	.w5(32'hbafda566),
	.w6(32'h38ca7916),
	.w7(32'hbb494c36),
	.w8(32'hbb9cee22),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dac436),
	.w1(32'h39c95d81),
	.w2(32'hbb3faa15),
	.w3(32'h3a70ac9a),
	.w4(32'h3a9efe83),
	.w5(32'hbb13c1c3),
	.w6(32'h3903cc33),
	.w7(32'h399e3ca2),
	.w8(32'hbb296be5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95c6a6),
	.w1(32'hbb382ed1),
	.w2(32'hbb9eb51b),
	.w3(32'hb9d63822),
	.w4(32'hbb1ea05d),
	.w5(32'hbbac86b1),
	.w6(32'hb959a821),
	.w7(32'hbaef7b53),
	.w8(32'hbbbf5b7a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952a222),
	.w1(32'h3a4147a3),
	.w2(32'h39961312),
	.w3(32'h396d2c8e),
	.w4(32'h3a335cd3),
	.w5(32'h3a1c38db),
	.w6(32'h390842d7),
	.w7(32'h3a1a5bf4),
	.w8(32'h3a050285),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a010),
	.w1(32'hbb21f560),
	.w2(32'hbb56ad0f),
	.w3(32'hb97b22f4),
	.w4(32'hbace02b1),
	.w5(32'hbaebcd1b),
	.w6(32'h38b85189),
	.w7(32'hba7bb1ef),
	.w8(32'hbab3a53f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a150c5),
	.w1(32'hb5ae7350),
	.w2(32'hb737bae3),
	.w3(32'hb833435d),
	.w4(32'hb7c21d2c),
	.w5(32'hb7bd55a3),
	.w6(32'h37b62f15),
	.w7(32'hb80e9b16),
	.w8(32'h382f96df),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f07b7),
	.w1(32'hba846caf),
	.w2(32'hbaaafdfe),
	.w3(32'hb9cd8c01),
	.w4(32'hbaa1ef57),
	.w5(32'hbadfc01b),
	.w6(32'hba0b2b3c),
	.w7(32'hba89c770),
	.w8(32'hbaef8ee0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3c477),
	.w1(32'hba148d20),
	.w2(32'hb8879732),
	.w3(32'hb97682ac),
	.w4(32'hba467a03),
	.w5(32'hb9c6dba4),
	.w6(32'hb9ef934c),
	.w7(32'hba180408),
	.w8(32'hb9e0aa7e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911eddf),
	.w1(32'hbab1c6fa),
	.w2(32'hbb39dca8),
	.w3(32'hba9949fc),
	.w4(32'hbab3b0c2),
	.w5(32'hbae3ff29),
	.w6(32'hba8be9d5),
	.w7(32'hbaf3d47a),
	.w8(32'hbb42fd3b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736f2bb),
	.w1(32'h38b5fea4),
	.w2(32'h38f2edb1),
	.w3(32'h364848c3),
	.w4(32'h392a287a),
	.w5(32'h38e20eda),
	.w6(32'h3916a77e),
	.w7(32'h391c4f00),
	.w8(32'h38f59994),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39029fd4),
	.w1(32'h392e1d4f),
	.w2(32'hb82e077b),
	.w3(32'h3935f267),
	.w4(32'h3981aaa8),
	.w5(32'h387735a3),
	.w6(32'h3990f290),
	.w7(32'h39969c68),
	.w8(32'h391ba2ab),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d067ce),
	.w1(32'h39871e1d),
	.w2(32'h38610b01),
	.w3(32'h3a27efa1),
	.w4(32'h39f33766),
	.w5(32'h393136d4),
	.w6(32'h38fe4074),
	.w7(32'h383146af),
	.w8(32'hb9e6c010),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f3fc0),
	.w1(32'h3aa56468),
	.w2(32'hbb8026a6),
	.w3(32'h3ad20d45),
	.w4(32'h3ab7c453),
	.w5(32'hbb6875f4),
	.w6(32'hb8910158),
	.w7(32'hbaaae86a),
	.w8(32'hbb80816e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b506b2),
	.w1(32'h3a612801),
	.w2(32'hbb203a56),
	.w3(32'hba91eac6),
	.w4(32'h3a8e124c),
	.w5(32'hbaf3f0fe),
	.w6(32'h3a6e8cd4),
	.w7(32'h3b084b78),
	.w8(32'hba990fde),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9217a3b),
	.w1(32'h3506b049),
	.w2(32'h39c14d50),
	.w3(32'hba1a04f2),
	.w4(32'hb88f06ee),
	.w5(32'h39d8abe7),
	.w6(32'hba30d5b3),
	.w7(32'hb9ef92d9),
	.w8(32'hb80d3729),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be19638),
	.w1(32'h3b339ae4),
	.w2(32'hbbaf2a0c),
	.w3(32'h3c2efdb3),
	.w4(32'h3b82caa9),
	.w5(32'hbbd9f578),
	.w6(32'h3beb840b),
	.w7(32'h3b1e7f94),
	.w8(32'hbc0e6954),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf62704),
	.w1(32'hbb12cd1f),
	.w2(32'hbb7735b3),
	.w3(32'h37d42674),
	.w4(32'h3b089d94),
	.w5(32'h3afe2ace),
	.w6(32'hbadd772d),
	.w7(32'h3a8c94fa),
	.w8(32'h3adaf9e9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a5ba),
	.w1(32'h39c558e1),
	.w2(32'hba8ada0f),
	.w3(32'h3a5c077a),
	.w4(32'h39ad0261),
	.w5(32'hba56425e),
	.w6(32'h3a5fe0c6),
	.w7(32'h3a2287b1),
	.w8(32'hb9d883f5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cc99e),
	.w1(32'hb96fa193),
	.w2(32'hb96db946),
	.w3(32'h38b4560d),
	.w4(32'hb983527e),
	.w5(32'hb91e2b0f),
	.w6(32'hb8f0aa76),
	.w7(32'hb99904b8),
	.w8(32'hb9910e31),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9405618),
	.w1(32'h3869ff87),
	.w2(32'h3819cb85),
	.w3(32'hb8661584),
	.w4(32'h3865e64e),
	.w5(32'hb90303ab),
	.w6(32'h398be7db),
	.w7(32'hb8f2d267),
	.w8(32'h38498eb4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875cd3d),
	.w1(32'hb847c5e6),
	.w2(32'h383959e1),
	.w3(32'h38a6ccf8),
	.w4(32'hb5f78bed),
	.w5(32'h381a6cdc),
	.w6(32'h37be2f38),
	.w7(32'h37bc4f2a),
	.w8(32'h390ad8ee),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd0d3a),
	.w1(32'h3985d47d),
	.w2(32'hbb0652a6),
	.w3(32'h3a5dcbf4),
	.w4(32'h37ad66c0),
	.w5(32'hbb08519a),
	.w6(32'h39bb8ed9),
	.w7(32'h39f52f97),
	.w8(32'hba993d41),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73e69b),
	.w1(32'hbaf713ae),
	.w2(32'hbb0ad816),
	.w3(32'hba5bb79b),
	.w4(32'h39bf52ba),
	.w5(32'hbaad8bf6),
	.w6(32'hbb06393c),
	.w7(32'hbb21ec6d),
	.w8(32'hbb5b6a1c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1b976),
	.w1(32'h38ccf58f),
	.w2(32'hbb37645e),
	.w3(32'hb92e28ff),
	.w4(32'h3a8ad843),
	.w5(32'hbabc24f1),
	.w6(32'hbab2a1c0),
	.w7(32'hb9ee88a5),
	.w8(32'hbb4af433),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba123932),
	.w1(32'hb91583c2),
	.w2(32'hb905c793),
	.w3(32'hb9c13344),
	.w4(32'hb9d795c8),
	.w5(32'hba4a1d28),
	.w6(32'hb915cb46),
	.w7(32'hb5fcb2fb),
	.w8(32'hba09645e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7d6ba),
	.w1(32'h3b1abcf3),
	.w2(32'hbba74a63),
	.w3(32'h3ad2c07a),
	.w4(32'h3b0dc31c),
	.w5(32'hbb9cb75a),
	.w6(32'h39071d25),
	.w7(32'h397f21e8),
	.w8(32'hbbbbb07e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c67bb),
	.w1(32'h3968244e),
	.w2(32'hba4e7005),
	.w3(32'h39b5503b),
	.w4(32'hb921245e),
	.w5(32'hba6c25f0),
	.w6(32'h3a266366),
	.w7(32'hba3a7691),
	.w8(32'hbaf8eb9e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948e7e6),
	.w1(32'h389eb264),
	.w2(32'h38a6f799),
	.w3(32'h396e961f),
	.w4(32'h389d97af),
	.w5(32'h38b1e4e3),
	.w6(32'h38cbde95),
	.w7(32'h38936421),
	.w8(32'h390be882),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bba2fd),
	.w1(32'hba0b2bfd),
	.w2(32'hba4a97d7),
	.w3(32'hb9825512),
	.w4(32'hba05a381),
	.w5(32'h37932710),
	.w6(32'h3a0496fd),
	.w7(32'hb9076e11),
	.w8(32'hb75b629e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da3b57),
	.w1(32'h3710e032),
	.w2(32'h3810f5f0),
	.w3(32'hb7b6c78a),
	.w4(32'h385bfa3e),
	.w5(32'h38b9a64e),
	.w6(32'h38994a0b),
	.w7(32'hb8161df9),
	.w8(32'h3898804b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fcfcd),
	.w1(32'h3afbc7fe),
	.w2(32'hbb1f0d97),
	.w3(32'h3b309c73),
	.w4(32'h3b2d7776),
	.w5(32'hbac6deb6),
	.w6(32'h3ac231fa),
	.w7(32'h3a54f09f),
	.w8(32'hbb492d17),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51e591),
	.w1(32'h39cf100d),
	.w2(32'h39d8bbd3),
	.w3(32'hbb389294),
	.w4(32'h3ab12eb6),
	.w5(32'h3b02beb9),
	.w6(32'hbb91df69),
	.w7(32'hb9f7e32c),
	.w8(32'h3a0d26cb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20651c),
	.w1(32'h3996b193),
	.w2(32'hbb1d4330),
	.w3(32'h3a0ecf22),
	.w4(32'h3ada1177),
	.w5(32'hbae0382b),
	.w6(32'hb99dc071),
	.w7(32'h3a5c586d),
	.w8(32'hbb0e9ea8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a400478),
	.w1(32'h3a7276fe),
	.w2(32'h390bd001),
	.w3(32'h3a3c3188),
	.w4(32'h3a3e63a9),
	.w5(32'h39862ff0),
	.w6(32'h3990a5df),
	.w7(32'h3a180045),
	.w8(32'h39b18e74),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980f3f2),
	.w1(32'h3a31619b),
	.w2(32'hbaf283fe),
	.w3(32'h3affe8f1),
	.w4(32'h3b0f13bd),
	.w5(32'hba032aab),
	.w6(32'h398cc318),
	.w7(32'h3a5c89a7),
	.w8(32'hbb30f3f0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e29d1f),
	.w1(32'h39638434),
	.w2(32'hbb38250e),
	.w3(32'h3a81f073),
	.w4(32'h3a6234bb),
	.w5(32'hbb1b33ee),
	.w6(32'h3944e45e),
	.w7(32'h3a0d2d49),
	.w8(32'hbb26f10c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8c9f8),
	.w1(32'h3ab1f606),
	.w2(32'hbad8152d),
	.w3(32'h3b06f66a),
	.w4(32'h3a30abfb),
	.w5(32'hbb4f5354),
	.w6(32'hbac487fb),
	.w7(32'hbb0d0010),
	.w8(32'hbbc17a8d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9099f99),
	.w1(32'h395ea468),
	.w2(32'h395fece1),
	.w3(32'hb8fa43ef),
	.w4(32'h398b4171),
	.w5(32'h39a7fb22),
	.w6(32'h396f8798),
	.w7(32'h39112972),
	.w8(32'h39939ac5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb6867),
	.w1(32'h38a88d47),
	.w2(32'hb82bbf84),
	.w3(32'h397d18f0),
	.w4(32'hb6e9ebf9),
	.w5(32'hb92f2308),
	.w6(32'h3851a152),
	.w7(32'hb706a8d1),
	.w8(32'hb74d8103),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7460a1),
	.w1(32'h3ad34bda),
	.w2(32'hbb624684),
	.w3(32'h3ab28350),
	.w4(32'h3b30dd20),
	.w5(32'hbafb11d4),
	.w6(32'hba890ef3),
	.w7(32'hb904adf8),
	.w8(32'hbb69d673),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ba2f7),
	.w1(32'hb981b6a0),
	.w2(32'hbba824cc),
	.w3(32'h3ab97bb1),
	.w4(32'h3a80d54e),
	.w5(32'hbba43089),
	.w6(32'hb992f107),
	.w7(32'hba97ba8d),
	.w8(32'hbbf0a650),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4117a4),
	.w1(32'hb9e27d62),
	.w2(32'hbb5586e9),
	.w3(32'h3a9fb1b9),
	.w4(32'h3ac32f37),
	.w5(32'hbb154b9b),
	.w6(32'hba72dd30),
	.w7(32'hb99ed338),
	.w8(32'hbb738e30),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5d0b3),
	.w1(32'hba6eb7e4),
	.w2(32'hbb290457),
	.w3(32'hb9d27fda),
	.w4(32'hbad68864),
	.w5(32'hbb3e15af),
	.w6(32'h3af22855),
	.w7(32'h38eee85b),
	.w8(32'hbaa69449),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8945922),
	.w1(32'hb8bf9713),
	.w2(32'hb976ffe3),
	.w3(32'hb91d99eb),
	.w4(32'hb8bf5797),
	.w5(32'hb8ac70b7),
	.w6(32'h3823d5de),
	.w7(32'hb8a0dab2),
	.w8(32'hb8ad9c18),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39419c59),
	.w1(32'hb96381c1),
	.w2(32'hba07dba4),
	.w3(32'h39d4e4b2),
	.w4(32'h37cfbd96),
	.w5(32'hba089edb),
	.w6(32'h39a9bdd8),
	.w7(32'hb846ca06),
	.w8(32'hb9e628c2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aa3dc),
	.w1(32'h3b3101f3),
	.w2(32'hbbd4f919),
	.w3(32'hba8b80d0),
	.w4(32'h39cd24a3),
	.w5(32'hbbb4d924),
	.w6(32'hba523a13),
	.w7(32'h39a9cd98),
	.w8(32'hbb85f693),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac07f2),
	.w1(32'h3af7781c),
	.w2(32'hbb31d94f),
	.w3(32'h3af5db85),
	.w4(32'h3a80199d),
	.w5(32'hbb46572f),
	.w6(32'h3aa8d7b5),
	.w7(32'hba341a02),
	.w8(32'hbbb0811a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11d24e),
	.w1(32'hba44c986),
	.w2(32'hbba9d06d),
	.w3(32'hba5f129d),
	.w4(32'hba42d5c2),
	.w5(32'hbb2fe289),
	.w6(32'hb90d9fb4),
	.w7(32'hba143ce9),
	.w8(32'hbb0c8ad6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1854c0),
	.w1(32'h3b05cdc6),
	.w2(32'h3a5098f7),
	.w3(32'h3a31983f),
	.w4(32'h3b194bfd),
	.w5(32'h3ad7e136),
	.w6(32'hbabb321b),
	.w7(32'h39d6ff90),
	.w8(32'h39f0fce0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacebf36),
	.w1(32'hbaa3fa82),
	.w2(32'hbb53f754),
	.w3(32'h399cb80b),
	.w4(32'h3a54ac66),
	.w5(32'hbb1599f2),
	.w6(32'hba701586),
	.w7(32'hb912d813),
	.w8(32'hbb5da0b6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eaf0d2),
	.w1(32'h391f1b0d),
	.w2(32'h38f0467b),
	.w3(32'hb8d32092),
	.w4(32'h393efd4c),
	.w5(32'h392da433),
	.w6(32'h3895ded2),
	.w7(32'h37da5008),
	.w8(32'h38ce8a47),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df9ef6),
	.w1(32'h396c4aa9),
	.w2(32'h39689487),
	.w3(32'h391c8474),
	.w4(32'h3989f66a),
	.w5(32'h3906c642),
	.w6(32'h39849549),
	.w7(32'h397b6dbf),
	.w8(32'h3942ea10),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4780f0),
	.w1(32'h392dd887),
	.w2(32'hb979b750),
	.w3(32'h3a3fe483),
	.w4(32'hb9b88ee6),
	.w5(32'hb9c5e031),
	.w6(32'h3943f36e),
	.w7(32'hb94388ab),
	.w8(32'hb9aad09f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388365f6),
	.w1(32'hb9952d96),
	.w2(32'hb91043a8),
	.w3(32'h3886241d),
	.w4(32'hb977a0a9),
	.w5(32'hb903f36d),
	.w6(32'hb904f06b),
	.w7(32'hb942e424),
	.w8(32'hb90eb39c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d1e64),
	.w1(32'hb8dba631),
	.w2(32'hbab626da),
	.w3(32'hb89e16ce),
	.w4(32'hb9a391e1),
	.w5(32'hba7d1b01),
	.w6(32'h38d43e53),
	.w7(32'hb9e1041f),
	.w8(32'hba55b8b8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d804d4),
	.w1(32'hbacb765d),
	.w2(32'hbba1fa23),
	.w3(32'h3acbf623),
	.w4(32'h39c234ac),
	.w5(32'hbb7d06e6),
	.w6(32'h3947f656),
	.w7(32'hb932bf35),
	.w8(32'hbba5f3ca),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3f2f4),
	.w1(32'hb99de5cd),
	.w2(32'hbb1eff3e),
	.w3(32'h398f2fde),
	.w4(32'h39fe826f),
	.w5(32'hbb35cfbd),
	.w6(32'hb995aa35),
	.w7(32'hb8a015a3),
	.w8(32'hbb4b7e3e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b83348),
	.w1(32'h39ebd01f),
	.w2(32'h3a4d8d13),
	.w3(32'h39211bf9),
	.w4(32'h39de14b5),
	.w5(32'h39bcef3a),
	.w6(32'h39cf1f7c),
	.w7(32'h39f0a921),
	.w8(32'h39cfa993),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af66eab),
	.w1(32'h3a4e75f2),
	.w2(32'hbbe26000),
	.w3(32'hb88423dc),
	.w4(32'h3abaee68),
	.w5(32'hbba40fc2),
	.w6(32'h3a58555c),
	.w7(32'h3a596cb6),
	.w8(32'hbb8855eb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b23982),
	.w1(32'hba3c4f57),
	.w2(32'hbb02170f),
	.w3(32'h3993771e),
	.w4(32'hba2d1370),
	.w5(32'hbaf1c941),
	.w6(32'hb99c8917),
	.w7(32'hbaa94986),
	.w8(32'hbb153f70),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8014f5e),
	.w1(32'hb9d9d733),
	.w2(32'hba1df962),
	.w3(32'hb8dbf6c7),
	.w4(32'hba36674a),
	.w5(32'hba3ba17b),
	.w6(32'h38196690),
	.w7(32'hba04cca0),
	.w8(32'hba2952d5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac34fb),
	.w1(32'h3a5c420e),
	.w2(32'hbb0615a7),
	.w3(32'h3a0b327f),
	.w4(32'h39d1a3d6),
	.w5(32'hbadb8e6b),
	.w6(32'h3a1c60c7),
	.w7(32'h39462f47),
	.w8(32'hbabe5990),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d365e),
	.w1(32'h3926d981),
	.w2(32'h3948a6e7),
	.w3(32'h388e8fdc),
	.w4(32'h39714cd5),
	.w5(32'h39320809),
	.w6(32'h391e4185),
	.w7(32'h379af3de),
	.w8(32'h38c8476d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d35a65),
	.w1(32'hb952aa3d),
	.w2(32'hb90dec1b),
	.w3(32'hb8bb710c),
	.w4(32'hb8bfd6de),
	.w5(32'hb8025046),
	.w6(32'hb81ee909),
	.w7(32'hb99ebae0),
	.w8(32'hb9b4166b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dea7fd),
	.w1(32'h3895a833),
	.w2(32'h388636ff),
	.w3(32'hb65049bd),
	.w4(32'h37ab97d0),
	.w5(32'h3706ceff),
	.w6(32'h38667cac),
	.w7(32'h387e870b),
	.w8(32'h38aba1fa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3821e8dd),
	.w1(32'hb7e7f590),
	.w2(32'h38776d5e),
	.w3(32'h3882df01),
	.w4(32'h39288ad2),
	.w5(32'h39340f84),
	.w6(32'hb891fd8c),
	.w7(32'hb8e2f6e3),
	.w8(32'h381a7d04),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a621c3d),
	.w1(32'h3aa9c463),
	.w2(32'hb914029e),
	.w3(32'h39c11841),
	.w4(32'h3a9462ef),
	.w5(32'h37fc2923),
	.w6(32'hba8c0573),
	.w7(32'hb7a25823),
	.w8(32'h38e938fd),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeec82),
	.w1(32'hbb81e882),
	.w2(32'hbbf3a43a),
	.w3(32'h38bbfc51),
	.w4(32'hbb369d67),
	.w5(32'hbbbbdeb2),
	.w6(32'hb94d7d88),
	.w7(32'hbb3a92af),
	.w8(32'hbbd37ef1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cadf6c),
	.w1(32'h36c860d1),
	.w2(32'hbb7b334b),
	.w3(32'h3af026c3),
	.w4(32'h3a5f88f6),
	.w5(32'hbb3dddd0),
	.w6(32'h3af65b8e),
	.w7(32'h3a4179d6),
	.w8(32'hbb297623),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804f21),
	.w1(32'hba95a773),
	.w2(32'hbb861c83),
	.w3(32'h3a80c61f),
	.w4(32'hba35e908),
	.w5(32'hbb3f413e),
	.w6(32'h39049d93),
	.w7(32'hbaa7ec83),
	.w8(32'hbb941220),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f03224),
	.w1(32'hb7930ac1),
	.w2(32'hb78d571a),
	.w3(32'hb8fd2649),
	.w4(32'h3797d4fe),
	.w5(32'h38410b89),
	.w6(32'hb820d489),
	.w7(32'h37b68990),
	.w8(32'h39189922),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2dbc7),
	.w1(32'hb8f0fee1),
	.w2(32'hb9134c75),
	.w3(32'h3985234a),
	.w4(32'hb8c7e773),
	.w5(32'hb8d63dfe),
	.w6(32'h392cbca5),
	.w7(32'hb6b07bda),
	.w8(32'hb8205fc3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1f1f8),
	.w1(32'h38ad5973),
	.w2(32'h385ec848),
	.w3(32'h38851ff0),
	.w4(32'h37414e33),
	.w5(32'h372e5331),
	.w6(32'h38bdf0f7),
	.w7(32'h382a4919),
	.w8(32'h38301ab9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d634b6),
	.w1(32'h3909b41e),
	.w2(32'h3879d600),
	.w3(32'h37da94f8),
	.w4(32'h38a1b906),
	.w5(32'h383dae65),
	.w6(32'h3920f09c),
	.w7(32'h38cec45e),
	.w8(32'h38d1b5b0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94967df),
	.w1(32'hba9bb166),
	.w2(32'hbb3da0cf),
	.w3(32'h3a73cbee),
	.w4(32'hb9e05ab6),
	.w5(32'hbae8d25b),
	.w6(32'h3a08c307),
	.w7(32'hba85ce8f),
	.w8(32'hbb305dc7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9977435),
	.w1(32'hb9fbb391),
	.w2(32'hb9b2c8e9),
	.w3(32'h38561f31),
	.w4(32'hb9ab6c46),
	.w5(32'hb9e48708),
	.w6(32'h38bab963),
	.w7(32'h390ab49e),
	.w8(32'hb80bc10a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b92f1),
	.w1(32'h3a7c71af),
	.w2(32'h39297c19),
	.w3(32'h3984097d),
	.w4(32'h3a672770),
	.w5(32'h39ea8be7),
	.w6(32'h39650436),
	.w7(32'h3a4ef5c1),
	.w8(32'h3a03222f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37022a),
	.w1(32'hb9cbccd4),
	.w2(32'hb9a5ed3a),
	.w3(32'hb9f0ffdc),
	.w4(32'hba31ceb1),
	.w5(32'hb978f1aa),
	.w6(32'hb83f7859),
	.w7(32'hb89b9473),
	.w8(32'h3938154e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73b5045),
	.w1(32'h393b3168),
	.w2(32'h389df6c8),
	.w3(32'hb84a9e7b),
	.w4(32'h38345a85),
	.w5(32'h388b785a),
	.w6(32'h38aff8a0),
	.w7(32'hb7dd16aa),
	.w8(32'h38e1d52e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a041269),
	.w1(32'h3980041b),
	.w2(32'hba7583ed),
	.w3(32'h3a4fe78b),
	.w4(32'h3aa8c633),
	.w5(32'hb9c19b69),
	.w6(32'h37942cc0),
	.w7(32'h39212519),
	.w8(32'hba6add36),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc3249),
	.w1(32'h38167258),
	.w2(32'hb8977162),
	.w3(32'h396bd9b0),
	.w4(32'h38bf62d8),
	.w5(32'h378fc9df),
	.w6(32'h3985448c),
	.w7(32'h3888276a),
	.w8(32'h388cfa9b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d3c9),
	.w1(32'hbb7b8311),
	.w2(32'hbbbbd6c1),
	.w3(32'hb94839dc),
	.w4(32'hbb519434),
	.w5(32'hbb29c478),
	.w6(32'hba80c213),
	.w7(32'hbb046228),
	.w8(32'hbb488590),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b38d3b),
	.w1(32'hb74f6a68),
	.w2(32'hb7b6d942),
	.w3(32'h38814da1),
	.w4(32'hb820fcf7),
	.w5(32'hb726f802),
	.w6(32'h38a1d058),
	.w7(32'hb84bbe7f),
	.w8(32'h375841b8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bd98b),
	.w1(32'h3b0d5fc5),
	.w2(32'h3a15551f),
	.w3(32'hb9a5e949),
	.w4(32'h3a903190),
	.w5(32'h3a2b0d35),
	.w6(32'hbb6a0ea1),
	.w7(32'h374df79f),
	.w8(32'h3ae1bf9a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule