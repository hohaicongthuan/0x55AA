module layer_10_featuremap_206(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a773b),
	.w1(32'h3bb3e909),
	.w2(32'h3be38368),
	.w3(32'h3a85dc83),
	.w4(32'h3ae1d21f),
	.w5(32'h3ad71c38),
	.w6(32'h3b9ee40c),
	.w7(32'h3b6952d2),
	.w8(32'h3aed0985),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b49a1),
	.w1(32'hb98851c5),
	.w2(32'hb892e5d6),
	.w3(32'h3aece53b),
	.w4(32'hb9b7bc52),
	.w5(32'hb99b59c5),
	.w6(32'h389987ac),
	.w7(32'hb9aeb82d),
	.w8(32'h393cbc20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397034ec),
	.w1(32'h3a3006fc),
	.w2(32'h3b0182c8),
	.w3(32'h391ce509),
	.w4(32'hba0c8438),
	.w5(32'hb9eccab6),
	.w6(32'hba050ee8),
	.w7(32'hb94674e4),
	.w8(32'hb9d63e34),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cbc40),
	.w1(32'h39450ef5),
	.w2(32'hbad61e72),
	.w3(32'hb9c25729),
	.w4(32'h3aa18d1f),
	.w5(32'h3b0b3a77),
	.w6(32'hb97c9927),
	.w7(32'hba197462),
	.w8(32'h39311a72),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ca9f1),
	.w1(32'h3b3fe54b),
	.w2(32'h3a9e3a59),
	.w3(32'h3a1c78f3),
	.w4(32'h3b81b618),
	.w5(32'h3a9c987c),
	.w6(32'h3b3705f5),
	.w7(32'h3affa916),
	.w8(32'h3afcc85b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f45b2),
	.w1(32'h3aa850b0),
	.w2(32'h390a37a0),
	.w3(32'hb885f227),
	.w4(32'h3ad51362),
	.w5(32'h392e5394),
	.w6(32'h3abb4745),
	.w7(32'h3a3d521c),
	.w8(32'h3aa54200),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b4d12),
	.w1(32'h3aa8896c),
	.w2(32'h3a956686),
	.w3(32'h3aa60dcd),
	.w4(32'h3ad83481),
	.w5(32'h3a715ad3),
	.w6(32'h3acb36a3),
	.w7(32'h3aa78955),
	.w8(32'h3ac96d9e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9942f4),
	.w1(32'h39d3beba),
	.w2(32'hb94438c7),
	.w3(32'h3a22bf3d),
	.w4(32'h398b4c24),
	.w5(32'hb7a11072),
	.w6(32'h3a78adf4),
	.w7(32'h39c280dc),
	.w8(32'h3906ef74),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39661fec),
	.w1(32'hb882d67d),
	.w2(32'hb944fa63),
	.w3(32'h39fa2247),
	.w4(32'hb979f71c),
	.w5(32'hba28ed30),
	.w6(32'h398b7106),
	.w7(32'h393e5ab1),
	.w8(32'hb8dc5ed6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba096c80),
	.w1(32'h3a3a7395),
	.w2(32'hb9aee2cb),
	.w3(32'hb9859227),
	.w4(32'h3a5c7993),
	.w5(32'h39a7da16),
	.w6(32'h38b79c48),
	.w7(32'h38389fda),
	.w8(32'h3ac30b5b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f1c52),
	.w1(32'hb81cc9ef),
	.w2(32'h389bfcd7),
	.w3(32'h3ad55d48),
	.w4(32'h39a447a8),
	.w5(32'h3ae5a179),
	.w6(32'hbaeaa09f),
	.w7(32'hbaeafa51),
	.w8(32'hbab1ee1c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6949e5),
	.w1(32'h3a0808b7),
	.w2(32'hba132d36),
	.w3(32'h39f6180b),
	.w4(32'hba08624b),
	.w5(32'hba8ba97f),
	.w6(32'hb8c417bb),
	.w7(32'h3a8b497c),
	.w8(32'h3ac123fc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4d696),
	.w1(32'hba30d2cb),
	.w2(32'hb714c282),
	.w3(32'hb9d964e2),
	.w4(32'hb95e43d4),
	.w5(32'h395ebe01),
	.w6(32'hba48d7ec),
	.w7(32'hba543e78),
	.w8(32'hba7ffe2f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ab45f),
	.w1(32'hba883e39),
	.w2(32'hba55341c),
	.w3(32'h39743b8a),
	.w4(32'hbaae432f),
	.w5(32'hbaa58888),
	.w6(32'h379b4ae4),
	.w7(32'hba6da96f),
	.w8(32'hba89879b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12279),
	.w1(32'h3b02290d),
	.w2(32'h38159b7d),
	.w3(32'hba4921a9),
	.w4(32'h3b1f2a7e),
	.w5(32'hb9c571fd),
	.w6(32'h3a1a3ad5),
	.w7(32'h3b2b9987),
	.w8(32'h3b14873c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa922f9),
	.w1(32'h3a02ea7b),
	.w2(32'hb91782b6),
	.w3(32'hbac0bed5),
	.w4(32'h3a36fa9d),
	.w5(32'h39bcd3d3),
	.w6(32'h3a42dfd6),
	.w7(32'h3a35311b),
	.w8(32'h3a3a0668),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a73bc),
	.w1(32'h3aedce86),
	.w2(32'h3b34b8d2),
	.w3(32'h3a285f5d),
	.w4(32'hb922070b),
	.w5(32'hba0bcde4),
	.w6(32'h3a588f57),
	.w7(32'h3a6c3f4c),
	.w8(32'h3977a57c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8d5d0),
	.w1(32'h3a2564fb),
	.w2(32'h3a2faba4),
	.w3(32'h39470bc1),
	.w4(32'h3a1d23ec),
	.w5(32'h3a33bd9c),
	.w6(32'h39f51207),
	.w7(32'h3a96f0d9),
	.w8(32'h3a0867fd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e41d0),
	.w1(32'hb99f30bb),
	.w2(32'h391f6d2f),
	.w3(32'h3a78c80e),
	.w4(32'hb9a61b89),
	.w5(32'hb9c23f32),
	.w6(32'hb9bcfc87),
	.w7(32'h39606eb1),
	.w8(32'hb84a68aa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0c8a5),
	.w1(32'hb866ec83),
	.w2(32'hb971b6f2),
	.w3(32'hb9e97b31),
	.w4(32'hba05b715),
	.w5(32'hba396517),
	.w6(32'hb7fcd05b),
	.w7(32'hb8cfcddb),
	.w8(32'hb9a2b7a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3869e9),
	.w1(32'hba044433),
	.w2(32'hba992c57),
	.w3(32'hb9934dd0),
	.w4(32'hb9bcd7d1),
	.w5(32'hba1fe233),
	.w6(32'hba0e7135),
	.w7(32'hba052747),
	.w8(32'hb9d7f1ec),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ac9f5),
	.w1(32'h3ae5426f),
	.w2(32'h3be22c2d),
	.w3(32'h39153d35),
	.w4(32'h3a94c4af),
	.w5(32'h39a6efeb),
	.w6(32'h3a9d3b12),
	.w7(32'hbaeed12e),
	.w8(32'hbb3ea6be),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bfe46),
	.w1(32'hbadcfaf8),
	.w2(32'hb9d75a7b),
	.w3(32'hb9ca24f7),
	.w4(32'hba4edf42),
	.w5(32'hb99e074c),
	.w6(32'hba2fa379),
	.w7(32'h3a00df8e),
	.w8(32'hb8a47800),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39829097),
	.w1(32'h3a4447f4),
	.w2(32'h3a131ba1),
	.w3(32'h3a402e2d),
	.w4(32'h3a1869a5),
	.w5(32'h39be4d27),
	.w6(32'h3a87be98),
	.w7(32'h3a02bd3a),
	.w8(32'h39141038),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc278f),
	.w1(32'hbabad651),
	.w2(32'hbb0671bb),
	.w3(32'h3a1af3da),
	.w4(32'hba8163eb),
	.w5(32'hb973b0dc),
	.w6(32'hbae6422f),
	.w7(32'hba85a6c8),
	.w8(32'hba6b8f4e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082f74),
	.w1(32'hba359924),
	.w2(32'h3a37cc6c),
	.w3(32'h398bbd32),
	.w4(32'hbaa10789),
	.w5(32'hba8de729),
	.w6(32'h383f6d3f),
	.w7(32'h3a154185),
	.w8(32'h3a18227d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aded96),
	.w1(32'hb9c80e7d),
	.w2(32'hb9d2a5ac),
	.w3(32'hba8e19d0),
	.w4(32'hba20313b),
	.w5(32'hba624be1),
	.w6(32'hb9c92b8e),
	.w7(32'hb9d88eb6),
	.w8(32'hb992ff7d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e4eb5),
	.w1(32'h3987fb4b),
	.w2(32'hba85b35f),
	.w3(32'hb9d0f26e),
	.w4(32'hb884d2fb),
	.w5(32'h39e877a6),
	.w6(32'hba4cf69b),
	.w7(32'hb88985b7),
	.w8(32'hba0e6644),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990fcc4),
	.w1(32'hbb3e7051),
	.w2(32'hbb2851f5),
	.w3(32'h397883de),
	.w4(32'hbb3236dd),
	.w5(32'hbb00fe1b),
	.w6(32'hbb12eb9d),
	.w7(32'hbb23df76),
	.w8(32'hba412af7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9081427),
	.w1(32'hb8c4caba),
	.w2(32'h3a91e4c9),
	.w3(32'h3903d5ef),
	.w4(32'hbaafb683),
	.w5(32'hb8778a02),
	.w6(32'hba126e3e),
	.w7(32'hb8cc2069),
	.w8(32'h3930d2b4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e46c3c),
	.w1(32'hba016d43),
	.w2(32'hba57825d),
	.w3(32'h39e337b6),
	.w4(32'hb98ee183),
	.w5(32'hba38c68d),
	.w6(32'hb9bcdc39),
	.w7(32'hba223313),
	.w8(32'hb9d10f7b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba347486),
	.w1(32'hb9222dd5),
	.w2(32'h381534cc),
	.w3(32'hb9e1a2c8),
	.w4(32'h387623cf),
	.w5(32'hb8ee8d64),
	.w6(32'hb9b86267),
	.w7(32'hb9d503da),
	.w8(32'hb9c9f970),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8551d7c),
	.w1(32'h3a8a6854),
	.w2(32'hba180f39),
	.w3(32'h38fac776),
	.w4(32'h3a1e5b8f),
	.w5(32'hbac4920a),
	.w6(32'h3aadc3c7),
	.w7(32'hba07fe7c),
	.w8(32'hbaa6fd5b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac180ae),
	.w1(32'hba597ef9),
	.w2(32'hba6951b4),
	.w3(32'hbafdfe15),
	.w4(32'hbadd3cf1),
	.w5(32'hbb0a1ad9),
	.w6(32'hb98c48bd),
	.w7(32'hba726446),
	.w8(32'hbaa2a349),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c0255),
	.w1(32'hb9680bb0),
	.w2(32'hb9d49176),
	.w3(32'hba2da252),
	.w4(32'h391cdb87),
	.w5(32'hb95716c4),
	.w6(32'hb9bf0453),
	.w7(32'h38570d79),
	.w8(32'h3a369b7f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b3030),
	.w1(32'hba013ab6),
	.w2(32'hb9883aa6),
	.w3(32'h3a82d033),
	.w4(32'hba0f6c81),
	.w5(32'hba4f86b6),
	.w6(32'hba5a8826),
	.w7(32'hba38d2fb),
	.w8(32'hba4a17ec),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac36140),
	.w1(32'hb9584369),
	.w2(32'hb9d030b0),
	.w3(32'hba97b72a),
	.w4(32'h3a0cc738),
	.w5(32'h39946231),
	.w6(32'hba77244b),
	.w7(32'h388e8a6c),
	.w8(32'h38e1d746),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1880bc),
	.w1(32'h3a4600d9),
	.w2(32'h3a9740ef),
	.w3(32'h382ced5a),
	.w4(32'h39882d43),
	.w5(32'h3982edce),
	.w6(32'h39ff3a9a),
	.w7(32'h3999a53c),
	.w8(32'h39ba9e63),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947222),
	.w1(32'h3a6ac6db),
	.w2(32'h3a24fef8),
	.w3(32'h3a1f6bee),
	.w4(32'h3a28dd8c),
	.w5(32'h399a1d16),
	.w6(32'h3a94ec46),
	.w7(32'h39992512),
	.w8(32'hb8c45484),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d369),
	.w1(32'h39aa228e),
	.w2(32'h39e5da09),
	.w3(32'h3a32a114),
	.w4(32'h3a001b44),
	.w5(32'h394419ae),
	.w6(32'h39d3c765),
	.w7(32'h399d86bc),
	.w8(32'h392925a5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c6c194),
	.w1(32'h39116a80),
	.w2(32'h39bae56f),
	.w3(32'h390b9605),
	.w4(32'hb9c581ee),
	.w5(32'hb84acee2),
	.w6(32'h39c5104d),
	.w7(32'h3995c700),
	.w8(32'hb9f1cc8e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a50a8),
	.w1(32'hba223372),
	.w2(32'hba174d74),
	.w3(32'hb9debbfe),
	.w4(32'hbab1ba5c),
	.w5(32'hba4a41f9),
	.w6(32'hba786a25),
	.w7(32'hb9e22b2b),
	.w8(32'hbaac4405),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d335c),
	.w1(32'h384f0d7d),
	.w2(32'h3a1248a9),
	.w3(32'hba88e296),
	.w4(32'h38e05885),
	.w5(32'h3a300f7b),
	.w6(32'hb9b6f788),
	.w7(32'hb8cc7a00),
	.w8(32'h39191c72),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ec171),
	.w1(32'h3afbac3b),
	.w2(32'h395e55f0),
	.w3(32'h3a833efa),
	.w4(32'h3b206dec),
	.w5(32'h3ab53587),
	.w6(32'h3ae14906),
	.w7(32'h3a9e307b),
	.w8(32'h3b3e6b2e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b267545),
	.w1(32'h39be9f16),
	.w2(32'h3ad9f739),
	.w3(32'h3b28dfa5),
	.w4(32'hb92140c5),
	.w5(32'h3a3d5d4c),
	.w6(32'h396de168),
	.w7(32'hb9af4794),
	.w8(32'hba9130ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919ff86),
	.w1(32'h3a381c57),
	.w2(32'h3a013f21),
	.w3(32'h3aec3c4f),
	.w4(32'h3acdd23c),
	.w5(32'h3aa4e478),
	.w6(32'h3a4bb656),
	.w7(32'hb75d63bc),
	.w8(32'h398fb13a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62a4c6),
	.w1(32'h3b207d6e),
	.w2(32'h39742861),
	.w3(32'h3aaa4def),
	.w4(32'h3b3e0c26),
	.w5(32'h3ae42946),
	.w6(32'h3b0d877d),
	.w7(32'h3b8074f7),
	.w8(32'h3b8751fd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa2758),
	.w1(32'hb9d5edf4),
	.w2(32'h37d473e5),
	.w3(32'h3a6090b2),
	.w4(32'hba9aa525),
	.w5(32'hba66932f),
	.w6(32'hb9cfbc43),
	.w7(32'hb9caa4cc),
	.w8(32'hba64712d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2519e),
	.w1(32'hb9025ca5),
	.w2(32'h3a532b7c),
	.w3(32'hba51f102),
	.w4(32'hb98cf809),
	.w5(32'h399ca055),
	.w6(32'hba103ffc),
	.w7(32'hb97a2f4a),
	.w8(32'hb87b737a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7eba5),
	.w1(32'h3783672b),
	.w2(32'hba1c7d16),
	.w3(32'h3a342650),
	.w4(32'hb82433ee),
	.w5(32'hba096be7),
	.w6(32'h3a11b78c),
	.w7(32'hb9917f4e),
	.w8(32'hb9ebcf15),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba261588),
	.w1(32'h3a64761b),
	.w2(32'h38941560),
	.w3(32'hb949d5d5),
	.w4(32'h3a60d276),
	.w5(32'h3a5df393),
	.w6(32'hb8b15434),
	.w7(32'hb92dbcc1),
	.w8(32'h39b2ce78),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f95313),
	.w1(32'h3b318e20),
	.w2(32'hbac0ff2a),
	.w3(32'h3a0a1491),
	.w4(32'h3af18cc3),
	.w5(32'h3b43d1a6),
	.w6(32'h3b624b86),
	.w7(32'h3b87c4d8),
	.w8(32'h3b113f23),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa59a0),
	.w1(32'hb97623b5),
	.w2(32'hba9e5a93),
	.w3(32'h3b2dd3ab),
	.w4(32'hb90bfa29),
	.w5(32'hba9cf8bd),
	.w6(32'h39e0bd36),
	.w7(32'hb9fdf14c),
	.w8(32'hb93a7bac),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52faaf),
	.w1(32'h3ad8a74b),
	.w2(32'h3a25ce69),
	.w3(32'hb8612053),
	.w4(32'h3b80252f),
	.w5(32'h3a16643d),
	.w6(32'h3abfb9b0),
	.w7(32'h3adf0112),
	.w8(32'h3a93dfc0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88fe86c),
	.w1(32'hba24e1a8),
	.w2(32'h39ac1e10),
	.w3(32'hba7fe528),
	.w4(32'hba562082),
	.w5(32'hb99c4d61),
	.w6(32'hba2121df),
	.w7(32'hb89487c4),
	.w8(32'hb930559d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f4819),
	.w1(32'hbb0ef9c5),
	.w2(32'hba838d9f),
	.w3(32'h36b76373),
	.w4(32'hbab6409f),
	.w5(32'hbae63f65),
	.w6(32'hbac94c80),
	.w7(32'hba9d7293),
	.w8(32'hba716c7b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace27fc),
	.w1(32'hbab74a8d),
	.w2(32'hbb0c059c),
	.w3(32'hbac0302e),
	.w4(32'hbb013722),
	.w5(32'hbb0fad07),
	.w6(32'hbaa7d87a),
	.w7(32'hbb04d489),
	.w8(32'hbb060633),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332a90),
	.w1(32'h3b2c6cf3),
	.w2(32'hba428554),
	.w3(32'hbaca7579),
	.w4(32'h3b4e2098),
	.w5(32'h39fabec0),
	.w6(32'h3a577145),
	.w7(32'hb9cdad23),
	.w8(32'h3a8996fe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3f5d9),
	.w1(32'h399aa209),
	.w2(32'h3a2f83c2),
	.w3(32'hbaa8ac16),
	.w4(32'hb97ad5c2),
	.w5(32'h3958e5b9),
	.w6(32'h39e2a650),
	.w7(32'h38f94d6c),
	.w8(32'h392ffdcf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a4cd7),
	.w1(32'h3a3b63af),
	.w2(32'h3a2c2926),
	.w3(32'h3a73944b),
	.w4(32'h3a0b2463),
	.w5(32'h39a41ecb),
	.w6(32'h3a70bf98),
	.w7(32'h3a067a2d),
	.w8(32'h388885c2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b8e02),
	.w1(32'hb9c0e01b),
	.w2(32'h3a67fdf6),
	.w3(32'h3a1a4f13),
	.w4(32'hba1b06cb),
	.w5(32'hb9b4b60d),
	.w6(32'hb9ff75ee),
	.w7(32'h39809f40),
	.w8(32'h39118eed),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aeb64),
	.w1(32'hb9bc88ad),
	.w2(32'h36f9b953),
	.w3(32'h3986eeb4),
	.w4(32'hba1c0a05),
	.w5(32'hba29f896),
	.w6(32'hb954a488),
	.w7(32'hb9eaff6e),
	.w8(32'hba62999b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba422a99),
	.w1(32'h3aa62af6),
	.w2(32'h3b1f5997),
	.w3(32'hb9fdb6e0),
	.w4(32'hba9233f1),
	.w5(32'hbb2efa72),
	.w6(32'h3ae37e41),
	.w7(32'hbb001fac),
	.w8(32'hbb8170e4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080772),
	.w1(32'h3a8c2cd6),
	.w2(32'h38906d3e),
	.w3(32'hbad9ec73),
	.w4(32'h3abf361e),
	.w5(32'h3a6acd8a),
	.w6(32'h3a409ee5),
	.w7(32'h3a083c94),
	.w8(32'h3af41860),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2463f),
	.w1(32'hba45e822),
	.w2(32'hb9abe3a7),
	.w3(32'h3ada3c57),
	.w4(32'hb9ac5203),
	.w5(32'hb91e954f),
	.w6(32'hba013a3d),
	.w7(32'hb972debe),
	.w8(32'hb7aad9c3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b91cb),
	.w1(32'hbac700b0),
	.w2(32'hbadfb158),
	.w3(32'h394fa311),
	.w4(32'hb97a400e),
	.w5(32'h39baf957),
	.w6(32'hbac331d0),
	.w7(32'hbad094d0),
	.w8(32'hba8d2493),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dc91d),
	.w1(32'h3a0fbdf0),
	.w2(32'h3ad4df59),
	.w3(32'hba988ca8),
	.w4(32'hb9ee9f18),
	.w5(32'h36722df8),
	.w6(32'hb5a59fc1),
	.w7(32'h39e891e1),
	.w8(32'hb9178c55),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd8e27),
	.w1(32'h388414e4),
	.w2(32'hba928067),
	.w3(32'hb8ee48a5),
	.w4(32'h39e41465),
	.w5(32'hba446da3),
	.w6(32'h3a0ad30d),
	.w7(32'hb91ae632),
	.w8(32'hb9e6cb25),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf516),
	.w1(32'h39fbb16a),
	.w2(32'hba54451e),
	.w3(32'hb9e1560f),
	.w4(32'h3a6e2d95),
	.w5(32'h3816dd21),
	.w6(32'h3a92a723),
	.w7(32'h3a3ec1ab),
	.w8(32'h3a04995d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a16f),
	.w1(32'h3a54dd71),
	.w2(32'hba675ef6),
	.w3(32'h3a5aac23),
	.w4(32'h3abab604),
	.w5(32'h3a95b93a),
	.w6(32'hb998ad7e),
	.w7(32'hba4e73fa),
	.w8(32'h3a39e60a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f37407),
	.w1(32'h399cac40),
	.w2(32'h3a355e34),
	.w3(32'h39a21037),
	.w4(32'hb9534e1f),
	.w5(32'hb833d20a),
	.w6(32'h383d5333),
	.w7(32'h38f12588),
	.w8(32'hb9fb8605),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39117f73),
	.w1(32'h398c1155),
	.w2(32'h37f2f5fc),
	.w3(32'h3979bd21),
	.w4(32'h39c051b0),
	.w5(32'hb951e182),
	.w6(32'h3a00c7d4),
	.w7(32'h388bb316),
	.w8(32'hb8ff629a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388aa2bb),
	.w1(32'h3a3f6786),
	.w2(32'h3a0b1291),
	.w3(32'h39532704),
	.w4(32'h3a28d8c9),
	.w5(32'h39c253aa),
	.w6(32'h3a66b0fa),
	.w7(32'h3a087491),
	.w8(32'h3942d100),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965992c),
	.w1(32'hb9f27b13),
	.w2(32'hb9cbcd22),
	.w3(32'h3a1c475c),
	.w4(32'hb9838fc4),
	.w5(32'hb9909041),
	.w6(32'hba213250),
	.w7(32'hba3ed897),
	.w8(32'hba3f2b34),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb2024),
	.w1(32'hba959505),
	.w2(32'hba9c60bb),
	.w3(32'hb7dd48df),
	.w4(32'hba66a3be),
	.w5(32'h3839c695),
	.w6(32'hba087ead),
	.w7(32'hb7999da4),
	.w8(32'hb94b5b9f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02edcd),
	.w1(32'hb9beaffd),
	.w2(32'hba9d55dc),
	.w3(32'h39c634fc),
	.w4(32'hbacc2463),
	.w5(32'hba536a2d),
	.w6(32'h3a0dc6f0),
	.w7(32'h3a949e56),
	.w8(32'hb9827127),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961c0e7),
	.w1(32'h39b80312),
	.w2(32'hb9f8e5a2),
	.w3(32'hbb369325),
	.w4(32'h3a324883),
	.w5(32'hb9608d8e),
	.w6(32'h3a8690b1),
	.w7(32'h38d1b7f8),
	.w8(32'h39a95c05),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc2d3c),
	.w1(32'hba9acaf4),
	.w2(32'h3a1ea627),
	.w3(32'h3a006f56),
	.w4(32'hbaecb3d2),
	.w5(32'hbab0e9de),
	.w6(32'hba531bfb),
	.w7(32'hba90234a),
	.w8(32'hbadf88fd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9e940),
	.w1(32'hb7a8dceb),
	.w2(32'h3a85cf5f),
	.w3(32'hb8ee6d02),
	.w4(32'h3943d1d4),
	.w5(32'h3a840b08),
	.w6(32'h37c4e37b),
	.w7(32'h39e3d198),
	.w8(32'h3a43316d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b8777),
	.w1(32'hb9b191c2),
	.w2(32'hbab3c96c),
	.w3(32'h3a3fd4ca),
	.w4(32'hb640439a),
	.w5(32'hba51a39e),
	.w6(32'hb96c5fbc),
	.w7(32'hba603567),
	.w8(32'hba467ed5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba893ca7),
	.w1(32'hba035490),
	.w2(32'hbad3adb0),
	.w3(32'hb9f06b15),
	.w4(32'hba6a0a88),
	.w5(32'hbaed6fae),
	.w6(32'hb8abcb31),
	.w7(32'hba39743b),
	.w8(32'hba691e54),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b5b9),
	.w1(32'hb92ab841),
	.w2(32'hb9c2003f),
	.w3(32'hbabf89ce),
	.w4(32'hb9c16bd3),
	.w5(32'hba278460),
	.w6(32'h3902fdab),
	.w7(32'hb9a2246c),
	.w8(32'h3970a2ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d14fa6),
	.w1(32'hba8876f8),
	.w2(32'hba30f13d),
	.w3(32'hb9aee662),
	.w4(32'hbabaaee3),
	.w5(32'hbaa4ef72),
	.w6(32'hba96e23a),
	.w7(32'hba93bde4),
	.w8(32'hbaabe16b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f4dbb),
	.w1(32'h395e9d17),
	.w2(32'h3a91973f),
	.w3(32'hba5bedae),
	.w4(32'hba2fb62d),
	.w5(32'hb9897fb6),
	.w6(32'h399b8e68),
	.w7(32'h3933dbf1),
	.w8(32'h393a9434),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c98e2),
	.w1(32'h38a924b9),
	.w2(32'h3a977a24),
	.w3(32'h3a064984),
	.w4(32'hb90373ed),
	.w5(32'h3a4c2b2e),
	.w6(32'h3a569c07),
	.w7(32'h3a3e9b2b),
	.w8(32'h3a44c985),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399685db),
	.w1(32'hba37513e),
	.w2(32'h392b7c24),
	.w3(32'hb828d5cb),
	.w4(32'hba8adb49),
	.w5(32'hba4696d1),
	.w6(32'hba822947),
	.w7(32'hba8de911),
	.w8(32'hba9bedcf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a844f),
	.w1(32'hba4fa970),
	.w2(32'hb9d0ea4e),
	.w3(32'hba88a310),
	.w4(32'hbae4271e),
	.w5(32'hba76d7a5),
	.w6(32'hba2dc666),
	.w7(32'hba06f6ce),
	.w8(32'hbaaebfc7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa96820),
	.w1(32'hb9ae34f4),
	.w2(32'hba675c86),
	.w3(32'hbb082523),
	.w4(32'hb953f058),
	.w5(32'hb9ddd99c),
	.w6(32'hb95fdf7c),
	.w7(32'hb9e72a85),
	.w8(32'hb9983091),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba127803),
	.w1(32'hba30873f),
	.w2(32'hb9ba121c),
	.w3(32'hb907bb39),
	.w4(32'hba34148f),
	.w5(32'hba44d0f6),
	.w6(32'hb9f37bd5),
	.w7(32'h38e6a592),
	.w8(32'h392e1411),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2ded0),
	.w1(32'hb972e8a8),
	.w2(32'hba522a44),
	.w3(32'hb97506d5),
	.w4(32'h38829f9f),
	.w5(32'hb9f2cf22),
	.w6(32'hb8c400c1),
	.w7(32'hb93f6cd6),
	.w8(32'hb9fb7f73),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a5c8b),
	.w1(32'hb997c782),
	.w2(32'hba16c5c6),
	.w3(32'hb9213997),
	.w4(32'hb7eeffbe),
	.w5(32'hb9a935af),
	.w6(32'hba2d13c8),
	.w7(32'hba8938de),
	.w8(32'hba0c24e8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa9395),
	.w1(32'h3988c8c4),
	.w2(32'h39300320),
	.w3(32'h38554c51),
	.w4(32'h39ace890),
	.w5(32'h38515cf3),
	.w6(32'hb81315ee),
	.w7(32'h39efeaac),
	.w8(32'h3a7f81be),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f4ecd),
	.w1(32'hbad5be07),
	.w2(32'hba859505),
	.w3(32'h3a34cdd9),
	.w4(32'hbb1fc08d),
	.w5(32'hbb1b8a1e),
	.w6(32'hba67e22c),
	.w7(32'hba558d2c),
	.w8(32'hb9b7f0d3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39e90b),
	.w1(32'hbacccb86),
	.w2(32'hbb330aeb),
	.w3(32'hba933f78),
	.w4(32'hbabdc667),
	.w5(32'hbb13a6fe),
	.w6(32'hba6e5cb1),
	.w7(32'hbaa7aca2),
	.w8(32'hba2a917a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f4072),
	.w1(32'h38c6afec),
	.w2(32'h3ac1d3f9),
	.w3(32'hba1aabe8),
	.w4(32'hb784b97d),
	.w5(32'hb9036b8a),
	.w6(32'hb937472d),
	.w7(32'h399cf266),
	.w8(32'hb73fae47),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09101a),
	.w1(32'h3ae62dcf),
	.w2(32'h3b179f0a),
	.w3(32'h35ea6a87),
	.w4(32'h3adde3be),
	.w5(32'hba52ebf2),
	.w6(32'h3b2181f3),
	.w7(32'h3ac2d02f),
	.w8(32'h3aa8fd62),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2607e4),
	.w1(32'hba7f5e9a),
	.w2(32'h3a8de59c),
	.w3(32'hba358b9b),
	.w4(32'hba5e4637),
	.w5(32'h3a1b486a),
	.w6(32'hba71c02f),
	.w7(32'h3a1d00cd),
	.w8(32'h3886c991),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba383a57),
	.w1(32'hb9403874),
	.w2(32'hba93792c),
	.w3(32'hb9d8a28c),
	.w4(32'hba975944),
	.w5(32'hba2e37c5),
	.w6(32'hb7d7c472),
	.w7(32'hbaa0ecff),
	.w8(32'hbabafbcd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bdf74f),
	.w1(32'hba3f238a),
	.w2(32'hb8ab579f),
	.w3(32'h3a07af9c),
	.w4(32'hba8b7f6a),
	.w5(32'hbad3daeb),
	.w6(32'h39522cf4),
	.w7(32'hb9c90a1f),
	.w8(32'hbaba7828),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f6c7),
	.w1(32'hbad9c913),
	.w2(32'hbb1c146d),
	.w3(32'hbad3cbcd),
	.w4(32'hbaae0cb4),
	.w5(32'hbad75208),
	.w6(32'hbab6b6b7),
	.w7(32'hba21fee2),
	.w8(32'hba122bae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab854d5),
	.w1(32'h3b14ac1e),
	.w2(32'hbae55f71),
	.w3(32'hba437a6d),
	.w4(32'h3b4b873c),
	.w5(32'hba5823cc),
	.w6(32'h3a94b3d9),
	.w7(32'hba190498),
	.w8(32'h3b1a6283),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8978e),
	.w1(32'h3b0336bd),
	.w2(32'h3a0cb1c5),
	.w3(32'hba8cec12),
	.w4(32'h3b8a5875),
	.w5(32'h3b72f41c),
	.w6(32'h3b5a224e),
	.w7(32'h39e6c60d),
	.w8(32'h3a849acd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574a3a),
	.w1(32'h39d12124),
	.w2(32'hba0fa682),
	.w3(32'h3a23b0dc),
	.w4(32'h3a94b639),
	.w5(32'hb98fa97a),
	.w6(32'h3ab7b245),
	.w7(32'h38bb588b),
	.w8(32'h39c357c7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ebcbad),
	.w1(32'h3a42a8f5),
	.w2(32'hb94675f6),
	.w3(32'h3a2ae10a),
	.w4(32'h3a50aeb0),
	.w5(32'hb9a45e9e),
	.w6(32'h3a4d2985),
	.w7(32'h39737d0d),
	.w8(32'h389c609d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5dd6d),
	.w1(32'h391f2bec),
	.w2(32'hba24b9b3),
	.w3(32'hb8e70017),
	.w4(32'h3a15bf84),
	.w5(32'hb97078c4),
	.w6(32'h3a2758f5),
	.w7(32'h38fc1924),
	.w8(32'h3952fb0b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9036029),
	.w1(32'h387b070d),
	.w2(32'h36bdbdce),
	.w3(32'h399a7d26),
	.w4(32'hba15c1e7),
	.w5(32'hba5fd169),
	.w6(32'hb88359e3),
	.w7(32'hb85423da),
	.w8(32'hb9500059),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dc5e1),
	.w1(32'h38a0f2e3),
	.w2(32'h3ad1fe55),
	.w3(32'hba179751),
	.w4(32'hba919331),
	.w5(32'hba89f7d8),
	.w6(32'hb998ebe1),
	.w7(32'hb9e83728),
	.w8(32'hba094b7a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a398155),
	.w1(32'hb9f8b5a2),
	.w2(32'hba727ac2),
	.w3(32'hba2c87ed),
	.w4(32'hb9b2f2b7),
	.w5(32'hba222ae5),
	.w6(32'hba4df0e0),
	.w7(32'hba6dc2c6),
	.w8(32'hba3cbf6f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d29b2),
	.w1(32'h39b2f40a),
	.w2(32'hb928f075),
	.w3(32'h38430a40),
	.w4(32'h3a2eb02c),
	.w5(32'hb8b0ec1d),
	.w6(32'h3a613d5c),
	.w7(32'h389ab216),
	.w8(32'h398d41bd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f3605),
	.w1(32'h3a19a34e),
	.w2(32'h3b1cd4b3),
	.w3(32'h39afc26e),
	.w4(32'h3891bd08),
	.w5(32'h3aa2fbc0),
	.w6(32'h39670105),
	.w7(32'h3a256a01),
	.w8(32'h3986c9d2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb972a),
	.w1(32'h3a7c5f03),
	.w2(32'h398784ff),
	.w3(32'h3b152121),
	.w4(32'h3a03adbc),
	.w5(32'h39fc9f74),
	.w6(32'h3a9e3779),
	.w7(32'h3a96e560),
	.w8(32'h3a2691fc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fdd3e),
	.w1(32'h3b13672e),
	.w2(32'h3b967b71),
	.w3(32'h3a8aa0e5),
	.w4(32'hba74ec40),
	.w5(32'h3ab84992),
	.w6(32'h3ae4b1cf),
	.w7(32'h3a979d62),
	.w8(32'hbaf095ae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8c60c),
	.w1(32'h3aca916e),
	.w2(32'h39b50887),
	.w3(32'h3ab39190),
	.w4(32'h3ab0318e),
	.w5(32'h3a74e22c),
	.w6(32'h3ab2da57),
	.w7(32'h3ab65289),
	.w8(32'h3aa94a67),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccb595),
	.w1(32'hb8937d64),
	.w2(32'h3a368090),
	.w3(32'h3a7e0f32),
	.w4(32'h3807794d),
	.w5(32'h3a83e7af),
	.w6(32'hba981585),
	.w7(32'hb945d9a6),
	.w8(32'hb8a0442f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10ada9),
	.w1(32'hb920459e),
	.w2(32'hb9084908),
	.w3(32'h3a80519e),
	.w4(32'h38fa309c),
	.w5(32'hb93c378f),
	.w6(32'h39b25570),
	.w7(32'hba5fa170),
	.w8(32'hba88f90e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e8c7f),
	.w1(32'h39c0d261),
	.w2(32'hb9b1d710),
	.w3(32'hb9c217f1),
	.w4(32'h3a500cad),
	.w5(32'hb9544b5a),
	.w6(32'h3a8c6633),
	.w7(32'hb9033f2a),
	.w8(32'h3991920a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a90f20),
	.w1(32'h39f88363),
	.w2(32'h39b3b6a3),
	.w3(32'h39fe6936),
	.w4(32'h3a09f066),
	.w5(32'h393b5304),
	.w6(32'h3a46e20b),
	.w7(32'h3964bc76),
	.w8(32'h394ebd7d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6f574),
	.w1(32'h399b49ed),
	.w2(32'hb83093a7),
	.w3(32'h3a20e557),
	.w4(32'h3a06d478),
	.w5(32'h37f57013),
	.w6(32'h3a299b0e),
	.w7(32'h37fe8e7d),
	.w8(32'h39855cbf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab6036),
	.w1(32'h399f581a),
	.w2(32'h3b347e76),
	.w3(32'h3a1b6f2a),
	.w4(32'hba1ee09a),
	.w5(32'hb97372b6),
	.w6(32'hba2f91ce),
	.w7(32'hbaeccc06),
	.w8(32'hbb097657),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59ea3d),
	.w1(32'h3ab3812b),
	.w2(32'h3a29e54f),
	.w3(32'h3a894844),
	.w4(32'h3ab67040),
	.w5(32'h3a7d2d89),
	.w6(32'h3a1273ee),
	.w7(32'h39fb8d7b),
	.w8(32'hb9713da4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a84f77),
	.w1(32'hb9991106),
	.w2(32'hba9ad173),
	.w3(32'hba1b8efb),
	.w4(32'h3a4a5d38),
	.w5(32'hbaa282f5),
	.w6(32'h3907d76f),
	.w7(32'hba3eff5c),
	.w8(32'hba59edaa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab86dc6),
	.w1(32'hb9f7a9c5),
	.w2(32'hba66f0c6),
	.w3(32'hb99c596c),
	.w4(32'hb9e31bb4),
	.w5(32'hba986e14),
	.w6(32'h3980bfc6),
	.w7(32'hb7a789e4),
	.w8(32'hb9218cc5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e51ab7),
	.w1(32'h3a2486d8),
	.w2(32'h39ff2561),
	.w3(32'h390c399d),
	.w4(32'h3a109528),
	.w5(32'h39b7602d),
	.w6(32'h3a817334),
	.w7(32'h39963345),
	.w8(32'h3874b4db),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963dfa9),
	.w1(32'h3b7eb1ea),
	.w2(32'h3bb3d999),
	.w3(32'h3a268a06),
	.w4(32'h3b09504b),
	.w5(32'hba2d9fdc),
	.w6(32'h3ba91eb9),
	.w7(32'h3b39d583),
	.w8(32'h3aa6bb4c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95ba26),
	.w1(32'h3a7f149d),
	.w2(32'hba0cc363),
	.w3(32'h3ad96a80),
	.w4(32'h3a2831e7),
	.w5(32'hbad006e2),
	.w6(32'h3b13f0f7),
	.w7(32'h39d67b06),
	.w8(32'h39c7dc57),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffc76c),
	.w1(32'hba86cf90),
	.w2(32'hbaf1049a),
	.w3(32'hba2058fb),
	.w4(32'hba782b0d),
	.w5(32'hbabd7264),
	.w6(32'hba3748cd),
	.w7(32'hbaae52c9),
	.w8(32'hba53e852),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819609),
	.w1(32'h39788f0c),
	.w2(32'h379eeb7c),
	.w3(32'hb9c5128a),
	.w4(32'h399951b7),
	.w5(32'hb902176d),
	.w6(32'h390e1772),
	.w7(32'h39ab4907),
	.w8(32'hb7b313e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933c85a),
	.w1(32'h3a517127),
	.w2(32'h3a399bb6),
	.w3(32'hb6b170d8),
	.w4(32'h3a6c3649),
	.w5(32'h3a129b71),
	.w6(32'h3a140082),
	.w7(32'h3a4d7f4f),
	.w8(32'h3a09a052),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a377b32),
	.w1(32'h39e5dd37),
	.w2(32'hb8d2553c),
	.w3(32'h3a150b28),
	.w4(32'h3a9d596f),
	.w5(32'h3a3a955f),
	.w6(32'h3842efd6),
	.w7(32'hb8baa343),
	.w8(32'hba325f7b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807ee02),
	.w1(32'h3a18d572),
	.w2(32'h39eefb4c),
	.w3(32'h3a0dc061),
	.w4(32'h3a5cc434),
	.w5(32'h3a189cca),
	.w6(32'h39e64559),
	.w7(32'h3a1c8b5c),
	.w8(32'h3a467d50),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a409881),
	.w1(32'h37d13704),
	.w2(32'hb99ffda3),
	.w3(32'h3a84a910),
	.w4(32'h3a0c8d1d),
	.w5(32'h3931535b),
	.w6(32'h395f50ba),
	.w7(32'h39cb34e7),
	.w8(32'h3a301cb9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ca228),
	.w1(32'hb9d2cc42),
	.w2(32'hb95f00aa),
	.w3(32'h3a2e6a4c),
	.w4(32'hb89fb8e6),
	.w5(32'h39431b70),
	.w6(32'hb91f7098),
	.w7(32'hba31817f),
	.w8(32'h389758c3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9301b5e),
	.w1(32'h3a140201),
	.w2(32'h39a8a374),
	.w3(32'h3976c3b0),
	.w4(32'h3a986340),
	.w5(32'h398a23a4),
	.w6(32'hb88ca463),
	.w7(32'h3a8bd82f),
	.w8(32'h39ef7e1d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2e3a2),
	.w1(32'h3a0ece18),
	.w2(32'h39fecd0d),
	.w3(32'hb9aa24b0),
	.w4(32'h3a61f77e),
	.w5(32'h3a550896),
	.w6(32'h3a038815),
	.w7(32'h3a0d7a76),
	.w8(32'h3a3bfc07),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e0b07),
	.w1(32'h3a3d61e8),
	.w2(32'h3a2abeb4),
	.w3(32'h3a27fc8c),
	.w4(32'h3aa4393e),
	.w5(32'h3a6ee15f),
	.w6(32'h3a242cd8),
	.w7(32'h3a8e9a14),
	.w8(32'h3a4b70a4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ce29a),
	.w1(32'h39933347),
	.w2(32'h399c3b94),
	.w3(32'h3aca814f),
	.w4(32'h39851c5a),
	.w5(32'h39107680),
	.w6(32'h37bdf67b),
	.w7(32'hb923c741),
	.w8(32'hb982f898),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38478a87),
	.w1(32'h382eb38a),
	.w2(32'hb87df87c),
	.w3(32'hb788546c),
	.w4(32'hb8a8d814),
	.w5(32'hb99302f5),
	.w6(32'h394689cf),
	.w7(32'h39c859de),
	.w8(32'h38f0e8f4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9298ed6),
	.w1(32'h3a18c88a),
	.w2(32'h384d2a07),
	.w3(32'hb92da6c5),
	.w4(32'h3a9e9370),
	.w5(32'h3a64af1b),
	.w6(32'h39e814fa),
	.w7(32'h3a09c238),
	.w8(32'h3a4783c1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bb65b),
	.w1(32'hba054cea),
	.w2(32'hb8c7b669),
	.w3(32'h3ac67838),
	.w4(32'hb940ef78),
	.w5(32'hb99cd788),
	.w6(32'hb9c82a2e),
	.w7(32'hba182cbe),
	.w8(32'h398e8566),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39154dd5),
	.w1(32'hb9602e0b),
	.w2(32'h3a498a12),
	.w3(32'hb9e71f27),
	.w4(32'h3a1232ee),
	.w5(32'h3a89f98a),
	.w6(32'hb91270be),
	.w7(32'hb980fae6),
	.w8(32'h39a7c710),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c69e41),
	.w1(32'h39817cd5),
	.w2(32'h39737eb6),
	.w3(32'h3a4555d8),
	.w4(32'h39abc41e),
	.w5(32'h3910d5b1),
	.w6(32'h3829631e),
	.w7(32'hb8e4bb02),
	.w8(32'hb97fbd9e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a62423),
	.w1(32'h399a4ba4),
	.w2(32'h39ecbe06),
	.w3(32'h38831cc7),
	.w4(32'h3905d165),
	.w5(32'h3896119e),
	.w6(32'h38fa9b9c),
	.w7(32'hb924c294),
	.w8(32'hb93e5eb7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab941a),
	.w1(32'h3a2d8869),
	.w2(32'h3ae1ed21),
	.w3(32'hb92758f7),
	.w4(32'h3a80ed3f),
	.w5(32'h3a98f104),
	.w6(32'hba18e7a0),
	.w7(32'hb98cea86),
	.w8(32'h3a50098a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a382c38),
	.w1(32'h3a0f381e),
	.w2(32'h39594ebf),
	.w3(32'h398ca034),
	.w4(32'h39c9d6a2),
	.w5(32'h39741bea),
	.w6(32'h3a08b5bb),
	.w7(32'h3a037ed6),
	.w8(32'h39b6112b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39606850),
	.w1(32'hb9637eb4),
	.w2(32'h383e9763),
	.w3(32'h390cd627),
	.w4(32'hb9bdc235),
	.w5(32'hba72f7fb),
	.w6(32'hb9d9888b),
	.w7(32'h392605b2),
	.w8(32'h39162a62),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dead0a),
	.w1(32'h3a1c9850),
	.w2(32'h39ada947),
	.w3(32'hba957fc2),
	.w4(32'h3a4a4e4e),
	.w5(32'h39e075f4),
	.w6(32'h3a315c70),
	.w7(32'h3a4f244b),
	.w8(32'h3a5fa2ba),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f37c),
	.w1(32'h39e5a51c),
	.w2(32'h39764776),
	.w3(32'h3a95ce05),
	.w4(32'h3a20e989),
	.w5(32'h394efa7e),
	.w6(32'h38b99955),
	.w7(32'h39cae16e),
	.w8(32'h3a0b8bc1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e5b86),
	.w1(32'h389509d8),
	.w2(32'hb914cff7),
	.w3(32'h3a4a86ce),
	.w4(32'hb806465f),
	.w5(32'hb9642f28),
	.w6(32'h38cf0065),
	.w7(32'h389cc89e),
	.w8(32'hb8dde515),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914bc4b),
	.w1(32'h39fc22fe),
	.w2(32'h37fadef3),
	.w3(32'hb955de9b),
	.w4(32'h3a21355b),
	.w5(32'h3a126c19),
	.w6(32'h3a192a0a),
	.w7(32'h39dbedc8),
	.w8(32'h39508be0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38142417),
	.w1(32'hbaa32ef8),
	.w2(32'hba0883f7),
	.w3(32'h39debd2a),
	.w4(32'h3a939f48),
	.w5(32'h3a785b6f),
	.w6(32'hb9acb331),
	.w7(32'hb9728406),
	.w8(32'h3a8fc52c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39595010),
	.w1(32'hba20ef71),
	.w2(32'hba8a0282),
	.w3(32'h3a64dea3),
	.w4(32'hba5413a6),
	.w5(32'hbae3a23e),
	.w6(32'hb8d5e8ff),
	.w7(32'h3993914d),
	.w8(32'h379089dd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba576161),
	.w1(32'h39bff913),
	.w2(32'h39b91e36),
	.w3(32'hba163a3e),
	.w4(32'h3a1bccd1),
	.w5(32'h3999ce99),
	.w6(32'h39b06a63),
	.w7(32'h39cced17),
	.w8(32'h382e428e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04d784),
	.w1(32'h39f520a0),
	.w2(32'h395fb2bb),
	.w3(32'h39857663),
	.w4(32'h398d742f),
	.w5(32'hb8f53732),
	.w6(32'hb8301703),
	.w7(32'hb998ecd7),
	.w8(32'h395323f8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6fa04),
	.w1(32'hba732251),
	.w2(32'hba04e585),
	.w3(32'h38a6998f),
	.w4(32'hb9af6756),
	.w5(32'hb9f16128),
	.w6(32'hba93af8b),
	.w7(32'hba934a57),
	.w8(32'hba1c41a6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8213e3),
	.w1(32'hb9314ebe),
	.w2(32'hb9886e95),
	.w3(32'hb998682a),
	.w4(32'hb771c1a4),
	.w5(32'hb8986935),
	.w6(32'hb9848c7d),
	.w7(32'hb9dbb98c),
	.w8(32'hba0f4144),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9773200),
	.w1(32'hba1dd832),
	.w2(32'hba30f516),
	.w3(32'hb90055f0),
	.w4(32'hba29ba65),
	.w5(32'hba119049),
	.w6(32'hba42d736),
	.w7(32'hba5cc42e),
	.w8(32'hba17fd19),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d645a6),
	.w1(32'h3952e200),
	.w2(32'hba07fa10),
	.w3(32'hba20f90c),
	.w4(32'h38e5f41a),
	.w5(32'hba602098),
	.w6(32'hb899a6b4),
	.w7(32'hb9c5c96f),
	.w8(32'hb90c8cf9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995f60d),
	.w1(32'h391d80f6),
	.w2(32'h394dc657),
	.w3(32'hba0eb849),
	.w4(32'hb93328c1),
	.w5(32'hb92e277b),
	.w6(32'h39394a71),
	.w7(32'h39c55a91),
	.w8(32'h39e0caf4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c59ea2),
	.w1(32'h39a207a7),
	.w2(32'hb6e4243b),
	.w3(32'hb9b3bcc4),
	.w4(32'h39d4ad3f),
	.w5(32'h390d1475),
	.w6(32'h39a1e83b),
	.w7(32'h39861fbc),
	.w8(32'h37b3a25c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1330c),
	.w1(32'h3896078e),
	.w2(32'hb8babcb4),
	.w3(32'h3823e726),
	.w4(32'h398c4b13),
	.w5(32'hb7d055f3),
	.w6(32'h3784b327),
	.w7(32'hb9699d94),
	.w8(32'hb9ea3987),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e5230),
	.w1(32'hb971db9c),
	.w2(32'hba449a4e),
	.w3(32'hb8d22502),
	.w4(32'hb98cb1a4),
	.w5(32'hba5480e5),
	.w6(32'hb994248e),
	.w7(32'hba3a9beb),
	.w8(32'hba6f72dc),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810435),
	.w1(32'h385e4e91),
	.w2(32'hb9c4d20e),
	.w3(32'hba9fd831),
	.w4(32'hb9e49e19),
	.w5(32'hba12fb65),
	.w6(32'h3a1fe455),
	.w7(32'hb6afa7f6),
	.w8(32'hba8a9bf4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba451b31),
	.w1(32'h3aa6d0db),
	.w2(32'h3a6a2145),
	.w3(32'hba83b31a),
	.w4(32'h3ae52e44),
	.w5(32'h3ac68012),
	.w6(32'h3a8e2e11),
	.w7(32'h3a696d5a),
	.w8(32'h3aae0674),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe8af8),
	.w1(32'hb9665bbd),
	.w2(32'hb9b535ab),
	.w3(32'h3b082a17),
	.w4(32'hb75e015e),
	.w5(32'hb98be3eb),
	.w6(32'hba117dd5),
	.w7(32'hba32bc97),
	.w8(32'hba3e9c21),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d26ee0),
	.w1(32'h3a469cf7),
	.w2(32'h3a5aa1c3),
	.w3(32'hb9a30aae),
	.w4(32'h3a593854),
	.w5(32'h39fd226f),
	.w6(32'h39d039ac),
	.w7(32'h3a4783a4),
	.w8(32'h3a08f33d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e316d),
	.w1(32'h3a19af77),
	.w2(32'h39c77d33),
	.w3(32'h3a495afc),
	.w4(32'h3a62e674),
	.w5(32'h39f9afe6),
	.w6(32'h3a2cd72d),
	.w7(32'h3a63fca9),
	.w8(32'h3a77d3da),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47b454),
	.w1(32'h3a149a19),
	.w2(32'h3a34f9d5),
	.w3(32'h3a7e0471),
	.w4(32'h3a2d03cb),
	.w5(32'h3a158ad2),
	.w6(32'h39f4131b),
	.w7(32'h39f4cc49),
	.w8(32'h39956688),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2758fd),
	.w1(32'h39fdf342),
	.w2(32'h3a027b53),
	.w3(32'h3a04fed5),
	.w4(32'h3a19bbe3),
	.w5(32'h3a003be6),
	.w6(32'h39acb1b8),
	.w7(32'h39e6c161),
	.w8(32'h39d7a99b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0faf52),
	.w1(32'h3a1d06be),
	.w2(32'h39d5de5a),
	.w3(32'h3a3df5be),
	.w4(32'h39a042ef),
	.w5(32'h3994659e),
	.w6(32'h3a045db3),
	.w7(32'h3a5179a5),
	.w8(32'h3975cdb3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f4ba08),
	.w1(32'hb9120402),
	.w2(32'h37f8e88a),
	.w3(32'h38b9e818),
	.w4(32'hb9782cc1),
	.w5(32'hb80d9136),
	.w6(32'h38c34155),
	.w7(32'hb9a30071),
	.w8(32'h390e7abd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f60af0),
	.w1(32'h38b0800e),
	.w2(32'hb6002af1),
	.w3(32'h38ffd022),
	.w4(32'hb71b71ed),
	.w5(32'hb9178a75),
	.w6(32'hb8c4a26c),
	.w7(32'hb9af6767),
	.w8(32'hb9dee8c9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb50e47d6),
	.w1(32'h39c0925c),
	.w2(32'h3804dee3),
	.w3(32'hb88e4057),
	.w4(32'h3a60e5f6),
	.w5(32'h3a6cfe0b),
	.w6(32'h3912d783),
	.w7(32'h391fb2cb),
	.w8(32'h3a5e924d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42cb0c),
	.w1(32'h399ddfcd),
	.w2(32'hb8d22e20),
	.w3(32'h3aca1ab1),
	.w4(32'h3a3c37c1),
	.w5(32'h39aa21a2),
	.w6(32'h3a116f8a),
	.w7(32'h3a18a726),
	.w8(32'h3a2ba40d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2aae6),
	.w1(32'h3952fd00),
	.w2(32'h398685db),
	.w3(32'h396e807f),
	.w4(32'h3a29461f),
	.w5(32'h3a1457ea),
	.w6(32'h39d64ad7),
	.w7(32'h3a575472),
	.w8(32'h3a4d85ee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8273ad),
	.w1(32'h3a10c704),
	.w2(32'h3a6b9b02),
	.w3(32'h3a9408d6),
	.w4(32'h3aa52d06),
	.w5(32'h3aaba1f1),
	.w6(32'hb7eda347),
	.w7(32'hbaa9d83a),
	.w8(32'hb8bef981),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b03a7e),
	.w1(32'hb98d332e),
	.w2(32'hba3a0cd0),
	.w3(32'h3a0db054),
	.w4(32'hba53996f),
	.w5(32'hbb04f525),
	.w6(32'hb9008e16),
	.w7(32'h3a218fd6),
	.w8(32'h3989cbad),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe2d16),
	.w1(32'hb9733cc6),
	.w2(32'hb9b952a9),
	.w3(32'hbaae5cfb),
	.w4(32'hb90527ef),
	.w5(32'hb9d7847d),
	.w6(32'hb99fe168),
	.w7(32'hb9f333cf),
	.w8(32'hba01c68f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9895845),
	.w1(32'h390d573e),
	.w2(32'h3953e16a),
	.w3(32'hb93ab384),
	.w4(32'h380f344c),
	.w5(32'hb72e698d),
	.w6(32'h3795cb97),
	.w7(32'hb8dabc9b),
	.w8(32'hb992f059),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e34257),
	.w1(32'h3a02e26f),
	.w2(32'h3a6d0f8b),
	.w3(32'hb983ab3c),
	.w4(32'h3a0d76ab),
	.w5(32'h39f9448b),
	.w6(32'hb99474d4),
	.w7(32'h38b94189),
	.w8(32'hb6969ae7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18c3fa),
	.w1(32'hb9f53b45),
	.w2(32'hbaa74106),
	.w3(32'h3a77fee3),
	.w4(32'hba95375c),
	.w5(32'hbab62d8c),
	.w6(32'h39c7a564),
	.w7(32'hba9ea7d3),
	.w8(32'hba165f8d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cedd0),
	.w1(32'h3a1c8090),
	.w2(32'h3931b046),
	.w3(32'hba81938c),
	.w4(32'h3a4c8660),
	.w5(32'h39c0d64f),
	.w6(32'h3966e3fa),
	.w7(32'h397aab03),
	.w8(32'h394d134c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac556f),
	.w1(32'h3a78b1e3),
	.w2(32'h3a8dc8ae),
	.w3(32'h39a59568),
	.w4(32'h3a9c5ca4),
	.w5(32'h3a91b4c4),
	.w6(32'h398edc19),
	.w7(32'h3a9a20cb),
	.w8(32'h39d330b1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9b0b7),
	.w1(32'h3a337e5d),
	.w2(32'h39ab77df),
	.w3(32'h3a4713a5),
	.w4(32'h3a283943),
	.w5(32'h394a4303),
	.w6(32'h39cc995c),
	.w7(32'h39eb735b),
	.w8(32'h3a566628),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ad8b3),
	.w1(32'hb95eefc9),
	.w2(32'h386367d2),
	.w3(32'h39a83b07),
	.w4(32'h38d3265c),
	.w5(32'hb91a4903),
	.w6(32'hb99eb6ab),
	.w7(32'hb93987f6),
	.w8(32'hba120903),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f9ce1e),
	.w1(32'hba2232fb),
	.w2(32'hba2be5c8),
	.w3(32'h38bb5253),
	.w4(32'hba249ae4),
	.w5(32'hba2ee2f6),
	.w6(32'hb9eb08ef),
	.w7(32'hb97459a9),
	.w8(32'h3781c797),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c75267),
	.w1(32'h3a0aa8c8),
	.w2(32'h39a08856),
	.w3(32'hb9d1e967),
	.w4(32'h3a81e014),
	.w5(32'h3a116fbe),
	.w6(32'hb9c3e692),
	.w7(32'h3a302c25),
	.w8(32'h3a01e030),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a600e71),
	.w1(32'h3a2954d9),
	.w2(32'h39b4a8db),
	.w3(32'h3a4e14fc),
	.w4(32'h3a820c66),
	.w5(32'h3a376c28),
	.w6(32'h39954bf9),
	.w7(32'h397e98ac),
	.w8(32'h3a08ee31),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a331abd),
	.w1(32'h3a1c2b9d),
	.w2(32'h3a13255b),
	.w3(32'h3a90db15),
	.w4(32'h3a4696c5),
	.w5(32'h39e0175e),
	.w6(32'h3a38a2e1),
	.w7(32'h3a3957eb),
	.w8(32'h3984d5b5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39dbc2),
	.w1(32'h3a19ec44),
	.w2(32'h39bba53e),
	.w3(32'h39f4460d),
	.w4(32'h3a2695f4),
	.w5(32'h3a366d91),
	.w6(32'h39d25289),
	.w7(32'h38ec6875),
	.w8(32'h3a0aa239),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a260f4e),
	.w1(32'h396eee78),
	.w2(32'h38df62ff),
	.w3(32'h3a87fe10),
	.w4(32'h3859fe17),
	.w5(32'h3899eac1),
	.w6(32'h399b1157),
	.w7(32'h39ab0ae0),
	.w8(32'hb814266b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb832c25e),
	.w1(32'h3a220ca3),
	.w2(32'hb997b6a7),
	.w3(32'hb8f6938c),
	.w4(32'h3a2380f0),
	.w5(32'h39bb6010),
	.w6(32'h3a597ad9),
	.w7(32'h398c92c6),
	.w8(32'hb7ba0014),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f18e4),
	.w1(32'h398ce4b0),
	.w2(32'h382e875c),
	.w3(32'hba25e5ae),
	.w4(32'h3a3240a5),
	.w5(32'h3a2e270a),
	.w6(32'h387d11a1),
	.w7(32'h38bd7219),
	.w8(32'h3a10d14a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08d1a1),
	.w1(32'h38958b36),
	.w2(32'hb8daa01a),
	.w3(32'h3a91f1b1),
	.w4(32'h39a7121d),
	.w5(32'h387b82e1),
	.w6(32'hb9b80226),
	.w7(32'hb8a318c3),
	.w8(32'h39920def),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a50347),
	.w1(32'h3750ad27),
	.w2(32'h38cdcd31),
	.w3(32'h39b824f2),
	.w4(32'h38dd8eee),
	.w5(32'hb92da392),
	.w6(32'h381c0693),
	.w7(32'h3a88594b),
	.w8(32'h3a2db49e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914d4b8),
	.w1(32'h39a24cfc),
	.w2(32'h3a0fe761),
	.w3(32'h38fee3ec),
	.w4(32'h399601a9),
	.w5(32'h3a3ffc62),
	.w6(32'h3a0c4e58),
	.w7(32'h3a1f6c90),
	.w8(32'h3a308e0c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f4eef),
	.w1(32'h3942289e),
	.w2(32'hb9afc107),
	.w3(32'h3a36a408),
	.w4(32'hb989093a),
	.w5(32'hba85a9d9),
	.w6(32'h39c50f02),
	.w7(32'h3a302f04),
	.w8(32'h3821f8ae),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd6fd6),
	.w1(32'h3a823705),
	.w2(32'h3a330a8f),
	.w3(32'hb9ee4c80),
	.w4(32'h3a625e4c),
	.w5(32'h3a31030e),
	.w6(32'h3a375c68),
	.w7(32'h3a0ea3ad),
	.w8(32'h39b18d6f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d67bd),
	.w1(32'h3a896a75),
	.w2(32'h3a787d7a),
	.w3(32'h3a019109),
	.w4(32'h3a41f7ad),
	.w5(32'h3a08f39e),
	.w6(32'h394d352d),
	.w7(32'h3a4ccf2a),
	.w8(32'h399dc3b6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a183324),
	.w1(32'h39d2e023),
	.w2(32'h39a663f8),
	.w3(32'h3a6b1bce),
	.w4(32'h3a081d7d),
	.w5(32'h39ab32a2),
	.w6(32'h3a03557d),
	.w7(32'h3a405e15),
	.w8(32'h3a723451),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48bfd4),
	.w1(32'h3a25f3b6),
	.w2(32'h3a0d024a),
	.w3(32'h3a3e0225),
	.w4(32'h3a237536),
	.w5(32'h39e2e94b),
	.w6(32'h3a06e073),
	.w7(32'h39e3af4f),
	.w8(32'h3946ad6c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a20e93),
	.w1(32'h39e67947),
	.w2(32'h3a04b072),
	.w3(32'h396b46dc),
	.w4(32'h39ef324c),
	.w5(32'h39cddba2),
	.w6(32'h3a08b9fe),
	.w7(32'h39d47217),
	.w8(32'h39459ef2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08deeb),
	.w1(32'h37f40924),
	.w2(32'hb941b919),
	.w3(32'h39ed56ae),
	.w4(32'h3977c790),
	.w5(32'hb836d21f),
	.w6(32'hb983a7f0),
	.w7(32'hba096b9a),
	.w8(32'hba201bb2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c93b4),
	.w1(32'h39bab3a7),
	.w2(32'h37f4834d),
	.w3(32'hb91eb788),
	.w4(32'h39cf1f2b),
	.w5(32'h38188402),
	.w6(32'hb90cfc2f),
	.w7(32'hb92b362a),
	.w8(32'h394988fb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e5ce3),
	.w1(32'hbab91c7f),
	.w2(32'h39cdb2bf),
	.w3(32'h38fc90a8),
	.w4(32'hba82eef0),
	.w5(32'hba208e78),
	.w6(32'hba9627f5),
	.w7(32'hbb18be80),
	.w8(32'hba6dece7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9997e85),
	.w1(32'hb8449a86),
	.w2(32'hb8ebd10a),
	.w3(32'hb8da3ccb),
	.w4(32'hb91cb122),
	.w5(32'hb9ad00f6),
	.w6(32'h37ad53fd),
	.w7(32'h36d99708),
	.w8(32'hb95961f8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98aa08c),
	.w1(32'h3a4ec1e8),
	.w2(32'h39c966cb),
	.w3(32'hb9ee5b29),
	.w4(32'h3a4cb0d2),
	.w5(32'h39dab1dc),
	.w6(32'h3a98e0d9),
	.w7(32'h3a6d64f9),
	.w8(32'h3a5c6e6d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22f3f7),
	.w1(32'hb920871a),
	.w2(32'hb7c9c291),
	.w3(32'h3a054559),
	.w4(32'hba0b7a24),
	.w5(32'hba720171),
	.w6(32'hb986c9d5),
	.w7(32'h3885b7c8),
	.w8(32'h393bdb61),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f283ee),
	.w1(32'h3a131521),
	.w2(32'h392babfa),
	.w3(32'hb9e385ba),
	.w4(32'h3a10a262),
	.w5(32'h39ab88bc),
	.w6(32'h3a07b4ba),
	.w7(32'h3a0240e8),
	.w8(32'h39404c7f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ec3d86),
	.w1(32'h39c53e0b),
	.w2(32'hb8939a85),
	.w3(32'h38ade9fd),
	.w4(32'hb93240d9),
	.w5(32'hba361075),
	.w6(32'h39d63e8d),
	.w7(32'h3a5a464a),
	.w8(32'hb818c255),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967f4dc),
	.w1(32'h3a0df507),
	.w2(32'h3a25d2dc),
	.w3(32'hb9dd125e),
	.w4(32'h3a5b96e1),
	.w5(32'h3a36cd36),
	.w6(32'h3936f20b),
	.w7(32'h399148ad),
	.w8(32'h39f27103),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4535e2),
	.w1(32'h389abafd),
	.w2(32'hb91e85dd),
	.w3(32'h3a5361aa),
	.w4(32'hb966f577),
	.w5(32'hba0c04e7),
	.w6(32'hb987b564),
	.w7(32'hb913547f),
	.w8(32'hb8cae546),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a36ff2),
	.w1(32'h3a49416f),
	.w2(32'h39a9d6dd),
	.w3(32'hb92e5fa5),
	.w4(32'h3a940cb5),
	.w5(32'h3a61a146),
	.w6(32'h39e02828),
	.w7(32'h3a19661d),
	.w8(32'h3a136f5b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c000fa),
	.w1(32'hb8aef023),
	.w2(32'h394daf73),
	.w3(32'h3a540a4c),
	.w4(32'hba1ea00f),
	.w5(32'hbaad4e70),
	.w6(32'h3a830af2),
	.w7(32'h3ae21385),
	.w8(32'h3a615787),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6820),
	.w1(32'h390576d6),
	.w2(32'h399bade0),
	.w3(32'hba3fc685),
	.w4(32'h3856167c),
	.w5(32'h38af1ff8),
	.w6(32'h3974bfbf),
	.w7(32'h3a01136e),
	.w8(32'h3a340d4f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986d834),
	.w1(32'hba1d65f7),
	.w2(32'h393f7550),
	.w3(32'h38c0c582),
	.w4(32'hba6f777c),
	.w5(32'hb99d3996),
	.w6(32'hba15051d),
	.w7(32'hba48f1b0),
	.w8(32'hba022700),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905a854),
	.w1(32'h39978041),
	.w2(32'h38729c0a),
	.w3(32'hb8250e94),
	.w4(32'h399af0ce),
	.w5(32'h39702830),
	.w6(32'h3992346e),
	.w7(32'h393eca3b),
	.w8(32'hb63a9986),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b860a6),
	.w1(32'h3a7a349f),
	.w2(32'h39fdbc39),
	.w3(32'h3920a3b9),
	.w4(32'h3a8895a1),
	.w5(32'h3a3022ed),
	.w6(32'h3a1f3150),
	.w7(32'h3a1be4c9),
	.w8(32'h3a7cc795),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a9f44),
	.w1(32'h3a2bfb3d),
	.w2(32'h39a796a2),
	.w3(32'h39ceb08d),
	.w4(32'h3a09c041),
	.w5(32'h39b22782),
	.w6(32'h39c45e54),
	.w7(32'h39eb93fe),
	.w8(32'h39be7141),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912f3c3),
	.w1(32'h39d181b4),
	.w2(32'h375f96c7),
	.w3(32'h391c0b23),
	.w4(32'h3a1f533a),
	.w5(32'h392e3a60),
	.w6(32'h3a15d8d7),
	.w7(32'h3a01a008),
	.w8(32'hb5bf24b7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a364e0),
	.w1(32'h39f7feee),
	.w2(32'hb8df82e7),
	.w3(32'h384b2e53),
	.w4(32'h3a39a58a),
	.w5(32'h39ce0fcb),
	.w6(32'h3a26c365),
	.w7(32'h3a8871de),
	.w8(32'h3a958a10),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7725),
	.w1(32'h39ce1572),
	.w2(32'h3955cbd2),
	.w3(32'h3a5e4cf7),
	.w4(32'h3a0e826d),
	.w5(32'h38bf090e),
	.w6(32'h39200a2a),
	.w7(32'h396cd62e),
	.w8(32'h39db6472),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3c3da),
	.w1(32'h38be7d93),
	.w2(32'hb9f0e021),
	.w3(32'h395d0444),
	.w4(32'hb99d612c),
	.w5(32'hba53122a),
	.w6(32'h39052702),
	.w7(32'h37189182),
	.w8(32'hb99dd700),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9920077),
	.w1(32'h38965306),
	.w2(32'h3801f420),
	.w3(32'hb9a1a418),
	.w4(32'h3a041e08),
	.w5(32'h39b140d5),
	.w6(32'h3955668b),
	.w7(32'h399e9533),
	.w8(32'h39f251cd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992feb6),
	.w1(32'h391cd1ea),
	.w2(32'h3a8fd9ee),
	.w3(32'h3a3200e9),
	.w4(32'h3a1173d7),
	.w5(32'h3a922823),
	.w6(32'hb91f3666),
	.w7(32'h3610ffb9),
	.w8(32'hb9a4882c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779d3f),
	.w1(32'hb952317a),
	.w2(32'hba2cb848),
	.w3(32'h3aa30cfb),
	.w4(32'hba699757),
	.w5(32'hbab64572),
	.w6(32'h38841990),
	.w7(32'h39c8bc7d),
	.w8(32'hb9b7f099),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aced4),
	.w1(32'hba2aad3d),
	.w2(32'hba66d458),
	.w3(32'hb79d1e66),
	.w4(32'hba35910c),
	.w5(32'hba80b711),
	.w6(32'h39aa15ea),
	.w7(32'hb97f334a),
	.w8(32'hba02903c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081a81),
	.w1(32'h3a1f6838),
	.w2(32'h3a08c363),
	.w3(32'hb9f2f28f),
	.w4(32'h3a69225f),
	.w5(32'h3a096b42),
	.w6(32'h39bf29d0),
	.w7(32'h3a1f1303),
	.w8(32'h3a08f5c0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a6c3),
	.w1(32'h39955b8c),
	.w2(32'hb968eba3),
	.w3(32'h3a8803ba),
	.w4(32'h38bd187b),
	.w5(32'hba3d7a53),
	.w6(32'hb893dcb0),
	.w7(32'h39656dc0),
	.w8(32'h3997f87e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899d43a),
	.w1(32'hb9c35bde),
	.w2(32'h393f41bf),
	.w3(32'hb9b551e9),
	.w4(32'h38ab407c),
	.w5(32'h371ea391),
	.w6(32'hba1d7f2b),
	.w7(32'h3a0c8433),
	.w8(32'hb7b26959),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a078297),
	.w1(32'h3a9d735e),
	.w2(32'h3ad5118a),
	.w3(32'h3a265680),
	.w4(32'h3a8aed77),
	.w5(32'h3aa48f03),
	.w6(32'h3a056f8c),
	.w7(32'h3aa09547),
	.w8(32'h3a948436),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e45dd),
	.w1(32'hb822cdd2),
	.w2(32'hb9bcad96),
	.w3(32'h3a9872a0),
	.w4(32'hb8a0caf3),
	.w5(32'hba19d3fe),
	.w6(32'h38598e65),
	.w7(32'h39ee89c4),
	.w8(32'hb9580f87),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1796c),
	.w1(32'h3a41c4a9),
	.w2(32'h3a1ac4c0),
	.w3(32'hba2c65ff),
	.w4(32'h3a5b9591),
	.w5(32'h3a11fa2d),
	.w6(32'h3a19fc67),
	.w7(32'h3a0d0173),
	.w8(32'h399e0b9b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2d178),
	.w1(32'hb871837d),
	.w2(32'hb8ef50d7),
	.w3(32'h398ab7f2),
	.w4(32'hb8e3d65a),
	.w5(32'hb992d137),
	.w6(32'h37b62ac9),
	.w7(32'hb669f9a8),
	.w8(32'hb94b0877),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946ba68),
	.w1(32'hb92c8ab2),
	.w2(32'hb9ade92d),
	.w3(32'hb99c9658),
	.w4(32'hb94d59fe),
	.w5(32'hb97b8035),
	.w6(32'hb85763a9),
	.w7(32'hb8babce3),
	.w8(32'hb9a8602d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6aad9),
	.w1(32'h39cef70b),
	.w2(32'h38d18c93),
	.w3(32'hb9367ba4),
	.w4(32'h3a82711c),
	.w5(32'h3a4deaa3),
	.w6(32'h39ef0e65),
	.w7(32'h3a0e1ce2),
	.w8(32'h3a8ac47e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb3bcf),
	.w1(32'h3a007d8e),
	.w2(32'h38e74854),
	.w3(32'h3a40d13b),
	.w4(32'h3a1b3e0a),
	.w5(32'h39c15b0a),
	.w6(32'h3a02eec3),
	.w7(32'h39e8b701),
	.w8(32'h38b0a0f6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377b72ed),
	.w1(32'hb7dd524b),
	.w2(32'hb8d28946),
	.w3(32'h39b7271d),
	.w4(32'hb8aa4fc1),
	.w5(32'hb98285cf),
	.w6(32'h388eb1ce),
	.w7(32'h389f043a),
	.w8(32'hb91aa423),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93da980),
	.w1(32'h3a690cbe),
	.w2(32'h3a51c9eb),
	.w3(32'hb9a83f6e),
	.w4(32'h3aad7c80),
	.w5(32'h3a7895f2),
	.w6(32'h3a2097d6),
	.w7(32'h39de8e73),
	.w8(32'h3a5b0bcc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a1391),
	.w1(32'h39ef6bb5),
	.w2(32'h3982f178),
	.w3(32'h3a8aad66),
	.w4(32'h39ce318f),
	.w5(32'h3938cae4),
	.w6(32'h39de4786),
	.w7(32'h392acdf8),
	.w8(32'h3936de01),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e96e2c),
	.w1(32'h390b8583),
	.w2(32'hb9ffc71c),
	.w3(32'h39d2ec6b),
	.w4(32'h39a64865),
	.w5(32'h379c0533),
	.w6(32'h3a4c39be),
	.w7(32'hb9ae5b0a),
	.w8(32'hb9b6867b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4faeb7),
	.w1(32'h3a07cf2f),
	.w2(32'h39232ad8),
	.w3(32'h38d6988a),
	.w4(32'h3a125d21),
	.w5(32'h397bc3db),
	.w6(32'h3a1d866d),
	.w7(32'h3a07fd2c),
	.w8(32'h39d404b8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1139e),
	.w1(32'h39c338b9),
	.w2(32'h3a0e29e9),
	.w3(32'h3992f884),
	.w4(32'h3a3e2369),
	.w5(32'h3a74da74),
	.w6(32'hb7d4b897),
	.w7(32'hb8f82a42),
	.w8(32'h39c038be),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b9be1),
	.w1(32'h39a7622c),
	.w2(32'h39fe1641),
	.w3(32'h3a9d4cdd),
	.w4(32'h3946e36c),
	.w5(32'h38890496),
	.w6(32'h383df729),
	.w7(32'hb9073769),
	.w8(32'hb9250434),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a3ef0),
	.w1(32'hb8afaef3),
	.w2(32'hb9484b46),
	.w3(32'hb8bc1877),
	.w4(32'hb933f98d),
	.w5(32'hb9de557f),
	.w6(32'h388a18c1),
	.w7(32'h387db361),
	.w8(32'hb96c0a2e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d4a42),
	.w1(32'h3987543f),
	.w2(32'h3973acc8),
	.w3(32'hba05a250),
	.w4(32'h39974a20),
	.w5(32'h39104726),
	.w6(32'h397aa232),
	.w7(32'h395f3508),
	.w8(32'h380744d2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992c742),
	.w1(32'h394b0805),
	.w2(32'h39176ced),
	.w3(32'h390062fc),
	.w4(32'h39849baf),
	.w5(32'h384b20e8),
	.w6(32'h3939e0d6),
	.w7(32'h391e46f6),
	.w8(32'hb8742e27),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d9986),
	.w1(32'h39758c35),
	.w2(32'h39c66329),
	.w3(32'hb7b80f42),
	.w4(32'h3a67625e),
	.w5(32'h3a7f52a6),
	.w6(32'h3926514f),
	.w7(32'hb92975f5),
	.w8(32'hb9a91b7b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01d5b1),
	.w1(32'hb9046298),
	.w2(32'hb98baf8f),
	.w3(32'h3a437ad6),
	.w4(32'hb93094b0),
	.w5(32'hba568019),
	.w6(32'hb9675c1a),
	.w7(32'h3a2bb018),
	.w8(32'h3966b5a6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1b7f8),
	.w1(32'h38882e05),
	.w2(32'hb9080c7c),
	.w3(32'h3a130543),
	.w4(32'h3a19964f),
	.w5(32'h3a04bf49),
	.w6(32'hb8dbe1e9),
	.w7(32'hb97b4bef),
	.w8(32'hb9a7a364),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be75cd),
	.w1(32'h3a0cde2b),
	.w2(32'h39805c94),
	.w3(32'h3937042f),
	.w4(32'h3a3db752),
	.w5(32'h3a04ae0c),
	.w6(32'h3992f5fe),
	.w7(32'h399e5912),
	.w8(32'h38083b29),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6e6b7),
	.w1(32'h39e899f6),
	.w2(32'h3a026529),
	.w3(32'h3a007218),
	.w4(32'h39ffab41),
	.w5(32'h39cb895d),
	.w6(32'h3997423d),
	.w7(32'h396bbc5b),
	.w8(32'h381044a8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b405f8),
	.w1(32'h3a83f6f7),
	.w2(32'h3ab47751),
	.w3(32'h398ad87e),
	.w4(32'h3b0d39ae),
	.w5(32'h3b349de3),
	.w6(32'h3a62f8cc),
	.w7(32'h397c6cf7),
	.w8(32'h39afa945),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1ab18),
	.w1(32'h3925afed),
	.w2(32'h3a0819f3),
	.w3(32'h3b43d5ee),
	.w4(32'h3a1d2825),
	.w5(32'h39d58f29),
	.w6(32'hb9473fe6),
	.w7(32'h392e3fbb),
	.w8(32'hb84dbcf4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b425),
	.w1(32'h3925770a),
	.w2(32'hb911cb7f),
	.w3(32'h39aebd37),
	.w4(32'h397a0a72),
	.w5(32'h385b185e),
	.w6(32'h38b95545),
	.w7(32'h33f864ae),
	.w8(32'hb9c8ff64),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950d8bf),
	.w1(32'hb877c9df),
	.w2(32'hbbf09140),
	.w3(32'h37f55d9a),
	.w4(32'hba2b958c),
	.w5(32'hbb021379),
	.w6(32'h37eddc58),
	.w7(32'hbb930f9d),
	.w8(32'h3b01ba63),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d01b1),
	.w1(32'h3aaac11e),
	.w2(32'h3a88d60e),
	.w3(32'hbab27a52),
	.w4(32'hbaa483fe),
	.w5(32'hbae3d79b),
	.w6(32'h3ad5335c),
	.w7(32'h3a34a879),
	.w8(32'h38a91a3d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule