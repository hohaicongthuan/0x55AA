module layer_10_featuremap_489(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fca93),
	.w1(32'hba14e11a),
	.w2(32'h3b4291dd),
	.w3(32'h3b84129f),
	.w4(32'h3b6b3375),
	.w5(32'h3bf0844f),
	.w6(32'h3bd8908b),
	.w7(32'hba15646c),
	.w8(32'h3bbe4898),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855512),
	.w1(32'h3b75513e),
	.w2(32'hba68adea),
	.w3(32'h3bccc5d0),
	.w4(32'h3be32193),
	.w5(32'h3c042b43),
	.w6(32'h3beaf0dc),
	.w7(32'h3c2d3363),
	.w8(32'h3b9a1c8f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a51b0f),
	.w1(32'hba9527e7),
	.w2(32'hbbe2c313),
	.w3(32'hbb1cf611),
	.w4(32'h3afbc690),
	.w5(32'hbaea5aff),
	.w6(32'h3b2db2d7),
	.w7(32'hbb844b41),
	.w8(32'h3933c429),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4735e),
	.w1(32'h3c031814),
	.w2(32'h3c491517),
	.w3(32'hb6f99622),
	.w4(32'h3b0e6f8b),
	.w5(32'h3a85f1e4),
	.w6(32'h3b589739),
	.w7(32'h3b611934),
	.w8(32'h3a377dc2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d747),
	.w1(32'hbba921b1),
	.w2(32'hbb474c25),
	.w3(32'hbc3dbc18),
	.w4(32'hbbf1da8b),
	.w5(32'hbc0101da),
	.w6(32'hbb02c51d),
	.w7(32'h3b682975),
	.w8(32'hbbd0f2d6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9abbb6),
	.w1(32'hbbbf341f),
	.w2(32'hbb445079),
	.w3(32'hbba90b2a),
	.w4(32'hbb1ba256),
	.w5(32'h39fbce0f),
	.w6(32'hbb4356e0),
	.w7(32'hbb840cd2),
	.w8(32'hbb4dac57),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11fe38),
	.w1(32'hbc2f8342),
	.w2(32'hbc353dcd),
	.w3(32'h3b8a9422),
	.w4(32'hbc24210f),
	.w5(32'hbc1d9331),
	.w6(32'hbabed83c),
	.w7(32'hbc650bed),
	.w8(32'hbc1e7e27),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61db48),
	.w1(32'hbb127bf6),
	.w2(32'hbb43470b),
	.w3(32'h3a2ba3b2),
	.w4(32'h3aa98554),
	.w5(32'hbbb3e2fd),
	.w6(32'hbbbb3e9b),
	.w7(32'h3bc03ff7),
	.w8(32'hbb4a7af7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae44132),
	.w1(32'h39ccccdf),
	.w2(32'h3bb31df9),
	.w3(32'h3ae7db3e),
	.w4(32'hbbae7b2f),
	.w5(32'h3c18a4fb),
	.w6(32'h3b7f00a3),
	.w7(32'hbbe181c3),
	.w8(32'hbba4d739),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0fe4),
	.w1(32'hba4c6122),
	.w2(32'h3a49ba1b),
	.w3(32'hbb243ac5),
	.w4(32'hbb8e745e),
	.w5(32'hbb20db3b),
	.w6(32'hbc030f4b),
	.w7(32'hbb43de7e),
	.w8(32'hb981c6e4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914585),
	.w1(32'hbaf2d9ce),
	.w2(32'hbbcd8e91),
	.w3(32'h3b28c70a),
	.w4(32'hbaa87991),
	.w5(32'hbb97f353),
	.w6(32'h3b0dff74),
	.w7(32'h3b7113fe),
	.w8(32'hbb986082),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bae84),
	.w1(32'h3a7c2cc7),
	.w2(32'hbab27078),
	.w3(32'hbab4ddaa),
	.w4(32'hb8e33138),
	.w5(32'h39e6d7ef),
	.w6(32'h39291cc2),
	.w7(32'h3ac76b54),
	.w8(32'hbac4ffd6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6f20e),
	.w1(32'h3bb0a202),
	.w2(32'h3c81632d),
	.w3(32'hb9223328),
	.w4(32'h3b0f7388),
	.w5(32'h3c8e682c),
	.w6(32'hba777566),
	.w7(32'hbb63203c),
	.w8(32'h3c38556e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0642b),
	.w1(32'hbb5042e6),
	.w2(32'h3b203dd4),
	.w3(32'h3abc6c68),
	.w4(32'h3b15ce83),
	.w5(32'h3c256e13),
	.w6(32'h3bff4513),
	.w7(32'hbb038a2b),
	.w8(32'h3c2b844d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e2a9),
	.w1(32'h3a8d50dd),
	.w2(32'hbc2cd5f7),
	.w3(32'hbaabf773),
	.w4(32'hba294f64),
	.w5(32'hbc0f5e05),
	.w6(32'h3b3c14b2),
	.w7(32'h3b63dc85),
	.w8(32'hbc42d797),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43939c),
	.w1(32'hbb6772bf),
	.w2(32'hba633d1b),
	.w3(32'hbc0fc044),
	.w4(32'hbb1e55af),
	.w5(32'hbb21f62a),
	.w6(32'hbbb728ff),
	.w7(32'hbc051508),
	.w8(32'hbadbdd7e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d47ae),
	.w1(32'h3ab61ea8),
	.w2(32'hbbe4b06c),
	.w3(32'hbbb4795f),
	.w4(32'h3956b4bb),
	.w5(32'hbbe7b41c),
	.w6(32'hbc1e7e14),
	.w7(32'h3b928d8f),
	.w8(32'hba55b6b6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba038ef),
	.w1(32'hb96d7066),
	.w2(32'h3b1ad007),
	.w3(32'hbc1166e9),
	.w4(32'h3b59bd83),
	.w5(32'h3a31a9c3),
	.w6(32'hbb635abb),
	.w7(32'h3b96d1b7),
	.w8(32'h3bc75984),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213635),
	.w1(32'hbb3d3b04),
	.w2(32'hbba92055),
	.w3(32'h3bcb3b39),
	.w4(32'h3a41a41b),
	.w5(32'hba72e903),
	.w6(32'h3bc52138),
	.w7(32'h3b1fa34e),
	.w8(32'hbbb58022),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3224d),
	.w1(32'hbbc4b579),
	.w2(32'h3b17d256),
	.w3(32'hbbbf90ff),
	.w4(32'h3be0bd8c),
	.w5(32'h3ab3aabc),
	.w6(32'hbc01780d),
	.w7(32'h3bc38b88),
	.w8(32'h3bb0afd8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b145191),
	.w1(32'h3833d47f),
	.w2(32'hbb53ecb1),
	.w3(32'h3afdce6f),
	.w4(32'h3b2d2dbc),
	.w5(32'hbb73d493),
	.w6(32'h3ad3b051),
	.w7(32'hbb10abae),
	.w8(32'hbb6949f8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2161),
	.w1(32'hbb4cea87),
	.w2(32'hbbc858ed),
	.w3(32'h3a207313),
	.w4(32'hbb45f2b9),
	.w5(32'hbc05fce6),
	.w6(32'hbb0b6f13),
	.w7(32'hbb58a443),
	.w8(32'hbba2cc2a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf45b30),
	.w1(32'hba9b6cf5),
	.w2(32'h3b11df34),
	.w3(32'hbbd354f6),
	.w4(32'hbbb7770a),
	.w5(32'hbbc7cec3),
	.w6(32'hbbb3c4f1),
	.w7(32'hbbea54d6),
	.w8(32'hbb8ab59c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfec1f),
	.w1(32'hbbe01f6c),
	.w2(32'h3c8df635),
	.w3(32'hbb473d34),
	.w4(32'hbbaca867),
	.w5(32'h3cbb11cf),
	.w6(32'hbba4a001),
	.w7(32'hbc66143e),
	.w8(32'h3c683f2c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0edd45),
	.w1(32'hba328509),
	.w2(32'hbb8aff9a),
	.w3(32'hbbb9fd6a),
	.w4(32'hbac2d22f),
	.w5(32'hbb4cd848),
	.w6(32'hbc81b5dc),
	.w7(32'hbbebbd61),
	.w8(32'hbbe4d239),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe3ac4),
	.w1(32'hbb39c00e),
	.w2(32'hbba72ecc),
	.w3(32'hbbb773de),
	.w4(32'hbba8699b),
	.w5(32'hbbefcefd),
	.w6(32'hbc3b90c2),
	.w7(32'hbbf911f5),
	.w8(32'hbc49e531),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab4fde),
	.w1(32'hbbacba53),
	.w2(32'hbad13f71),
	.w3(32'h3b58b26e),
	.w4(32'hbb198340),
	.w5(32'hbb402756),
	.w6(32'hb9d8fc52),
	.w7(32'hb9f0ef8e),
	.w8(32'hbb89c6ce),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0125bf),
	.w1(32'hba11b68c),
	.w2(32'hbbc5d901),
	.w3(32'h3b7b5a25),
	.w4(32'h3a13f371),
	.w5(32'hbb842dad),
	.w6(32'h3bb764ec),
	.w7(32'hbb9a9d3a),
	.w8(32'hbbb01b6e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbe264),
	.w1(32'hbba16472),
	.w2(32'h39a5cbea),
	.w3(32'h3b348d7b),
	.w4(32'hbc1d33f8),
	.w5(32'hbb8c0b9c),
	.w6(32'hba53052b),
	.w7(32'hbbd4376a),
	.w8(32'hbb4f41e2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb3d5),
	.w1(32'h3ae1dddc),
	.w2(32'h3ba8c2ee),
	.w3(32'hba5098f9),
	.w4(32'h3b1801c3),
	.w5(32'h3c23027d),
	.w6(32'hba901d53),
	.w7(32'h3bdc622d),
	.w8(32'h3c2aa014),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf349da),
	.w1(32'hba9e51ce),
	.w2(32'hbaab720d),
	.w3(32'h3c2068eb),
	.w4(32'h3b1ece19),
	.w5(32'h3b6822be),
	.w6(32'h3c44deab),
	.w7(32'hba0de455),
	.w8(32'h3a971de7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fac3d7),
	.w1(32'h3b7b3a8e),
	.w2(32'h3b13d9e5),
	.w3(32'h38c5566a),
	.w4(32'h3b41bc7d),
	.w5(32'h3c09f990),
	.w6(32'h3b5f887b),
	.w7(32'hbae6daf1),
	.w8(32'h3b8d0aa7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c408),
	.w1(32'h3ba5bde8),
	.w2(32'h3bcce643),
	.w3(32'h3a0e8eb2),
	.w4(32'h3bee56f3),
	.w5(32'h3bef7109),
	.w6(32'h3b83bf4e),
	.w7(32'h3b918268),
	.w8(32'h3b9cb317),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafddf0),
	.w1(32'h3aba07db),
	.w2(32'hbb1b123a),
	.w3(32'h3c0e4ebf),
	.w4(32'h3bd75542),
	.w5(32'h39d58b13),
	.w6(32'h3bcb167c),
	.w7(32'h3a220f85),
	.w8(32'hba836ac6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c19a1),
	.w1(32'h3a5eb2a4),
	.w2(32'h39f03700),
	.w3(32'h3a8ad6d7),
	.w4(32'h3b1c8f11),
	.w5(32'h3bcd9ef7),
	.w6(32'hbb6d75cb),
	.w7(32'hbba2cd55),
	.w8(32'hbb3d2bea),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa540),
	.w1(32'h3b9f176c),
	.w2(32'h3be38f54),
	.w3(32'h3b188bc5),
	.w4(32'h3b895f41),
	.w5(32'h3beb95d9),
	.w6(32'h3ac5f322),
	.w7(32'h3bb1b3aa),
	.w8(32'h3c0f564c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6396a),
	.w1(32'hbc1b5b9c),
	.w2(32'hbc52ffa1),
	.w3(32'h3c24053c),
	.w4(32'hbc160062),
	.w5(32'hbb769030),
	.w6(32'h3bf34373),
	.w7(32'hbc3fc6ea),
	.w8(32'hbc09e97b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2d70),
	.w1(32'h3b2c202f),
	.w2(32'h3b5df883),
	.w3(32'hbbe2414c),
	.w4(32'h3bd7dac2),
	.w5(32'h3c5dbbf4),
	.w6(32'hbbc28965),
	.w7(32'h39c9ad67),
	.w8(32'h3c155eea),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba67e36),
	.w1(32'h3a12bdd4),
	.w2(32'hbc1b15f3),
	.w3(32'h3bc93450),
	.w4(32'hbb860f5f),
	.w5(32'hbbd72ec5),
	.w6(32'h3c12ddee),
	.w7(32'hbbe47dc7),
	.w8(32'hbbd85195),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996067),
	.w1(32'h3ba4de4d),
	.w2(32'h3b8480ad),
	.w3(32'hbb22334f),
	.w4(32'h3b63adf9),
	.w5(32'h3b3914f6),
	.w6(32'h3abbcaff),
	.w7(32'h3a6edf27),
	.w8(32'hbaa7dd5f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0b575),
	.w1(32'hbb89a523),
	.w2(32'h3b7c35c5),
	.w3(32'h3bf4c520),
	.w4(32'hbc4e95f7),
	.w5(32'hbbcb3653),
	.w6(32'h3bdb3dde),
	.w7(32'hbc3c8520),
	.w8(32'hbb0b63c6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55260c),
	.w1(32'hbb736bd2),
	.w2(32'hbc3e2985),
	.w3(32'hbc345861),
	.w4(32'hbbb67128),
	.w5(32'hbc4bc8af),
	.w6(32'hbb76ba13),
	.w7(32'hbacbe364),
	.w8(32'hbc43bbe6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9795a),
	.w1(32'h3bd1ac2b),
	.w2(32'h3c3e065e),
	.w3(32'hbb63e34d),
	.w4(32'h3c09604a),
	.w5(32'h3c819310),
	.w6(32'h3ab347f4),
	.w7(32'h3c012e0f),
	.w8(32'h3c51e1c6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7059df),
	.w1(32'h3a497f87),
	.w2(32'h38bb424d),
	.w3(32'hbaf5bcae),
	.w4(32'h3a468735),
	.w5(32'hbb0c051c),
	.w6(32'h3bde1a59),
	.w7(32'hbaca6877),
	.w8(32'hbba4cfcf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb094),
	.w1(32'h3b68462c),
	.w2(32'h39d89ede),
	.w3(32'hbbd9acf4),
	.w4(32'h3ba98f50),
	.w5(32'h3a6021c0),
	.w6(32'hbb6dbfe7),
	.w7(32'h3b359967),
	.w8(32'hb8c510bb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59df00),
	.w1(32'hbaa964d8),
	.w2(32'h3b8aa944),
	.w3(32'hbb4493a7),
	.w4(32'hbaa4ccde),
	.w5(32'h3b110588),
	.w6(32'hbb9841d9),
	.w7(32'hbc02aa9f),
	.w8(32'hbac46fd1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c9332),
	.w1(32'h3af6b343),
	.w2(32'hbb6563c7),
	.w3(32'h39c53326),
	.w4(32'hba01208e),
	.w5(32'hbb787300),
	.w6(32'hbb7cd9bb),
	.w7(32'hbb67a34c),
	.w8(32'hba832bc6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdee54d),
	.w1(32'hbb3aa7a0),
	.w2(32'h39a2b867),
	.w3(32'hbc097583),
	.w4(32'hbad264f9),
	.w5(32'h3b4f6425),
	.w6(32'hbb24c23a),
	.w7(32'hbb512da3),
	.w8(32'h3a7e3fc6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21bea1),
	.w1(32'h3b0a0626),
	.w2(32'hbb636bb6),
	.w3(32'h3b72fd70),
	.w4(32'h3a82e00f),
	.w5(32'hbb38f50c),
	.w6(32'hbb5f3ad4),
	.w7(32'h3b78d5f9),
	.w8(32'h384c7aba),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb629afe),
	.w1(32'h3b0c83eb),
	.w2(32'h3b0a61b8),
	.w3(32'h3a0a9a58),
	.w4(32'hbb04df0e),
	.w5(32'h3a75644a),
	.w6(32'hbb868a59),
	.w7(32'h3a484a6c),
	.w8(32'h3a325c22),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b7b8),
	.w1(32'h3b31c016),
	.w2(32'hbabf9e09),
	.w3(32'h3abbb3dd),
	.w4(32'hba19a8b4),
	.w5(32'h3a30617d),
	.w6(32'hbb531870),
	.w7(32'h3b598509),
	.w8(32'hbb4f0ac7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ab33),
	.w1(32'hbae574b7),
	.w2(32'h3c2612c4),
	.w3(32'hbbc569e3),
	.w4(32'hbb0a315d),
	.w5(32'h3cbc1d7d),
	.w6(32'hbc182e8a),
	.w7(32'hbaf00337),
	.w8(32'h3bfdb9ef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d3f1),
	.w1(32'h3be302a2),
	.w2(32'hba41e2f0),
	.w3(32'h3c2985c1),
	.w4(32'h3bd77d3e),
	.w5(32'h3ae3cbd9),
	.w6(32'h3bcca95c),
	.w7(32'h3bb93d2c),
	.w8(32'h3acf1bc9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ea11),
	.w1(32'h3c7c7f1b),
	.w2(32'h3c84bb32),
	.w3(32'h3b0c7952),
	.w4(32'h3c83ca85),
	.w5(32'h3ca2dff9),
	.w6(32'h3a8cdaf9),
	.w7(32'h3c070160),
	.w8(32'h3c0b9de4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86de7b),
	.w1(32'hb911b751),
	.w2(32'h3b4f0049),
	.w3(32'h3c70701b),
	.w4(32'h397e9ba8),
	.w5(32'hb8abe986),
	.w6(32'h3bc8ddb8),
	.w7(32'hbb14af0d),
	.w8(32'h3b8fc78a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f26d7),
	.w1(32'h3c197cb6),
	.w2(32'h3c3a229c),
	.w3(32'h3b402787),
	.w4(32'h3c8dbf78),
	.w5(32'h3cd567c7),
	.w6(32'h3ba72fc0),
	.w7(32'h3c010dd8),
	.w8(32'h3cc62376),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9401f8),
	.w1(32'hbb871f34),
	.w2(32'h3a0db803),
	.w3(32'h3c394073),
	.w4(32'hbbad8f52),
	.w5(32'h39b9bb5d),
	.w6(32'h3c4e61f8),
	.w7(32'h3aa49328),
	.w8(32'hb9e29e55),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02264a),
	.w1(32'h3b64a7e4),
	.w2(32'hbaee8599),
	.w3(32'h3b2edfe9),
	.w4(32'h3bef9d7e),
	.w5(32'hba8c0847),
	.w6(32'h3b8bd688),
	.w7(32'h3bb06654),
	.w8(32'hbbb77d60),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c1f9),
	.w1(32'h3b97e193),
	.w2(32'h3bd35f27),
	.w3(32'hbb140d06),
	.w4(32'h3b90aea3),
	.w5(32'hba55b9c7),
	.w6(32'hbb79db30),
	.w7(32'h3b67052b),
	.w8(32'h3b7c07d4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2961a),
	.w1(32'h3b1a406f),
	.w2(32'hba3e0adb),
	.w3(32'h3987769e),
	.w4(32'h3ba5758e),
	.w5(32'hbbd21e81),
	.w6(32'h3bb436bc),
	.w7(32'h3c0e4e35),
	.w8(32'hbb6acbe8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff4fd),
	.w1(32'hba40ce4b),
	.w2(32'hbbf49fee),
	.w3(32'h3bdfde2d),
	.w4(32'hba58830f),
	.w5(32'hbbe32f22),
	.w6(32'h3ad0d0bf),
	.w7(32'h3aada5dd),
	.w8(32'h3a0f0523),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d6495),
	.w1(32'hbba10563),
	.w2(32'hbc58cef5),
	.w3(32'h3bf93572),
	.w4(32'hbb478e33),
	.w5(32'hbc123c00),
	.w6(32'h3bc93b16),
	.w7(32'hba9c6107),
	.w8(32'hbc2f3a0f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade113),
	.w1(32'h3c15be32),
	.w2(32'h3bb160a2),
	.w3(32'hbc224126),
	.w4(32'h3bdeab56),
	.w5(32'h3bbf18b1),
	.w6(32'hbbb87cbf),
	.w7(32'h3c1f8e4b),
	.w8(32'h3c2745cd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe25501),
	.w1(32'hbad47179),
	.w2(32'h3a876b02),
	.w3(32'hbc3258e0),
	.w4(32'hbb3122e7),
	.w5(32'hbb6b9b13),
	.w6(32'hbaa6f5d3),
	.w7(32'hb9c7dfd5),
	.w8(32'hbb48dda8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4633),
	.w1(32'hbb6295b9),
	.w2(32'h3b7baa81),
	.w3(32'hbba2eed8),
	.w4(32'h3afbc9ea),
	.w5(32'h3c32936d),
	.w6(32'hbb4e0914),
	.w7(32'h3b65acc8),
	.w8(32'h3c262c30),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0915),
	.w1(32'hbc06321a),
	.w2(32'hbc45dc50),
	.w3(32'h3b52c390),
	.w4(32'hbc2077da),
	.w5(32'hbc6542e0),
	.w6(32'h3aadfa08),
	.w7(32'hbc22f9c0),
	.w8(32'hbc88c333),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dbe91),
	.w1(32'hba188738),
	.w2(32'hbc01154c),
	.w3(32'hbbc4d1b5),
	.w4(32'h3b96ab27),
	.w5(32'hbb995ae3),
	.w6(32'hbc02baf7),
	.w7(32'h3bd3862e),
	.w8(32'h3afbe5f1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39228d06),
	.w1(32'h39d59c94),
	.w2(32'hbb516d27),
	.w3(32'hbafe6233),
	.w4(32'h3baa2802),
	.w5(32'h3b5cc980),
	.w6(32'h3b4d9172),
	.w7(32'h3b958ae9),
	.w8(32'h3c02a2d8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149ebb),
	.w1(32'h3b0428d2),
	.w2(32'hbbce7b54),
	.w3(32'hbbda3f99),
	.w4(32'h3c025213),
	.w5(32'hbb80af89),
	.w6(32'hbbfd71e7),
	.w7(32'h3bb75c7a),
	.w8(32'hbabe7018),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16c2a1),
	.w1(32'hbbe981ee),
	.w2(32'hbc145078),
	.w3(32'hbbe88a1d),
	.w4(32'hbb78bd22),
	.w5(32'hbc4d6613),
	.w6(32'hbc2ab525),
	.w7(32'hbbb7fe78),
	.w8(32'hbb6725e3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe31430),
	.w1(32'h3ba624bd),
	.w2(32'hba8266d4),
	.w3(32'hbbae8e9c),
	.w4(32'h3b676af0),
	.w5(32'hbb96f7b9),
	.w6(32'hbb55d9b2),
	.w7(32'h3b16bd5f),
	.w8(32'hb8c1b948),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7827b9),
	.w1(32'hbb11f374),
	.w2(32'hbbad712d),
	.w3(32'h3adf8000),
	.w4(32'hba736336),
	.w5(32'hbbfa0138),
	.w6(32'hb944d4d8),
	.w7(32'h39d338b8),
	.w8(32'hbb970b55),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946806d),
	.w1(32'hbb48f237),
	.w2(32'h3b05ddc7),
	.w3(32'h3c075b95),
	.w4(32'hbbb70023),
	.w5(32'hbae4c95c),
	.w6(32'h3ba3663a),
	.w7(32'hba21476a),
	.w8(32'hbacc0ff9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933f1e),
	.w1(32'hbac01c57),
	.w2(32'hbb6b14e7),
	.w3(32'h39ce6791),
	.w4(32'hbba7d85d),
	.w5(32'h3a7378e6),
	.w6(32'hbc18760c),
	.w7(32'hb91fdd9c),
	.w8(32'hba39776b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2d8ee),
	.w1(32'h3c0d5717),
	.w2(32'hbba223da),
	.w3(32'hbb18a60f),
	.w4(32'h3c56a89e),
	.w5(32'hbbae7d22),
	.w6(32'hbba05890),
	.w7(32'h3afd1d41),
	.w8(32'hbbce81f9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dc8d1),
	.w1(32'h3afca8c0),
	.w2(32'h3c57abd4),
	.w3(32'h3b6732c1),
	.w4(32'h3a871628),
	.w5(32'h3bca1213),
	.w6(32'hba3736c4),
	.w7(32'h3b45be79),
	.w8(32'hba8f070a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c726709),
	.w1(32'hbb81653e),
	.w2(32'hbb80a47a),
	.w3(32'h3c021867),
	.w4(32'hbbfdeb95),
	.w5(32'hbbe110f5),
	.w6(32'hbabc0568),
	.w7(32'hbbf95dac),
	.w8(32'hbc0c6a52),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061329),
	.w1(32'hba447213),
	.w2(32'hba0f055b),
	.w3(32'hbc24f026),
	.w4(32'hbaddcf3c),
	.w5(32'hbb37000f),
	.w6(32'hbc278fd6),
	.w7(32'h3b6f3684),
	.w8(32'hbb8c1753),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8870),
	.w1(32'hbb91b83a),
	.w2(32'hbbf0103b),
	.w3(32'hba8ce268),
	.w4(32'hbb9f70d6),
	.w5(32'hba5daba3),
	.w6(32'hbb13dc82),
	.w7(32'hbb344dd2),
	.w8(32'hbbdfa461),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d91c),
	.w1(32'h3bed9b35),
	.w2(32'h3b165054),
	.w3(32'hbbc0d939),
	.w4(32'h3cb57d36),
	.w5(32'h3bbd5138),
	.w6(32'hbb1aeff8),
	.w7(32'h3c2d11ab),
	.w8(32'h3c9c9aca),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d2bd),
	.w1(32'hbc56b431),
	.w2(32'hbc1f31ad),
	.w3(32'hbb26b9a3),
	.w4(32'hbc0d0f63),
	.w5(32'h3be79fdd),
	.w6(32'h3bafb66d),
	.w7(32'hbc336ac0),
	.w8(32'hbc134a08),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c8b0b),
	.w1(32'hb9452db0),
	.w2(32'h3a5cae16),
	.w3(32'hbc83c59e),
	.w4(32'hbb5bbc9c),
	.w5(32'hbb5a7429),
	.w6(32'hbc8e5428),
	.w7(32'hbb7b5ae1),
	.w8(32'hbb08b305),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3be6c3),
	.w1(32'h3ababeb8),
	.w2(32'h3afd8e79),
	.w3(32'h382170f2),
	.w4(32'hbae89495),
	.w5(32'h3b594c57),
	.w6(32'h3a79c850),
	.w7(32'hbb8acf50),
	.w8(32'hbac2c7a7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49ebe6),
	.w1(32'h3b300522),
	.w2(32'h3b9feb82),
	.w3(32'h3b871f25),
	.w4(32'hba807e2b),
	.w5(32'h3b013815),
	.w6(32'h3b4e1aae),
	.w7(32'h3b1a453f),
	.w8(32'h3ba17985),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2ccd8),
	.w1(32'h3a2db605),
	.w2(32'h3b097226),
	.w3(32'h3bd1c5ea),
	.w4(32'hb927ae2c),
	.w5(32'hba214a7c),
	.w6(32'h3a40d3bb),
	.w7(32'h3ab0a991),
	.w8(32'h3a9eff37),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1f25),
	.w1(32'h39e4552b),
	.w2(32'hbc086507),
	.w3(32'h3b377899),
	.w4(32'hbb5bee59),
	.w5(32'hbc1116fb),
	.w6(32'hba0929e2),
	.w7(32'h3a7e9fd4),
	.w8(32'h3b31c0ac),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc035),
	.w1(32'h3b891f84),
	.w2(32'h3b4b1627),
	.w3(32'h3bdd37a0),
	.w4(32'h3b27654f),
	.w5(32'h3b7b7a56),
	.w6(32'h3c08b3bf),
	.w7(32'hbbeedb32),
	.w8(32'h3a73cd3e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7adf4b),
	.w1(32'h3ad2a2bf),
	.w2(32'h39cb01d4),
	.w3(32'h3aedfeb8),
	.w4(32'hbbc8ba53),
	.w5(32'hb7aa6bb1),
	.w6(32'h3b25f912),
	.w7(32'hbc0007dc),
	.w8(32'hbb44d4e5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b240bdb),
	.w1(32'h3be3fcf0),
	.w2(32'h3bb74dc5),
	.w3(32'h3b63eefa),
	.w4(32'hbb3916ea),
	.w5(32'hbbc19347),
	.w6(32'hbaa0b15c),
	.w7(32'hb9fbeed2),
	.w8(32'h3b2d550e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f2c2),
	.w1(32'hba60b50f),
	.w2(32'h3ab5f804),
	.w3(32'hbb328593),
	.w4(32'hbbd1755f),
	.w5(32'hbc0779c6),
	.w6(32'h3c1caa58),
	.w7(32'hbb4388c3),
	.w8(32'hbb925ac6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a692683),
	.w1(32'h3bbd52d8),
	.w2(32'h3b9425e9),
	.w3(32'hbb3215e8),
	.w4(32'h3b855a87),
	.w5(32'hbc20d578),
	.w6(32'hb97ea17e),
	.w7(32'h3a94efff),
	.w8(32'hbb47b922),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0a9af),
	.w1(32'h3b68f34d),
	.w2(32'hbba5da64),
	.w3(32'hbbbb18ac),
	.w4(32'hbb2c5f34),
	.w5(32'hbbfde4b7),
	.w6(32'h3acbce3b),
	.w7(32'hba4271d9),
	.w8(32'hbbca7f9f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab913f8),
	.w1(32'hbbf3fd45),
	.w2(32'hbc03aa16),
	.w3(32'hbb4eebe7),
	.w4(32'hbb8e9e3b),
	.w5(32'h3b98639b),
	.w6(32'hbbf055ee),
	.w7(32'hbb83e100),
	.w8(32'hbad4d13e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf992c0),
	.w1(32'hba8772ab),
	.w2(32'h3b5ed4be),
	.w3(32'hbb0ce416),
	.w4(32'hbbb63a48),
	.w5(32'h3bddaabb),
	.w6(32'hbbc84a3f),
	.w7(32'hbb47d960),
	.w8(32'h3ac159b4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba046b10),
	.w1(32'hba80c843),
	.w2(32'hbb04a743),
	.w3(32'hbaf9db9c),
	.w4(32'h3c12a809),
	.w5(32'h39db667d),
	.w6(32'hbbc99ffd),
	.w7(32'h3c2d1bb0),
	.w8(32'h3bb2ae56),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37673f),
	.w1(32'h38db89da),
	.w2(32'h3b95d661),
	.w3(32'hba830c67),
	.w4(32'h3a82479e),
	.w5(32'h3a8cf619),
	.w6(32'h3b84731c),
	.w7(32'h3b83aed6),
	.w8(32'h3bc8d550),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8569e7),
	.w1(32'h3ba0b14a),
	.w2(32'hbad69619),
	.w3(32'hb9cc814e),
	.w4(32'h3a2dad4a),
	.w5(32'hbb3ee762),
	.w6(32'hbb41a45d),
	.w7(32'h3a96f160),
	.w8(32'h3b7677f0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd023),
	.w1(32'hbb087e5f),
	.w2(32'hbbbbf68d),
	.w3(32'hb9d0ab08),
	.w4(32'hbb458cff),
	.w5(32'hbbedb10d),
	.w6(32'h3a4a2cd5),
	.w7(32'hbb0ae1a3),
	.w8(32'hbb8faa5f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8569),
	.w1(32'hbb29e498),
	.w2(32'hbbabc99d),
	.w3(32'hbbac9b44),
	.w4(32'hbb7d313b),
	.w5(32'hbcb2ff48),
	.w6(32'hbbe7832e),
	.w7(32'hbc43193d),
	.w8(32'hbbc9379b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cde85),
	.w1(32'hbac9f133),
	.w2(32'hbb9f0417),
	.w3(32'hbbf18113),
	.w4(32'hbb9efeff),
	.w5(32'hbc1f118a),
	.w6(32'hbbbb2a8e),
	.w7(32'hbadfcbde),
	.w8(32'hbb95b394),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca343),
	.w1(32'h3bd18f36),
	.w2(32'h3b444765),
	.w3(32'h3b14d9ee),
	.w4(32'h3bb619df),
	.w5(32'hbae76903),
	.w6(32'hbb20dd64),
	.w7(32'h3bd7660c),
	.w8(32'h3ac0b8dc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba035074),
	.w1(32'hbb554660),
	.w2(32'hbc0a76ef),
	.w3(32'h3940c5b0),
	.w4(32'hbbfaf3ed),
	.w5(32'hbbc08a78),
	.w6(32'hb83489cf),
	.w7(32'hbbebbf03),
	.w8(32'hbc176e2a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda4b0),
	.w1(32'hbb5fa073),
	.w2(32'h3a22ad96),
	.w3(32'h3baaf938),
	.w4(32'hbbd026df),
	.w5(32'hbb05a513),
	.w6(32'hbaa14172),
	.w7(32'hbaebe37b),
	.w8(32'hbb9cd618),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66166c),
	.w1(32'hbc1a2be4),
	.w2(32'hbb919a1a),
	.w3(32'hba4e2fc7),
	.w4(32'hbb87709f),
	.w5(32'hb9c16cc0),
	.w6(32'hbafe0f4c),
	.w7(32'hbb0d81c3),
	.w8(32'hbae645b3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af80a71),
	.w1(32'h39a859ef),
	.w2(32'hbb231eae),
	.w3(32'h3b49ea33),
	.w4(32'hb9b07d5d),
	.w5(32'h39cfb4fe),
	.w6(32'hbaefb8b0),
	.w7(32'hbb87f05b),
	.w8(32'hbb9e31f4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac4f1),
	.w1(32'h3bf6cb7b),
	.w2(32'h3a380b31),
	.w3(32'h3b1718a1),
	.w4(32'h3be0968e),
	.w5(32'h39f2ada9),
	.w6(32'h3aefe1e3),
	.w7(32'h3c17788c),
	.w8(32'h3be13de1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b4ce),
	.w1(32'hbb09af52),
	.w2(32'hba0933b4),
	.w3(32'hba60cb1d),
	.w4(32'hb988a497),
	.w5(32'h3b8befb4),
	.w6(32'h3b80fd32),
	.w7(32'hb9f6a05e),
	.w8(32'h3b216d13),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f7a8),
	.w1(32'hbbd6db62),
	.w2(32'hbbad00ad),
	.w3(32'h3a6d6240),
	.w4(32'hbb16b280),
	.w5(32'hbba53139),
	.w6(32'h39b8788f),
	.w7(32'hbb13c8d8),
	.w8(32'h36dc316a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98963),
	.w1(32'hbaf1b9a6),
	.w2(32'hbb2fa050),
	.w3(32'hbc426f49),
	.w4(32'hbb3f7796),
	.w5(32'h3b7a0860),
	.w6(32'hbc1b1bc0),
	.w7(32'hbbcaf2b5),
	.w8(32'hbb6a3638),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16b0c8),
	.w1(32'h3b8a0a99),
	.w2(32'hbb9b8a8f),
	.w3(32'hb99ab68c),
	.w4(32'h3b302ae1),
	.w5(32'h3b4e8a59),
	.w6(32'hbb92ce59),
	.w7(32'hbbc7eb3c),
	.w8(32'h3919eaf4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0996eb),
	.w1(32'h3c0fe6ef),
	.w2(32'hba5f0a34),
	.w3(32'hbafa5560),
	.w4(32'hbb8eaba8),
	.w5(32'hbc389eb8),
	.w6(32'h3a87d314),
	.w7(32'hbb3c0bc2),
	.w8(32'hbbb9bd16),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad8a8),
	.w1(32'h3c22cff8),
	.w2(32'h3b8b5af7),
	.w3(32'hbc0c7431),
	.w4(32'h3c01613c),
	.w5(32'hbbd91505),
	.w6(32'hbbbe3c21),
	.w7(32'h3c158505),
	.w8(32'hbaa196b9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba815f78),
	.w1(32'hbaffa9f7),
	.w2(32'h3ad4021d),
	.w3(32'h3bdb62af),
	.w4(32'hbbae5717),
	.w5(32'h3b2cf4f2),
	.w6(32'h3b0aa0c0),
	.w7(32'h3af914dd),
	.w8(32'h3b8a901a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae448b),
	.w1(32'hbbfe8116),
	.w2(32'hbbbbbf9d),
	.w3(32'h3ac01ecb),
	.w4(32'hbba008fe),
	.w5(32'h3c45f9ae),
	.w6(32'h3b11e866),
	.w7(32'h3abd9d79),
	.w8(32'h3b475f94),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16c5be),
	.w1(32'hbb54fcf9),
	.w2(32'hbc230576),
	.w3(32'h3b1fc470),
	.w4(32'hbbc4682c),
	.w5(32'hbb97be7b),
	.w6(32'h396307c0),
	.w7(32'h3a337faf),
	.w8(32'hbb02cbc2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60cc64),
	.w1(32'hbb65449d),
	.w2(32'h3aea364a),
	.w3(32'hbbe4716a),
	.w4(32'hbb4f00ba),
	.w5(32'hbb707d81),
	.w6(32'hbb97c1eb),
	.w7(32'h3a12f362),
	.w8(32'h3a1a3deb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac79774),
	.w1(32'h3a6c0e12),
	.w2(32'h390ad149),
	.w3(32'h39e5ae0e),
	.w4(32'h3b39dc79),
	.w5(32'h3aaa1935),
	.w6(32'h3a0d8f90),
	.w7(32'h3c126605),
	.w8(32'h3b9016d1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256088),
	.w1(32'h3a14c82c),
	.w2(32'hbaf22619),
	.w3(32'hb9ce56e2),
	.w4(32'hbb7f5d71),
	.w5(32'hb93887d1),
	.w6(32'h39147dca),
	.w7(32'h3acf94c6),
	.w8(32'hbaed5538),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad23b38),
	.w1(32'hb999aeec),
	.w2(32'h3afd400b),
	.w3(32'hbc133d55),
	.w4(32'hbb9dcada),
	.w5(32'hb9205c25),
	.w6(32'hbbd7c9f8),
	.w7(32'hba8a8bd0),
	.w8(32'hba76a067),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c196e),
	.w1(32'hbb5ecc5a),
	.w2(32'hbb877f53),
	.w3(32'h3bc2890d),
	.w4(32'hbb85ad16),
	.w5(32'h3a66cf06),
	.w6(32'h3b2bb4a9),
	.w7(32'hbad6f881),
	.w8(32'h3b9f48ab),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba724db3),
	.w1(32'hbafad003),
	.w2(32'hba4bf706),
	.w3(32'h3a93e598),
	.w4(32'hbb92b116),
	.w5(32'h39eec2a4),
	.w6(32'h389873aa),
	.w7(32'hbb65c501),
	.w8(32'hbaf95546),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ce2e),
	.w1(32'h3b6b7730),
	.w2(32'h3b89a66b),
	.w3(32'hbad4481f),
	.w4(32'h3c435bf7),
	.w5(32'h3aeda198),
	.w6(32'hba9513c5),
	.w7(32'h3b2543da),
	.w8(32'hbb27d8ec),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cce4d1),
	.w1(32'h3ba070a0),
	.w2(32'h3b8eb615),
	.w3(32'hbbb13ec6),
	.w4(32'h3bb3f4cf),
	.w5(32'h3bff8a10),
	.w6(32'hbb150eca),
	.w7(32'h3b9c9a4c),
	.w8(32'h3bad2d3b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aa541),
	.w1(32'h3aa9a761),
	.w2(32'hbafa33b8),
	.w3(32'h3c395fa0),
	.w4(32'hbb6ed6f3),
	.w5(32'hb6d4925a),
	.w6(32'h3bcf30e6),
	.w7(32'hbae53b0b),
	.w8(32'hbb812bb3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb0f18),
	.w1(32'hbb239234),
	.w2(32'hbb99dd2b),
	.w3(32'hbc06624a),
	.w4(32'hba1e1f17),
	.w5(32'h3a474cab),
	.w6(32'hbbcb2f2d),
	.w7(32'hba3654f7),
	.w8(32'hbbb58ad2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0627e),
	.w1(32'h3c0485bd),
	.w2(32'h3a02dfae),
	.w3(32'hb9592141),
	.w4(32'h3b1bd8de),
	.w5(32'hb9ba3b1f),
	.w6(32'hbb867740),
	.w7(32'h3af3a9a7),
	.w8(32'hbacd313d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb909),
	.w1(32'h3c303e0a),
	.w2(32'hbabf538c),
	.w3(32'h3a4d4e70),
	.w4(32'h3c402f81),
	.w5(32'hbca7774f),
	.w6(32'h3b6d7fb1),
	.w7(32'h3c1313f4),
	.w8(32'hbbf7d9c8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef4850),
	.w1(32'hbaafa72a),
	.w2(32'hbb7c6fba),
	.w3(32'hbc83fdc8),
	.w4(32'hbaea398e),
	.w5(32'hbc02d6f9),
	.w6(32'hbc1b92ff),
	.w7(32'h3b64e74b),
	.w8(32'h3b934fa2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fb075),
	.w1(32'h3c2e36cc),
	.w2(32'h3afe74f8),
	.w3(32'h3bebc16a),
	.w4(32'h3c024a41),
	.w5(32'hbae6c86a),
	.w6(32'h3bf4895b),
	.w7(32'h3b784961),
	.w8(32'h3bd5cc8b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfd203),
	.w1(32'h3ba768d1),
	.w2(32'hb838f373),
	.w3(32'hbc1a2a68),
	.w4(32'hba069d9a),
	.w5(32'hbc061874),
	.w6(32'h3aeed217),
	.w7(32'h3b3cf940),
	.w8(32'hbbaa5726),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea46f0),
	.w1(32'hbb8408a2),
	.w2(32'h3b431e01),
	.w3(32'h3bfdb381),
	.w4(32'hbb43cb1f),
	.w5(32'hbb85850a),
	.w6(32'h3bd89e57),
	.w7(32'h3b38bf46),
	.w8(32'h3b8740c2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1663e5),
	.w1(32'hbb78f2d7),
	.w2(32'h3a6574a5),
	.w3(32'hbab7211b),
	.w4(32'h3a65e43b),
	.w5(32'hba8fbe7b),
	.w6(32'hbba0c89b),
	.w7(32'h3becfc24),
	.w8(32'hbaeca88b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29f072),
	.w1(32'h3a4a3e87),
	.w2(32'hbaebda73),
	.w3(32'hbb01a631),
	.w4(32'h3b25fef1),
	.w5(32'h3ba29140),
	.w6(32'h3bb4fbdb),
	.w7(32'hb7e28ec8),
	.w8(32'h3a9f71d5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9367e4),
	.w1(32'hba8fc94d),
	.w2(32'hba9543aa),
	.w3(32'h3a1d1f5b),
	.w4(32'hbb9cc8ba),
	.w5(32'hba802335),
	.w6(32'hba993cd5),
	.w7(32'h352189f0),
	.w8(32'hbb8e905f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c88549),
	.w1(32'hbb882730),
	.w2(32'h3a81ad11),
	.w3(32'h3acd2644),
	.w4(32'hbb864601),
	.w5(32'hbb04dbc7),
	.w6(32'h3abee2c1),
	.w7(32'hbb1feab0),
	.w8(32'hbb160a21),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393914a6),
	.w1(32'hbafc964a),
	.w2(32'hb9d76161),
	.w3(32'h3b130c8b),
	.w4(32'hbbc90ba4),
	.w5(32'h3bb85dc3),
	.w6(32'hbaf77764),
	.w7(32'hbb20fb54),
	.w8(32'hb9fff53b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a3570),
	.w1(32'hb9895b82),
	.w2(32'hbb2964d3),
	.w3(32'hbc100750),
	.w4(32'h3b080d6a),
	.w5(32'h3bdfc9b9),
	.w6(32'hbbee3282),
	.w7(32'h3bd7490f),
	.w8(32'h3b8757e1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b81e),
	.w1(32'hba9b1d24),
	.w2(32'h3a0d3aa3),
	.w3(32'h3bbd40ac),
	.w4(32'h39f73936),
	.w5(32'h3ab7ac8b),
	.w6(32'h3bbbca5a),
	.w7(32'hb9d85962),
	.w8(32'h3b170653),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc6b62),
	.w1(32'hbb1562bd),
	.w2(32'hbb4808d3),
	.w3(32'hba0c58cb),
	.w4(32'h3b153dbc),
	.w5(32'hb6b0f721),
	.w6(32'h3b8ed484),
	.w7(32'h3b4e4add),
	.w8(32'h3b9d523c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074103),
	.w1(32'hbc0ab469),
	.w2(32'hbb02aa92),
	.w3(32'hb8aedd64),
	.w4(32'hbc0d06d1),
	.w5(32'hb9ea48f6),
	.w6(32'h3b1a2fc9),
	.w7(32'hbc1ac710),
	.w8(32'hbbbfdfea),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f929a),
	.w1(32'h3bfb50ac),
	.w2(32'h3a0a9877),
	.w3(32'hbae448f0),
	.w4(32'h3b879170),
	.w5(32'hbbcdefd6),
	.w6(32'hbbc7021c),
	.w7(32'h3bf1ea03),
	.w8(32'hbb5f25f5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b8f3b),
	.w1(32'hba8d3f77),
	.w2(32'h3ba025e3),
	.w3(32'h3ac89e94),
	.w4(32'h3a65ab9c),
	.w5(32'h3b911ec0),
	.w6(32'hbadb6e60),
	.w7(32'h3b7c9d0a),
	.w8(32'h3c3b2b88),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02f9bc),
	.w1(32'hba9d9140),
	.w2(32'h3a98910c),
	.w3(32'h3bb271e5),
	.w4(32'hba4a7f2d),
	.w5(32'h3b5747a6),
	.w6(32'h3c0a37a5),
	.w7(32'h3a41a094),
	.w8(32'h3a19b4c6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e6e11),
	.w1(32'hbb692284),
	.w2(32'hba4cff26),
	.w3(32'h3bf3a29b),
	.w4(32'hbb87459b),
	.w5(32'h3a38571d),
	.w6(32'h3b0c167b),
	.w7(32'hbb9c9a1a),
	.w8(32'hbaf54114),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf50f6),
	.w1(32'h3c127123),
	.w2(32'h3c7cfac8),
	.w3(32'hba5c4cec),
	.w4(32'h3a8ade67),
	.w5(32'h3b1cdd25),
	.w6(32'hbbb09555),
	.w7(32'hbb7b1a36),
	.w8(32'hbb34be5b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca328cc),
	.w1(32'h3bc90c37),
	.w2(32'h3bb17dea),
	.w3(32'h3c422f6c),
	.w4(32'h3b5e25e1),
	.w5(32'h3ba50563),
	.w6(32'hb9acbae8),
	.w7(32'h3b0faa09),
	.w8(32'h3ba28516),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ce715),
	.w1(32'h3a85cddb),
	.w2(32'h3adc360d),
	.w3(32'hbc0bd957),
	.w4(32'hba7e778c),
	.w5(32'h3b3f809f),
	.w6(32'hbb92c03b),
	.w7(32'hba16ba42),
	.w8(32'h3839abc9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5db7d),
	.w1(32'hbb1602ed),
	.w2(32'h3babab4d),
	.w3(32'h3ac0a239),
	.w4(32'hbc210257),
	.w5(32'hbc090042),
	.w6(32'h3b19dda1),
	.w7(32'hbc4b7d54),
	.w8(32'hbb86df7b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf2a93),
	.w1(32'hbb85a2eb),
	.w2(32'hbadb832f),
	.w3(32'h3c25f968),
	.w4(32'hb99e418f),
	.w5(32'h3ba470a9),
	.w6(32'h3a6801da),
	.w7(32'hbb64d45d),
	.w8(32'h3b4c6169),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ea43),
	.w1(32'h3a9a6750),
	.w2(32'hbbb4e593),
	.w3(32'hbb890681),
	.w4(32'h3ae440f2),
	.w5(32'hbbbd669a),
	.w6(32'hbab8d3e9),
	.w7(32'h3b9ea578),
	.w8(32'hbb03439c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9685be),
	.w1(32'h3bbb1462),
	.w2(32'h3b13e926),
	.w3(32'h3a63e307),
	.w4(32'h3c01ff94),
	.w5(32'hbbd37b60),
	.w6(32'h3b714516),
	.w7(32'h3b791a07),
	.w8(32'hbbc97426),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c006a),
	.w1(32'hb9bb9b1b),
	.w2(32'h3c4e726c),
	.w3(32'hbb045d32),
	.w4(32'h3bfb2136),
	.w5(32'h3cbf8bee),
	.w6(32'hba30ae69),
	.w7(32'h3a59060a),
	.w8(32'h3c32ce08),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d39c),
	.w1(32'h3ba2ac69),
	.w2(32'h3c026832),
	.w3(32'h3c0bcb17),
	.w4(32'h3b6fd4c2),
	.w5(32'hbb67fed7),
	.w6(32'h3bb8fc01),
	.w7(32'h3bf46255),
	.w8(32'h3b99be86),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb50b),
	.w1(32'hbb1b007d),
	.w2(32'hbbd292f5),
	.w3(32'hbc0e2bea),
	.w4(32'hbaef5806),
	.w5(32'hbb34590a),
	.w6(32'hbbc04425),
	.w7(32'h3a032fdd),
	.w8(32'hbb75e462),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc9da0),
	.w1(32'h3babda49),
	.w2(32'h35b5da80),
	.w3(32'hbbf8f69b),
	.w4(32'hbbb6a0ed),
	.w5(32'hbbff1bde),
	.w6(32'hbbeea0db),
	.w7(32'hbbaa7630),
	.w8(32'hbc1b1d27),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d456c),
	.w1(32'hbb8fe01f),
	.w2(32'hbb9904e9),
	.w3(32'hbb5e1025),
	.w4(32'hbb5da2c4),
	.w5(32'hbbf9a2dd),
	.w6(32'hbbea4742),
	.w7(32'hbb37ab35),
	.w8(32'hbbd3376c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14288e),
	.w1(32'h3cadab72),
	.w2(32'h3cb4fe88),
	.w3(32'hbb77f668),
	.w4(32'h3cd56db5),
	.w5(32'h39fe0281),
	.w6(32'hbb51f22f),
	.w7(32'h3b2f5c7a),
	.w8(32'hbb966727),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194b8e),
	.w1(32'h3a98530f),
	.w2(32'h3a96c447),
	.w3(32'hbb279fa1),
	.w4(32'hbb864129),
	.w5(32'hbaa5049a),
	.w6(32'hbb8bef36),
	.w7(32'hba9f2054),
	.w8(32'h3ad0e917),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3ba3b),
	.w1(32'hba6a7ba8),
	.w2(32'hba817c93),
	.w3(32'hbbced22f),
	.w4(32'hbb9ee1ab),
	.w5(32'hbbb73758),
	.w6(32'hbb428987),
	.w7(32'hbb5e32c2),
	.w8(32'hbb8a9bc7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5495e5),
	.w1(32'h3b4ca5cd),
	.w2(32'hb99bd7e8),
	.w3(32'h3acfc41d),
	.w4(32'h3afdfe85),
	.w5(32'h3ab7e147),
	.w6(32'hb990c21c),
	.w7(32'h3b941f67),
	.w8(32'h3b1d029e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3942d6),
	.w1(32'hbbccfb7f),
	.w2(32'hbba7605d),
	.w3(32'h3b2a6034),
	.w4(32'hbbda4ad0),
	.w5(32'hbb84dcf7),
	.w6(32'h3a2e9644),
	.w7(32'hbc022bb8),
	.w8(32'hbbf03d3b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9705df),
	.w1(32'h3ba933ef),
	.w2(32'hbb49a49f),
	.w3(32'h395e13d5),
	.w4(32'hba8c3b40),
	.w5(32'hbbcc3ca2),
	.w6(32'hbb8ee1e6),
	.w7(32'h3b9e2aae),
	.w8(32'h3b1df70f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a045),
	.w1(32'hba1bff94),
	.w2(32'h3b56274f),
	.w3(32'hbbd683c5),
	.w4(32'h3a9afb20),
	.w5(32'h3c0848c1),
	.w6(32'hbb3306d7),
	.w7(32'hbaccdbb4),
	.w8(32'h3bb60937),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e007f2),
	.w1(32'hbbcce244),
	.w2(32'hbbfbaf81),
	.w3(32'h3a84bdea),
	.w4(32'hbb8ae4ed),
	.w5(32'hbb1c4652),
	.w6(32'h3946f227),
	.w7(32'hbb9128ff),
	.w8(32'hbb713268),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9b83),
	.w1(32'h3b76945a),
	.w2(32'h3c2dd949),
	.w3(32'hbc00f94a),
	.w4(32'h3c453fea),
	.w5(32'h3bfce51a),
	.w6(32'hbb3feeb7),
	.w7(32'h3bc1e821),
	.w8(32'h3c1dbcac),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ad948),
	.w1(32'hbc0314b8),
	.w2(32'hbb4e46c9),
	.w3(32'h3baaa2c3),
	.w4(32'hbc462b4b),
	.w5(32'hbc2243f5),
	.w6(32'h3bc3d592),
	.w7(32'hbbdb8843),
	.w8(32'hbc2b9db8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba00438),
	.w1(32'hbbc7bc86),
	.w2(32'hbbda8135),
	.w3(32'h3bb12802),
	.w4(32'hbbbc9e5f),
	.w5(32'hbc1b8d7c),
	.w6(32'hba666185),
	.w7(32'hbbb2cc79),
	.w8(32'hbadebcfb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef6f5),
	.w1(32'hbbb19e10),
	.w2(32'hbb5b6970),
	.w3(32'hbbd25194),
	.w4(32'h3aa7e053),
	.w5(32'hb9283bfd),
	.w6(32'hbba4f177),
	.w7(32'hba18089f),
	.w8(32'hbb0654ac),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9374fe9),
	.w1(32'h3a9c567f),
	.w2(32'h3ba8baf1),
	.w3(32'hbb9823ed),
	.w4(32'h3b5c65ef),
	.w5(32'h3c1ea703),
	.w6(32'hbac8beaa),
	.w7(32'h36c6f6e3),
	.w8(32'hbb44b5cb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84f043),
	.w1(32'h3b7d289b),
	.w2(32'hbb495fcf),
	.w3(32'h3bfb0715),
	.w4(32'hbb250fa9),
	.w5(32'h3a55e502),
	.w6(32'hbb995c4f),
	.w7(32'h3b09f1c4),
	.w8(32'h3aac608a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5bf27),
	.w1(32'h3bb455ba),
	.w2(32'h3bad89e9),
	.w3(32'h3b625707),
	.w4(32'h3b1a69fb),
	.w5(32'h3b0df781),
	.w6(32'h3bc03ada),
	.w7(32'h3bc93c88),
	.w8(32'h3b266574),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942d8d2),
	.w1(32'hbbaf12e4),
	.w2(32'hbbef4e6e),
	.w3(32'hbbbf08ce),
	.w4(32'hbadc80bf),
	.w5(32'hbba1a79e),
	.w6(32'h3b07f87d),
	.w7(32'h3a660306),
	.w8(32'hba8779a6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacca831),
	.w1(32'hbb765a6a),
	.w2(32'hbae2a12a),
	.w3(32'hbbf1291e),
	.w4(32'hbb5e66be),
	.w5(32'hbb09a743),
	.w6(32'hbbfd4204),
	.w7(32'hbb56f02f),
	.w8(32'hbb9e3202),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1470e),
	.w1(32'hb9a04b06),
	.w2(32'h3bbb3296),
	.w3(32'hbb473fa0),
	.w4(32'hba62ec7d),
	.w5(32'h3a92fa58),
	.w6(32'hbbe52c57),
	.w7(32'hbb0584f9),
	.w8(32'h3a82e5ed),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba763a1d),
	.w1(32'h3a9435c0),
	.w2(32'hbb890b23),
	.w3(32'h3b739a9a),
	.w4(32'hba6496af),
	.w5(32'hbbaa8372),
	.w6(32'hbb308c8f),
	.w7(32'hba87b293),
	.w8(32'hba3afcc1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9073),
	.w1(32'h3bf1a35e),
	.w2(32'h3bf27474),
	.w3(32'hbaab4e05),
	.w4(32'h3c1102fa),
	.w5(32'h393c2d78),
	.w6(32'hba2c2330),
	.w7(32'h3c32360f),
	.w8(32'h3c262b9f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c341841),
	.w1(32'h3bf26739),
	.w2(32'h3a289964),
	.w3(32'h3c1b1f5e),
	.w4(32'h3c15cf9a),
	.w5(32'h3c185441),
	.w6(32'h3c2f9917),
	.w7(32'h3bb220c8),
	.w8(32'hba39d07a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8f3ca),
	.w1(32'hb8d6d031),
	.w2(32'hbb7f331d),
	.w3(32'hbbe35436),
	.w4(32'hbb120472),
	.w5(32'h3bb4ece3),
	.w6(32'hbbac6a6d),
	.w7(32'hbb2d4b5a),
	.w8(32'hbac0739e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5e3db),
	.w1(32'h3c46f66c),
	.w2(32'h3af4d44c),
	.w3(32'hbbc57dd2),
	.w4(32'h3c1fc7f7),
	.w5(32'hbb21bee2),
	.w6(32'hba222ce2),
	.w7(32'h3bb57a14),
	.w8(32'h3b5054b6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a136ce6),
	.w1(32'h3bbcf482),
	.w2(32'h3bcfe96f),
	.w3(32'hba37b3b9),
	.w4(32'h3aa62a6a),
	.w5(32'h3bb73057),
	.w6(32'h3bc9a66d),
	.w7(32'hbbe7e760),
	.w8(32'h3ab36183),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c34fb),
	.w1(32'hbb826a34),
	.w2(32'hbb2b3d30),
	.w3(32'h3ad4842c),
	.w4(32'hbbb21114),
	.w5(32'h3b758529),
	.w6(32'h3b8ca1ea),
	.w7(32'h3a0c2afb),
	.w8(32'h3b3e8d92),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a4604),
	.w1(32'hbb2e3d78),
	.w2(32'h3b06d7b3),
	.w3(32'hbb8768ea),
	.w4(32'hbb87419e),
	.w5(32'h3ba96ab0),
	.w6(32'hbb806c99),
	.w7(32'hbc147737),
	.w8(32'hbaae0882),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38249),
	.w1(32'hbb53d488),
	.w2(32'hb9c75486),
	.w3(32'hbbb2974d),
	.w4(32'hbb8d2271),
	.w5(32'hbb63f4cf),
	.w6(32'hbbb51295),
	.w7(32'hbb83a061),
	.w8(32'h39c74071),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cb233),
	.w1(32'hbb8354c5),
	.w2(32'hbbbab8d1),
	.w3(32'hb9cfe8c8),
	.w4(32'hbbf96fc2),
	.w5(32'hba8db3a6),
	.w6(32'hb890e175),
	.w7(32'hbb07aa2b),
	.w8(32'hbb3c0002),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf299d),
	.w1(32'h3b9864ba),
	.w2(32'hb9edaafe),
	.w3(32'hba4e5c2d),
	.w4(32'hbac6d922),
	.w5(32'hbb97b5e1),
	.w6(32'hbaac8eda),
	.w7(32'h3a691dc0),
	.w8(32'hbb13901a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a466d),
	.w1(32'hbbc5609d),
	.w2(32'h3b215814),
	.w3(32'hbb4924fa),
	.w4(32'hbb9d8622),
	.w5(32'hbba7f9a9),
	.w6(32'hba920388),
	.w7(32'h39ffd69e),
	.w8(32'hbba550d7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb214b64),
	.w1(32'h3bbdf536),
	.w2(32'h3c1d89fd),
	.w3(32'hba033f0e),
	.w4(32'hbb496ce3),
	.w5(32'hbacf430f),
	.w6(32'hbbc7d068),
	.w7(32'hbb5835e8),
	.w8(32'h3b3f190b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeed1b),
	.w1(32'hbb3617cc),
	.w2(32'hbba0a729),
	.w3(32'hbbed8a8b),
	.w4(32'h3c070057),
	.w5(32'hbb9c7ebc),
	.w6(32'hbbd94eb9),
	.w7(32'hb98208da),
	.w8(32'h3b99afa2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9949f8),
	.w1(32'hbc0bd4e0),
	.w2(32'hbaa18dc8),
	.w3(32'hbbc4cb90),
	.w4(32'hbc2cf231),
	.w5(32'hbc84088a),
	.w6(32'hbc10b4d6),
	.w7(32'hbc6257de),
	.w8(32'hbc3e5c22),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef2eee),
	.w1(32'h3abbcf9d),
	.w2(32'hb93f8cb3),
	.w3(32'hbc60a282),
	.w4(32'hb9b05dc0),
	.w5(32'h3b5c4b2b),
	.w6(32'hbc6c9fab),
	.w7(32'h3b082e1f),
	.w8(32'h3ac8b61d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c7cdd),
	.w1(32'h3ba1d373),
	.w2(32'h3c15976a),
	.w3(32'hbbb5c1a6),
	.w4(32'h3bcc6e19),
	.w5(32'h3c102d10),
	.w6(32'hbb27e71c),
	.w7(32'h39c05ae9),
	.w8(32'h3bd75652),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d69d),
	.w1(32'hb994cf26),
	.w2(32'h3b20dda6),
	.w3(32'hbb312a54),
	.w4(32'hbaaa4049),
	.w5(32'hbb17dac7),
	.w6(32'h3af0848a),
	.w7(32'h3a40b152),
	.w8(32'h39fd867d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd4d9a),
	.w1(32'h3aaf95be),
	.w2(32'h3a100e12),
	.w3(32'hba907bc1),
	.w4(32'h3b828114),
	.w5(32'h3c05e7b2),
	.w6(32'h3a94d317),
	.w7(32'hbb418c1f),
	.w8(32'hbbfbf077),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17498b),
	.w1(32'hbbb3c4ff),
	.w2(32'hba8e3ebe),
	.w3(32'hbc47c4f7),
	.w4(32'hbb985c30),
	.w5(32'h3b403b69),
	.w6(32'hbc885505),
	.w7(32'hbaf1260d),
	.w8(32'hbb09e678),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6516e),
	.w1(32'h3c03de74),
	.w2(32'hbb8f1dff),
	.w3(32'hbaaf57fa),
	.w4(32'h3c048c2b),
	.w5(32'hbc1cfd5c),
	.w6(32'hbbb76907),
	.w7(32'h3c727c74),
	.w8(32'h3bfc93c6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b158f),
	.w1(32'h3c5890e6),
	.w2(32'h3c05f763),
	.w3(32'hbbdcb0a9),
	.w4(32'h3c32fa3f),
	.w5(32'hbaf6258f),
	.w6(32'h3bdbac6a),
	.w7(32'h3b8b19c4),
	.w8(32'h3baa1bf2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9699d8),
	.w1(32'h3be122ce),
	.w2(32'h3b40a8cb),
	.w3(32'hbc4e8d56),
	.w4(32'h3bedb31b),
	.w5(32'hbc26f94c),
	.w6(32'hbb213f27),
	.w7(32'h3b88dbea),
	.w8(32'h3ae14aea),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913a1b),
	.w1(32'h3b16ae27),
	.w2(32'hbbedf17e),
	.w3(32'hb710f392),
	.w4(32'hbb65496e),
	.w5(32'hbc05e9cd),
	.w6(32'h3b5a43c2),
	.w7(32'h3b0f86cf),
	.w8(32'hbbbb16bb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeef02),
	.w1(32'h3b0f57ba),
	.w2(32'h3c496e9b),
	.w3(32'h3b5953c0),
	.w4(32'h3c0291ec),
	.w5(32'h3ccde1a7),
	.w6(32'h3c4948fe),
	.w7(32'h3bab8ce3),
	.w8(32'hbb752b99),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46a467),
	.w1(32'h3ac02cf8),
	.w2(32'hbc1b6eca),
	.w3(32'h3c04d860),
	.w4(32'hbb95dbb5),
	.w5(32'h3b43778b),
	.w6(32'hba58f977),
	.w7(32'h3b91e6ec),
	.w8(32'h3bf25cab),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9feb538),
	.w1(32'h3a976039),
	.w2(32'hbc04e29e),
	.w3(32'h3c146778),
	.w4(32'hbb273505),
	.w5(32'hbc40a7d5),
	.w6(32'h3bd7c9c5),
	.w7(32'h3b0a9a3d),
	.w8(32'hbbf9bfea),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221521),
	.w1(32'hbb18377c),
	.w2(32'hbba81659),
	.w3(32'hbb44f784),
	.w4(32'hbaf53b69),
	.w5(32'h39c116b3),
	.w6(32'h3ac102bb),
	.w7(32'h3aa028d1),
	.w8(32'h3bcb6e5b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1624a8),
	.w1(32'hbba3afb3),
	.w2(32'hbc6cc018),
	.w3(32'h3b13b7d1),
	.w4(32'hbc362bcc),
	.w5(32'hbc293b28),
	.w6(32'h3af0c851),
	.w7(32'hbc3785d1),
	.w8(32'hbc09ab0b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5b635),
	.w1(32'hbb6975dc),
	.w2(32'h3b017529),
	.w3(32'hbc6761e5),
	.w4(32'hbaf65eb0),
	.w5(32'h3afedaa7),
	.w6(32'hba6b8b79),
	.w7(32'h3af4d21a),
	.w8(32'hba373ba9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c9c3a),
	.w1(32'hbaeb1b19),
	.w2(32'hbc1200a4),
	.w3(32'h3b6c1016),
	.w4(32'h3a803b43),
	.w5(32'hba651114),
	.w6(32'h3baae041),
	.w7(32'h3b5f331b),
	.w8(32'h3bb548be),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0375df),
	.w1(32'hbb4e04cc),
	.w2(32'hbbcdf9b5),
	.w3(32'h3c3903b0),
	.w4(32'hbb9ff955),
	.w5(32'hbce261eb),
	.w6(32'h3bc5aff2),
	.w7(32'hbb8becdc),
	.w8(32'hbbf60f12),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25bde2),
	.w1(32'h3b5adb97),
	.w2(32'h3bc3e538),
	.w3(32'hbca261d3),
	.w4(32'h3a9a0606),
	.w5(32'h3c046fc5),
	.w6(32'hb909e0d6),
	.w7(32'h3baf89f7),
	.w8(32'h3aac3ecc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0b69),
	.w1(32'hb8d4b8a6),
	.w2(32'h38d0f5d6),
	.w3(32'h3bb5c078),
	.w4(32'h3b05206c),
	.w5(32'hbb574e88),
	.w6(32'hbb42817e),
	.w7(32'hbaece7be),
	.w8(32'hbabee4a4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62c1e),
	.w1(32'hbb9fe2de),
	.w2(32'hbc016bf8),
	.w3(32'h3c29c211),
	.w4(32'hbb955abe),
	.w5(32'h3ad50875),
	.w6(32'h3c38e18c),
	.w7(32'h3b968fd3),
	.w8(32'hb7eaa678),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af17e01),
	.w1(32'hbbb854e0),
	.w2(32'h3b22513a),
	.w3(32'h3b6c88bb),
	.w4(32'h3b9767a1),
	.w5(32'h39ae1009),
	.w6(32'hbb7abe71),
	.w7(32'h3b414a60),
	.w8(32'hbacf727f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf59065),
	.w1(32'hbba05d15),
	.w2(32'hbb440ab9),
	.w3(32'h3af566bb),
	.w4(32'h3b64ba27),
	.w5(32'h3bcd2289),
	.w6(32'hbbb14593),
	.w7(32'h3bf5f062),
	.w8(32'h3bc7e1f3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafb47c),
	.w1(32'hbb615fa2),
	.w2(32'h3b5cff0c),
	.w3(32'h3c10e618),
	.w4(32'hbb71c958),
	.w5(32'h3bf18b1f),
	.w6(32'hb9f6e8b4),
	.w7(32'hbbf90434),
	.w8(32'hb9477cec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8ab9c),
	.w1(32'hbaf89c5c),
	.w2(32'hbad1797e),
	.w3(32'h3bdbd5d8),
	.w4(32'hbb8405bc),
	.w5(32'hbc8d1a2d),
	.w6(32'h3b92d554),
	.w7(32'hbba1ecd4),
	.w8(32'hbc10bb0b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a983ba),
	.w1(32'hbaf3465a),
	.w2(32'h3bcfeaa8),
	.w3(32'hbb8b306f),
	.w4(32'h3c36195b),
	.w5(32'h3c519729),
	.w6(32'h3b35dfb2),
	.w7(32'h3af3f9c9),
	.w8(32'h3b10d788),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e416),
	.w1(32'hbb1b9b3b),
	.w2(32'hbb963126),
	.w3(32'h3b7f13d2),
	.w4(32'hbc4d5647),
	.w5(32'hbcb0fec7),
	.w6(32'h3b60a60b),
	.w7(32'hbc186a03),
	.w8(32'hbc677331),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeedf02),
	.w1(32'hbc20712c),
	.w2(32'h39101063),
	.w3(32'hbc46a550),
	.w4(32'hba5261fe),
	.w5(32'h3c85faaf),
	.w6(32'hb89cd6b2),
	.w7(32'h3b92b1a0),
	.w8(32'hbb069ba9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175dd8),
	.w1(32'h3a1ea044),
	.w2(32'hbc03d793),
	.w3(32'h3b2b0a72),
	.w4(32'hbbbc912e),
	.w5(32'h3aadff39),
	.w6(32'hbb4baa41),
	.w7(32'hbbb6241e),
	.w8(32'h3b5dc523),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b471060),
	.w1(32'h3c0ae6cf),
	.w2(32'h3baa422f),
	.w3(32'h3bcee7c2),
	.w4(32'h3bdb3b0f),
	.w5(32'hbc35e49e),
	.w6(32'h39a19185),
	.w7(32'hb9d2a40a),
	.w8(32'hbbe28ed3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf122dd),
	.w1(32'hbab849ce),
	.w2(32'hbc2ce2d4),
	.w3(32'hbabe6074),
	.w4(32'hbb17aeb3),
	.w5(32'hbc72bf94),
	.w6(32'hbb9f1048),
	.w7(32'hbc295b3a),
	.w8(32'hbbcbb2f9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab401c),
	.w1(32'h3a32017a),
	.w2(32'h3bba82af),
	.w3(32'hbbf85167),
	.w4(32'h3b85002d),
	.w5(32'h3a438227),
	.w6(32'hbb61840c),
	.w7(32'hbc72b7f8),
	.w8(32'hbb0b8a27),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349305),
	.w1(32'hbb1a94c4),
	.w2(32'hbacebfef),
	.w3(32'hbc28a130),
	.w4(32'hbb72ab47),
	.w5(32'h3bbbb9ff),
	.w6(32'h39f07c2d),
	.w7(32'hbb35196d),
	.w8(32'hbaad3e01),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e71c),
	.w1(32'h3a6faabb),
	.w2(32'hbac47fa9),
	.w3(32'hb9a18280),
	.w4(32'h3baf96a1),
	.w5(32'h3bbe999a),
	.w6(32'h3b9fe6f0),
	.w7(32'h3a8fd17c),
	.w8(32'hba3913ae),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5b754),
	.w1(32'hbacb8f63),
	.w2(32'h3b509913),
	.w3(32'h3bcfe45a),
	.w4(32'h3a8f56f8),
	.w5(32'h3b06eee8),
	.w6(32'hba8f7e8a),
	.w7(32'hbc1891e1),
	.w8(32'hbc2397bc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d789),
	.w1(32'h3c1a5604),
	.w2(32'hbc00c59a),
	.w3(32'hbbfc2bef),
	.w4(32'hba28e508),
	.w5(32'hbbc9fd84),
	.w6(32'hbb9949e0),
	.w7(32'hbb643e82),
	.w8(32'hbb167ebd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2258a3),
	.w1(32'hbc53df76),
	.w2(32'h3b94cbcb),
	.w3(32'h38acd360),
	.w4(32'h3b1f036a),
	.w5(32'h3cbb6d48),
	.w6(32'h3b5a750a),
	.w7(32'h3b161020),
	.w8(32'h3ae897a9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982697),
	.w1(32'hbb10993a),
	.w2(32'hbb54541b),
	.w3(32'h3be304fd),
	.w4(32'hb893b977),
	.w5(32'hbc57c70d),
	.w6(32'hbba1d05a),
	.w7(32'hba87a87a),
	.w8(32'hbbbc6d59),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88024d),
	.w1(32'h3c3b05f5),
	.w2(32'h3b9a6295),
	.w3(32'h3a435fb6),
	.w4(32'hbaa1a79e),
	.w5(32'hbb548e5a),
	.w6(32'h3b708c80),
	.w7(32'hbada0dc8),
	.w8(32'h3b875e72),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613bca),
	.w1(32'h3c485fb6),
	.w2(32'h3b4bbccf),
	.w3(32'hbb0c6fff),
	.w4(32'hbbe9c279),
	.w5(32'hbc2e2554),
	.w6(32'h3b1c28b6),
	.w7(32'hbb9b5e60),
	.w8(32'h3b9f5c0f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12c332),
	.w1(32'hbb617353),
	.w2(32'h3b40bfc2),
	.w3(32'hb8fb5881),
	.w4(32'h3b33d0f7),
	.w5(32'h3c8aabe9),
	.w6(32'h3bcb08a5),
	.w7(32'h3aff1000),
	.w8(32'h3aaf0a45),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff48cd),
	.w1(32'hbbb824c9),
	.w2(32'h3b82132d),
	.w3(32'h3b421bc0),
	.w4(32'hbbc4bcc5),
	.w5(32'hbc2e90e7),
	.w6(32'hbbdbc5eb),
	.w7(32'hbb943a86),
	.w8(32'hbb8f7ad8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a7bd),
	.w1(32'h3b6a51f8),
	.w2(32'h3b139b81),
	.w3(32'hbbedc832),
	.w4(32'h3a4435f1),
	.w5(32'hbb94c23a),
	.w6(32'hbb76b5aa),
	.w7(32'hbaa5b330),
	.w8(32'hbb4b4897),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6698b4),
	.w1(32'hba732c98),
	.w2(32'h3bd59fe8),
	.w3(32'hbb62b6b0),
	.w4(32'hbafb4eee),
	.w5(32'hbc2e11fc),
	.w6(32'h3b361515),
	.w7(32'hb986c121),
	.w8(32'hbc0e4330),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898e4a),
	.w1(32'hbb983d8b),
	.w2(32'h3b1e10c2),
	.w3(32'hbb4f4f45),
	.w4(32'h3c3c2f8d),
	.w5(32'h3d18cd36),
	.w6(32'h3b1ddda9),
	.w7(32'h3c0dc22d),
	.w8(32'h3be0ae6d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c520383),
	.w1(32'h3a1738f4),
	.w2(32'h3af321f9),
	.w3(32'h3bf73f4d),
	.w4(32'h3b3f3e59),
	.w5(32'h3bfe75cf),
	.w6(32'hbc0bb37f),
	.w7(32'h3b814a03),
	.w8(32'h39cfbc27),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc146ee),
	.w1(32'hba951955),
	.w2(32'h3c0c0035),
	.w3(32'h3bb74028),
	.w4(32'h3c5bb7c8),
	.w5(32'h3c4f8d45),
	.w6(32'hbb98d451),
	.w7(32'h3bfca718),
	.w8(32'hbbb99d61),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beef88c),
	.w1(32'hbb73ed45),
	.w2(32'h3b35b7f6),
	.w3(32'h3b9b08c1),
	.w4(32'hbba54990),
	.w5(32'hbc43b359),
	.w6(32'hbbf97f60),
	.w7(32'hbba9c455),
	.w8(32'hbb74fea4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ea8b),
	.w1(32'h3ae6d116),
	.w2(32'hbb4d6da2),
	.w3(32'hbc3b725d),
	.w4(32'hbaf294ff),
	.w5(32'hbbe35bca),
	.w6(32'hba0d8ba1),
	.w7(32'h3a46a586),
	.w8(32'hbb9b55ca),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bb286),
	.w1(32'hbb8ece7b),
	.w2(32'hbc2167cd),
	.w3(32'hba344dcb),
	.w4(32'h3bd2ff91),
	.w5(32'hbbcd34cf),
	.w6(32'h3ba8e9ba),
	.w7(32'hbbe7e428),
	.w8(32'hbc6e2e0b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cde79),
	.w1(32'h3cb726cd),
	.w2(32'h3cb90ccc),
	.w3(32'hbc2416f1),
	.w4(32'h3c28a9b3),
	.w5(32'hbc70ac93),
	.w6(32'hbbb496ac),
	.w7(32'hbbcf4455),
	.w8(32'h3a411b66),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc2882),
	.w1(32'hbbb0c29d),
	.w2(32'hbbd08e96),
	.w3(32'hbaf132d8),
	.w4(32'hbbb18a2f),
	.w5(32'hbc1b41eb),
	.w6(32'h3b0fa639),
	.w7(32'hbb81699b),
	.w8(32'hbabd7a79),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f152),
	.w1(32'hbb6fc9e0),
	.w2(32'hbbb331f9),
	.w3(32'hbb9278db),
	.w4(32'hbb7c63b8),
	.w5(32'hbb5135fc),
	.w6(32'hbb493ce3),
	.w7(32'hbab9a388),
	.w8(32'h39e5f43a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc017961),
	.w1(32'h3a902844),
	.w2(32'hbc0fb7d6),
	.w3(32'hbb78bb7d),
	.w4(32'hbb328386),
	.w5(32'h3c45c0a7),
	.w6(32'hbac5ec6a),
	.w7(32'h367222d5),
	.w8(32'hbb08ebf2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe675c),
	.w1(32'h39fa1541),
	.w2(32'hbc1d9fb2),
	.w3(32'hbabfc6d0),
	.w4(32'hbc4135ca),
	.w5(32'hbbf6c7e8),
	.w6(32'h3abd017c),
	.w7(32'hbb067c62),
	.w8(32'h3affb9fc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9765dfe),
	.w1(32'h3b546fb5),
	.w2(32'h3bed3f20),
	.w3(32'h3b6fd904),
	.w4(32'h3bcb327d),
	.w5(32'h3b8a3715),
	.w6(32'h3b88a567),
	.w7(32'h3c30ca65),
	.w8(32'h3b090938),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1deeac),
	.w1(32'h3b915dde),
	.w2(32'hbb989b39),
	.w3(32'h3aae33d5),
	.w4(32'h3ab9eac5),
	.w5(32'hbc182e15),
	.w6(32'h394f3959),
	.w7(32'hbbc4b70d),
	.w8(32'h3a6b36d4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecd06e),
	.w1(32'h38b41e80),
	.w2(32'hbc35b0ed),
	.w3(32'hbac3e23f),
	.w4(32'h3ab74b13),
	.w5(32'hbc29b175),
	.w6(32'h3c3af5a6),
	.w7(32'hba75a2d6),
	.w8(32'h3ba74521),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11991c),
	.w1(32'hbbb9d7a0),
	.w2(32'hbbd5250c),
	.w3(32'h3b52c81e),
	.w4(32'hbaebe75d),
	.w5(32'hbbff0a0d),
	.w6(32'h3b5466ee),
	.w7(32'hbbbae7a0),
	.w8(32'hbb851a4b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d79b),
	.w1(32'h3b66ab7c),
	.w2(32'hbb24cfda),
	.w3(32'hbbcb7ad6),
	.w4(32'hbb2fac87),
	.w5(32'hbc2e9e8c),
	.w6(32'hbb802ad9),
	.w7(32'hbb590de8),
	.w8(32'hbc0c4991),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcde6e),
	.w1(32'hbbde9964),
	.w2(32'hbbed791e),
	.w3(32'hbb9ed390),
	.w4(32'hb9118371),
	.w5(32'h3b778115),
	.w6(32'hba4f9690),
	.w7(32'h3ae5eb16),
	.w8(32'h3b945886),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8e8d),
	.w1(32'hbb0e88cb),
	.w2(32'h3a490d16),
	.w3(32'h3c0e087d),
	.w4(32'h3b524b6e),
	.w5(32'h3c080225),
	.w6(32'h3b8574e5),
	.w7(32'h3b3aee98),
	.w8(32'hbbf93695),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c925a),
	.w1(32'hbbc0846f),
	.w2(32'h3bddd88e),
	.w3(32'hbc06c71d),
	.w4(32'h3aef7452),
	.w5(32'h3d0374d6),
	.w6(32'hbb9e18b5),
	.w7(32'h3bc72c6f),
	.w8(32'h3b86f41d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdcfa7),
	.w1(32'hbbc8226b),
	.w2(32'h3c180822),
	.w3(32'h3bf33dd3),
	.w4(32'h3b556021),
	.w5(32'h3beed3c4),
	.w6(32'hba84cecd),
	.w7(32'h3adce682),
	.w8(32'hba2e4f47),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e72e5),
	.w1(32'hbad5885a),
	.w2(32'hbba9415d),
	.w3(32'hbaced528),
	.w4(32'hbc0f5217),
	.w5(32'hbc61b1bf),
	.w6(32'hbb73dc10),
	.w7(32'hba8ea53a),
	.w8(32'hbb281bc5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f89ca7),
	.w1(32'hbb6de84c),
	.w2(32'h3a8ec1c5),
	.w3(32'h393eb7fc),
	.w4(32'hb92d43bc),
	.w5(32'h3c36c917),
	.w6(32'h3bece3f8),
	.w7(32'h3a6b4543),
	.w8(32'h3b350462),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cc651),
	.w1(32'h3bdb981e),
	.w2(32'h3a471c55),
	.w3(32'hbbaf8021),
	.w4(32'h3994667f),
	.w5(32'hbbb32f4e),
	.w6(32'hbb6e2e37),
	.w7(32'hbc12e84a),
	.w8(32'hbabbb822),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6e06),
	.w1(32'hba8974b3),
	.w2(32'hbb39adea),
	.w3(32'hbc0a72f3),
	.w4(32'hbbe7582e),
	.w5(32'hbba95d33),
	.w6(32'h3b9c9121),
	.w7(32'hbbe49afa),
	.w8(32'hbbddb4ae),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule