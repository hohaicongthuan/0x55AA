module layer_8_featuremap_60(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab06ae2),
	.w1(32'hbb9079f3),
	.w2(32'hbbb8e87d),
	.w3(32'hba66846e),
	.w4(32'hbb88d66d),
	.w5(32'hbbd38f4d),
	.w6(32'hbaa52c1a),
	.w7(32'hbb5e3cbf),
	.w8(32'hbba52b86),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6874d),
	.w1(32'h3b3a5f74),
	.w2(32'h3bbf526d),
	.w3(32'h3b2f5c4f),
	.w4(32'h3b57f349),
	.w5(32'h3ba21773),
	.w6(32'h3b354de3),
	.w7(32'h3b2c0c02),
	.w8(32'h3b7d9ed3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4675c7),
	.w1(32'h3b6d1901),
	.w2(32'h3b9edc35),
	.w3(32'h3b48bcd6),
	.w4(32'h3b822771),
	.w5(32'h3b8b7dc2),
	.w6(32'h3b3f5011),
	.w7(32'h3b247459),
	.w8(32'h3b3539cf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c94f4),
	.w1(32'hbb3230b4),
	.w2(32'hbb4fa084),
	.w3(32'hbad78246),
	.w4(32'hbb911689),
	.w5(32'hbb70b10e),
	.w6(32'hbac1549c),
	.w7(32'hbb5d2d7c),
	.w8(32'hbb3a9480),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e9bd0),
	.w1(32'h3a9c4778),
	.w2(32'h3b59b2df),
	.w3(32'hb9bf40be),
	.w4(32'h3afc5600),
	.w5(32'h3b2ad9ca),
	.w6(32'hb90921ae),
	.w7(32'h3aafef4a),
	.w8(32'h3b1adf63),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2a43),
	.w1(32'h3b175adb),
	.w2(32'h3866a616),
	.w3(32'h3b22d2aa),
	.w4(32'h3b906465),
	.w5(32'h3ab2ade4),
	.w6(32'h3b1b8aa3),
	.w7(32'h3b9209d9),
	.w8(32'hba4017c5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec661d),
	.w1(32'h3964a1c0),
	.w2(32'h397170be),
	.w3(32'h3a055a4d),
	.w4(32'h3a186116),
	.w5(32'h39b38a4e),
	.w6(32'h39cf4a69),
	.w7(32'h39c0e107),
	.w8(32'hb69f9eba),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b309e7c),
	.w1(32'h3b5c336a),
	.w2(32'h3bfd2e55),
	.w3(32'h3926b849),
	.w4(32'h3a0ff054),
	.w5(32'h3b84fd4c),
	.w6(32'h3aa27772),
	.w7(32'h391963c1),
	.w8(32'h3b819de4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f3440),
	.w1(32'h3b85e965),
	.w2(32'h3bc75bea),
	.w3(32'h3ad4483e),
	.w4(32'h3b5595bd),
	.w5(32'h3b8f5002),
	.w6(32'h39ff934e),
	.w7(32'h3ae983fc),
	.w8(32'hb9d0fa58),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae76eb),
	.w1(32'hba92268e),
	.w2(32'h3af497ad),
	.w3(32'h3a98c88e),
	.w4(32'hbaf3dec9),
	.w5(32'hba180201),
	.w6(32'h3b09bfd4),
	.w7(32'h3a815269),
	.w8(32'h3ad6615e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddf659),
	.w1(32'hbb5062c2),
	.w2(32'hbb5adab7),
	.w3(32'hb9c835c4),
	.w4(32'hbb711a51),
	.w5(32'hbb8334c3),
	.w6(32'hba23f68c),
	.w7(32'hbb2851d8),
	.w8(32'hbb528b81),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8b9a6),
	.w1(32'hb9b670da),
	.w2(32'hbb16f421),
	.w3(32'h3ac8ead8),
	.w4(32'hb9328b6f),
	.w5(32'hbb478f28),
	.w6(32'h3b44efd6),
	.w7(32'h3b1fdc8a),
	.w8(32'hb9893104),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fc673),
	.w1(32'h3b4b98df),
	.w2(32'h3b80be60),
	.w3(32'h3afde5a2),
	.w4(32'h3b5f66c3),
	.w5(32'h3b5cfa2e),
	.w6(32'h3b0b9e66),
	.w7(32'h3b2877ff),
	.w8(32'h3b7400da),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a659077),
	.w1(32'h39fe882b),
	.w2(32'h3a6dd57a),
	.w3(32'h3aca7a79),
	.w4(32'h3ab16059),
	.w5(32'h3aaa26d1),
	.w6(32'h3a2cf83f),
	.w7(32'h3aa10083),
	.w8(32'h39abe9a3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00a5d2),
	.w1(32'h399f47bd),
	.w2(32'h3a5d333c),
	.w3(32'h3a42b334),
	.w4(32'h3a3c3b56),
	.w5(32'h3a52b47e),
	.w6(32'h3a1f1a0b),
	.w7(32'h3a889473),
	.w8(32'hb8ab6bff),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9351c50),
	.w1(32'hb8f8d656),
	.w2(32'hb9d1d683),
	.w3(32'hb86febb8),
	.w4(32'h388ddfed),
	.w5(32'hb9e4aff8),
	.w6(32'hb8c8a1ca),
	.w7(32'hb9c126d2),
	.w8(32'hba7998af),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad35607),
	.w1(32'hba803e09),
	.w2(32'hbaaa465b),
	.w3(32'h3ae999ed),
	.w4(32'hba0beebc),
	.w5(32'hbafff1a1),
	.w6(32'hba506bd9),
	.w7(32'hbad609c5),
	.w8(32'hba3253d3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe46a),
	.w1(32'hbb4520c3),
	.w2(32'hba93c66e),
	.w3(32'h376c290b),
	.w4(32'hba42c26e),
	.w5(32'hba366ae9),
	.w6(32'h3aaaa370),
	.w7(32'h3a003fba),
	.w8(32'hb9d9c9ce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd89c64),
	.w1(32'hbbf8c74d),
	.w2(32'hbc028e6d),
	.w3(32'h3ba46753),
	.w4(32'hbc14c431),
	.w5(32'hbc0827df),
	.w6(32'h3c1c65c7),
	.w7(32'h3b098b9b),
	.w8(32'h3b38800b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4667f),
	.w1(32'hbbd84166),
	.w2(32'hbc027416),
	.w3(32'hbb8ef6ea),
	.w4(32'hbb80bbef),
	.w5(32'hbc17fd5a),
	.w6(32'hbb9a91f7),
	.w7(32'hbba46c69),
	.w8(32'hbb437677),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054a27),
	.w1(32'h3b31f915),
	.w2(32'hbafef430),
	.w3(32'h3b83d718),
	.w4(32'h3b9b8a44),
	.w5(32'hba75887d),
	.w6(32'h3baaaf8d),
	.w7(32'h3bc776c1),
	.w8(32'h3a0d83f2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10eb34),
	.w1(32'h3b8c1a27),
	.w2(32'h3bd63fba),
	.w3(32'h3b3611e6),
	.w4(32'h3b993e8d),
	.w5(32'h3bc72ae3),
	.w6(32'h3b4d5251),
	.w7(32'h3b88d3b5),
	.w8(32'h3bb85fad),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16dbfa),
	.w1(32'hbb3c1803),
	.w2(32'hbb771aba),
	.w3(32'h3c2ceb9a),
	.w4(32'hbbfd809a),
	.w5(32'hbbf7df1e),
	.w6(32'h3a95010d),
	.w7(32'hbbce1a82),
	.w8(32'hbb85c615),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37142),
	.w1(32'hbb8f1b0d),
	.w2(32'hbaa026f2),
	.w3(32'hbb6cb7fe),
	.w4(32'hbac5385b),
	.w5(32'hba279bb0),
	.w6(32'hbb1d973a),
	.w7(32'hbaae5f0a),
	.w8(32'hbb2c467f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928d7fc),
	.w1(32'h39d6fd20),
	.w2(32'hb8a8331e),
	.w3(32'hba020aa6),
	.w4(32'hba5bb5bc),
	.w5(32'hba6e7989),
	.w6(32'hb9067285),
	.w7(32'hba8a8f0a),
	.w8(32'h38803376),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df90b8),
	.w1(32'hbb852915),
	.w2(32'hbb8c9978),
	.w3(32'hb99d713d),
	.w4(32'hbbb77934),
	.w5(32'hbc0a9a39),
	.w6(32'hbb1c0162),
	.w7(32'hbb9e8903),
	.w8(32'hbbb3bef9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a14dd),
	.w1(32'hb9059493),
	.w2(32'hb95936ab),
	.w3(32'h3a832409),
	.w4(32'h3962c594),
	.w5(32'h3a03c9a5),
	.w6(32'hb9f0484a),
	.w7(32'hb9ce7158),
	.w8(32'h3a5a6075),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82e95),
	.w1(32'hbbf3b54b),
	.w2(32'hbc773a15),
	.w3(32'hbc07adb8),
	.w4(32'hbd140cb2),
	.w5(32'hbd0b62ad),
	.w6(32'hbd070799),
	.w7(32'hbc688e21),
	.w8(32'hbbdc8485),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92cbfa),
	.w1(32'h3ab2d38f),
	.w2(32'h39538bcb),
	.w3(32'h39dea5de),
	.w4(32'hbb16d3f1),
	.w5(32'hbb0b7a28),
	.w6(32'h3ab3b66d),
	.w7(32'hba73ce51),
	.w8(32'hba6136e5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d9c58),
	.w1(32'h3a8ad71a),
	.w2(32'h3acaa05d),
	.w3(32'h3a6449df),
	.w4(32'h3a93d69c),
	.w5(32'h3a9d5891),
	.w6(32'h3a3be9ef),
	.w7(32'h3a2de11c),
	.w8(32'hb9ab9389),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d83f2),
	.w1(32'hbabf6f09),
	.w2(32'hb9aaf1f7),
	.w3(32'hbad7953f),
	.w4(32'hbb0a2b17),
	.w5(32'hba09a4e6),
	.w6(32'hbaecfb85),
	.w7(32'hbb1f2c05),
	.w8(32'h3b0499ca),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28f783),
	.w1(32'h3b62c7b3),
	.w2(32'h3b0abf77),
	.w3(32'h3b41e67c),
	.w4(32'h3b75783e),
	.w5(32'h3ad8760f),
	.w6(32'h3b0b37d0),
	.w7(32'h3b310d7b),
	.w8(32'h39ba1c3d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2b8d4),
	.w1(32'hbb111b7a),
	.w2(32'hba1b292b),
	.w3(32'hba898b33),
	.w4(32'hbaa044e0),
	.w5(32'hb9e912eb),
	.w6(32'hbad4f4a2),
	.w7(32'hba6e2e52),
	.w8(32'h39c4872b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3daf0d),
	.w1(32'hbae46959),
	.w2(32'hba6eebb9),
	.w3(32'hba9cd8b8),
	.w4(32'hbb15fe09),
	.w5(32'hba85fe2d),
	.w6(32'h3671fbb6),
	.w7(32'hbae0f859),
	.w8(32'h3a3822ab),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25d6b4),
	.w1(32'h39ea2163),
	.w2(32'h3b0f942d),
	.w3(32'h3b55baf2),
	.w4(32'h3bc418a4),
	.w5(32'h3be357ed),
	.w6(32'h3b374d18),
	.w7(32'h3b98fe0e),
	.w8(32'h3b8e2457),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219cd5),
	.w1(32'hbb2fc3f5),
	.w2(32'hbb57e693),
	.w3(32'hbb6d20e8),
	.w4(32'hbb89b324),
	.w5(32'hbba58897),
	.w6(32'hbb537075),
	.w7(32'hba8b58bb),
	.w8(32'hbb31fa38),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a6855),
	.w1(32'h3a3d3613),
	.w2(32'h380165e6),
	.w3(32'hba0116f5),
	.w4(32'hb9a5ecf5),
	.w5(32'hba07f8ea),
	.w6(32'hb8ef9ee0),
	.w7(32'hb9775041),
	.w8(32'h3914a0c5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b561a5f),
	.w1(32'h3b6c91d0),
	.w2(32'h3bb18476),
	.w3(32'h3b3ea2c3),
	.w4(32'h3b452453),
	.w5(32'h3b89f9a8),
	.w6(32'h3b372aec),
	.w7(32'h3b3452bf),
	.w8(32'h3b945800),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7066c0),
	.w1(32'h39cf2752),
	.w2(32'h3af4dee2),
	.w3(32'h3ac88689),
	.w4(32'h3aaed2d3),
	.w5(32'h3adb7b88),
	.w6(32'h3a95b641),
	.w7(32'h3b0f47a1),
	.w8(32'h39b4517b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56394f),
	.w1(32'h399b1bf3),
	.w2(32'h37c6ec82),
	.w3(32'h3acbb1d8),
	.w4(32'h3896e263),
	.w5(32'h36b832b4),
	.w6(32'h3a5da9f2),
	.w7(32'h390e1506),
	.w8(32'h398617c9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eaafa),
	.w1(32'hbbe1d23f),
	.w2(32'hbc5b6496),
	.w3(32'hbb7cd3ba),
	.w4(32'hbc3c5260),
	.w5(32'hbc7e1c93),
	.w6(32'hbb3bb302),
	.w7(32'hbbc7acac),
	.w8(32'hbbf98a78),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28526e),
	.w1(32'h3b86e4be),
	.w2(32'hbc09de4f),
	.w3(32'h3b85499a),
	.w4(32'h3a996418),
	.w5(32'hbab5ac7f),
	.w6(32'h3bb4f845),
	.w7(32'h3a845ad9),
	.w8(32'hbb95f977),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafaf67),
	.w1(32'hbc5b4ab2),
	.w2(32'hbcbc9093),
	.w3(32'hbc6e496e),
	.w4(32'hbd14fcf5),
	.w5(32'hbcc214f8),
	.w6(32'hbcdc206d),
	.w7(32'hbc80828e),
	.w8(32'h38b23357),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ea28),
	.w1(32'hbb3e8dde),
	.w2(32'hbc85401a),
	.w3(32'h3a6f5f19),
	.w4(32'hbbc9e1c1),
	.w5(32'hbc2d0933),
	.w6(32'hba8b2bb2),
	.w7(32'hbbb0e15f),
	.w8(32'h3abc1e8f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c835e78),
	.w1(32'h3ad71924),
	.w2(32'hbc87193b),
	.w3(32'h3c2804e1),
	.w4(32'hbbb9f3ff),
	.w5(32'hbc7e6e7f),
	.w6(32'h3c0e4813),
	.w7(32'hbb86edb1),
	.w8(32'hbb97fe0c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d9e58),
	.w1(32'hbba519c9),
	.w2(32'hbc6d1d86),
	.w3(32'hbaa94cdd),
	.w4(32'hbb9c43eb),
	.w5(32'hbc643ca3),
	.w6(32'hbaa1ce73),
	.w7(32'hbbb9a98f),
	.w8(32'hbb86968a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe383b),
	.w1(32'hbb8646c9),
	.w2(32'hbc4f916a),
	.w3(32'h3c06fef1),
	.w4(32'hbb150283),
	.w5(32'h3a85dce6),
	.w6(32'hbc948bf5),
	.w7(32'hbadb6378),
	.w8(32'h3bccf84f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd32d),
	.w1(32'h3ac99435),
	.w2(32'hbca41a4e),
	.w3(32'hbb8eb528),
	.w4(32'hbbf42015),
	.w5(32'hbc410e56),
	.w6(32'h3c01e5be),
	.w7(32'hbbf913e9),
	.w8(32'hbc6b85bb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb83418),
	.w1(32'hbad09a7c),
	.w2(32'h3d17181e),
	.w3(32'hbc1b5f61),
	.w4(32'hba01b01e),
	.w5(32'h3cca5e75),
	.w6(32'hbc3d56c9),
	.w7(32'h3c4102da),
	.w8(32'h3bb1673f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82ad04),
	.w1(32'h3b8d1cae),
	.w2(32'hbc934aea),
	.w3(32'h3bdbda76),
	.w4(32'hbb1a8858),
	.w5(32'hbc95044f),
	.w6(32'h3bf25de2),
	.w7(32'hbbaee957),
	.w8(32'h39e8fedc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c887324),
	.w1(32'h3c0762cc),
	.w2(32'h3b977a2e),
	.w3(32'h3c51a6bf),
	.w4(32'h3c083034),
	.w5(32'h3bcd0115),
	.w6(32'h3c4bdd0a),
	.w7(32'h3c324142),
	.w8(32'h3c852bfd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf8250),
	.w1(32'hbb8cc128),
	.w2(32'hbca20c9c),
	.w3(32'h3c24d8b7),
	.w4(32'hbc55cfad),
	.w5(32'hbc5d87f1),
	.w6(32'h3c331c03),
	.w7(32'hbbe53eca),
	.w8(32'hbbfa4819),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e638a),
	.w1(32'hbaab275d),
	.w2(32'hbb2b361d),
	.w3(32'h3b85236a),
	.w4(32'hbbf291da),
	.w5(32'hbc9ec868),
	.w6(32'hbcae23ea),
	.w7(32'hbc5ef5ac),
	.w8(32'hbba6540c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe6707),
	.w1(32'hbb86700d),
	.w2(32'h3ba8fa6e),
	.w3(32'h3bce9edf),
	.w4(32'h3a1e6805),
	.w5(32'h3a81c084),
	.w6(32'hb98740ad),
	.w7(32'hbae2c764),
	.w8(32'hbcb54f40),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4cd7a),
	.w1(32'hbc2cbd84),
	.w2(32'hbc908694),
	.w3(32'hbd0c7897),
	.w4(32'hbce7461b),
	.w5(32'hbca2f9b5),
	.w6(32'hbccbe23b),
	.w7(32'hbc487944),
	.w8(32'hbc165838),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4bc50),
	.w1(32'h3ae368d9),
	.w2(32'hbc8e8cd4),
	.w3(32'h3c838215),
	.w4(32'h3b02da68),
	.w5(32'hbc2d67e4),
	.w6(32'hbbe082a4),
	.w7(32'h3b82286f),
	.w8(32'hbc1575ed),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceea7f),
	.w1(32'h3b9209ac),
	.w2(32'hbad62070),
	.w3(32'hbb6ab2e1),
	.w4(32'h37d19c74),
	.w5(32'hbbd8a79f),
	.w6(32'hbc1b34df),
	.w7(32'hba4c9ffa),
	.w8(32'hbb871e66),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcade5c3),
	.w1(32'hbb1cb941),
	.w2(32'hbc3ce723),
	.w3(32'hbbdf6685),
	.w4(32'hbbb122b6),
	.w5(32'hbb859e38),
	.w6(32'h3c19454e),
	.w7(32'h3bdc70cb),
	.w8(32'h3b94f9dd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c763ae7),
	.w1(32'hbafff445),
	.w2(32'h3b61dbeb),
	.w3(32'h3b7a9aa1),
	.w4(32'hbc22ad8e),
	.w5(32'h3ae26b02),
	.w6(32'hbbe57343),
	.w7(32'h3a1f2856),
	.w8(32'hbb93514f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e376a),
	.w1(32'h3a6201aa),
	.w2(32'hbc08d466),
	.w3(32'hbb642783),
	.w4(32'hbc283ea1),
	.w5(32'hbc66c871),
	.w6(32'hbae64c67),
	.w7(32'hbc6d2829),
	.w8(32'hbb819918),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3eec),
	.w1(32'hbb678025),
	.w2(32'hbaf56499),
	.w3(32'hbd0306d5),
	.w4(32'hbc862971),
	.w5(32'hbc7e1901),
	.w6(32'hbc9a23b1),
	.w7(32'hbc210947),
	.w8(32'h3ae9293c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf65397),
	.w1(32'hbb6b8da7),
	.w2(32'hbcbdba0d),
	.w3(32'hbaebc703),
	.w4(32'hba831026),
	.w5(32'hbba27d63),
	.w6(32'h3abd18a2),
	.w7(32'hbc348261),
	.w8(32'h3cad2007),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2ef4c),
	.w1(32'h3b25c06d),
	.w2(32'hbc981518),
	.w3(32'h3ca1c768),
	.w4(32'hba787b0c),
	.w5(32'hbca45efa),
	.w6(32'h3c7db82a),
	.w7(32'hbacb157f),
	.w8(32'hbc6fdfbf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0f719),
	.w1(32'hbcb80c7f),
	.w2(32'hbc4645a5),
	.w3(32'h3b56a11e),
	.w4(32'h3c0c07fb),
	.w5(32'h3d156432),
	.w6(32'h3c814237),
	.w7(32'h3bf3c846),
	.w8(32'h3b2b0979),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c181d2c),
	.w1(32'h3b2ffb69),
	.w2(32'hbbda9a67),
	.w3(32'h3b4d164a),
	.w4(32'hb9356363),
	.w5(32'hbbace5f0),
	.w6(32'h3b144fa5),
	.w7(32'hbaff15f0),
	.w8(32'hba6ed8c9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c3b78),
	.w1(32'hb926f39b),
	.w2(32'hbb76df67),
	.w3(32'hb94497cc),
	.w4(32'hbb0be532),
	.w5(32'hbb283243),
	.w6(32'h39b328a0),
	.w7(32'hba27d4fd),
	.w8(32'h3ad9b4ad),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfdd1d),
	.w1(32'h3a8bab3d),
	.w2(32'hbb90bca3),
	.w3(32'h3b8a9714),
	.w4(32'h3aa1f309),
	.w5(32'hbb2a21f6),
	.w6(32'h3b74eada),
	.w7(32'h392ff7cc),
	.w8(32'h3ba34577),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3cfe3),
	.w1(32'hbc1ef346),
	.w2(32'hbc61261d),
	.w3(32'h3c01ae4d),
	.w4(32'hbb075f8f),
	.w5(32'hbbd2a9d5),
	.w6(32'h3bfda6c4),
	.w7(32'h3c0cf28e),
	.w8(32'h3b340f82),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0de4ba),
	.w1(32'h3b395f51),
	.w2(32'hbc51121d),
	.w3(32'h3b5e9238),
	.w4(32'hbac46140),
	.w5(32'hbc4c6278),
	.w6(32'h3b855b92),
	.w7(32'hbb9cb874),
	.w8(32'h3cbe3d22),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4c7771),
	.w1(32'hbadef800),
	.w2(32'hbd21dbcd),
	.w3(32'h3c85cfe1),
	.w4(32'hbc9427ef),
	.w5(32'hbd021281),
	.w6(32'hba774382),
	.w7(32'hbc27f8c4),
	.w8(32'hbb586dd0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c540f),
	.w1(32'h3b90aa35),
	.w2(32'hbbf029af),
	.w3(32'h3bc7b37d),
	.w4(32'h3b032e62),
	.w5(32'hbb47365b),
	.w6(32'h3b9c9596),
	.w7(32'hba90af1d),
	.w8(32'h3b03b345),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be11aa7),
	.w1(32'h3b2769d4),
	.w2(32'hbc713c9b),
	.w3(32'hbabd5fff),
	.w4(32'hbbaf7b18),
	.w5(32'hbc8d49e1),
	.w6(32'h3b0778e1),
	.w7(32'hbc0530cf),
	.w8(32'hbabaaa3a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3b700),
	.w1(32'h3b93e3ac),
	.w2(32'hbc11564d),
	.w3(32'h3b1ae3fc),
	.w4(32'h37b9c653),
	.w5(32'hbbc4e2a9),
	.w6(32'h3b8482d6),
	.w7(32'hba83e3a3),
	.w8(32'hbc61c728),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f5ee0),
	.w1(32'hbc56f7d1),
	.w2(32'h3cbe67e0),
	.w3(32'h3c580e10),
	.w4(32'hbc07f225),
	.w5(32'hbc603e35),
	.w6(32'hbb42b704),
	.w7(32'h3c9115fd),
	.w8(32'h3ab00a08),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8cdd),
	.w1(32'hbbbff728),
	.w2(32'hbc855e64),
	.w3(32'hbb4eea3d),
	.w4(32'hbc10ba42),
	.w5(32'hbc4eab53),
	.w6(32'h3b053f35),
	.w7(32'hbbe3e894),
	.w8(32'h3b0c3db8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36bd39),
	.w1(32'h3bbf0d73),
	.w2(32'hbba50674),
	.w3(32'h3bb863f4),
	.w4(32'h3a7592c1),
	.w5(32'hbb0ff493),
	.w6(32'h3b255535),
	.w7(32'hbb311e10),
	.w8(32'h3a7c91a4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd68d2),
	.w1(32'hbb24c139),
	.w2(32'hbc581555),
	.w3(32'h3b120d29),
	.w4(32'hbb2533f7),
	.w5(32'hbb8c82bd),
	.w6(32'h3a9d21c1),
	.w7(32'hbb9d8436),
	.w8(32'h3cd53e0b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5ce69b),
	.w1(32'hbb7d368b),
	.w2(32'hbd13b440),
	.w3(32'h3c5e2c98),
	.w4(32'hbcb18647),
	.w5(32'hbce364d5),
	.w6(32'hbb163475),
	.w7(32'hbc3c27ec),
	.w8(32'h3c1d2cd8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0bbfc),
	.w1(32'hb9a41e6b),
	.w2(32'hbcd02d85),
	.w3(32'h3c486787),
	.w4(32'hbbdfa632),
	.w5(32'hbca6b8f1),
	.w6(32'h3bbd3b2c),
	.w7(32'hbbdeb9df),
	.w8(32'h3a37f538),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb07dad),
	.w1(32'hbb0607d9),
	.w2(32'hbb85e4d8),
	.w3(32'hb99ca89c),
	.w4(32'hbb319413),
	.w5(32'h397818e5),
	.w6(32'h3a18e4c3),
	.w7(32'h39a9e779),
	.w8(32'h3b2087f6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca01607),
	.w1(32'hbc1bce34),
	.w2(32'h3cde9c4f),
	.w3(32'h3a0fb963),
	.w4(32'hbbfcadae),
	.w5(32'h399ce2fb),
	.w6(32'hb997e863),
	.w7(32'h3b88e0fa),
	.w8(32'h398eadd7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ecc1c),
	.w1(32'hbb522c42),
	.w2(32'hbc67fa52),
	.w3(32'h39ec56fa),
	.w4(32'hbab2e221),
	.w5(32'hbbd179c0),
	.w6(32'h3a45ebad),
	.w7(32'hbbb0ef08),
	.w8(32'hbc2236ba),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eda3eb),
	.w1(32'hbc2154dd),
	.w2(32'hbcd09910),
	.w3(32'hbc0bc077),
	.w4(32'hbc7a8751),
	.w5(32'hbcb8c74a),
	.w6(32'hbb9a2d44),
	.w7(32'hbc209cbd),
	.w8(32'hbc97ef43),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c7619),
	.w1(32'hbb7e618d),
	.w2(32'hbd05723e),
	.w3(32'hbcc0fd6d),
	.w4(32'hbcc0b0c6),
	.w5(32'hbcf9ffe6),
	.w6(32'hbc53a27e),
	.w7(32'hbc50a657),
	.w8(32'hbb59d7ba),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2db608),
	.w1(32'hbb5e8335),
	.w2(32'hbc08834b),
	.w3(32'hbb66bd40),
	.w4(32'hbc32b171),
	.w5(32'hbca11695),
	.w6(32'hba7eb40e),
	.w7(32'hbc11716e),
	.w8(32'h3b90ef58),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e087f),
	.w1(32'hba92a739),
	.w2(32'hbca954bd),
	.w3(32'h3c17465e),
	.w4(32'hbbbf59d4),
	.w5(32'hbcac47cc),
	.w6(32'h3c151278),
	.w7(32'hbc147da2),
	.w8(32'hbccde573),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf266e9),
	.w1(32'hbb3a8e5d),
	.w2(32'h3d46781b),
	.w3(32'hbc4b6ad7),
	.w4(32'hbae04464),
	.w5(32'h3d02b1d2),
	.w6(32'hbc863f84),
	.w7(32'h3c64f805),
	.w8(32'hbb743fae),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be17dc8),
	.w1(32'h3b9d588a),
	.w2(32'hbbebaac1),
	.w3(32'hbc000224),
	.w4(32'hbbd4b879),
	.w5(32'hbc100e44),
	.w6(32'hba62a5b5),
	.w7(32'hbb0ea3d2),
	.w8(32'h3bd90248),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cbfd),
	.w1(32'hb95ac908),
	.w2(32'hbb0f303c),
	.w3(32'hbb85b433),
	.w4(32'hbba074cf),
	.w5(32'hbb9264b1),
	.w6(32'h3a21a1cd),
	.w7(32'hbbad4888),
	.w8(32'hbc882103),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5a52c),
	.w1(32'hbb0ee907),
	.w2(32'h3d3bc58b),
	.w3(32'hbc51ab3f),
	.w4(32'hbb38913b),
	.w5(32'h3ceb9b40),
	.w6(32'hbc8a5a1e),
	.w7(32'h3c4cb569),
	.w8(32'hbc8442db),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc77057),
	.w1(32'hbb7c41dd),
	.w2(32'h3d160283),
	.w3(32'hbc1a46ac),
	.w4(32'hbb36fbd7),
	.w5(32'h3cbe48fd),
	.w6(32'hbc412aa3),
	.w7(32'h3c2b5abc),
	.w8(32'hba4ba558),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed686),
	.w1(32'h3b023278),
	.w2(32'h3b9133fa),
	.w3(32'h3b7dea10),
	.w4(32'hbb46b7a5),
	.w5(32'hbbaf581a),
	.w6(32'hba4df3a3),
	.w7(32'hbb9123c0),
	.w8(32'hbc1df7bc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cf7b1),
	.w1(32'h3c39f257),
	.w2(32'hbb0220d4),
	.w3(32'hbc04bb40),
	.w4(32'hbc030c5b),
	.w5(32'hbc33f2c1),
	.w6(32'hbbba0419),
	.w7(32'hbb86c9db),
	.w8(32'h3b0944e3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbccc29),
	.w1(32'hbaec65a4),
	.w2(32'hbbb5b359),
	.w3(32'h3b205662),
	.w4(32'hbafa82b1),
	.w5(32'hbb72a556),
	.w6(32'h3ada81ea),
	.w7(32'hbab1fb8a),
	.w8(32'h3b92ee37),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a3bf1),
	.w1(32'h3b53cef2),
	.w2(32'hbb7d7605),
	.w3(32'hbccb587b),
	.w4(32'h3c1d7154),
	.w5(32'h3d159ca0),
	.w6(32'h3b77cf4d),
	.w7(32'hbc54f41d),
	.w8(32'h3c07836b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5415),
	.w1(32'h3ad11627),
	.w2(32'hbba14dc8),
	.w3(32'h3bb89c2d),
	.w4(32'hb91ee122),
	.w5(32'hbc5908d0),
	.w6(32'h3baa17f6),
	.w7(32'hbbe2bb6e),
	.w8(32'hba51aebf),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d165d33),
	.w1(32'h3c1b6cc2),
	.w2(32'hbca2e6ea),
	.w3(32'hbc1ddf87),
	.w4(32'hbc45fcc6),
	.w5(32'hbbf7cffc),
	.w6(32'hbae1d35b),
	.w7(32'hbc126417),
	.w8(32'h3bb4baf9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc516f19),
	.w1(32'h3bad735d),
	.w2(32'h3b33a920),
	.w3(32'hbbe4529e),
	.w4(32'hba45601a),
	.w5(32'h3b44754e),
	.w6(32'h3b4125c0),
	.w7(32'hbbfb0ef7),
	.w8(32'h3cbaea81),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3faaf2),
	.w1(32'hb9f278e6),
	.w2(32'hbcdecb22),
	.w3(32'h3c5ec849),
	.w4(32'hbc54c8dc),
	.w5(32'hbc9430fb),
	.w6(32'h3a7d400d),
	.w7(32'hbbdd498b),
	.w8(32'hbb590868),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6b6c7),
	.w1(32'h3b715359),
	.w2(32'hbc4467c7),
	.w3(32'hba77da0e),
	.w4(32'hbb5799f4),
	.w5(32'hbbf89784),
	.w6(32'hba6edb5d),
	.w7(32'hbb75c480),
	.w8(32'h3a09507f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfacc45),
	.w1(32'hbbb0f580),
	.w2(32'hbb9a72ec),
	.w3(32'hba517a05),
	.w4(32'hbc0e876a),
	.w5(32'hbc1ffb58),
	.w6(32'hbae54868),
	.w7(32'hbbf53a43),
	.w8(32'h3b683d2c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8271),
	.w1(32'h3a1caf30),
	.w2(32'hbb9a3951),
	.w3(32'h3bc527ef),
	.w4(32'h3ab78090),
	.w5(32'hbb56dc95),
	.w6(32'h3b8fe308),
	.w7(32'h3a851b9b),
	.w8(32'h3ccea7dd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6ea2a4),
	.w1(32'h3c18a969),
	.w2(32'hbd470749),
	.w3(32'h3cc702fc),
	.w4(32'hbc0464df),
	.w5(32'hbd1b4e23),
	.w6(32'h3c40bfe5),
	.w7(32'hbc66f3a3),
	.w8(32'h3aa59e65),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec71b3),
	.w1(32'h3acd7d91),
	.w2(32'h3afb6512),
	.w3(32'hb96bb053),
	.w4(32'hbb3641fd),
	.w5(32'hbb20e54d),
	.w6(32'hbb19a5be),
	.w7(32'hbb8bd0c5),
	.w8(32'hbbb150e8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50af8d),
	.w1(32'hb9d15cae),
	.w2(32'h3c9d3d2d),
	.w3(32'hbb91be7a),
	.w4(32'h3ae1fea0),
	.w5(32'h3c6445bc),
	.w6(32'hbbb67444),
	.w7(32'h3bd28a9a),
	.w8(32'h3b3a5880),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac6ed3),
	.w1(32'hbac7177a),
	.w2(32'hbc24e28e),
	.w3(32'hbb76812e),
	.w4(32'hbbe36664),
	.w5(32'hbc03261e),
	.w6(32'hbaab8023),
	.w7(32'hbb59efd5),
	.w8(32'hbc82635e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc554333),
	.w1(32'hbb848956),
	.w2(32'hbbe9e8aa),
	.w3(32'hbc9bb226),
	.w4(32'hbc5c4bd7),
	.w5(32'hbc0130c1),
	.w6(32'hbc461243),
	.w7(32'hbc620e3e),
	.w8(32'hba440d20),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe085b),
	.w1(32'hba80ae34),
	.w2(32'hbc24c626),
	.w3(32'h3b0ce123),
	.w4(32'hb8fd96da),
	.w5(32'hbb18791e),
	.w6(32'hba3f3be8),
	.w7(32'hbb88c0f7),
	.w8(32'hb8e4a6f4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07e71b),
	.w1(32'h3acb1261),
	.w2(32'hbb81f307),
	.w3(32'h39776f17),
	.w4(32'h3aeba0f6),
	.w5(32'h3a0abd2d),
	.w6(32'h3af629a9),
	.w7(32'hba868fc1),
	.w8(32'hbbef6aed),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6c028),
	.w1(32'h3ae3708a),
	.w2(32'h3b35adb1),
	.w3(32'hbba935a1),
	.w4(32'h3b5a5672),
	.w5(32'h3bb2c8e0),
	.w6(32'h3bbaf1ab),
	.w7(32'h3c040a16),
	.w8(32'hbaffc6b2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f61fe),
	.w1(32'hbb985e13),
	.w2(32'hbc23bb44),
	.w3(32'h3b1e685e),
	.w4(32'hbaf8d496),
	.w5(32'hb9b17b82),
	.w6(32'h3b318b4b),
	.w7(32'h3bf74273),
	.w8(32'hbc0e9004),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3f0e),
	.w1(32'hb99b456c),
	.w2(32'hbb736138),
	.w3(32'hbc84e2be),
	.w4(32'hbba3f42d),
	.w5(32'h3a9adb93),
	.w6(32'hba4f4440),
	.w7(32'h3b284203),
	.w8(32'hbc708afe),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc28bbc),
	.w1(32'h3b217e20),
	.w2(32'h3d1ece25),
	.w3(32'hbc68d84f),
	.w4(32'hbae4ee44),
	.w5(32'h3cc3ea75),
	.w6(32'hbb49cca5),
	.w7(32'h3ca3fc15),
	.w8(32'h3b8548bc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59e308),
	.w1(32'h3b2658df),
	.w2(32'hbbb002c6),
	.w3(32'h3851c431),
	.w4(32'h3b1d68cf),
	.w5(32'h39da91d9),
	.w6(32'h3b9a2289),
	.w7(32'h3911ed43),
	.w8(32'h3b1df153),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e5eb),
	.w1(32'hba80d6af),
	.w2(32'hbbc4e3d8),
	.w3(32'h3b15e1b8),
	.w4(32'h38acce35),
	.w5(32'hbb5a4408),
	.w6(32'h3a71fadb),
	.w7(32'hbae88d35),
	.w8(32'h3b70ba3a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c238c51),
	.w1(32'hbac362f8),
	.w2(32'hbc22d459),
	.w3(32'h3b9addab),
	.w4(32'h3a4ff440),
	.w5(32'hbac8fd70),
	.w6(32'hb9371e5f),
	.w7(32'hbb321fe4),
	.w8(32'h3bae7ebd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884adf),
	.w1(32'h3964c1a7),
	.w2(32'hbb193727),
	.w3(32'hbba406ea),
	.w4(32'hbad9abc4),
	.w5(32'hbbee0864),
	.w6(32'hbc168109),
	.w7(32'hbb987a8f),
	.w8(32'hbc8cb0c7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc0a17),
	.w1(32'hb9b50d25),
	.w2(32'h3cc85279),
	.w3(32'hbc59dd21),
	.w4(32'hbad190fc),
	.w5(32'h3c648700),
	.w6(32'h3ac04190),
	.w7(32'h3c94b643),
	.w8(32'hbc7b4d6e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc944c6c),
	.w1(32'hb9e8b957),
	.w2(32'hbc5348c1),
	.w3(32'hbcbf3208),
	.w4(32'hbc44f7ba),
	.w5(32'hbc333857),
	.w6(32'hbb9dd3a2),
	.w7(32'hbc0a06c6),
	.w8(32'h3c81e1cb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9818de),
	.w1(32'h3c27ddc6),
	.w2(32'hbc27f220),
	.w3(32'h3c5436e3),
	.w4(32'h3c558c08),
	.w5(32'h3bdf94f9),
	.w6(32'h3c47049e),
	.w7(32'h3c11e80f),
	.w8(32'h3aadc1b4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a356),
	.w1(32'h3bd07798),
	.w2(32'h3ba919a5),
	.w3(32'h3b8f0018),
	.w4(32'h3bb108c9),
	.w5(32'h39b46269),
	.w6(32'hb95bb0ff),
	.w7(32'hbb2fd48c),
	.w8(32'hbbe77fa6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d4690),
	.w1(32'hbc4ceead),
	.w2(32'hbba56030),
	.w3(32'hbc1af4bc),
	.w4(32'h3a98157d),
	.w5(32'h3be3e7e2),
	.w6(32'hbb8f0322),
	.w7(32'hbacb2990),
	.w8(32'h3c2a21c0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d02f7),
	.w1(32'h3a2dc785),
	.w2(32'hbbc10ad6),
	.w3(32'h3c29a9af),
	.w4(32'hbb74ee98),
	.w5(32'hbb70a65c),
	.w6(32'hbbc349cb),
	.w7(32'hbc15ac7f),
	.w8(32'hbc1877cd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8316aa),
	.w1(32'h3b9aeac9),
	.w2(32'h3c326907),
	.w3(32'hbc1baa9d),
	.w4(32'hbb169e2b),
	.w5(32'hbb845771),
	.w6(32'h380521c3),
	.w7(32'hb9580eb7),
	.w8(32'h3c15acf8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baddefe),
	.w1(32'h3bffe7af),
	.w2(32'h3c42af71),
	.w3(32'hbc7d81d9),
	.w4(32'h3b2b1814),
	.w5(32'hbbbf20e9),
	.w6(32'h3c378bfa),
	.w7(32'h3c8aee80),
	.w8(32'h380af62a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be227b3),
	.w1(32'h3c0a44ad),
	.w2(32'h3a2a6ff2),
	.w3(32'hbbae32bc),
	.w4(32'h3be0114c),
	.w5(32'h3c158a85),
	.w6(32'h3c0a2197),
	.w7(32'h3bafb205),
	.w8(32'h3c5a8556),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ea72b),
	.w1(32'h3c0fad0b),
	.w2(32'hbb7b46db),
	.w3(32'h3c4f8e79),
	.w4(32'h3c297444),
	.w5(32'h3a1f6d1c),
	.w6(32'h3c08568b),
	.w7(32'hba9a06b8),
	.w8(32'hbc064dfb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68829d),
	.w1(32'hbbb119fd),
	.w2(32'h3c3b4677),
	.w3(32'h3af2448c),
	.w4(32'hbabb931a),
	.w5(32'h3c90178c),
	.w6(32'h3b7b6ce4),
	.w7(32'h37f747ec),
	.w8(32'h3a9cd41f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule