module layer_6_featuremap_119(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ecf58),
	.w1(32'hbb0316c9),
	.w2(32'hbac85837),
	.w3(32'hbb416b6b),
	.w4(32'hbb729916),
	.w5(32'hbb47d102),
	.w6(32'hbb6c2f3e),
	.w7(32'hbb77d415),
	.w8(32'hbb71c153),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21cb4),
	.w1(32'hbad7a14e),
	.w2(32'hbab07d66),
	.w3(32'h3a1ef1ab),
	.w4(32'h3a33cc62),
	.w5(32'h39a33bdb),
	.w6(32'h3a91d0a7),
	.w7(32'h3aa4585f),
	.w8(32'h3a8fd465),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8ef13),
	.w1(32'h3a81d02b),
	.w2(32'hb91c7578),
	.w3(32'hbb7da607),
	.w4(32'h3a4e85c7),
	.w5(32'h39e47f62),
	.w6(32'h3a5fbbdd),
	.w7(32'h3abeec09),
	.w8(32'hbb0a65db),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20544b),
	.w1(32'hb8830eb4),
	.w2(32'hb9ba1d52),
	.w3(32'h3ad6cf12),
	.w4(32'h3b012152),
	.w5(32'h3aed855a),
	.w6(32'h3a97ac02),
	.w7(32'h3a9c0154),
	.w8(32'h3aaf81e2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e2cbd),
	.w1(32'h3aa82362),
	.w2(32'hba009972),
	.w3(32'h3b810780),
	.w4(32'h3afef51d),
	.w5(32'h3b34cf2c),
	.w6(32'h3b4d413b),
	.w7(32'h3983b05e),
	.w8(32'hba2aa4b6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39572525),
	.w1(32'hbb086186),
	.w2(32'hbb014930),
	.w3(32'hbbaa451a),
	.w4(32'hbbb921c8),
	.w5(32'hbbae4059),
	.w6(32'hbb8316d2),
	.w7(32'hbb897b2a),
	.w8(32'hbb87725d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8218e),
	.w1(32'h3aa6c3cb),
	.w2(32'h3a31c669),
	.w3(32'h3be23626),
	.w4(32'h3be8c6ec),
	.w5(32'h3bd23e2b),
	.w6(32'h3b8b3aa5),
	.w7(32'h3b83c4ec),
	.w8(32'h3b838e08),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82de30),
	.w1(32'h3ad1457a),
	.w2(32'h3b109d01),
	.w3(32'h3b001d2c),
	.w4(32'hb9f617c3),
	.w5(32'hb93ad2cd),
	.w6(32'h392aa1b7),
	.w7(32'h3afb508d),
	.w8(32'h3a38468c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a827f),
	.w1(32'h3b2c3196),
	.w2(32'hbab051fc),
	.w3(32'h3aae53e0),
	.w4(32'h3a9ff532),
	.w5(32'h3abb31c0),
	.w6(32'h3b83627c),
	.w7(32'h3b1cde25),
	.w8(32'h3a2fee54),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f4c2),
	.w1(32'h394424e1),
	.w2(32'h39b119ec),
	.w3(32'hbb1bfc2c),
	.w4(32'hbb281fbb),
	.w5(32'hbb064e75),
	.w6(32'hbab2508b),
	.w7(32'hbaa7f89e),
	.w8(32'hba815b5f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54f4d5),
	.w1(32'hb89a7a42),
	.w2(32'hbb1c8e8e),
	.w3(32'hb9c4ffee),
	.w4(32'hbb50c8f3),
	.w5(32'hb9a00918),
	.w6(32'hbae8a75e),
	.w7(32'hbb23e5ef),
	.w8(32'hbb2ed970),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5b5d6),
	.w1(32'hba8361c6),
	.w2(32'hba3d9278),
	.w3(32'hba13582a),
	.w4(32'hba1aa4ea),
	.w5(32'hb9875688),
	.w6(32'hbaf3a625),
	.w7(32'hbaea757f),
	.w8(32'hba8c1c14),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f847bb),
	.w1(32'h39df2ef2),
	.w2(32'h3a187f3d),
	.w3(32'h3a912456),
	.w4(32'h3acea38c),
	.w5(32'h3a8e76c3),
	.w6(32'h3a775ce0),
	.w7(32'h3aae6366),
	.w8(32'h3a7607da),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35e543),
	.w1(32'h3ba0796f),
	.w2(32'h3b8e6f89),
	.w3(32'h3aec9af5),
	.w4(32'h3b2cb3e9),
	.w5(32'h3b0b2fe7),
	.w6(32'h3b8262d9),
	.w7(32'h3ae7ce4c),
	.w8(32'hba18ee7d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27dfd7),
	.w1(32'hb863d41c),
	.w2(32'hb83aaaca),
	.w3(32'h3ae856b9),
	.w4(32'h3ada30eb),
	.w5(32'h3ae37e53),
	.w6(32'h3a4e0c5e),
	.w7(32'h3a826287),
	.w8(32'h3a18c295),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9390d40),
	.w1(32'hb95c309a),
	.w2(32'hba77e164),
	.w3(32'hbad95621),
	.w4(32'hbae92136),
	.w5(32'hbaf6bebc),
	.w6(32'hbad5799c),
	.w7(32'hbb00b16c),
	.w8(32'hbb24d2b1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4bb38),
	.w1(32'h3b8423cc),
	.w2(32'h3ac64fe1),
	.w3(32'h39603259),
	.w4(32'h385e6558),
	.w5(32'hb9c3d535),
	.w6(32'h3b2b476d),
	.w7(32'h3a0edcde),
	.w8(32'hba4878ba),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964c02b),
	.w1(32'h3a2d24eb),
	.w2(32'h3a1ba8ee),
	.w3(32'hba3be852),
	.w4(32'hba928ce5),
	.w5(32'hba99b27b),
	.w6(32'hba8339ae),
	.w7(32'hba93560d),
	.w8(32'hba8f016b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c1265),
	.w1(32'hbaa27356),
	.w2(32'hbab4ae99),
	.w3(32'h38a8f698),
	.w4(32'h393fef14),
	.w5(32'hb5ae5015),
	.w6(32'hba4c3710),
	.w7(32'hba3d1be7),
	.w8(32'hba1ea1c3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba718a0c),
	.w1(32'hb94cfbff),
	.w2(32'hb98745fd),
	.w3(32'hba6d5df0),
	.w4(32'hbac5aed8),
	.w5(32'h3a98b682),
	.w6(32'hbad38db8),
	.w7(32'hbaa8ef20),
	.w8(32'hb8f55146),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d5306),
	.w1(32'hb9f72cb9),
	.w2(32'hba244bd8),
	.w3(32'h39b9490c),
	.w4(32'h39c1b2d0),
	.w5(32'h39757634),
	.w6(32'h391cd209),
	.w7(32'h391ce4b4),
	.w8(32'h38a2a2e8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a856760),
	.w1(32'h3b4383dd),
	.w2(32'hba32e607),
	.w3(32'hbb0037b0),
	.w4(32'hbab949f3),
	.w5(32'hba4c43fa),
	.w6(32'h3a566585),
	.w7(32'hbb01f6a7),
	.w8(32'hbb293647),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c0c55),
	.w1(32'hba68d7e1),
	.w2(32'hba73e24c),
	.w3(32'hb98c5b39),
	.w4(32'h37953d23),
	.w5(32'hbb05bd28),
	.w6(32'h3a1bfeba),
	.w7(32'h398945d9),
	.w8(32'hba65f66a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2623c7),
	.w1(32'h3adc5070),
	.w2(32'h3a59d36c),
	.w3(32'hbb3767dc),
	.w4(32'hbb7a3f48),
	.w5(32'hb9d28f67),
	.w6(32'hba3e0b49),
	.w7(32'hbb67dac5),
	.w8(32'hbb33eb8a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658ff3),
	.w1(32'h3ad05d51),
	.w2(32'h3a4dc121),
	.w3(32'hbaf75c78),
	.w4(32'h3a754a9d),
	.w5(32'h3b10c992),
	.w6(32'hba162a8c),
	.w7(32'hba660f73),
	.w8(32'hbb27eb7e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b76cc),
	.w1(32'h3a793949),
	.w2(32'hb9504b66),
	.w3(32'h39b9b210),
	.w4(32'h3a3b8149),
	.w5(32'h3a1bb250),
	.w6(32'h3a1c3588),
	.w7(32'h3a58d863),
	.w8(32'h3a9fc9ca),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39993cb1),
	.w1(32'h3b3f6c04),
	.w2(32'h3acfcc34),
	.w3(32'h3a4398d8),
	.w4(32'h3919bc75),
	.w5(32'h3b11915e),
	.w6(32'h39653cbf),
	.w7(32'hbaa36c2b),
	.w8(32'hba64ee69),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2708b1),
	.w1(32'h3a933f5e),
	.w2(32'hb93793c2),
	.w3(32'h3b847fca),
	.w4(32'h3ba8ae0c),
	.w5(32'h3b94e0e0),
	.w6(32'h3b292915),
	.w7(32'h3b3574ce),
	.w8(32'h3b2f7c0d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d829a8),
	.w1(32'h390bfc62),
	.w2(32'h39383214),
	.w3(32'h39132b4b),
	.w4(32'h398f4d07),
	.w5(32'h3a0993e7),
	.w6(32'h3807cd63),
	.w7(32'hb6e990ed),
	.w8(32'h3951311e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb30ca8),
	.w1(32'hbadd35e9),
	.w2(32'hbbaaa1b2),
	.w3(32'h3c31a1d2),
	.w4(32'hba537240),
	.w5(32'hbb67284c),
	.w6(32'hbbe6bdde),
	.w7(32'hbbe4a1c7),
	.w8(32'hbaf49e75),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2812),
	.w1(32'hbb47a6a2),
	.w2(32'hbbc41366),
	.w3(32'hbaa6aae1),
	.w4(32'hbb2fef06),
	.w5(32'hbb502ac1),
	.w6(32'hbb3bb1a4),
	.w7(32'hbbdb15b2),
	.w8(32'hbbc356e8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75315),
	.w1(32'hb9353257),
	.w2(32'hbb0be722),
	.w3(32'hbab0835b),
	.w4(32'hbb14f584),
	.w5(32'hbaf2752f),
	.w6(32'hb9572188),
	.w7(32'hbad2c192),
	.w8(32'hbadc045e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c9fa4),
	.w1(32'hba02f35d),
	.w2(32'hba8ab96a),
	.w3(32'hba478b9e),
	.w4(32'hbaa90db3),
	.w5(32'hbb381e1f),
	.w6(32'hba08b31e),
	.w7(32'h3a283b29),
	.w8(32'hbae8ec9a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4f6f0),
	.w1(32'h3a9d8855),
	.w2(32'hbb1870ca),
	.w3(32'hbabd8d4a),
	.w4(32'hbb4c8611),
	.w5(32'hba4c6c1f),
	.w6(32'hb9bfe1b6),
	.w7(32'hb969f026),
	.w8(32'hbb258c61),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba966aa0),
	.w1(32'hba8f31ce),
	.w2(32'hbaa829b1),
	.w3(32'hbb7e04a0),
	.w4(32'hbb8548b1),
	.w5(32'hbb7ab026),
	.w6(32'hbb07f620),
	.w7(32'hbb120f58),
	.w8(32'hbb042547),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38716738),
	.w1(32'hb8356ffa),
	.w2(32'h3b1976d1),
	.w3(32'hb8973651),
	.w4(32'h3b7c534f),
	.w5(32'h3a776952),
	.w6(32'hbb3ad0be),
	.w7(32'hba04ff72),
	.w8(32'hb9dded1b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872739),
	.w1(32'hb9823a8b),
	.w2(32'hb9c6730f),
	.w3(32'hba425b09),
	.w4(32'hbab18613),
	.w5(32'hba6a79df),
	.w6(32'hba8dfc88),
	.w7(32'hbae6a6a9),
	.w8(32'hbac87d7f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3c5cd),
	.w1(32'hba06648d),
	.w2(32'hba45618a),
	.w3(32'h3aea6067),
	.w4(32'h3ab942c9),
	.w5(32'h3a0b31b9),
	.w6(32'hb994a597),
	.w7(32'hb88ddf84),
	.w8(32'h3a1803d1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b89c5),
	.w1(32'h3a503d98),
	.w2(32'h3a7eb1a2),
	.w3(32'h3a157678),
	.w4(32'h3b157df2),
	.w5(32'h3969836f),
	.w6(32'h3ac7305e),
	.w7(32'hb98ed435),
	.w8(32'h398db666),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5751f),
	.w1(32'h3bbc61c5),
	.w2(32'h3b1bef70),
	.w3(32'hbabad566),
	.w4(32'h3b1def1f),
	.w5(32'h3bc989af),
	.w6(32'h3b311ab2),
	.w7(32'hba8bec2d),
	.w8(32'hbaa29af9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa619),
	.w1(32'hbb40fe46),
	.w2(32'hbb388e35),
	.w3(32'hbb0b382b),
	.w4(32'h39fea231),
	.w5(32'h3b27dfaa),
	.w6(32'hbab24d0f),
	.w7(32'hba07456b),
	.w8(32'h3b2cf4e8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac75ac2),
	.w1(32'hba4a5df0),
	.w2(32'hba816dc0),
	.w3(32'h3aff419a),
	.w4(32'h3b085d8f),
	.w5(32'h3ac4fff9),
	.w6(32'h38c9be88),
	.w7(32'h3a262944),
	.w8(32'h3aa5f44e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9bc22),
	.w1(32'h3adb4550),
	.w2(32'h3a88e0ff),
	.w3(32'h3a4b9e9f),
	.w4(32'hb8fdf1a3),
	.w5(32'hb8af1e70),
	.w6(32'h3aa29ac1),
	.w7(32'h3a67a45e),
	.w8(32'h3a0e66c1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d6dd),
	.w1(32'hbae8a1c7),
	.w2(32'hbb9f4701),
	.w3(32'h3c01623e),
	.w4(32'hb8bdc457),
	.w5(32'hbbbd5c65),
	.w6(32'hbc10b1e0),
	.w7(32'hbbfa6a5a),
	.w8(32'hba5d8d3e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad069e1),
	.w1(32'h3b793944),
	.w2(32'h3ae6d87d),
	.w3(32'h38e4189c),
	.w4(32'h3b1e3ea4),
	.w5(32'h3b55337c),
	.w6(32'h3af1c49d),
	.w7(32'hb8e42057),
	.w8(32'hbada9105),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d0847),
	.w1(32'hbab8f439),
	.w2(32'h39b809f3),
	.w3(32'h39f03602),
	.w4(32'h37a09258),
	.w5(32'hbadf4589),
	.w6(32'h3b03f847),
	.w7(32'h3a552cdd),
	.w8(32'h39c006ef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba829461),
	.w1(32'hbb464b0c),
	.w2(32'hbb6b82b6),
	.w3(32'h395345f6),
	.w4(32'hb84c1ea2),
	.w5(32'h3b475f20),
	.w6(32'h3a2388e9),
	.w7(32'h3941b821),
	.w8(32'h3a5a0d7b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9bdae),
	.w1(32'hbae86fe6),
	.w2(32'hbbce33a9),
	.w3(32'hba5b3852),
	.w4(32'hbbce8f40),
	.w5(32'hbb976e7b),
	.w6(32'hba386590),
	.w7(32'hbbd0abcf),
	.w8(32'hbba26eaf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592c4b),
	.w1(32'hbaaf913d),
	.w2(32'hba6473cf),
	.w3(32'hbac836cb),
	.w4(32'hba9b8c18),
	.w5(32'hba9e4f74),
	.w6(32'hba8e41a5),
	.w7(32'hba51952c),
	.w8(32'hba68cbc9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb616b62),
	.w1(32'hbb3d272c),
	.w2(32'hbb2560e2),
	.w3(32'hba994835),
	.w4(32'hbae06b8e),
	.w5(32'h3a7b3a69),
	.w6(32'hbb8d5d6f),
	.w7(32'hbbd135fd),
	.w8(32'hbba8c028),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeda3a6),
	.w1(32'h39437262),
	.w2(32'hbab3ba07),
	.w3(32'h3aadf6e7),
	.w4(32'h3ae57460),
	.w5(32'h3ade7d97),
	.w6(32'h3accc52b),
	.w7(32'h3aada6f0),
	.w8(32'h3b018ed5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3c0b5),
	.w1(32'h39c35bc8),
	.w2(32'h3afe5f9b),
	.w3(32'h3a893c3b),
	.w4(32'h3b792ad5),
	.w5(32'h3b8c3ebd),
	.w6(32'h3a8e3598),
	.w7(32'h3b547f9f),
	.w8(32'h3b817112),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34017c),
	.w1(32'h3ba099b7),
	.w2(32'h3afbad80),
	.w3(32'h3b6efeed),
	.w4(32'h3bb2cb95),
	.w5(32'h3b8c1e0a),
	.w6(32'h3b8cfd18),
	.w7(32'h3b65dac4),
	.w8(32'h3a0a95fa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afc012),
	.w1(32'hba8095e8),
	.w2(32'hbaae26b1),
	.w3(32'h3bd4fc98),
	.w4(32'h3bbecad0),
	.w5(32'h3ba6bc52),
	.w6(32'h3b619d22),
	.w7(32'h3b3ed5e1),
	.w8(32'h3ac7ef27),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2abd88),
	.w1(32'h38e71b06),
	.w2(32'hba3393f6),
	.w3(32'h3aae5d26),
	.w4(32'h3b003c32),
	.w5(32'h3adbe7ce),
	.w6(32'h3b2df38a),
	.w7(32'h3b3878c1),
	.w8(32'h3b384ce3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f9088),
	.w1(32'hbbebe549),
	.w2(32'hbc448cd5),
	.w3(32'h3c5297af),
	.w4(32'h3cda06eb),
	.w5(32'h3cb4458e),
	.w6(32'h3cc56ff3),
	.w7(32'h3cbc9587),
	.w8(32'h3b896703),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15246d),
	.w1(32'hbaec7b40),
	.w2(32'h3b095905),
	.w3(32'hbc8bc55d),
	.w4(32'hbc62014c),
	.w5(32'hbc1ffac8),
	.w6(32'hbbb23bc1),
	.w7(32'h3b6406bf),
	.w8(32'h3b29f6a8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12b080),
	.w1(32'hbae478f0),
	.w2(32'hbc68f63d),
	.w3(32'hbbbe9cfb),
	.w4(32'hbc80156c),
	.w5(32'hbc97e42b),
	.w6(32'hbae229f5),
	.w7(32'h3b1f2c62),
	.w8(32'h3a9af3fc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb940c3),
	.w1(32'hbbfce04f),
	.w2(32'hbc06f624),
	.w3(32'h3b4acf2f),
	.w4(32'hb9d24d5f),
	.w5(32'hbadb6dcc),
	.w6(32'hbb7f7d5e),
	.w7(32'hbbc6cd25),
	.w8(32'hbbf0ba2c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdce147),
	.w1(32'h3c5e9cc5),
	.w2(32'h3caa2b28),
	.w3(32'hbcdc360c),
	.w4(32'h39ef721c),
	.w5(32'h3c1420c5),
	.w6(32'h3d16ecea),
	.w7(32'h3cefdf25),
	.w8(32'h3a418b91),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38274e),
	.w1(32'hbaf52d4f),
	.w2(32'hbc43612c),
	.w3(32'h3bfe8455),
	.w4(32'h3b361d50),
	.w5(32'hbadb5a96),
	.w6(32'h3b2be586),
	.w7(32'hbbcf598d),
	.w8(32'hbc2add7b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf65925),
	.w1(32'hbbb5b035),
	.w2(32'hba34c2f3),
	.w3(32'hbb5d1a72),
	.w4(32'hbc17442c),
	.w5(32'h3aea5f36),
	.w6(32'h3b7aa877),
	.w7(32'h3c821435),
	.w8(32'h3c680fa5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe40877),
	.w1(32'h3c345b60),
	.w2(32'h3cfe4743),
	.w3(32'hbc54b125),
	.w4(32'hbcb34738),
	.w5(32'hbce5d3e0),
	.w6(32'h3b127202),
	.w7(32'h3c21d836),
	.w8(32'h3c963b78),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbce4c),
	.w1(32'hbbd683f7),
	.w2(32'hbc653971),
	.w3(32'h3cb2e5f6),
	.w4(32'h3c9f7426),
	.w5(32'h3c688e62),
	.w6(32'h39c3181c),
	.w7(32'hbc462777),
	.w8(32'hbc17c6b1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule