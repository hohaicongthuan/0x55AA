module layer_8_featuremap_17(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1173ac),
	.w1(32'h3b154431),
	.w2(32'h3b84916d),
	.w3(32'hbbdcb97d),
	.w4(32'h3bed5c3e),
	.w5(32'h3c242d75),
	.w6(32'hbb434772),
	.w7(32'h3bf3e405),
	.w8(32'h3904c9c8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c1d8),
	.w1(32'hbae49918),
	.w2(32'hbb327e94),
	.w3(32'h3ba74877),
	.w4(32'hbbcf9148),
	.w5(32'hbb80d66d),
	.w6(32'h3bf3bbc3),
	.w7(32'hbba00d11),
	.w8(32'h3b00bab7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a9e15),
	.w1(32'hbb951f00),
	.w2(32'hbc47fb1f),
	.w3(32'h3a81f2b6),
	.w4(32'hb94f9192),
	.w5(32'hbbd781d9),
	.w6(32'h3bd1d003),
	.w7(32'h3bb6151b),
	.w8(32'hbb88256d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67728a),
	.w1(32'h3c595f4f),
	.w2(32'h3bce9efc),
	.w3(32'h3c401e7c),
	.w4(32'h3c5fcdcf),
	.w5(32'h3be12945),
	.w6(32'h3aea0f6e),
	.w7(32'h3ca10969),
	.w8(32'h3beb92ce),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bef08),
	.w1(32'hbb262497),
	.w2(32'hbaa7db22),
	.w3(32'h3b004377),
	.w4(32'hbb2d8682),
	.w5(32'hba07e8d2),
	.w6(32'h3a15cef1),
	.w7(32'hbb298f10),
	.w8(32'h3b241be9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b9582),
	.w1(32'hbc852b74),
	.w2(32'hbb2ae490),
	.w3(32'h3c2001e0),
	.w4(32'hbc01d00c),
	.w5(32'hbb1e38b2),
	.w6(32'h3aff937f),
	.w7(32'hbb699b1f),
	.w8(32'h3b44bd6b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1522),
	.w1(32'hbb3dfea8),
	.w2(32'h3ab527f7),
	.w3(32'hbb70d0ba),
	.w4(32'hbab26d9e),
	.w5(32'hbba305a4),
	.w6(32'h3b966393),
	.w7(32'h3b82ddfb),
	.w8(32'h3a3ca5e4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba63d0e),
	.w1(32'hbc483125),
	.w2(32'hbc1f0564),
	.w3(32'h3cb61f70),
	.w4(32'h3c27f8a1),
	.w5(32'h3ba83bbd),
	.w6(32'h3b76bbc7),
	.w7(32'h3c0cd183),
	.w8(32'h3be1799d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb313f6d),
	.w1(32'hbbad0a64),
	.w2(32'hbbe6b896),
	.w3(32'hba0bd86f),
	.w4(32'hbb9816f3),
	.w5(32'hbb7d9fab),
	.w6(32'h3b659bb8),
	.w7(32'h3bc5503c),
	.w8(32'h3bbfa3b2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d0e5),
	.w1(32'h3c044d99),
	.w2(32'h3b990265),
	.w3(32'hbb5ebfb5),
	.w4(32'h3bd4a517),
	.w5(32'h3b8b73df),
	.w6(32'hbb3366cf),
	.w7(32'h3c14819b),
	.w8(32'h3b1cb58e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e324),
	.w1(32'h3c08e5ff),
	.w2(32'hbb874341),
	.w3(32'h3aa284e3),
	.w4(32'h3c8ced79),
	.w5(32'h3c854dff),
	.w6(32'h3c870be8),
	.w7(32'h3b7d0045),
	.w8(32'h3cac5e5e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e87b01),
	.w1(32'h3b928fe8),
	.w2(32'h3be0fbdb),
	.w3(32'h398333fa),
	.w4(32'h3c652256),
	.w5(32'h3c367dd3),
	.w6(32'hbbc0b42f),
	.w7(32'hbbbae18a),
	.w8(32'h3b8e5001),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d30ee),
	.w1(32'hbb50f7a3),
	.w2(32'h3b83cc4f),
	.w3(32'h3ba49a3b),
	.w4(32'hba807273),
	.w5(32'hbbc0bf63),
	.w6(32'h3bc06d26),
	.w7(32'h3bd3e465),
	.w8(32'hbb94c48b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2255e0),
	.w1(32'h3b7ed6e7),
	.w2(32'hbb06dda0),
	.w3(32'h3adfb237),
	.w4(32'h3b8caaa4),
	.w5(32'hbbf8dd5f),
	.w6(32'hbb008f06),
	.w7(32'h3ca76464),
	.w8(32'h3afaedfc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4de8c0),
	.w1(32'hba267dcc),
	.w2(32'hbc157407),
	.w3(32'hbb4b558e),
	.w4(32'hbb8bcddf),
	.w5(32'h3b9c756d),
	.w6(32'h3c97c595),
	.w7(32'h3b006c7d),
	.w8(32'hbba727bd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fbaa1),
	.w1(32'h3b4241cb),
	.w2(32'h3c108cb7),
	.w3(32'hbba4d8ea),
	.w4(32'hbbf7a596),
	.w5(32'hbc0869d6),
	.w6(32'hbaf8b574),
	.w7(32'h3b17f2d6),
	.w8(32'h3b250a64),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa1c4),
	.w1(32'hbb2ece6f),
	.w2(32'hbb0914d5),
	.w3(32'h3ba10727),
	.w4(32'h3bc5b128),
	.w5(32'h3c8a124e),
	.w6(32'h3bbd8752),
	.w7(32'h391fb68c),
	.w8(32'h3c13128a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e2dec),
	.w1(32'h3c33e4c8),
	.w2(32'hbab0bc7b),
	.w3(32'h3b3cd788),
	.w4(32'h3b92d2dc),
	.w5(32'h3c857b14),
	.w6(32'hbbec8ab4),
	.w7(32'hbb8fac79),
	.w8(32'hbb9a8efa),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b258ffd),
	.w1(32'h3b842681),
	.w2(32'hba7b6d29),
	.w3(32'hbc69b2c9),
	.w4(32'h3d9433bb),
	.w5(32'h3d289e85),
	.w6(32'hbc90652b),
	.w7(32'h3b2e4517),
	.w8(32'hbbf76d78),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bddf6),
	.w1(32'h3b5e5eed),
	.w2(32'h3cc6ad8f),
	.w3(32'hbc10eeae),
	.w4(32'h3bf8dce6),
	.w5(32'h3bfa9920),
	.w6(32'hbc496e93),
	.w7(32'hbc5ca9dc),
	.w8(32'h3c610a73),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35fb22),
	.w1(32'h3c819467),
	.w2(32'h3c590dd3),
	.w3(32'hbc564c24),
	.w4(32'h3b5808af),
	.w5(32'h3cc074e8),
	.w6(32'hbca88c0a),
	.w7(32'hbc4f5820),
	.w8(32'h3c628914),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab9239),
	.w1(32'h3c1ff6c8),
	.w2(32'hbb7ab74c),
	.w3(32'hba89313d),
	.w4(32'hbc1cfd64),
	.w5(32'hbc36a9ae),
	.w6(32'h3c54d73e),
	.w7(32'hbb1702d9),
	.w8(32'hbb6c67b9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc903c82),
	.w1(32'hbc4c44a0),
	.w2(32'h39dc8c66),
	.w3(32'hbd434e67),
	.w4(32'h3cd09ea1),
	.w5(32'h3d1abc29),
	.w6(32'hbcc2cd5a),
	.w7(32'h3c59128c),
	.w8(32'h3cad992a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0acb),
	.w1(32'hbb4925b9),
	.w2(32'h3b34db0e),
	.w3(32'hbbc967d9),
	.w4(32'hbbb9cd78),
	.w5(32'hbbf2dd68),
	.w6(32'hb9b39fec),
	.w7(32'h38b99836),
	.w8(32'h3b3d36e7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc72d2e),
	.w1(32'h3bcd5132),
	.w2(32'hbb889578),
	.w3(32'h3a7e59aa),
	.w4(32'h3c8f4fcf),
	.w5(32'hbc4a5c36),
	.w6(32'hb94e8b53),
	.w7(32'h3c654b00),
	.w8(32'h3b6bfdb7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd227e5),
	.w1(32'hbb30669e),
	.w2(32'hbace563f),
	.w3(32'hbc8518c6),
	.w4(32'h3b4bd798),
	.w5(32'h3cf7872e),
	.w6(32'hbc1a7ce9),
	.w7(32'hbb30d2c1),
	.w8(32'h3c8a0cc1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45eeeb),
	.w1(32'hbb60244c),
	.w2(32'hbbc39176),
	.w3(32'h3c067be2),
	.w4(32'h3b523b9d),
	.w5(32'h3af2a9e6),
	.w6(32'h3b5de110),
	.w7(32'h39d244f6),
	.w8(32'hbaec09b0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e0e1f52),
	.w1(32'h3d0857b8),
	.w2(32'hbda172fc),
	.w3(32'hbd89b334),
	.w4(32'h3cafdf0d),
	.w5(32'h3e745215),
	.w6(32'hbcc50e8e),
	.w7(32'h3d593ca1),
	.w8(32'h3d55fbf8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad7e01),
	.w1(32'h3a3ec06f),
	.w2(32'hbacae024),
	.w3(32'h3ade65a9),
	.w4(32'h3ccc4e67),
	.w5(32'h3c659b44),
	.w6(32'h3bb0d0df),
	.w7(32'h3bc4800b),
	.w8(32'h3c47461f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8420b),
	.w1(32'hbb1d9c1d),
	.w2(32'hbb340b4c),
	.w3(32'hbb65d415),
	.w4(32'hbb04da51),
	.w5(32'hba9895bc),
	.w6(32'hbb0a0640),
	.w7(32'h3be3d928),
	.w8(32'h39864099),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c4407),
	.w1(32'h3bd8886c),
	.w2(32'hb936e7ed),
	.w3(32'h3972c400),
	.w4(32'hbb34b3b0),
	.w5(32'h3a397104),
	.w6(32'hbb003a80),
	.w7(32'hbaf4cf29),
	.w8(32'hbaa4d963),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36ac0),
	.w1(32'hbbc50027),
	.w2(32'hba92a313),
	.w3(32'hbc2901fe),
	.w4(32'hbc527f51),
	.w5(32'h3aa1442c),
	.w6(32'hbb84cefc),
	.w7(32'hbb18eeb7),
	.w8(32'hbc1b8503),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88db53),
	.w1(32'hbb9ae113),
	.w2(32'hbbbe816b),
	.w3(32'hb9f53cae),
	.w4(32'hbb626040),
	.w5(32'h39f97be0),
	.w6(32'hbbbc1130),
	.w7(32'h39a9a201),
	.w8(32'hbb367e9c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bcab2),
	.w1(32'h3bc14235),
	.w2(32'h3bdd56c9),
	.w3(32'hb91f19de),
	.w4(32'hbb58db75),
	.w5(32'hbc0609c8),
	.w6(32'h3a8013fc),
	.w7(32'h3c1fa8ed),
	.w8(32'h3b77dba8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e93be1),
	.w1(32'h3b85360a),
	.w2(32'h3c1a9e4c),
	.w3(32'hbc1d74da),
	.w4(32'hbc818a05),
	.w5(32'hbc6191ad),
	.w6(32'hbbc0f0e3),
	.w7(32'hbc802db0),
	.w8(32'hbc5e2921),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5580e0),
	.w1(32'h3c222c17),
	.w2(32'h3ab3b8e0),
	.w3(32'h3c2f42aa),
	.w4(32'h3cf76aa4),
	.w5(32'h3c58c2cb),
	.w6(32'h3c682c15),
	.w7(32'h3ce2c44e),
	.w8(32'h3b581c41),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70f49a),
	.w1(32'hbb2baf7b),
	.w2(32'h39e5197e),
	.w3(32'hba5c3939),
	.w4(32'h3a608224),
	.w5(32'hbb42fec0),
	.w6(32'h3a84a58f),
	.w7(32'hb90e894d),
	.w8(32'hbb0bb19d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53aa05),
	.w1(32'hbb8d21ca),
	.w2(32'hbc8d7bb9),
	.w3(32'hbbc447c3),
	.w4(32'hba388583),
	.w5(32'hbb7be800),
	.w6(32'hbb4a5926),
	.w7(32'h3a31a559),
	.w8(32'h3aa7df14),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71885c),
	.w1(32'h3b64da2d),
	.w2(32'h3cacfe58),
	.w3(32'hbc4a1f2f),
	.w4(32'hbb1d1c86),
	.w5(32'h3c46a262),
	.w6(32'h3bb0258f),
	.w7(32'hbc25f2b3),
	.w8(32'h3a9b3ba6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734824),
	.w1(32'h3a70ac25),
	.w2(32'hbc029aa3),
	.w3(32'hbb1b9925),
	.w4(32'hbb878219),
	.w5(32'hbbb2fb31),
	.w6(32'h3b5ef48f),
	.w7(32'h3b73c2ef),
	.w8(32'h3b982ed9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b787d46),
	.w1(32'h3c9f16d8),
	.w2(32'h3c8a8f3c),
	.w3(32'h3ca9b045),
	.w4(32'h3cac3558),
	.w5(32'h3d06f26a),
	.w6(32'h3c9a232d),
	.w7(32'h3cc0e55e),
	.w8(32'h3ca7e85d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2463c2),
	.w1(32'hbc7c0a4a),
	.w2(32'h3a115a6b),
	.w3(32'h3d15ff84),
	.w4(32'hbcc9ab79),
	.w5(32'hbb3c19f8),
	.w6(32'h3b1ee43e),
	.w7(32'hbbeec2dc),
	.w8(32'hbc00781c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16e197),
	.w1(32'hbbfe4dcc),
	.w2(32'hb88940dd),
	.w3(32'h3d4711cc),
	.w4(32'hbc5e675b),
	.w5(32'hbb7111b0),
	.w6(32'hbb2fbbc4),
	.w7(32'h3d1ae167),
	.w8(32'hbc14f817),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bcc18),
	.w1(32'h3a2bb6e2),
	.w2(32'hbc35dfc5),
	.w3(32'h3814b13b),
	.w4(32'h3b55a8e8),
	.w5(32'h3b855451),
	.w6(32'hbb7517fb),
	.w7(32'hbc8bd9b8),
	.w8(32'h3c4c6dc0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1b2b5),
	.w1(32'hbc8c025d),
	.w2(32'h3c33cae6),
	.w3(32'hbd110131),
	.w4(32'h3d849d35),
	.w5(32'h3cf287a7),
	.w6(32'hbc2e4b71),
	.w7(32'hbb8f82fd),
	.w8(32'h39df9154),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65c94b),
	.w1(32'hbb8e9c5b),
	.w2(32'h3c9b5e79),
	.w3(32'h3b3a795c),
	.w4(32'h3c13a6dd),
	.w5(32'h3aadb8df),
	.w6(32'h3b276d9d),
	.w7(32'h396267e8),
	.w8(32'hbcaf5b97),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae70b9),
	.w1(32'hbc9810c4),
	.w2(32'h3c101a97),
	.w3(32'hbc1a81cc),
	.w4(32'hbcc1e117),
	.w5(32'hbb804fa7),
	.w6(32'hba11556a),
	.w7(32'hbc679ef3),
	.w8(32'hbb1b239b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6ec85),
	.w1(32'hbc85c150),
	.w2(32'hbb259c9e),
	.w3(32'h3cdffe4a),
	.w4(32'h3c830992),
	.w5(32'h3c363b8a),
	.w6(32'hbc202f41),
	.w7(32'h3bc9c4dc),
	.w8(32'hbcabb1ac),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9691f),
	.w1(32'hb989bd4d),
	.w2(32'h3cb44bd3),
	.w3(32'hba0785ea),
	.w4(32'hbbe2d0a9),
	.w5(32'hbc8160ae),
	.w6(32'h3bbcaf4f),
	.w7(32'h3c3cfd83),
	.w8(32'h3c19ffdd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca85ff0),
	.w1(32'hbb1da968),
	.w2(32'h3bf1cc23),
	.w3(32'h3c2cc63a),
	.w4(32'hb9e6e744),
	.w5(32'h3d0bdce6),
	.w6(32'hbbd6ea0f),
	.w7(32'hb9d957bc),
	.w8(32'h3a97aae5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31d92),
	.w1(32'hbc98fab7),
	.w2(32'hbc00df2b),
	.w3(32'h3ba0ea6c),
	.w4(32'h3c63e0eb),
	.w5(32'hbd1c6fd9),
	.w6(32'hbca1a5b2),
	.w7(32'hbc48116b),
	.w8(32'hbc28a626),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30c2c6),
	.w1(32'hbd1d05fd),
	.w2(32'hbcec558d),
	.w3(32'hbc65780e),
	.w4(32'h3d2b2903),
	.w5(32'h3b66b41f),
	.w6(32'hbc0197c6),
	.w7(32'h3d52d04a),
	.w8(32'h3c1e4032),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd229f81),
	.w1(32'hbcfb14db),
	.w2(32'hbb1631cb),
	.w3(32'hbcad689d),
	.w4(32'h3ce6afb0),
	.w5(32'h3b43dade),
	.w6(32'h3cf82d8c),
	.w7(32'h3d5f20a8),
	.w8(32'h3ceefe92),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bfc99),
	.w1(32'h3c724178),
	.w2(32'h3c482b61),
	.w3(32'h3bfea68e),
	.w4(32'h3bcedc84),
	.w5(32'h3cc87cdc),
	.w6(32'hbc15c3d7),
	.w7(32'h3c918cd9),
	.w8(32'hbc454b0a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d09f2),
	.w1(32'hb9ff1990),
	.w2(32'h3b4dfbb5),
	.w3(32'h3c56126f),
	.w4(32'h3c5f1066),
	.w5(32'h3c862535),
	.w6(32'h3b43efcc),
	.w7(32'h3d5959d2),
	.w8(32'h3d12827e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd73bb9),
	.w1(32'h3ce26092),
	.w2(32'h3d0596cb),
	.w3(32'hbcf9e817),
	.w4(32'h3c6d7a1d),
	.w5(32'h3d4a6c1d),
	.w6(32'hba0cd396),
	.w7(32'h3b046d45),
	.w8(32'h3c10af28),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89414),
	.w1(32'hbb66001f),
	.w2(32'h3b920498),
	.w3(32'hbb180502),
	.w4(32'hbc3caa35),
	.w5(32'hbc481d9a),
	.w6(32'h3c23c26f),
	.w7(32'hbc01f1d7),
	.w8(32'h3c55660d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80abdf),
	.w1(32'hbc035b40),
	.w2(32'hbcddb4b5),
	.w3(32'h3c26f234),
	.w4(32'h3cf59ea1),
	.w5(32'hbb7cd918),
	.w6(32'h3ca75c9c),
	.w7(32'h3c670173),
	.w8(32'h3839dcb0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ddf50),
	.w1(32'hbb07fa4e),
	.w2(32'hbaf1dcfd),
	.w3(32'hbbe3e1b3),
	.w4(32'h39972428),
	.w5(32'h3ce8d54f),
	.w6(32'hbc014018),
	.w7(32'h3bc1a846),
	.w8(32'h3c3db9f4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8101),
	.w1(32'h3acec882),
	.w2(32'h3b91ccfd),
	.w3(32'h394c08e6),
	.w4(32'h3c531db7),
	.w5(32'h3c3d5c62),
	.w6(32'h3bbdff4b),
	.w7(32'h3bd0f1fc),
	.w8(32'hbb86ce7d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78b7b),
	.w1(32'hbb1ad129),
	.w2(32'h3b2a98bf),
	.w3(32'h3b1aab23),
	.w4(32'h3c189a6a),
	.w5(32'h3c0e69d2),
	.w6(32'hbb3e0d4d),
	.w7(32'h3b59dfb2),
	.w8(32'h3b2d41ac),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66cb9c),
	.w1(32'h3b554aab),
	.w2(32'h3afb101a),
	.w3(32'hbc2f85d5),
	.w4(32'h3b76f98b),
	.w5(32'h3c084cfc),
	.w6(32'hbc13cecc),
	.w7(32'h3b26ce58),
	.w8(32'hbabcbff5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2944b),
	.w1(32'h3cb76759),
	.w2(32'h3b31d72c),
	.w3(32'h3c5857ec),
	.w4(32'h3c9cc86c),
	.w5(32'h3cfae75c),
	.w6(32'hbc97abfe),
	.w7(32'h3bc749cf),
	.w8(32'h3c542598),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ac4f6),
	.w1(32'h3ae8d9ff),
	.w2(32'hbbaf7e85),
	.w3(32'h3b17fc2d),
	.w4(32'h3b1376ca),
	.w5(32'hb971bc9d),
	.w6(32'h3ac66738),
	.w7(32'h3b9edaba),
	.w8(32'h3c5a9fcc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2898da),
	.w1(32'h3add372a),
	.w2(32'h3be4b5b3),
	.w3(32'hba1a2805),
	.w4(32'h3a1fb2e7),
	.w5(32'h3b45485e),
	.w6(32'hba707929),
	.w7(32'hbabc01c7),
	.w8(32'h3b17c304),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eeb6cf),
	.w1(32'hbbdd5ce4),
	.w2(32'hbc1f88de),
	.w3(32'h3b77cf1a),
	.w4(32'h3b851496),
	.w5(32'h3c890ded),
	.w6(32'h3c0f3e0e),
	.w7(32'hbb774703),
	.w8(32'h3b23cf51),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf20fa),
	.w1(32'h3a4ac708),
	.w2(32'h3bab55d6),
	.w3(32'hbc09f7de),
	.w4(32'hbb91d391),
	.w5(32'h3b826a2d),
	.w6(32'hbbe8fddd),
	.w7(32'hbb3a32f4),
	.w8(32'hbb63a78c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc897a),
	.w1(32'hbbb46f8d),
	.w2(32'h3c5a61ca),
	.w3(32'h3c2e0e7d),
	.w4(32'hbbc84da4),
	.w5(32'hbcad6f20),
	.w6(32'h3c4de068),
	.w7(32'hbc14d30a),
	.w8(32'hbb80efde),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc63c0f),
	.w1(32'hbcab56e5),
	.w2(32'h3b9701f4),
	.w3(32'hbbcbdc5d),
	.w4(32'hbb2508be),
	.w5(32'h3c217958),
	.w6(32'hbbcc41b4),
	.w7(32'h3923b06f),
	.w8(32'hbb96d914),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd91fb5),
	.w1(32'hbcb4f4f0),
	.w2(32'hbb89f54f),
	.w3(32'hbcb0adcf),
	.w4(32'h3cdafd89),
	.w5(32'h3d4cef7c),
	.w6(32'h3b85dd35),
	.w7(32'h3ccc7d8a),
	.w8(32'h3d09c718),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba1ef7),
	.w1(32'hbac80613),
	.w2(32'hb9a40998),
	.w3(32'hbb621693),
	.w4(32'h3c8de212),
	.w5(32'hbb047b88),
	.w6(32'hbb211cf9),
	.w7(32'h3a044d80),
	.w8(32'h3bd411a3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fa99e),
	.w1(32'h37339a7f),
	.w2(32'h3a709de9),
	.w3(32'h3a81d6a5),
	.w4(32'hbb507fdd),
	.w5(32'h3bbc8cce),
	.w6(32'h3a7f43d4),
	.w7(32'h3aeefb83),
	.w8(32'h3c0bf3b0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245410),
	.w1(32'h3ab3ebec),
	.w2(32'hbbf7a171),
	.w3(32'h3b88a940),
	.w4(32'h3a958f73),
	.w5(32'h3b820602),
	.w6(32'h3addb401),
	.w7(32'h3b07da10),
	.w8(32'hbb077c1a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0d12c),
	.w1(32'h3cb56a06),
	.w2(32'h3c385fd7),
	.w3(32'h3c35e70b),
	.w4(32'h3bd03fc0),
	.w5(32'h3bed6612),
	.w6(32'h3c2905cb),
	.w7(32'h3ab919c4),
	.w8(32'hb93f54c8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195c28),
	.w1(32'hbad4edbf),
	.w2(32'h3ba268d0),
	.w3(32'hbbd7819b),
	.w4(32'h3befd148),
	.w5(32'hb9af013d),
	.w6(32'hbac97912),
	.w7(32'hbb406bd0),
	.w8(32'hbb1e0962),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9785),
	.w1(32'hbb384629),
	.w2(32'hbc157959),
	.w3(32'hbbb46d53),
	.w4(32'h3a375f7e),
	.w5(32'hbad9af6f),
	.w6(32'hb95bdcbe),
	.w7(32'h3bb40d07),
	.w8(32'h3c105435),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0a6be),
	.w1(32'h3be3fa5d),
	.w2(32'h38b62f33),
	.w3(32'hb92a4afd),
	.w4(32'hbc0b5538),
	.w5(32'hba1786f5),
	.w6(32'h3bdfc942),
	.w7(32'h3a5d7fd3),
	.w8(32'h3bd97e83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c36ec),
	.w1(32'h3b44c210),
	.w2(32'h3aa7a369),
	.w3(32'hbae7fe6a),
	.w4(32'h3cd1af09),
	.w5(32'h3cfd09a6),
	.w6(32'h3b52f67e),
	.w7(32'h3c2a4272),
	.w8(32'h3c0c5345),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c650730),
	.w1(32'h3c9417cb),
	.w2(32'h3c31ac2c),
	.w3(32'h3ba34cbc),
	.w4(32'h3bd2baa3),
	.w5(32'h3c52951e),
	.w6(32'h3c5221f9),
	.w7(32'h3b2572f2),
	.w8(32'h3b0f1423),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7009a),
	.w1(32'h3a326ce8),
	.w2(32'hba14453b),
	.w3(32'h39c752ff),
	.w4(32'hbbb55e8c),
	.w5(32'hbb40a54d),
	.w6(32'hbbe03d93),
	.w7(32'hbb6383de),
	.w8(32'hbb167d19),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71249a),
	.w1(32'hbb079dc1),
	.w2(32'h3b3b8ad3),
	.w3(32'h3a0ba6a9),
	.w4(32'hbb53d9d7),
	.w5(32'h3a4812d5),
	.w6(32'hbaa5a928),
	.w7(32'hbb61cb3d),
	.w8(32'h3ada03a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d8b1),
	.w1(32'h3bddf889),
	.w2(32'hbbf316a8),
	.w3(32'hbbac2cc6),
	.w4(32'h3b8fa526),
	.w5(32'hbb33e539),
	.w6(32'h3b25972a),
	.w7(32'h3b912c52),
	.w8(32'h3c61959f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072e05),
	.w1(32'hbb8ec0c0),
	.w2(32'hb9dea43e),
	.w3(32'hba933780),
	.w4(32'h3cb3d0e2),
	.w5(32'h3cc0d965),
	.w6(32'hba6060b4),
	.w7(32'h3c2ddb3c),
	.w8(32'h3c6c88dd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d0c20),
	.w1(32'h3c00fa14),
	.w2(32'h3d21c471),
	.w3(32'h3d0a8717),
	.w4(32'h3cc97be2),
	.w5(32'h3ca4e9b4),
	.w6(32'h3ccdbd9b),
	.w7(32'h3c6f9e29),
	.w8(32'h3c62621a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3809f8),
	.w1(32'hbbe2a227),
	.w2(32'h3c6619e1),
	.w3(32'h3bdf0fbf),
	.w4(32'h3d398a27),
	.w5(32'h3d3b59d8),
	.w6(32'h3c442b3c),
	.w7(32'h3c96e98c),
	.w8(32'h3cc6becb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f35c),
	.w1(32'h3bb4d7b3),
	.w2(32'hbb1d9d8c),
	.w3(32'h3b1d9ff8),
	.w4(32'h3bead026),
	.w5(32'h3bc786ab),
	.w6(32'hbc241f39),
	.w7(32'h3c2eaf17),
	.w8(32'h3cfed0d1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f9925),
	.w1(32'hba7f5d6c),
	.w2(32'hba5c45d8),
	.w3(32'hba0eba20),
	.w4(32'h3b4fba24),
	.w5(32'hbb4937d4),
	.w6(32'h3b83d9d9),
	.w7(32'hbb1db887),
	.w8(32'hbbe7b8c0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9bcd),
	.w1(32'h3b7e13b2),
	.w2(32'hbb43c20d),
	.w3(32'hb8e5cf6b),
	.w4(32'hb9c95b32),
	.w5(32'h3a84849f),
	.w6(32'h3bac17ab),
	.w7(32'h3b9e4f62),
	.w8(32'h3bcb7eb4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096fd0),
	.w1(32'hbbd7a1ee),
	.w2(32'h3bbf3e28),
	.w3(32'hbae64fc2),
	.w4(32'h3ae9df3e),
	.w5(32'hbb3b9091),
	.w6(32'hba3e2f15),
	.w7(32'hba51ccf6),
	.w8(32'h3c409371),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4afc),
	.w1(32'hba6a585d),
	.w2(32'h3a2f4f05),
	.w3(32'h38f2b5cb),
	.w4(32'h3b810ffa),
	.w5(32'h3c05fd05),
	.w6(32'h3a86d5c5),
	.w7(32'h3ba4947b),
	.w8(32'h3bfbb40a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba19252),
	.w1(32'h3be27568),
	.w2(32'hbb385c03),
	.w3(32'h39132193),
	.w4(32'h3c78c63e),
	.w5(32'h3c1abacc),
	.w6(32'hb8d536de),
	.w7(32'h3c7228ab),
	.w8(32'h3bdb34bf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9871e),
	.w1(32'h3b4103f2),
	.w2(32'h3b1b7415),
	.w3(32'hb9682662),
	.w4(32'h3b56e448),
	.w5(32'hbadc55e1),
	.w6(32'hbb115710),
	.w7(32'h3bc35a1a),
	.w8(32'h3bb9fd4b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a901bfc),
	.w1(32'hba3bea2f),
	.w2(32'hbb9fc046),
	.w3(32'hbb9844de),
	.w4(32'h3bdced25),
	.w5(32'hbc0c38e1),
	.w6(32'h3bc6ca90),
	.w7(32'h3c03627c),
	.w8(32'h3c187784),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d35d84),
	.w1(32'h3a8dca6a),
	.w2(32'h3a58107e),
	.w3(32'h3bddb989),
	.w4(32'h3be54b80),
	.w5(32'h3bedb81d),
	.w6(32'hbaa424af),
	.w7(32'h3b97ad59),
	.w8(32'h3bb636c6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8577e0),
	.w1(32'h3b14fd72),
	.w2(32'hbb2fb950),
	.w3(32'hbbe772f4),
	.w4(32'hba690c58),
	.w5(32'hba131c0b),
	.w6(32'hbbf6add8),
	.w7(32'hbc311226),
	.w8(32'hbbaead20),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f9fbb),
	.w1(32'hbbfe4719),
	.w2(32'h3c9a78f8),
	.w3(32'hbc26ee22),
	.w4(32'hbbb4775b),
	.w5(32'h3b9f43e5),
	.w6(32'hbbe44006),
	.w7(32'h3c086b39),
	.w8(32'hbb8eb2be),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257365),
	.w1(32'hba90b8f7),
	.w2(32'h3c0d3196),
	.w3(32'h3b82b447),
	.w4(32'h3ca0ce73),
	.w5(32'h3afcabd5),
	.w6(32'hbc457761),
	.w7(32'h3c201001),
	.w8(32'h3ca4597f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119e23),
	.w1(32'hbab61e7e),
	.w2(32'hbb0e9e73),
	.w3(32'h3b03bc65),
	.w4(32'hbc370b77),
	.w5(32'hbb692792),
	.w6(32'h3b3fd456),
	.w7(32'h3c0e39b5),
	.w8(32'h3d7e0c7d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62f3e),
	.w1(32'hbc97b4fe),
	.w2(32'h3c4ecc39),
	.w3(32'h3b9ad90a),
	.w4(32'h3c8db2d1),
	.w5(32'h3b0721de),
	.w6(32'h3c0f2e7c),
	.w7(32'h3c8aba7d),
	.w8(32'h3db76951),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8827),
	.w1(32'h3b68d24f),
	.w2(32'h3b23f3c3),
	.w3(32'hbccf14ca),
	.w4(32'h3b13c066),
	.w5(32'hbac987bb),
	.w6(32'h3bb987d1),
	.w7(32'h3d4276a3),
	.w8(32'h3c299732),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00db44),
	.w1(32'hba582859),
	.w2(32'hbc499dcb),
	.w3(32'h3d0a8ff9),
	.w4(32'h3c1de303),
	.w5(32'h3b453e02),
	.w6(32'hba8778a2),
	.w7(32'h3a00dca8),
	.w8(32'h3b0da9f7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6edfe),
	.w1(32'hbd39b7db),
	.w2(32'h3b9bdfcf),
	.w3(32'hbda7c15b),
	.w4(32'hbcebe00d),
	.w5(32'h3cbead7c),
	.w6(32'h3c2aa018),
	.w7(32'hbc25853c),
	.w8(32'h3b05ac18),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954b94),
	.w1(32'h3c13a0cb),
	.w2(32'hbc8033e3),
	.w3(32'h3d1cc991),
	.w4(32'hbbfd770b),
	.w5(32'h3be4e2e6),
	.w6(32'h3bba28d9),
	.w7(32'hbd8babb9),
	.w8(32'h3a8166e1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb910a),
	.w1(32'hbb22c373),
	.w2(32'hbb007ade),
	.w3(32'hbc81d506),
	.w4(32'hbb919bbb),
	.w5(32'h3b188aee),
	.w6(32'h3bca46cb),
	.w7(32'hbbf8dc90),
	.w8(32'h3b397249),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60b6b),
	.w1(32'h3b42ead6),
	.w2(32'h3b5b4112),
	.w3(32'hbbee043f),
	.w4(32'hbc8dc71a),
	.w5(32'h3d6f7935),
	.w6(32'h3b06f14b),
	.w7(32'hbba67661),
	.w8(32'hbced50b5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e315a),
	.w1(32'hbb9775f2),
	.w2(32'hbcc84a33),
	.w3(32'hbd2a87a4),
	.w4(32'h3c0a0d19),
	.w5(32'h3dce144c),
	.w6(32'h3c102e41),
	.w7(32'h3c93703a),
	.w8(32'h3c7a734b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd9ecb),
	.w1(32'hbc53ef81),
	.w2(32'h3c5a309d),
	.w3(32'h3c81b9cf),
	.w4(32'h3be52c4c),
	.w5(32'h3ba6c1e4),
	.w6(32'h3be8edfc),
	.w7(32'h3c07bca6),
	.w8(32'h397780e2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608a7e),
	.w1(32'hbc062392),
	.w2(32'hbd929b8d),
	.w3(32'h39b483c3),
	.w4(32'h391bbd39),
	.w5(32'h3ac38355),
	.w6(32'hbb8c8c95),
	.w7(32'h3bbc860d),
	.w8(32'h3be72091),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65ad2c),
	.w1(32'hbcb71e79),
	.w2(32'h3c27d4e9),
	.w3(32'h3b846beb),
	.w4(32'hbc19a421),
	.w5(32'hbc4cdc04),
	.w6(32'hbc81c2e1),
	.w7(32'h3b094632),
	.w8(32'hba425acc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1187cc),
	.w1(32'hbadadd0e),
	.w2(32'hbc8a191e),
	.w3(32'h3be55977),
	.w4(32'h3accbd15),
	.w5(32'h3bdfe002),
	.w6(32'h3c620110),
	.w7(32'h3bfaf3d2),
	.w8(32'h3c713ea9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd4a7),
	.w1(32'hbcb1e250),
	.w2(32'hbc1b2aab),
	.w3(32'hbc6de675),
	.w4(32'h3bf1146b),
	.w5(32'hbc848ea7),
	.w6(32'hbb5ccdce),
	.w7(32'hba93fb9a),
	.w8(32'h3c299234),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f2021),
	.w1(32'h392a6e0d),
	.w2(32'h3c179b10),
	.w3(32'h3c1a6214),
	.w4(32'h3bd71577),
	.w5(32'hbb46bffd),
	.w6(32'h3bc79eed),
	.w7(32'hbc8f03a7),
	.w8(32'hbb497883),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0e93),
	.w1(32'hbaaea9db),
	.w2(32'h3b47757a),
	.w3(32'h3d095a86),
	.w4(32'hbc66c074),
	.w5(32'hbc2cda06),
	.w6(32'h3b6e37a8),
	.w7(32'hbc598379),
	.w8(32'hbb515f80),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ab46a),
	.w1(32'hbc876bf0),
	.w2(32'hbb92c5ac),
	.w3(32'h3d404a15),
	.w4(32'h3ba9ebad),
	.w5(32'h3ced5995),
	.w6(32'h3ba0694b),
	.w7(32'hba05eb4a),
	.w8(32'h3b069316),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3188b1),
	.w1(32'h3c73ffd7),
	.w2(32'h3b20c8d1),
	.w3(32'hbbc328d8),
	.w4(32'h3b906ee2),
	.w5(32'h3b08287a),
	.w6(32'hbc0e2cf7),
	.w7(32'h3ac7c9cc),
	.w8(32'hb98859bf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25304),
	.w1(32'hbd1d3748),
	.w2(32'hbcdce398),
	.w3(32'h387b9821),
	.w4(32'h3c1aec0f),
	.w5(32'h3beddeca),
	.w6(32'h3a4a6538),
	.w7(32'hbc8c717d),
	.w8(32'h3beced2e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6812f7),
	.w1(32'h3cb9180d),
	.w2(32'hbc2d6437),
	.w3(32'hba74d432),
	.w4(32'hbc1c9594),
	.w5(32'hbd2cdab8),
	.w6(32'h395a50e6),
	.w7(32'h3b279564),
	.w8(32'hbbd5705c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e595),
	.w1(32'hbbf4c719),
	.w2(32'hbb70229e),
	.w3(32'h3bb3797e),
	.w4(32'h3c49e8fe),
	.w5(32'h3c19e15c),
	.w6(32'hba4df71c),
	.w7(32'h3b67bbf0),
	.w8(32'h3bf5f877),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d112c),
	.w1(32'hba511999),
	.w2(32'hbbed534d),
	.w3(32'h3a2a6638),
	.w4(32'h38955449),
	.w5(32'hb980dc9a),
	.w6(32'hbb164af6),
	.w7(32'h3aaf72e5),
	.w8(32'hbb9b40c6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10ab98),
	.w1(32'hbcaf27af),
	.w2(32'hbb7ac548),
	.w3(32'hbc7aac5b),
	.w4(32'h3aa4b3b7),
	.w5(32'hbb20f084),
	.w6(32'hbafa2a66),
	.w7(32'hbb5b7675),
	.w8(32'hbadd9bc0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3653c2),
	.w1(32'h3c9cd2fc),
	.w2(32'h3c1c3b0b),
	.w3(32'hbc1736ee),
	.w4(32'hbc34f518),
	.w5(32'hbc1b73ee),
	.w6(32'hbc30425c),
	.w7(32'h3bcfa962),
	.w8(32'h3c88857c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e540e),
	.w1(32'hb9177054),
	.w2(32'h3b093152),
	.w3(32'h3b8cf074),
	.w4(32'hba0b269b),
	.w5(32'hba2f7303),
	.w6(32'h3b2a97c6),
	.w7(32'h3ae06125),
	.w8(32'hbd415ba2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7634f1),
	.w1(32'h3aca5712),
	.w2(32'h3ade8539),
	.w3(32'h3a9913f8),
	.w4(32'hbc26eebc),
	.w5(32'h3ac0b481),
	.w6(32'h3a1be0f0),
	.w7(32'hbc4b88cd),
	.w8(32'h39998719),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32de74),
	.w1(32'h3a4e84e9),
	.w2(32'hbbba7b84),
	.w3(32'hbbd32399),
	.w4(32'hb992a0d2),
	.w5(32'hbbacb78e),
	.w6(32'hbc52cda9),
	.w7(32'hba6b13a3),
	.w8(32'hbc2665cd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fd6b),
	.w1(32'hbc3570c7),
	.w2(32'h3bee05fb),
	.w3(32'h3b8c58ec),
	.w4(32'hbb2d6a4b),
	.w5(32'h3aa2ace7),
	.w6(32'hb989a630),
	.w7(32'hbc94661f),
	.w8(32'hbbc73eb7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50bd69),
	.w1(32'hbb5ece3b),
	.w2(32'hbbe0d7f6),
	.w3(32'hb9e14fd6),
	.w4(32'hbae2f692),
	.w5(32'hbae5f16d),
	.w6(32'h3b4124b1),
	.w7(32'hba8a9790),
	.w8(32'h3c11556b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94146e6),
	.w1(32'hb9fa1a7f),
	.w2(32'hb913b548),
	.w3(32'h3b286580),
	.w4(32'h3b327358),
	.w5(32'hbac0200a),
	.w6(32'h3b77ac17),
	.w7(32'h3b342968),
	.w8(32'h3a8f06a6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000052),
	.w1(32'h3bed487a),
	.w2(32'h3c0f006e),
	.w3(32'hbbf46018),
	.w4(32'h3c00d716),
	.w5(32'h3c1b96b8),
	.w6(32'hbb806233),
	.w7(32'h3c34e82d),
	.w8(32'h3c1efb80),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule