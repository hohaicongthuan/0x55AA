module layer_10_featuremap_381(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58adb4),
	.w1(32'h3cbaf48b),
	.w2(32'h3add4e67),
	.w3(32'h3b4824c0),
	.w4(32'h3c8dd803),
	.w5(32'h3a1ce5f0),
	.w6(32'h3bccc279),
	.w7(32'h3c886c5d),
	.w8(32'h3baf6d72),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8015d4),
	.w1(32'hbbc9fdeb),
	.w2(32'hbba4f05d),
	.w3(32'hbca5f3e4),
	.w4(32'hbc226012),
	.w5(32'hbbd650d2),
	.w6(32'hbc05e18e),
	.w7(32'hbbee39b6),
	.w8(32'hbc1f52ae),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9736a),
	.w1(32'hbc526c89),
	.w2(32'h3c15b671),
	.w3(32'h3c57a063),
	.w4(32'hbcdd4a0f),
	.w5(32'h3c23e0e8),
	.w6(32'h3bade037),
	.w7(32'hbc9ac475),
	.w8(32'hbc649236),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3833c0),
	.w1(32'hbbd0df82),
	.w2(32'h3c28feff),
	.w3(32'h3c1219d4),
	.w4(32'hbbc6d278),
	.w5(32'hbc1b0e37),
	.w6(32'h39cdac9f),
	.w7(32'hbc396b80),
	.w8(32'h3bfefba0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad7d8),
	.w1(32'h3bee5fac),
	.w2(32'h3bade606),
	.w3(32'h3c6b7d7d),
	.w4(32'hbb9b1987),
	.w5(32'h3bc778d9),
	.w6(32'h3ca170cb),
	.w7(32'hbb61cec8),
	.w8(32'hbaafcb7a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbb7f2),
	.w1(32'h39ec7d92),
	.w2(32'hbb15e0a4),
	.w3(32'hbb8054c4),
	.w4(32'h3c132d32),
	.w5(32'h3c1a9c80),
	.w6(32'hbbbabeec),
	.w7(32'h3b0d426e),
	.w8(32'hbaeec3c7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75595f),
	.w1(32'h3c1ec657),
	.w2(32'h3b515e97),
	.w3(32'hbb7f9c46),
	.w4(32'h3b88559f),
	.w5(32'hbba65056),
	.w6(32'hbb9a3f4c),
	.w7(32'h3be987cb),
	.w8(32'h3b459891),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d5aaf),
	.w1(32'h3a4882dc),
	.w2(32'hba0360b8),
	.w3(32'h3aa61735),
	.w4(32'hb9faa709),
	.w5(32'hbb196bc5),
	.w6(32'h3bb777f5),
	.w7(32'hbbd75aee),
	.w8(32'hba5bab1a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda114a),
	.w1(32'hbca637bc),
	.w2(32'h3b84cb0f),
	.w3(32'hbbeff1dc),
	.w4(32'hbcd83f54),
	.w5(32'hbc6787f7),
	.w6(32'hbac3207d),
	.w7(32'hbc7b9ae1),
	.w8(32'hbb1d77ed),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca54de),
	.w1(32'hbbcbe6e4),
	.w2(32'hb92b26dd),
	.w3(32'h3c6efa69),
	.w4(32'hbc401a48),
	.w5(32'hbb081055),
	.w6(32'h3ca6bb1e),
	.w7(32'hbb2df578),
	.w8(32'h3be12cfd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bafdf),
	.w1(32'hbb57c6eb),
	.w2(32'h3989046a),
	.w3(32'h3bd00e92),
	.w4(32'hbc271f36),
	.w5(32'hbba87348),
	.w6(32'h3bf7f0a2),
	.w7(32'hbb0a41a4),
	.w8(32'hbc219934),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e436),
	.w1(32'h3bc7fb11),
	.w2(32'hbb2262bf),
	.w3(32'h3bcb405e),
	.w4(32'h3c4aef2f),
	.w5(32'h3bc220af),
	.w6(32'h3b2ed0ec),
	.w7(32'h3a4533a0),
	.w8(32'hbb0d00eb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc354a69),
	.w1(32'hbc010e8b),
	.w2(32'hbbc16b46),
	.w3(32'hbc802f31),
	.w4(32'hbc7bff22),
	.w5(32'hbcb73ad4),
	.w6(32'hbc6646cc),
	.w7(32'hbc1d5556),
	.w8(32'hbc212c01),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c269a3a),
	.w1(32'h3a0066a1),
	.w2(32'h3c4d6196),
	.w3(32'h3c9a2a5f),
	.w4(32'hbc167595),
	.w5(32'h3bd837dd),
	.w6(32'h3c51e911),
	.w7(32'hbc3789ff),
	.w8(32'hbb9c2551),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee9b88),
	.w1(32'hbc523938),
	.w2(32'hbae766fc),
	.w3(32'h39a69192),
	.w4(32'hbca7a3ce),
	.w5(32'hbc29eee7),
	.w6(32'h3adbe1c4),
	.w7(32'hbc19080a),
	.w8(32'hbc6dc320),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82598d),
	.w1(32'h3b02b590),
	.w2(32'hba8650ad),
	.w3(32'h3cc02576),
	.w4(32'hbc1702ea),
	.w5(32'h3afcca84),
	.w6(32'h3c3b5a47),
	.w7(32'hbb9cc69a),
	.w8(32'hbbb398be),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb15a4e),
	.w1(32'hbbfcff85),
	.w2(32'h3ba0ce86),
	.w3(32'h3c054fda),
	.w4(32'hbc271060),
	.w5(32'hbb3fe6bd),
	.w6(32'h3b945586),
	.w7(32'hbbfa40a7),
	.w8(32'hbbe7d41f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb20315),
	.w1(32'h3c1889be),
	.w2(32'h3834b1c0),
	.w3(32'h3bfdf88a),
	.w4(32'h3be4c092),
	.w5(32'h3c2fc743),
	.w6(32'hbbaa131a),
	.w7(32'h3c37e8df),
	.w8(32'h3bed4838),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc557275),
	.w1(32'hbbaa6d3f),
	.w2(32'hbb9d4795),
	.w3(32'hbc9011ba),
	.w4(32'hbc128ac8),
	.w5(32'hbc86d6f6),
	.w6(32'hbc441bfc),
	.w7(32'hbb0f1e61),
	.w8(32'hbc206a46),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86ea16),
	.w1(32'hba8e4ca0),
	.w2(32'hbbd46030),
	.w3(32'h3c4d7cfd),
	.w4(32'hbc0d2773),
	.w5(32'hbcb4092e),
	.w6(32'h3c07440e),
	.w7(32'hba5e6fd9),
	.w8(32'hbcc6eb66),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c377850),
	.w1(32'hba277a0c),
	.w2(32'hbb84ee0b),
	.w3(32'h3d025a74),
	.w4(32'h3c1a93ac),
	.w5(32'h3bfb4c63),
	.w6(32'h3b892fa6),
	.w7(32'hbb8b6a2a),
	.w8(32'hbc0487ee),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2347af),
	.w1(32'hbc3c6825),
	.w2(32'hbc4466f9),
	.w3(32'hbbe95795),
	.w4(32'hbb97e788),
	.w5(32'hbc8a1b11),
	.w6(32'hbbf8b49e),
	.w7(32'hbb9151c5),
	.w8(32'hbcc871be),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bf6e1),
	.w1(32'hbba6e190),
	.w2(32'hbb8bcac8),
	.w3(32'h3bb98fd6),
	.w4(32'hbc0e35da),
	.w5(32'h3c09c303),
	.w6(32'hbb517a30),
	.w7(32'h3b46e732),
	.w8(32'h3aac0d8d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1422a9),
	.w1(32'hbb82555d),
	.w2(32'hbc57706c),
	.w3(32'h3c12ac81),
	.w4(32'h39c03e74),
	.w5(32'hbbf3dd9f),
	.w6(32'h3b560644),
	.w7(32'hbbb9872d),
	.w8(32'hbc0f44ed),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e88eb),
	.w1(32'hbc846cac),
	.w2(32'hbb3245f1),
	.w3(32'h3c2f02bc),
	.w4(32'hbcffa5ab),
	.w5(32'h3b64bfbc),
	.w6(32'h3aae8b70),
	.w7(32'hbcd9f728),
	.w8(32'hbc620558),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81d223),
	.w1(32'h3cab3314),
	.w2(32'h3b4a0a05),
	.w3(32'h3cfb9015),
	.w4(32'h3c544177),
	.w5(32'hbbbe6a84),
	.w6(32'h3b6ab3fc),
	.w7(32'h3c44e675),
	.w8(32'hbc7ba3c0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d4a5),
	.w1(32'hbc20477e),
	.w2(32'hbc72b0ef),
	.w3(32'hbccc8f78),
	.w4(32'hbc25b0ed),
	.w5(32'hbc81b70e),
	.w6(32'hbc8a64bf),
	.w7(32'hbb7da10d),
	.w8(32'h3bba8e48),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7daa),
	.w1(32'hbc32375f),
	.w2(32'hbc1f4526),
	.w3(32'h3bed1495),
	.w4(32'hbc5809e2),
	.w5(32'hbc523249),
	.w6(32'h3c628e50),
	.w7(32'h3af6f9f0),
	.w8(32'h3b1c62f4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9a735),
	.w1(32'hbbf48b22),
	.w2(32'hbc1312cf),
	.w3(32'h3bc059f4),
	.w4(32'hbc8922c5),
	.w5(32'hbc00cca5),
	.w6(32'h3c1ba689),
	.w7(32'h3b919a66),
	.w8(32'h3c7c3e24),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6c718),
	.w1(32'h3c3b9af9),
	.w2(32'h3b6c1c97),
	.w3(32'h3b388586),
	.w4(32'h3c304e36),
	.w5(32'h3c73c870),
	.w6(32'h3b8c0574),
	.w7(32'h3bf05c77),
	.w8(32'h3b08da1a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd7a7d),
	.w1(32'hb89f7aff),
	.w2(32'h3c233d85),
	.w3(32'hbc8ff57d),
	.w4(32'hbc6b77c1),
	.w5(32'h3b1e3009),
	.w6(32'hbc8d9472),
	.w7(32'hbac71243),
	.w8(32'h3a5f3aaa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf93fcf),
	.w1(32'hbc73f085),
	.w2(32'h3a8c2a68),
	.w3(32'hbb983c4b),
	.w4(32'hbcbe4465),
	.w5(32'h398f7f22),
	.w6(32'hbc73cc49),
	.w7(32'hbc7c1346),
	.w8(32'hbafb7b42),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16a9c),
	.w1(32'hbbc45bae),
	.w2(32'h3b28ee46),
	.w3(32'h3c28ceb7),
	.w4(32'hbb909785),
	.w5(32'h3bb11c9f),
	.w6(32'h3bd95e7e),
	.w7(32'hbc420018),
	.w8(32'hba197cc3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9b211),
	.w1(32'h3b838866),
	.w2(32'h3b11b17f),
	.w3(32'h3bae65b1),
	.w4(32'hba83165b),
	.w5(32'hbb43d18f),
	.w6(32'h3b9cc234),
	.w7(32'h3b30e7d4),
	.w8(32'hbb8921db),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177b70),
	.w1(32'hbb19a1a1),
	.w2(32'hbbe4f811),
	.w3(32'hbb0bfd83),
	.w4(32'h3c05768c),
	.w5(32'h397ca91c),
	.w6(32'h3b4a06bb),
	.w7(32'h3bb4467e),
	.w8(32'h3b5aed9e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc61aa3),
	.w1(32'h3c63e288),
	.w2(32'h3a1b619e),
	.w3(32'hbc33733a),
	.w4(32'h3cf2d2f8),
	.w5(32'hbb9f2fac),
	.w6(32'h3b0a0d57),
	.w7(32'h3c00554c),
	.w8(32'hbbd787ca),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fc730),
	.w1(32'h3b90901b),
	.w2(32'h3c1f28b6),
	.w3(32'hbc8e0166),
	.w4(32'hbc919c1e),
	.w5(32'hbb852b69),
	.w6(32'hbc86a3b1),
	.w7(32'hbc022752),
	.w8(32'hbc6266bb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5bf0f),
	.w1(32'h39d86f9e),
	.w2(32'h3b6ceea7),
	.w3(32'h3c9a2417),
	.w4(32'hbb861576),
	.w5(32'hba21e2b2),
	.w6(32'h3c0276bf),
	.w7(32'hbc02ab9c),
	.w8(32'hbb55446e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990e42),
	.w1(32'h3c222c3c),
	.w2(32'h38bf6ded),
	.w3(32'h3c0de2c8),
	.w4(32'h3bd21cb3),
	.w5(32'hbca27723),
	.w6(32'hbab686db),
	.w7(32'h3a60806a),
	.w8(32'hbbc7d6fb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35dbc1),
	.w1(32'hbb76432f),
	.w2(32'hbb57f874),
	.w3(32'h3b5284d4),
	.w4(32'hbb0fbd03),
	.w5(32'hbc315311),
	.w6(32'hbb014fcb),
	.w7(32'hbb66bd4a),
	.w8(32'hbbc2b8d3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910652),
	.w1(32'hbaad87c9),
	.w2(32'hba1674f8),
	.w3(32'hb9fc6275),
	.w4(32'hbbcb1886),
	.w5(32'hbb103c8c),
	.w6(32'hbbdda6b5),
	.w7(32'hbc09880d),
	.w8(32'h3b06a965),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167556),
	.w1(32'h3b138c36),
	.w2(32'hbb49a5b6),
	.w3(32'h3c5d99ea),
	.w4(32'h39f3690d),
	.w5(32'hbc30c8c9),
	.w6(32'h3c505a64),
	.w7(32'h3ab601ec),
	.w8(32'hbaea9379),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9257a0c),
	.w1(32'hbc2ad9e0),
	.w2(32'hbb860fe3),
	.w3(32'h3c4a625c),
	.w4(32'hbbb40032),
	.w5(32'hbbfe0f41),
	.w6(32'h3ae4671e),
	.w7(32'hbbbb3d2c),
	.w8(32'h3bbb7196),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12761),
	.w1(32'h3bafdefd),
	.w2(32'hbb169b81),
	.w3(32'h3b9e1abd),
	.w4(32'h3c49174f),
	.w5(32'hbc03cf08),
	.w6(32'hbc0823fa),
	.w7(32'h3c2b3389),
	.w8(32'hbb07f475),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15aaed),
	.w1(32'hbb4e1ea1),
	.w2(32'hbbf7d398),
	.w3(32'hbc0cb08d),
	.w4(32'hbb92f41a),
	.w5(32'hbbe7f16e),
	.w6(32'h3b2d14b9),
	.w7(32'h3b9eeff7),
	.w8(32'h3ba6f3a0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f5e44),
	.w1(32'hbc123d55),
	.w2(32'hbb80f8c4),
	.w3(32'hbb3cfe36),
	.w4(32'hbc561ed8),
	.w5(32'h3c038987),
	.w6(32'hbb9cf640),
	.w7(32'hbbed07a0),
	.w8(32'h399f1492),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ba96f),
	.w1(32'hbb2754f8),
	.w2(32'hbbac7b2f),
	.w3(32'h3bb6218c),
	.w4(32'h398b904f),
	.w5(32'hbbea6ee7),
	.w6(32'h3be87696),
	.w7(32'hbba3f702),
	.w8(32'hbb8ea332),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59d4ef),
	.w1(32'hbc0fb25c),
	.w2(32'hbc1795e3),
	.w3(32'h3c2a8f08),
	.w4(32'hbc8ecc4a),
	.w5(32'hbc8f0c67),
	.w6(32'h3c2001b9),
	.w7(32'hbc5735f3),
	.w8(32'hbbaff96e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68db8e),
	.w1(32'hbbae4646),
	.w2(32'h3bd5b00b),
	.w3(32'h3c6c6278),
	.w4(32'h3cf1b250),
	.w5(32'h3cefbc83),
	.w6(32'h3c8dab78),
	.w7(32'h3bac954f),
	.w8(32'h3bf1ce39),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb609b),
	.w1(32'h3c455c93),
	.w2(32'h3adf0abf),
	.w3(32'hbc98fdec),
	.w4(32'h3d3b6c84),
	.w5(32'h3ca968ce),
	.w6(32'hbc658236),
	.w7(32'h3c797e07),
	.w8(32'h3b3a7029),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82891a),
	.w1(32'hbc11db1e),
	.w2(32'h3b106f1b),
	.w3(32'hbc351bea),
	.w4(32'hbc490b66),
	.w5(32'h3a0f4ab3),
	.w6(32'hbc662843),
	.w7(32'hbbf8bac8),
	.w8(32'hba58bae3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9149f),
	.w1(32'hba83e1bb),
	.w2(32'hbc350ff9),
	.w3(32'h3bf6fee9),
	.w4(32'hbc48808b),
	.w5(32'hbce6b3e7),
	.w6(32'h3b96468c),
	.w7(32'hbc37f529),
	.w8(32'hbc577f53),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56b75e),
	.w1(32'h3c20ec16),
	.w2(32'h3b002fca),
	.w3(32'h3c7a85c5),
	.w4(32'h3cd41725),
	.w5(32'h3c71ed4d),
	.w6(32'h3c60683a),
	.w7(32'h3c898295),
	.w8(32'h3b3b4d26),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f1da9),
	.w1(32'hbbb0a70a),
	.w2(32'hbb58f8c3),
	.w3(32'hbcf58d13),
	.w4(32'h3c20d45a),
	.w5(32'h3b40b509),
	.w6(32'hbcd9b2fb),
	.w7(32'h3b91066c),
	.w8(32'h3bdbe5b6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc385421),
	.w1(32'hbc4bea31),
	.w2(32'h3bc12f38),
	.w3(32'hbc75a7b8),
	.w4(32'hbd062828),
	.w5(32'hbb3c01ca),
	.w6(32'hbb7b4646),
	.w7(32'hbcb711f1),
	.w8(32'hbbb333a9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04de89),
	.w1(32'hbb126d5f),
	.w2(32'h3babbcbe),
	.w3(32'h3c81743d),
	.w4(32'hbba8bc0e),
	.w5(32'hbbf00731),
	.w6(32'h3a2aa677),
	.w7(32'hbba6668f),
	.w8(32'hbc294f40),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27779),
	.w1(32'h3bc370b7),
	.w2(32'hbad08ed7),
	.w3(32'hba249caf),
	.w4(32'h3ab48f5c),
	.w5(32'h3c5e13f7),
	.w6(32'hbb22ee79),
	.w7(32'h3b2c65a0),
	.w8(32'h3b3df8d4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74149a),
	.w1(32'hbc5be813),
	.w2(32'hbc123f7f),
	.w3(32'hbb945df3),
	.w4(32'hbcb709ae),
	.w5(32'hbc7cd3da),
	.w6(32'hbb5d37fe),
	.w7(32'hbca3229c),
	.w8(32'hbc6f39c7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d899),
	.w1(32'hbc51257e),
	.w2(32'hbcaf1643),
	.w3(32'h3b9c57cd),
	.w4(32'hbc93c66b),
	.w5(32'hbced7b84),
	.w6(32'h3b6fd93a),
	.w7(32'hbc3bdbc2),
	.w8(32'hbcd5db11),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69cc00),
	.w1(32'hbafa4c08),
	.w2(32'h3c0fa69c),
	.w3(32'h3b48eeb9),
	.w4(32'hbc9188f9),
	.w5(32'hbb8eca5d),
	.w6(32'hbbee629c),
	.w7(32'hbc8bb78f),
	.w8(32'hbc8561f8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be98e23),
	.w1(32'hba7bfea9),
	.w2(32'h3b2a68c8),
	.w3(32'h3cef8fc7),
	.w4(32'hbc1ff2ae),
	.w5(32'hba62e4ba),
	.w6(32'hbc4ff8a7),
	.w7(32'hbbfaf065),
	.w8(32'hbbac70a6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8142fb),
	.w1(32'hbbaa397c),
	.w2(32'hbb876012),
	.w3(32'hbb0c61ec),
	.w4(32'hbbd75a6c),
	.w5(32'hbc41365e),
	.w6(32'hbbf172be),
	.w7(32'hbb84347e),
	.w8(32'hbbc1508d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9426e8),
	.w1(32'hbc28d973),
	.w2(32'hbc0f89af),
	.w3(32'h3b23b496),
	.w4(32'hbc9d61a4),
	.w5(32'hbc473d3c),
	.w6(32'hbb933951),
	.w7(32'hbc46d7b5),
	.w8(32'h3ba7071a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c249809),
	.w1(32'hbb7cd617),
	.w2(32'hbb26fba7),
	.w3(32'h3ccdbeea),
	.w4(32'hbc11b53f),
	.w5(32'h3b578e9e),
	.w6(32'h3c6ce3d8),
	.w7(32'h3b603277),
	.w8(32'h3bd866a7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1e14),
	.w1(32'h3d18fa79),
	.w2(32'h3b0a5d18),
	.w3(32'hbada7234),
	.w4(32'h3d4648de),
	.w5(32'hbb0f375b),
	.w6(32'h3a72aa6b),
	.w7(32'h3d18ce46),
	.w8(32'hbaead04d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb772b0),
	.w1(32'h3c0b4566),
	.w2(32'h3baac769),
	.w3(32'hbd19b1e4),
	.w4(32'h3cc9d7b1),
	.w5(32'h3bc98999),
	.w6(32'hbce755ab),
	.w7(32'h3bfec71d),
	.w8(32'h3b3bea56),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc474aaf),
	.w1(32'hbbd787e1),
	.w2(32'h3ba700f4),
	.w3(32'hbc35beae),
	.w4(32'hbc555ed9),
	.w5(32'h3bffec76),
	.w6(32'hbc8b8120),
	.w7(32'hbc46540f),
	.w8(32'hbbe285f4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d76e57),
	.w1(32'hbc9312a8),
	.w2(32'h3b543d63),
	.w3(32'hbb944362),
	.w4(32'hbc8d30af),
	.w5(32'h3b4c8114),
	.w6(32'hb9a1ed73),
	.w7(32'hbc8fea49),
	.w8(32'h3b3797e2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59ed84),
	.w1(32'hbc83b083),
	.w2(32'hbb93d176),
	.w3(32'h3c339d0b),
	.w4(32'hbd0a3c74),
	.w5(32'hbc864fd4),
	.w6(32'h3c1c60c3),
	.w7(32'hbc7eed59),
	.w8(32'h3b81acc5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84eea4),
	.w1(32'h382213bb),
	.w2(32'hb8fb2761),
	.w3(32'h3c7f2da4),
	.w4(32'h3791c6a7),
	.w5(32'hb918753e),
	.w6(32'h3ca9da18),
	.w7(32'h38822ca6),
	.w8(32'hb86abced),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36217708),
	.w1(32'h3538395f),
	.w2(32'h353820f8),
	.w3(32'h35ec23f1),
	.w4(32'hb440b2d3),
	.w5(32'hb39303b4),
	.w6(32'h36316f77),
	.w7(32'h35a99a52),
	.w8(32'h35863da0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367c82ac),
	.w1(32'h351d54f2),
	.w2(32'h34a306d8),
	.w3(32'h36000c9f),
	.w4(32'hb5f6a9cd),
	.w5(32'h349aaea8),
	.w6(32'h368ad806),
	.w7(32'h3551b6f1),
	.w8(32'h353ab5a0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368c2df8),
	.w1(32'hb5b24016),
	.w2(32'h367d25df),
	.w3(32'h36a3c516),
	.w4(32'hb5a263ba),
	.w5(32'h34865525),
	.w6(32'h361d31a4),
	.w7(32'hb5a2be32),
	.w8(32'hb52ac52a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377b701b),
	.w1(32'h371e5d96),
	.w2(32'h37be0c9a),
	.w3(32'h37c3408f),
	.w4(32'h376a03f4),
	.w5(32'h378de23e),
	.w6(32'h373629dc),
	.w7(32'hb7063cf0),
	.w8(32'hb6a9aa1c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362f1485),
	.w1(32'h36178643),
	.w2(32'hb65a4407),
	.w3(32'h36040446),
	.w4(32'h3596721c),
	.w5(32'hb6aa1919),
	.w6(32'h36a3d158),
	.w7(32'h36850f36),
	.w8(32'hb51d1971),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6220ead),
	.w1(32'hb7d22baa),
	.w2(32'hb7d87e2f),
	.w3(32'h354d3b8b),
	.w4(32'h37ef85b4),
	.w5(32'hb7aa08ae),
	.w6(32'h37c2de10),
	.w7(32'h36febbb4),
	.w8(32'hb6b626eb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9b785),
	.w1(32'hb91aa884),
	.w2(32'hb875758c),
	.w3(32'h385a6618),
	.w4(32'hb886f435),
	.w5(32'hb8de642e),
	.w6(32'h394c7143),
	.w7(32'hb829e0b9),
	.w8(32'hb8161f5a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823384b),
	.w1(32'hb68ea160),
	.w2(32'hb89ca323),
	.w3(32'hb82c5429),
	.w4(32'h36bddc94),
	.w5(32'hb86e8cd9),
	.w6(32'hb7b64036),
	.w7(32'h377da8d0),
	.w8(32'hb788627b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377e0b08),
	.w1(32'h38709c9a),
	.w2(32'hb860aac0),
	.w3(32'hb8879f40),
	.w4(32'h37f30dd5),
	.w5(32'hb8f24c2d),
	.w6(32'hb8b98daf),
	.w7(32'hb81d874e),
	.w8(32'hb9260bcc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37186f13),
	.w1(32'h3723f56a),
	.w2(32'hb694630c),
	.w3(32'h36c82221),
	.w4(32'h371b2fac),
	.w5(32'hb789ceba),
	.w6(32'hb798e3b6),
	.w7(32'hb706f8c6),
	.w8(32'hb74db7b8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fefd2c),
	.w1(32'hb790ffd5),
	.w2(32'hb8be66d1),
	.w3(32'hb88c80e2),
	.w4(32'hb7bc5449),
	.w5(32'hb88da131),
	.w6(32'hb7225ddd),
	.w7(32'h3840975c),
	.w8(32'hb7833631),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ea41a),
	.w1(32'h36a428dc),
	.w2(32'hb70a29b6),
	.w3(32'h36bdc20e),
	.w4(32'h376f16e1),
	.w5(32'hb73ce877),
	.w6(32'hb7272608),
	.w7(32'hb6f0101c),
	.w8(32'hb7fd3d3a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b94b3f),
	.w1(32'hb669f621),
	.w2(32'hb54eb4f3),
	.w3(32'hb69ae00e),
	.w4(32'hb58f3ca0),
	.w5(32'h34f8d48d),
	.w6(32'h33ec59be),
	.w7(32'h360ddc62),
	.w8(32'h3619453b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b4c1c5),
	.w1(32'h331a6741),
	.w2(32'hb5fab4c8),
	.w3(32'h363c8ac7),
	.w4(32'hb58d4d93),
	.w5(32'hb6a70968),
	.w6(32'h3687a47d),
	.w7(32'h363703e9),
	.w8(32'hb59d0c13),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3367d6c7),
	.w1(32'hb4eb2240),
	.w2(32'hb2b76333),
	.w3(32'hb4e84c00),
	.w4(32'h350cf5c0),
	.w5(32'h361e0617),
	.w6(32'h3626b1e0),
	.w7(32'h35fe9a94),
	.w8(32'h35d8c923),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35869cae),
	.w1(32'h35f43a20),
	.w2(32'h35d632db),
	.w3(32'h35bd73a6),
	.w4(32'h360b00d6),
	.w5(32'h360263b2),
	.w6(32'h35be979d),
	.w7(32'hb4bd94f2),
	.w8(32'h35cb84ca),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b81195),
	.w1(32'hb7bcf25d),
	.w2(32'h36186e64),
	.w3(32'h37d650b2),
	.w4(32'h38217b37),
	.w5(32'h38150580),
	.w6(32'h37107f53),
	.w7(32'h374f2b66),
	.w8(32'h3800af45),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64778a6),
	.w1(32'h377cb3c1),
	.w2(32'h37b7ddad),
	.w3(32'hb631c371),
	.w4(32'h36a404ca),
	.w5(32'h371bb6fc),
	.w6(32'h351cfb27),
	.w7(32'h3703c1c1),
	.w8(32'h37658b59),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80453de),
	.w1(32'hb81277da),
	.w2(32'hb8ce3928),
	.w3(32'hb86f1f1e),
	.w4(32'hb80637c2),
	.w5(32'hb8f74524),
	.w6(32'hb81e6b22),
	.w7(32'hb6921958),
	.w8(32'hb8ad7d73),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8312236),
	.w1(32'h3517a3f2),
	.w2(32'hb633b130),
	.w3(32'hb81c628c),
	.w4(32'hb6012da8),
	.w5(32'hb8072365),
	.w6(32'hb84fa1ed),
	.w7(32'hb87c473d),
	.w8(32'hb8264770),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372408f3),
	.w1(32'h38993de9),
	.w2(32'h3858f1ed),
	.w3(32'h3845ebd0),
	.w4(32'h389dfcea),
	.w5(32'h37fc011e),
	.w6(32'h364602ef),
	.w7(32'h37ea19f5),
	.w8(32'h3818a4a5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8762817),
	.w1(32'hb8739b5e),
	.w2(32'hb9624370),
	.w3(32'hb873b4c7),
	.w4(32'hb907f317),
	.w5(32'hb97bc1e7),
	.w6(32'hb8820a8d),
	.w7(32'hb793e9e7),
	.w8(32'hb95a60e0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37632e8e),
	.w1(32'h38a4725c),
	.w2(32'h38b6f1af),
	.w3(32'h383c71a8),
	.w4(32'h38914e18),
	.w5(32'h3855ca5b),
	.w6(32'h36f9dd42),
	.w7(32'h37c2f33d),
	.w8(32'h368bbe54),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e880ae),
	.w1(32'hb9050e8b),
	.w2(32'hb983e719),
	.w3(32'hb9099890),
	.w4(32'hb8b02317),
	.w5(32'hb932239a),
	.w6(32'hb8aa84a2),
	.w7(32'hb7d23e07),
	.w8(32'hb8ec8f4a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a740c6),
	.w1(32'hb851446b),
	.w2(32'hb98704d0),
	.w3(32'h388f1e75),
	.w4(32'hb867b552),
	.w5(32'hb94e651d),
	.w6(32'h3935e6b6),
	.w7(32'h390ac480),
	.w8(32'hb87165f1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e822e5),
	.w1(32'hb8036aa1),
	.w2(32'hb8854e1c),
	.w3(32'hb8446d47),
	.w4(32'hb76a5a9f),
	.w5(32'hb81a03b9),
	.w6(32'hb711a033),
	.w7(32'h383fd693),
	.w8(32'hb7336484),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3698934b),
	.w1(32'h380c0812),
	.w2(32'hb82492cb),
	.w3(32'hb7b6a838),
	.w4(32'h371c93d2),
	.w5(32'hb82a27e6),
	.w6(32'h351d7c49),
	.w7(32'h3798e578),
	.w8(32'hb8195f44),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9789410),
	.w1(32'hb9090158),
	.w2(32'hb98948d2),
	.w3(32'hb998ffb6),
	.w4(32'hb8c63b60),
	.w5(32'hb985a742),
	.w6(32'hb8c4f1eb),
	.w7(32'h38b86ba7),
	.w8(32'hb8e3890a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868e002),
	.w1(32'h38a36c5a),
	.w2(32'h38b4c62d),
	.w3(32'h38873e54),
	.w4(32'h38fef361),
	.w5(32'h38fafff4),
	.w6(32'hb8ae98a2),
	.w7(32'hb89bf7c0),
	.w8(32'hb790ad36),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e0cfae),
	.w1(32'hb6737c27),
	.w2(32'h370b4cc0),
	.w3(32'hb7daa0b3),
	.w4(32'hb4f7380c),
	.w5(32'hb81eda1a),
	.w6(32'hb7ff66fe),
	.w7(32'hb8a7d728),
	.w8(32'hb860a982),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975fc34),
	.w1(32'hb845a430),
	.w2(32'hb9b1a667),
	.w3(32'hb9e4847b),
	.w4(32'hb91a0bae),
	.w5(32'hb9ae1223),
	.w6(32'hb990510e),
	.w7(32'h3856d095),
	.w8(32'hb9729f45),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3efd3),
	.w1(32'hb930c1b0),
	.w2(32'hb9845af1),
	.w3(32'hb9a00501),
	.w4(32'hb91182f7),
	.w5(32'hb95f79a9),
	.w6(32'hb90ac5f3),
	.w7(32'h3907192f),
	.w8(32'hb8a533ad),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365f605b),
	.w1(32'h385342e9),
	.w2(32'hb91a62cd),
	.w3(32'hb9177629),
	.w4(32'hb7a8dd92),
	.w5(32'hb922fa8c),
	.w6(32'hb96b3bf5),
	.w7(32'hb7120a55),
	.w8(32'hb95863af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739a03c),
	.w1(32'h38ed8863),
	.w2(32'h37f0c911),
	.w3(32'hb80ca211),
	.w4(32'h38cf228d),
	.w5(32'h34a3555d),
	.w6(32'h381d7a64),
	.w7(32'h38e365e4),
	.w8(32'h381c8d6e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec178d),
	.w1(32'h38b62a40),
	.w2(32'hb8ca4b59),
	.w3(32'h37dca559),
	.w4(32'h38e5e96f),
	.w5(32'hb88c2684),
	.w6(32'h372a0d25),
	.w7(32'hb7544128),
	.w8(32'hb8f22fa7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fe5742),
	.w1(32'hb69d21fa),
	.w2(32'hb7a02f6e),
	.w3(32'hb7ef7303),
	.w4(32'h36e7fce9),
	.w5(32'h369d99c4),
	.w6(32'h379111d2),
	.w7(32'hb85177dd),
	.w8(32'hb72231ca),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ed00f8),
	.w1(32'h377e4b7e),
	.w2(32'h377ede82),
	.w3(32'h378d2f5e),
	.w4(32'h37c3878c),
	.w5(32'h37a0b2da),
	.w6(32'h30957980),
	.w7(32'h364ee1c6),
	.w8(32'h36185893),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eebcbd),
	.w1(32'h365f988b),
	.w2(32'hb7f92579),
	.w3(32'hb7344198),
	.w4(32'h36615185),
	.w5(32'hb725b384),
	.w6(32'hb7058258),
	.w7(32'h361d4da9),
	.w8(32'hb6e6a3f5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9163e52),
	.w1(32'hb8a498b8),
	.w2(32'hb901a07f),
	.w3(32'hb93e51c8),
	.w4(32'hb8b49741),
	.w5(32'hb90057d7),
	.w6(32'hb88bb0ff),
	.w7(32'h389e4e05),
	.w8(32'hb7ff6ab5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940e1fb),
	.w1(32'hb8f8a8f0),
	.w2(32'hb9609a77),
	.w3(32'hb938841a),
	.w4(32'hb8c1e559),
	.w5(32'hb94210fd),
	.w6(32'h386c5dea),
	.w7(32'h38f5d97f),
	.w8(32'hb7e05dfe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b75c92),
	.w1(32'hb71d6654),
	.w2(32'hb8abb97c),
	.w3(32'hb828aa67),
	.w4(32'h381e4d86),
	.w5(32'hb8df3a1c),
	.w6(32'h3808f979),
	.w7(32'h38be22eb),
	.w8(32'hb7fde936),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cd4d6),
	.w1(32'h36adb5cf),
	.w2(32'hb7b8f1f6),
	.w3(32'hb8d47965),
	.w4(32'hb7c26639),
	.w5(32'hb883fd27),
	.w6(32'hb8fbc32e),
	.w7(32'hb8427e78),
	.w8(32'hb8f96bcc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5ea9b),
	.w1(32'h3868c8a0),
	.w2(32'h385b348d),
	.w3(32'hb75d0506),
	.w4(32'h3874696c),
	.w5(32'h385bfc26),
	.w6(32'hb797442b),
	.w7(32'h37e783d0),
	.w8(32'h37a0effb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dc6f3e),
	.w1(32'hb7a0bb0d),
	.w2(32'hb7cb4ce1),
	.w3(32'hb71426ea),
	.w4(32'hb6d69adf),
	.w5(32'hb84a6387),
	.w6(32'hb7c3889f),
	.w7(32'hb7c574b6),
	.w8(32'hb87a33d2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81fcdef),
	.w1(32'hb743bf30),
	.w2(32'hb804dff3),
	.w3(32'hb83bb79d),
	.w4(32'hb7a91dd7),
	.w5(32'hb81563c1),
	.w6(32'hb7e6c461),
	.w7(32'h36690c5e),
	.w8(32'hb7db8f78),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366d2752),
	.w1(32'h371f0a9b),
	.w2(32'hb75aa45d),
	.w3(32'hb7868974),
	.w4(32'hb776851b),
	.w5(32'hb7dbaedd),
	.w6(32'hb6948fff),
	.w7(32'hb792ccfa),
	.w8(32'hb249b3ce),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d54251),
	.w1(32'hb5e3bf47),
	.w2(32'hb4d9916c),
	.w3(32'h35eb8f80),
	.w4(32'hb5f6a6d8),
	.w5(32'h35487483),
	.w6(32'h361d91ee),
	.w7(32'hb5aeea53),
	.w8(32'hb56688ab),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a46e10),
	.w1(32'hb2c754a3),
	.w2(32'hb4fc25d0),
	.w3(32'h365a2c95),
	.w4(32'h35895039),
	.w5(32'h35b91e9d),
	.w6(32'h35b69ec8),
	.w7(32'h35406414),
	.w8(32'h34682a43),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37825032),
	.w1(32'h38603105),
	.w2(32'hb7227b99),
	.w3(32'h37d44296),
	.w4(32'hb79d9925),
	.w5(32'hb7fe6ff8),
	.w6(32'h3808e373),
	.w7(32'hb79407d7),
	.w8(32'hb605ccae),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37921e3e),
	.w1(32'hb84f0c84),
	.w2(32'hb9286a6f),
	.w3(32'hb8056c86),
	.w4(32'h37954eaa),
	.w5(32'hb8eb75d3),
	.w6(32'h389de745),
	.w7(32'h38fc587e),
	.w8(32'hb74b00a0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a53664),
	.w1(32'h38ca027c),
	.w2(32'hb8111e2c),
	.w3(32'h36df795d),
	.w4(32'hb786579b),
	.w5(32'hb8944fe4),
	.w6(32'hb6f26645),
	.w7(32'hb8781e94),
	.w8(32'hb89037d7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7345fd0),
	.w1(32'hb804c83f),
	.w2(32'hb8f0c348),
	.w3(32'hb836999e),
	.w4(32'hb7cb8c82),
	.w5(32'hb88d2768),
	.w6(32'hb814777a),
	.w7(32'hb789ee30),
	.w8(32'hb86f6ca5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b8643b),
	.w1(32'h37e40148),
	.w2(32'h37928059),
	.w3(32'h36463eea),
	.w4(32'h37fa5610),
	.w5(32'h367be825),
	.w6(32'hb7a6fe24),
	.w7(32'h37dc4d90),
	.w8(32'hb53725f9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36073785),
	.w1(32'h360186f0),
	.w2(32'h352a901c),
	.w3(32'h35699a41),
	.w4(32'hb49ad34b),
	.w5(32'h3627761a),
	.w6(32'h365f85e1),
	.w7(32'hb509577f),
	.w8(32'h3405a255),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34cac88f),
	.w1(32'h3725111d),
	.w2(32'h36b4c19f),
	.w3(32'hb5873fa9),
	.w4(32'h33872cc9),
	.w5(32'h360be946),
	.w6(32'hb60a145b),
	.w7(32'h357de740),
	.w8(32'h36272fe5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356e01ae),
	.w1(32'h35b50b7b),
	.w2(32'h36678906),
	.w3(32'h3696f12e),
	.w4(32'h35e646ba),
	.w5(32'h361ff6ef),
	.w6(32'h3632f85e),
	.w7(32'h36446880),
	.w8(32'h35ec0163),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3516f3bc),
	.w1(32'h38645d9d),
	.w2(32'hb80722c7),
	.w3(32'h35b1aaa1),
	.w4(32'h389844af),
	.w5(32'hb6cfa8b1),
	.w6(32'h36849d59),
	.w7(32'h388b2697),
	.w8(32'hb74a9c63),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85149e0),
	.w1(32'hb74d9b53),
	.w2(32'hb79f441c),
	.w3(32'hb824013e),
	.w4(32'h384397bd),
	.w5(32'hb6161aa4),
	.w6(32'hb8429171),
	.w7(32'hb5abef81),
	.w8(32'hb88e9370),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3478be2b),
	.w1(32'hb8805c08),
	.w2(32'hb9158e0d),
	.w3(32'hb901f3be),
	.w4(32'hb8370ebd),
	.w5(32'hb9007744),
	.w6(32'hb875f9ff),
	.w7(32'h3825ab47),
	.w8(32'hb8c16986),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35656043),
	.w1(32'hb4a87cf0),
	.w2(32'h34c96c48),
	.w3(32'h36a2ffa8),
	.w4(32'h367a8fcc),
	.w5(32'h3503fd64),
	.w6(32'h36b5f67e),
	.w7(32'hb597c707),
	.w8(32'hb6365fd3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb796adf2),
	.w1(32'hb5be214c),
	.w2(32'h36b6bf26),
	.w3(32'hb783f2f8),
	.w4(32'h36d43a50),
	.w5(32'h373bf909),
	.w6(32'hb79b48a4),
	.w7(32'hb6c64a7e),
	.w8(32'h36153c56),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ee4869),
	.w1(32'h371cef60),
	.w2(32'h34ddf90b),
	.w3(32'h369b3c7d),
	.w4(32'h3731ffc4),
	.w5(32'hb601e6fa),
	.w6(32'h3655df67),
	.w7(32'h36b0caab),
	.w8(32'hb69b8ea4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859f91a),
	.w1(32'hb7cac0dd),
	.w2(32'hb8899488),
	.w3(32'hb88080f3),
	.w4(32'hb78206b4),
	.w5(32'hb8824d0c),
	.w6(32'hb714323d),
	.w7(32'h383907cb),
	.w8(32'hb78bbf49),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb754e6ab),
	.w1(32'hb8ab9ae6),
	.w2(32'hb8332fa7),
	.w3(32'hb7ff52e5),
	.w4(32'hb8aa6f2c),
	.w5(32'hb8854c6b),
	.w6(32'h382a3d1d),
	.w7(32'hb8456361),
	.w8(32'hb86b7816),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a99a7),
	.w1(32'hb72f993e),
	.w2(32'hb8de9409),
	.w3(32'hb880b0fa),
	.w4(32'h36e87f2b),
	.w5(32'hb87acc6f),
	.w6(32'hb8999f98),
	.w7(32'h381666c7),
	.w8(32'hb7a4f862),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d49435),
	.w1(32'hb4a879f0),
	.w2(32'hb8347c3a),
	.w3(32'hb8058efa),
	.w4(32'hb6a761b7),
	.w5(32'hb8042f9e),
	.w6(32'hb78b6490),
	.w7(32'h375e2360),
	.w8(32'hb78beda1),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3ea81),
	.w1(32'hb8283426),
	.w2(32'hb83bdb86),
	.w3(32'hb832b92a),
	.w4(32'h350c66ec),
	.w5(32'hb81329b5),
	.w6(32'hb876e5aa),
	.w7(32'h366046fd),
	.w8(32'hb824d4ec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b08612),
	.w1(32'h37d6908e),
	.w2(32'hb8952a33),
	.w3(32'hb772d0e6),
	.w4(32'h38a86fe8),
	.w5(32'hb8cf79f0),
	.w6(32'hb81550cf),
	.w7(32'h3814868b),
	.w8(32'hb896a6fb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b318c5),
	.w1(32'h378a669d),
	.w2(32'h378d9457),
	.w3(32'hb83e120c),
	.w4(32'hb783b48e),
	.w5(32'h36b7d2f3),
	.w6(32'hb78bb867),
	.w7(32'hb828c6e4),
	.w8(32'h36dc3877),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb780dac3),
	.w1(32'hb7b9ae40),
	.w2(32'hb926464d),
	.w3(32'hb8b9113d),
	.w4(32'hb821dff2),
	.w5(32'hb9198265),
	.w6(32'h371a4014),
	.w7(32'h38ca16f5),
	.w8(32'hb8583d5d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77250fa),
	.w1(32'hb699be41),
	.w2(32'hb82fc005),
	.w3(32'hb7f9c345),
	.w4(32'hb7257244),
	.w5(32'hb8282c53),
	.w6(32'hb720941f),
	.w7(32'h3748718b),
	.w8(32'hb7b015f6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ee342),
	.w1(32'hb76ca590),
	.w2(32'hb91b1bc4),
	.w3(32'h38083766),
	.w4(32'h372a8fe2),
	.w5(32'hb90a53cd),
	.w6(32'h379c9991),
	.w7(32'h37efce56),
	.w8(32'hb91209a7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880e7d1),
	.w1(32'h379f5bed),
	.w2(32'hb8ddc05c),
	.w3(32'h37e88bc5),
	.w4(32'hb81b4789),
	.w5(32'hb8b3bed0),
	.w6(32'h38553363),
	.w7(32'h373d9ef0),
	.w8(32'hb8166bff),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34eedcec),
	.w1(32'h359d1582),
	.w2(32'h352ec672),
	.w3(32'h360e6b75),
	.w4(32'h35fd263f),
	.w5(32'h351e2b34),
	.w6(32'h35fcf018),
	.w7(32'h359fd328),
	.w8(32'h358be580),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d3f779),
	.w1(32'hb5a791ca),
	.w2(32'hb46589fc),
	.w3(32'h34cf388b),
	.w4(32'h348a5eb6),
	.w5(32'h3591f35e),
	.w6(32'h363eb336),
	.w7(32'h364bdfed),
	.w8(32'h35ebfecb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7374392),
	.w1(32'hb6d4ccbd),
	.w2(32'h3647dbe8),
	.w3(32'hb48c4b87),
	.w4(32'hb56933ff),
	.w5(32'h370652eb),
	.w6(32'hb71339a6),
	.w7(32'hb7899745),
	.w8(32'h3595080e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c1d5e4),
	.w1(32'hb8798e8b),
	.w2(32'hb8dabfc2),
	.w3(32'hb92393ca),
	.w4(32'hb864f10e),
	.w5(32'hb81a73f8),
	.w6(32'hb7fe638a),
	.w7(32'h382ca686),
	.w8(32'hb80bc879),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b8fbb0),
	.w1(32'h380919cc),
	.w2(32'hb86dba07),
	.w3(32'hb662edb3),
	.w4(32'h3730fc68),
	.w5(32'hb879a4e5),
	.w6(32'hb811a68c),
	.w7(32'hb826c591),
	.w8(32'hb8b0c9ca),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e73d54),
	.w1(32'hb51c628b),
	.w2(32'hb4d43709),
	.w3(32'hb53dcb23),
	.w4(32'hb4cdd65d),
	.w5(32'h34e302f9),
	.w6(32'hb4c613b4),
	.w7(32'hb5647055),
	.w8(32'hb4162975),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a333df),
	.w1(32'hb8b9a08f),
	.w2(32'hb96f63bb),
	.w3(32'hb8db4737),
	.w4(32'hb8a3b342),
	.w5(32'hb94908f4),
	.w6(32'h388016b9),
	.w7(32'h3804e867),
	.w8(32'hb8974d4c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e68f4d),
	.w1(32'hb98d7fc8),
	.w2(32'hb94a82e4),
	.w3(32'hb879695b),
	.w4(32'hb967f0cf),
	.w5(32'hb90cc9ff),
	.w6(32'hb940ba44),
	.w7(32'hb8939870),
	.w8(32'hb8f57e13),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89dc06c),
	.w1(32'h36c4a774),
	.w2(32'hb85c4012),
	.w3(32'hb82739fd),
	.w4(32'h381d00f5),
	.w5(32'hb81bb344),
	.w6(32'hb821e771),
	.w7(32'h37cef212),
	.w8(32'hb860b32c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c808ff),
	.w1(32'hb7f12241),
	.w2(32'hb8fcd63e),
	.w3(32'hb7db58f8),
	.w4(32'hb833f323),
	.w5(32'hb8f2e66e),
	.w6(32'h375e1672),
	.w7(32'h38628ecd),
	.w8(32'hb84bb8ab),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c77700),
	.w1(32'hb80bac98),
	.w2(32'h38297214),
	.w3(32'h36bf5768),
	.w4(32'hb742f99e),
	.w5(32'h3793e494),
	.w6(32'h3789bc97),
	.w7(32'h377605ef),
	.w8(32'h37fead1c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b8efe9),
	.w1(32'h38035f91),
	.w2(32'h37c927e6),
	.w3(32'h370a45be),
	.w4(32'h37dd52e4),
	.w5(32'h384658b1),
	.w6(32'h382543d7),
	.w7(32'h38238e1e),
	.w8(32'h37d7683d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8459959),
	.w1(32'hb81ba043),
	.w2(32'hb92c5d72),
	.w3(32'hb8b1772c),
	.w4(32'hb85c4330),
	.w5(32'hb9139f41),
	.w6(32'h37135400),
	.w7(32'h387e2d4d),
	.w8(32'hb741a88b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84e0423),
	.w1(32'hb84bb54b),
	.w2(32'hb8f6f922),
	.w3(32'h384b446e),
	.w4(32'hb71c7b70),
	.w5(32'hb870b99c),
	.w6(32'hb7a06f63),
	.w7(32'hb8640d7f),
	.w8(32'hb80001f6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba0aea),
	.w1(32'h3834c0be),
	.w2(32'h3858d77f),
	.w3(32'h37e43889),
	.w4(32'h38151403),
	.w5(32'h3819a91b),
	.w6(32'h37738bbd),
	.w7(32'h37b44c3f),
	.w8(32'h37db4708),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb620a1ec),
	.w1(32'hb605690b),
	.w2(32'hb5317604),
	.w3(32'h34d2158e),
	.w4(32'hb515e267),
	.w5(32'hb6201092),
	.w6(32'hb69c9477),
	.w7(32'hb696b2d7),
	.w8(32'hb6cded20),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d3565b),
	.w1(32'hb61e12a8),
	.w2(32'hb5c99691),
	.w3(32'h36a60f8e),
	.w4(32'h364b1b0d),
	.w5(32'h34421f40),
	.w6(32'h366d70e5),
	.w7(32'h368a3efb),
	.w8(32'h35e2640a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8849f63),
	.w1(32'hb730eccd),
	.w2(32'hb9035390),
	.w3(32'hb91b1b42),
	.w4(32'hb77a72f5),
	.w5(32'hb8d7749e),
	.w6(32'hb89c5ba8),
	.w7(32'h386ac05b),
	.w8(32'hb7a1279e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37be19b5),
	.w1(32'h330e0a6f),
	.w2(32'hb74a9731),
	.w3(32'h3775c6fe),
	.w4(32'hb6d70fe3),
	.w5(32'hb7a6f3da),
	.w6(32'h3756cfc9),
	.w7(32'hb69e5f5c),
	.w8(32'hb74d3486),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37639cf0),
	.w1(32'h385584a3),
	.w2(32'hb90e0d05),
	.w3(32'hb8ab21ee),
	.w4(32'hb7cd17c6),
	.w5(32'hb8f85c06),
	.w6(32'hb7f4b8d9),
	.w7(32'h385ae71f),
	.w8(32'hb8803579),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787f987),
	.w1(32'hb63b39fd),
	.w2(32'hb61194b5),
	.w3(32'hb6ac8d39),
	.w4(32'hb616dc85),
	.w5(32'hb694bd6f),
	.w6(32'hb77badb9),
	.w7(32'hb69d94f0),
	.w8(32'hb69d1220),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38258f27),
	.w1(32'h37ff559f),
	.w2(32'h383c1015),
	.w3(32'h38c07cee),
	.w4(32'h38a63ffe),
	.w5(32'h3856b23b),
	.w6(32'h389c2526),
	.w7(32'h380d18d4),
	.w8(32'h3797a325),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3731b775),
	.w1(32'h362041dd),
	.w2(32'h3692d2c9),
	.w3(32'hb626813c),
	.w4(32'h36fba526),
	.w5(32'h3732e346),
	.w6(32'hb7a3ef9e),
	.w7(32'h36ed1a06),
	.w8(32'h369749c5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3714800f),
	.w1(32'hb732d204),
	.w2(32'hb6ecceda),
	.w3(32'hb6088bd4),
	.w4(32'hb7254452),
	.w5(32'hb7891116),
	.w6(32'hb8177a3c),
	.w7(32'hb81d0711),
	.w8(32'hb7f00054),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716a8f4),
	.w1(32'h38e30dc7),
	.w2(32'hb9150854),
	.w3(32'hb8c7980b),
	.w4(32'h3885ef97),
	.w5(32'hb8ddd030),
	.w6(32'hb6658b40),
	.w7(32'h390625f4),
	.w8(32'h36e87fe5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb838897d),
	.w1(32'hb921ead2),
	.w2(32'hb99096f8),
	.w3(32'hb907e2c8),
	.w4(32'hb92a0575),
	.w5(32'hb96db90c),
	.w6(32'hb8cff117),
	.w7(32'hb7df78d5),
	.w8(32'hb9207e7c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c1f248),
	.w1(32'h38915fe1),
	.w2(32'h38b5e1fe),
	.w3(32'h383d5c42),
	.w4(32'h386d7e0f),
	.w5(32'h386f3135),
	.w6(32'h3819a060),
	.w7(32'h38512f87),
	.w8(32'h386503a3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928e293),
	.w1(32'hb8a2ea29),
	.w2(32'hb911a76a),
	.w3(32'hb8ff8b18),
	.w4(32'hb8b7902a),
	.w5(32'hb8d379bc),
	.w6(32'hb8d6d350),
	.w7(32'hb79b94f0),
	.w8(32'hb8aae071),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3719b3a0),
	.w1(32'h3715fd2a),
	.w2(32'hb5a292f0),
	.w3(32'h371009cc),
	.w4(32'h370019d9),
	.w5(32'hb62bc419),
	.w6(32'h361e1374),
	.w7(32'h36c197b6),
	.w8(32'hb6618e62),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8da908b),
	.w1(32'h36c1ebe6),
	.w2(32'hb8ff118c),
	.w3(32'hb8a36b7a),
	.w4(32'h38591c4e),
	.w5(32'hb864aa93),
	.w6(32'hb8740c88),
	.w7(32'h38c74234),
	.w8(32'hb82d8a4f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8895fe1),
	.w1(32'hb74dcdc4),
	.w2(32'hb81813e3),
	.w3(32'hb84f62ae),
	.w4(32'h3588f51b),
	.w5(32'hb7e46928),
	.w6(32'hb871342d),
	.w7(32'h364a6c36),
	.w8(32'hb78b1f62),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9603f87),
	.w1(32'hb98a30f0),
	.w2(32'hb9a2919e),
	.w3(32'hb97f4f8c),
	.w4(32'hb9620fdd),
	.w5(32'hb9311576),
	.w6(32'hb8a9ef42),
	.w7(32'hb6fa4485),
	.w8(32'hb8504372),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2c5ef),
	.w1(32'h38416bc2),
	.w2(32'hb8004baf),
	.w3(32'h36d343a8),
	.w4(32'hb612b25c),
	.w5(32'hb850b0de),
	.w6(32'h369a5c7b),
	.w7(32'h36f6c5a3),
	.w8(32'hb7b435e0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3734974e),
	.w1(32'hb8933246),
	.w2(32'hb8eb50f1),
	.w3(32'hb84f7a13),
	.w4(32'hb875275b),
	.w5(32'hb8a97b34),
	.w6(32'hb706d7ee),
	.w7(32'h36ab2c61),
	.w8(32'hb7b3ab9a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c02154),
	.w1(32'h34e48415),
	.w2(32'h354547a7),
	.w3(32'h36026691),
	.w4(32'h35a901f8),
	.w5(32'h35694724),
	.w6(32'h35990b41),
	.w7(32'h360a97e2),
	.w8(32'h35aee800),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb716f3f3),
	.w1(32'h3792cb31),
	.w2(32'h37fa73ca),
	.w3(32'h36b9a777),
	.w4(32'h37960506),
	.w5(32'h370e49fb),
	.w6(32'hb70724f0),
	.w7(32'h372b39b2),
	.w8(32'hb6e636cf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7242de1),
	.w1(32'hb6822e10),
	.w2(32'h35248b1b),
	.w3(32'hb6e0bf4e),
	.w4(32'hb506111f),
	.w5(32'hb61e592c),
	.w6(32'hb6ae5c32),
	.w7(32'h35204e70),
	.w8(32'hb6a591ef),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8435c1e),
	.w1(32'hb7f77483),
	.w2(32'hb840142f),
	.w3(32'hb814ee02),
	.w4(32'hb7c06cf6),
	.w5(32'hb81d520f),
	.w6(32'hb82d7f8d),
	.w7(32'hb7a585ac),
	.w8(32'hb83cb955),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ca7c65),
	.w1(32'h34364e86),
	.w2(32'h358bb3e1),
	.w3(32'h35b735e1),
	.w4(32'h35a32547),
	.w5(32'h35adc89f),
	.w6(32'hb4acba24),
	.w7(32'hb520fe11),
	.w8(32'hb478cb21),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae0d17),
	.w1(32'hb74eabfb),
	.w2(32'hb732bd7b),
	.w3(32'hb7298176),
	.w4(32'hb5e9507a),
	.w5(32'hb6a789ea),
	.w6(32'hb71284c9),
	.w7(32'h370ea33d),
	.w8(32'hb679225c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b05d92),
	.w1(32'h370c6009),
	.w2(32'h37087437),
	.w3(32'h3717fa5f),
	.w4(32'h3716bc90),
	.w5(32'h35f5df40),
	.w6(32'hb3bf4d27),
	.w7(32'h34b6cfea),
	.w8(32'hb637ac4d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849a4ca),
	.w1(32'h3883fee9),
	.w2(32'h379d0fb0),
	.w3(32'h3776beaf),
	.w4(32'h38803295),
	.w5(32'h37827fca),
	.w6(32'hb7889e27),
	.w7(32'h37c36253),
	.w8(32'h36f64683),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38657aa7),
	.w1(32'h37b2c5b8),
	.w2(32'hb7e0b520),
	.w3(32'h368af1d1),
	.w4(32'h36e43e56),
	.w5(32'hb79aa894),
	.w6(32'hb82ef257),
	.w7(32'hb815422a),
	.w8(32'hb826d9b4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aeb616),
	.w1(32'h379aad98),
	.w2(32'h36b205d0),
	.w3(32'h38a9ae24),
	.w4(32'h365833e2),
	.w5(32'h36599cb1),
	.w6(32'h38985354),
	.w7(32'hb71070f8),
	.w8(32'h37332084),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884b083),
	.w1(32'hb926baaa),
	.w2(32'hb9ac41b5),
	.w3(32'hb84ec707),
	.w4(32'h36c2c04f),
	.w5(32'hb9a118ae),
	.w6(32'h38e5388c),
	.w7(32'h392aee54),
	.w8(32'hb93aed5b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb653c4c0),
	.w1(32'hb808a09e),
	.w2(32'hb8d3194d),
	.w3(32'h38c3c7fd),
	.w4(32'h380c87dd),
	.w5(32'hb8b8e6d7),
	.w6(32'h38bcd28d),
	.w7(32'h38c0deb8),
	.w8(32'hb750a10f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c3ce2f),
	.w1(32'h33e12281),
	.w2(32'h372b6215),
	.w3(32'hb606c2cf),
	.w4(32'h36f8a304),
	.w5(32'h36a7f780),
	.w6(32'h34a52693),
	.w7(32'h370a35b5),
	.w8(32'h378039ac),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d57438),
	.w1(32'hb35f7c2e),
	.w2(32'h35e4feaa),
	.w3(32'h348dbc4d),
	.w4(32'hb5a0486e),
	.w5(32'hb570606a),
	.w6(32'hb61caa82),
	.w7(32'hb56597b2),
	.w8(32'hb5b96050),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b2aba),
	.w1(32'hb7d62918),
	.w2(32'hb8309390),
	.w3(32'hb7e4cedf),
	.w4(32'hb77c440f),
	.w5(32'hb81750f8),
	.w6(32'hb63556d5),
	.w7(32'h37bedbb2),
	.w8(32'hb7e0d52d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3372a8d7),
	.w1(32'h35c43ab2),
	.w2(32'h35e1eddb),
	.w3(32'h351a70d3),
	.w4(32'h3574acce),
	.w5(32'h33b1c6af),
	.w6(32'h35aaa671),
	.w7(32'h3594e102),
	.w8(32'h34debef1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69ced63),
	.w1(32'h37595f78),
	.w2(32'hb802472e),
	.w3(32'hb79502fd),
	.w4(32'h373a419e),
	.w5(32'hb7daa918),
	.w6(32'h365efdb1),
	.w7(32'h37ef288e),
	.w8(32'hb6c28fc8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e77296),
	.w1(32'hb6268d9c),
	.w2(32'h373f95fc),
	.w3(32'h379bda86),
	.w4(32'h37d18e6b),
	.w5(32'hb79acb86),
	.w6(32'hb84a0317),
	.w7(32'hb827893e),
	.w8(32'hb879c0ff),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83333b9),
	.w1(32'hb850afda),
	.w2(32'hb8cc8dc4),
	.w3(32'hb7eee689),
	.w4(32'hb807ba09),
	.w5(32'hb8b8e2ab),
	.w6(32'h38037bc1),
	.w7(32'h3838352f),
	.w8(32'hb77e8a5d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a3f4e0),
	.w1(32'hb681bf5e),
	.w2(32'hb6914ed7),
	.w3(32'hb7325c73),
	.w4(32'h3708cf4f),
	.w5(32'h36e1a5ac),
	.w6(32'hb7743071),
	.w7(32'h36b91c56),
	.w8(32'h36754952),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70e2a3c),
	.w1(32'hbbad6fd1),
	.w2(32'hbb0cf09a),
	.w3(32'hb8b39bcb),
	.w4(32'hbb58d00b),
	.w5(32'h3a9f3520),
	.w6(32'hb79db279),
	.w7(32'h3afc9d7d),
	.w8(32'h3b9485d2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e134),
	.w1(32'hbaa8ce10),
	.w2(32'hbaecbca7),
	.w3(32'hbba12a3f),
	.w4(32'hbaaaddf2),
	.w5(32'h3c5a7a5d),
	.w6(32'h3bf25ac6),
	.w7(32'h3c0352df),
	.w8(32'h3bb7d7c4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d33d3),
	.w1(32'h3a9432ff),
	.w2(32'h3ab7a2b7),
	.w3(32'h3ba50e38),
	.w4(32'hbb4fdc91),
	.w5(32'h3bcd360f),
	.w6(32'h3ae6050d),
	.w7(32'hbb6129c1),
	.w8(32'h3992a632),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4ddb),
	.w1(32'hb93e420f),
	.w2(32'h3bdffba0),
	.w3(32'hbbb2b6cb),
	.w4(32'hbba1401c),
	.w5(32'h3b974e9a),
	.w6(32'h3b39494f),
	.w7(32'hbb038626),
	.w8(32'hbb86d923),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27ccaa),
	.w1(32'hbc058814),
	.w2(32'hbc0c11e3),
	.w3(32'hbbef4826),
	.w4(32'hbad25894),
	.w5(32'h3ca8ae7f),
	.w6(32'hbc119911),
	.w7(32'h3c04d4c7),
	.w8(32'h3b23ec5f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4941cb),
	.w1(32'h3c1ba415),
	.w2(32'h3c0571ee),
	.w3(32'h3a415604),
	.w4(32'h3affdad8),
	.w5(32'hbbb5defe),
	.w6(32'hbc1c94c6),
	.w7(32'hbc13b450),
	.w8(32'h39f2e91a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f85922),
	.w1(32'hb9c85c4e),
	.w2(32'hbb93a316),
	.w3(32'hbb8c5aa3),
	.w4(32'hbada3774),
	.w5(32'h3c704424),
	.w6(32'h3ae6c5de),
	.w7(32'h3bdab8ba),
	.w8(32'h3b19be6f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e321b),
	.w1(32'h3aa1557a),
	.w2(32'h3b2f0839),
	.w3(32'h3c787a71),
	.w4(32'h3b27ccc0),
	.w5(32'h3b723f35),
	.w6(32'hbb8ae8b8),
	.w7(32'h3b0f79c9),
	.w8(32'h3b95684c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08aae7),
	.w1(32'h3923f6b1),
	.w2(32'hba8a1370),
	.w3(32'h3b6caaec),
	.w4(32'hbb9694cc),
	.w5(32'hbc4091cc),
	.w6(32'hbb29a6fd),
	.w7(32'h3a848c1e),
	.w8(32'h3a98498f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5bca),
	.w1(32'h3b54f4b7),
	.w2(32'h3c05dbe3),
	.w3(32'hba701fce),
	.w4(32'hbb5e5694),
	.w5(32'h3c155c35),
	.w6(32'h3be593b4),
	.w7(32'hbbd360a8),
	.w8(32'hbc1f9f24),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd34dc),
	.w1(32'h3a9a60a4),
	.w2(32'hbb85d81c),
	.w3(32'hbbfc5a74),
	.w4(32'h3a7520cf),
	.w5(32'hbab7b66d),
	.w6(32'hbc10159b),
	.w7(32'hbabdad84),
	.w8(32'h3b93c124),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab20a3),
	.w1(32'h394144b9),
	.w2(32'hbbb7187c),
	.w3(32'h3b64691f),
	.w4(32'hbba1ff21),
	.w5(32'hbbf268e1),
	.w6(32'hb995b8c2),
	.w7(32'h3af0b075),
	.w8(32'h3c369ca6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9b25e),
	.w1(32'hbaf73704),
	.w2(32'hba1846b4),
	.w3(32'h3bd29bea),
	.w4(32'hb9a57248),
	.w5(32'h3b3e8ef3),
	.w6(32'h3c922c75),
	.w7(32'h3acb5613),
	.w8(32'hbb2565a5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad0ce8),
	.w1(32'hbb6ca33c),
	.w2(32'hbc4cc6c3),
	.w3(32'h3b816e8f),
	.w4(32'hbc38dd64),
	.w5(32'hbc512aae),
	.w6(32'h3aa5b269),
	.w7(32'hbc484ebf),
	.w8(32'hbc104915),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc635e15),
	.w1(32'hbb572647),
	.w2(32'h3b348179),
	.w3(32'hbbc742fc),
	.w4(32'hbbde7ab0),
	.w5(32'h3c633fb0),
	.w6(32'h3bba1975),
	.w7(32'h3a13a51e),
	.w8(32'hbbe2032e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a40c),
	.w1(32'hbb74ddac),
	.w2(32'h3b3066f4),
	.w3(32'hbbae418e),
	.w4(32'hbc2954c4),
	.w5(32'h3b0e9322),
	.w6(32'hbbf5ca57),
	.w7(32'hbb839d7d),
	.w8(32'hba04dab2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5eb93),
	.w1(32'hb9cd8e98),
	.w2(32'hbb5a1560),
	.w3(32'hbc4c7668),
	.w4(32'hbb41995b),
	.w5(32'h3bb66d35),
	.w6(32'hbc350faa),
	.w7(32'h3b599570),
	.w8(32'h3a928826),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a931933),
	.w1(32'hbb303c36),
	.w2(32'hbb9e0140),
	.w3(32'h3bc46900),
	.w4(32'hbae8fc38),
	.w5(32'hbbd2f1e3),
	.w6(32'h3aa8ea63),
	.w7(32'h3b8cf78f),
	.w8(32'hb9df771c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1177),
	.w1(32'h3aadaebf),
	.w2(32'hbb6c5bc2),
	.w3(32'hbc1700cf),
	.w4(32'hbb6dd055),
	.w5(32'h3c141070),
	.w6(32'hbb0098ea),
	.w7(32'hbbba583d),
	.w8(32'hbae513a8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ad9a),
	.w1(32'h3bc7f5fb),
	.w2(32'h3b3ed027),
	.w3(32'hbc14c424),
	.w4(32'hba469439),
	.w5(32'hbaf7baa2),
	.w6(32'hbacae362),
	.w7(32'hbab3e5fe),
	.w8(32'h3af78142),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973200),
	.w1(32'h3ac8e43e),
	.w2(32'hbb1ac9ae),
	.w3(32'h3b28e980),
	.w4(32'h3a3bac8b),
	.w5(32'h39201cc1),
	.w6(32'hbafc9d7b),
	.w7(32'hb888cba6),
	.w8(32'hbbddecb5),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3705c3),
	.w1(32'hbb1de0af),
	.w2(32'h3abe9300),
	.w3(32'hbb7e4e7b),
	.w4(32'hbb876481),
	.w5(32'h3b115a61),
	.w6(32'hbba7d46e),
	.w7(32'hba246bf7),
	.w8(32'hbb961cb1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d430c),
	.w1(32'h3b3ece22),
	.w2(32'hbb0b2566),
	.w3(32'hbbce07a5),
	.w4(32'h3c5e296c),
	.w5(32'h3b0082b5),
	.w6(32'h3b12612d),
	.w7(32'hbb84df31),
	.w8(32'hbc1a85c1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8697f2),
	.w1(32'h3a666e71),
	.w2(32'hbb247c1a),
	.w3(32'hbb8911d3),
	.w4(32'hbb10b856),
	.w5(32'hbbfc722e),
	.w6(32'h3b956f93),
	.w7(32'h3aa98ff4),
	.w8(32'hbbc62a82),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf0b45),
	.w1(32'h3bac0e27),
	.w2(32'h3c148170),
	.w3(32'hbbf36458),
	.w4(32'h3c53dc3d),
	.w5(32'h3c6755e2),
	.w6(32'h3b3c6aaf),
	.w7(32'h3bba8124),
	.w8(32'h3b946805),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12484c),
	.w1(32'hbad5f487),
	.w2(32'hb9ed84fb),
	.w3(32'h3aad44eb),
	.w4(32'hbbbe0ce9),
	.w5(32'h3b8a835e),
	.w6(32'hbbb79348),
	.w7(32'hbbb10a88),
	.w8(32'hbc041299),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac6b91),
	.w1(32'hba669df0),
	.w2(32'h3b2cbc18),
	.w3(32'h39b5ffab),
	.w4(32'hbb5c28a6),
	.w5(32'h3cb0da2d),
	.w6(32'hbc109ef7),
	.w7(32'h3b7a3b4d),
	.w8(32'h3ba5bf42),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0426ef),
	.w1(32'hbbe661ca),
	.w2(32'hbc1d9658),
	.w3(32'h3b0f2951),
	.w4(32'hbc2fb50d),
	.w5(32'h3cae9370),
	.w6(32'hbbad691f),
	.w7(32'h39c0e5d3),
	.w8(32'h3c1645fc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e16b3),
	.w1(32'hbb1eb719),
	.w2(32'h3babb0e3),
	.w3(32'h3bba5c23),
	.w4(32'hbbe2a6d4),
	.w5(32'h3b0f46e8),
	.w6(32'hbbe26ea3),
	.w7(32'h3b2c96bb),
	.w8(32'h3b1e992e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6e68),
	.w1(32'hbbd3df00),
	.w2(32'h3a180b16),
	.w3(32'hbae3fb58),
	.w4(32'hbc23ed29),
	.w5(32'hbb16c3e3),
	.w6(32'hba7e0275),
	.w7(32'hbbbb5c0a),
	.w8(32'hbbdd1d63),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a5bf),
	.w1(32'h3b38d1e0),
	.w2(32'hba81c9f8),
	.w3(32'hba147cfa),
	.w4(32'hbaf7d23d),
	.w5(32'hbc016b4b),
	.w6(32'hbae0760c),
	.w7(32'hbbdf542e),
	.w8(32'hbb006326),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856d96),
	.w1(32'hbc4b6f84),
	.w2(32'hbc657c63),
	.w3(32'hb8c07aca),
	.w4(32'hbbf01f3b),
	.w5(32'h3c34aca4),
	.w6(32'hbb3b5564),
	.w7(32'h3c015859),
	.w8(32'hb93e200a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be61f28),
	.w1(32'hbc29fba4),
	.w2(32'h3a7f7024),
	.w3(32'h398e85dd),
	.w4(32'hbc18542e),
	.w5(32'h3b477996),
	.w6(32'hbc2b8c11),
	.w7(32'hbc00b1fa),
	.w8(32'hbc09801b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3762),
	.w1(32'h3be1a502),
	.w2(32'h3baad737),
	.w3(32'hbc067bdf),
	.w4(32'hbb9e6f2b),
	.w5(32'h3bd872e5),
	.w6(32'hbc80085e),
	.w7(32'hbbe40b39),
	.w8(32'h3a2c9301),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e470d),
	.w1(32'hbb62592d),
	.w2(32'h3ca78122),
	.w3(32'hbb150549),
	.w4(32'hbbddd2a4),
	.w5(32'h3cbe7175),
	.w6(32'h3c0d06db),
	.w7(32'h398e637c),
	.w8(32'hbc27490b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a84b),
	.w1(32'hbbb343fc),
	.w2(32'hbc09a69a),
	.w3(32'hbc89bce9),
	.w4(32'hbbb4f483),
	.w5(32'h3b6ec671),
	.w6(32'hbcac7c92),
	.w7(32'h3b17f782),
	.w8(32'h3c00677b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aea14),
	.w1(32'hbb9aca36),
	.w2(32'hbc053792),
	.w3(32'hbafaf5a9),
	.w4(32'hbb8fcb2f),
	.w5(32'hbc33dc49),
	.w6(32'h3c42581c),
	.w7(32'hbb971821),
	.w8(32'hbba55903),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdae09),
	.w1(32'hb9e08043),
	.w2(32'hbc17cf5c),
	.w3(32'hb9fea207),
	.w4(32'hbb62edf9),
	.w5(32'hbb30c59e),
	.w6(32'h39cd6a5e),
	.w7(32'h3a83d773),
	.w8(32'h3a9c339a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf2ad),
	.w1(32'h3a32795e),
	.w2(32'h3b7ecdab),
	.w3(32'h3b8cd614),
	.w4(32'h3ae9a7fd),
	.w5(32'hbc2e9de6),
	.w6(32'h3ae8e655),
	.w7(32'hbb99b2d9),
	.w8(32'hbbb4e8c3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd09610),
	.w1(32'hbb152010),
	.w2(32'hbb335cf4),
	.w3(32'hbaeeaeed),
	.w4(32'h38dc0c1e),
	.w5(32'hbbd0376e),
	.w6(32'h3b2d6ee2),
	.w7(32'h3a9ac54f),
	.w8(32'hba8077a1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac7da),
	.w1(32'hbc0d0d85),
	.w2(32'h3b8d1ce3),
	.w3(32'hbac2ce6e),
	.w4(32'hbaa39215),
	.w5(32'hbb5739f8),
	.w6(32'hbb50a9ea),
	.w7(32'hb9efe123),
	.w8(32'h3b00f009),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64bb47),
	.w1(32'h3bbca51f),
	.w2(32'h3a9b062c),
	.w3(32'hba42c7bf),
	.w4(32'h3b373cf3),
	.w5(32'h3bbfaeee),
	.w6(32'hba045744),
	.w7(32'h3b0387f8),
	.w8(32'hbb287eab),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d75f),
	.w1(32'h3aab255f),
	.w2(32'hbbfa27db),
	.w3(32'h3ac13ce0),
	.w4(32'hbb7520c8),
	.w5(32'hbbd2d125),
	.w6(32'hbace16a9),
	.w7(32'hbae67938),
	.w8(32'h3bb01dd1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e8d4),
	.w1(32'h3b848c06),
	.w2(32'hbbd6baad),
	.w3(32'h3b5fd87f),
	.w4(32'h3b7c2eb8),
	.w5(32'h3c36cf52),
	.w6(32'h3b1ecdc2),
	.w7(32'h3b4cf07e),
	.w8(32'h3b3e4d23),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3269a2),
	.w1(32'hbc26e0d3),
	.w2(32'hbcb35b83),
	.w3(32'h3b87db19),
	.w4(32'hbca1eeb8),
	.w5(32'h3c34e721),
	.w6(32'h3c018b1d),
	.w7(32'h3c067d96),
	.w8(32'h3c7dd1b6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94a500),
	.w1(32'h3a5bed58),
	.w2(32'hba8f85d7),
	.w3(32'h3bb0a1ff),
	.w4(32'hbbc8bf7c),
	.w5(32'hbb8ef0b7),
	.w6(32'hbc68d5f3),
	.w7(32'hbb8a2ce1),
	.w8(32'hbc0375ca),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4026b4),
	.w1(32'hbb3f43d3),
	.w2(32'hbba38723),
	.w3(32'h3beaeb07),
	.w4(32'hbab88f55),
	.w5(32'h3b5a765b),
	.w6(32'h3be881de),
	.w7(32'hbb834d19),
	.w8(32'h3bd9c37a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32d94a),
	.w1(32'h3b363986),
	.w2(32'hb9f5fdad),
	.w3(32'h3b73034c),
	.w4(32'h3b82f8ea),
	.w5(32'hbb84e097),
	.w6(32'h3bc4a08f),
	.w7(32'hbb6a99d2),
	.w8(32'hbbbd75da),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba631b46),
	.w1(32'h39454284),
	.w2(32'h3b658a88),
	.w3(32'h3bf5b756),
	.w4(32'h3b9c328b),
	.w5(32'h3b595176),
	.w6(32'h3aa5634b),
	.w7(32'h3b0ecf3f),
	.w8(32'hba425fb5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae18741),
	.w1(32'hbb3fb929),
	.w2(32'hbb1f3f6a),
	.w3(32'hba82958f),
	.w4(32'hba92abc6),
	.w5(32'h3bfa0ca0),
	.w6(32'h3b7cf4d0),
	.w7(32'h3af36ed5),
	.w8(32'hbb951ac4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18717f),
	.w1(32'hbbee1981),
	.w2(32'hbc4f2213),
	.w3(32'hbbf623e2),
	.w4(32'h3b241444),
	.w5(32'hbb9207bf),
	.w6(32'hbbb34320),
	.w7(32'hbbf72be8),
	.w8(32'hbc00b3cb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901713),
	.w1(32'hbb481fe9),
	.w2(32'h3938882f),
	.w3(32'h3a7c160b),
	.w4(32'hbb9adecc),
	.w5(32'h3b1dcc77),
	.w6(32'h3c0011c5),
	.w7(32'hb98372a2),
	.w8(32'h3bb94b26),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d16a),
	.w1(32'hb930c1f6),
	.w2(32'hbba858c6),
	.w3(32'h3bcc548b),
	.w4(32'hbb737145),
	.w5(32'hbb65f6d2),
	.w6(32'h3b1887b1),
	.w7(32'h3b78de1e),
	.w8(32'h3b2ab9e2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f9f8),
	.w1(32'h3b63a615),
	.w2(32'hbb5d47b7),
	.w3(32'hbaee352a),
	.w4(32'hbb215780),
	.w5(32'h3c10a61e),
	.w6(32'h3c4168ad),
	.w7(32'hbb44ad75),
	.w8(32'h3baf18d9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9b81),
	.w1(32'h3a2ceddf),
	.w2(32'hbba6b649),
	.w3(32'h3abc095b),
	.w4(32'h3ba716c0),
	.w5(32'h3a0944e0),
	.w6(32'h3c4540a7),
	.w7(32'h3b3c69d5),
	.w8(32'h3ad42387),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba4354),
	.w1(32'hbbad35f7),
	.w2(32'hbb18df00),
	.w3(32'h3ae86775),
	.w4(32'hba2a7140),
	.w5(32'hbac32aff),
	.w6(32'h3baf6836),
	.w7(32'h3b082930),
	.w8(32'h3b236530),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e36a9),
	.w1(32'h39f1d8f5),
	.w2(32'h3bea2791),
	.w3(32'h3b801eb6),
	.w4(32'h3b968762),
	.w5(32'h3d010345),
	.w6(32'h3abf4fa5),
	.w7(32'h3c006738),
	.w8(32'hbb05f850),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001ab4),
	.w1(32'hbbebac06),
	.w2(32'hbbc5698f),
	.w3(32'hb9e43358),
	.w4(32'hbbfc326d),
	.w5(32'hbc12885b),
	.w6(32'hba443a6e),
	.w7(32'hbb8dfc3b),
	.w8(32'hbc5d5825),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad114),
	.w1(32'hbb288543),
	.w2(32'hbc28abc6),
	.w3(32'hbc340596),
	.w4(32'hbc29994b),
	.w5(32'hbc8675d0),
	.w6(32'hbc291dd7),
	.w7(32'hbbb6362f),
	.w8(32'hbb94df95),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule