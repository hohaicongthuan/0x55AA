module layer_8_featuremap_43(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c991849),
	.w1(32'h3bbde4da),
	.w2(32'h3c312e2e),
	.w3(32'h3c8d2f53),
	.w4(32'h3c113269),
	.w5(32'h3bda1586),
	.w6(32'h3c6116ff),
	.w7(32'h3ca23bfb),
	.w8(32'hbb3cebff),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc479cae),
	.w1(32'h391d811d),
	.w2(32'h3c226b22),
	.w3(32'hbc314ff8),
	.w4(32'hb9d6ef5e),
	.w5(32'h3b2fbf92),
	.w6(32'h3a9ed197),
	.w7(32'h3b9af481),
	.w8(32'hbc365d3f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc669341),
	.w1(32'h3a8a8964),
	.w2(32'h3c6b80a7),
	.w3(32'hbc4191cc),
	.w4(32'h3aec85fe),
	.w5(32'h3beef870),
	.w6(32'hbb41997f),
	.w7(32'h3b8dda06),
	.w8(32'hb8e1322e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042081),
	.w1(32'h3a798cb2),
	.w2(32'h3c986cdf),
	.w3(32'hbbeb8774),
	.w4(32'h3c680264),
	.w5(32'h3c439a4e),
	.w6(32'h394e17de),
	.w7(32'hbc3de142),
	.w8(32'hbc279426),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaad4cd),
	.w1(32'h3a80a5e1),
	.w2(32'h3cde732c),
	.w3(32'hbc96e4b0),
	.w4(32'h39255ab2),
	.w5(32'h3c90bca6),
	.w6(32'h3bbb578f),
	.w7(32'h3cb06d18),
	.w8(32'hbce3ca24),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd413a5a),
	.w1(32'h3a625de8),
	.w2(32'h3db78269),
	.w3(32'hbd0f202f),
	.w4(32'h3b1ae19b),
	.w5(32'h3d259312),
	.w6(32'hbbd223dd),
	.w7(32'h3d537ef1),
	.w8(32'hbb0f1d51),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6a03),
	.w1(32'h3b8077a2),
	.w2(32'h3cb4a07a),
	.w3(32'hbc14305b),
	.w4(32'h3b79cf61),
	.w5(32'h3c64bc0c),
	.w6(32'h3ba9676d),
	.w7(32'h3c7bf499),
	.w8(32'hbc5c5af6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfae6a),
	.w1(32'hbc5d70ce),
	.w2(32'h3c992f3a),
	.w3(32'hbcce16dc),
	.w4(32'hbc8505e9),
	.w5(32'h3a31a53a),
	.w6(32'h3b5c004b),
	.w7(32'h3c5125fc),
	.w8(32'hbc92f85f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc698ac4),
	.w1(32'h3be787f1),
	.w2(32'h3cbcaef6),
	.w3(32'hbc74023e),
	.w4(32'h3ada82af),
	.w5(32'h3c0bfcfa),
	.w6(32'h3c04fc53),
	.w7(32'h3c5d3ebb),
	.w8(32'hbc03e724),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9749db),
	.w1(32'hbc3fcaf0),
	.w2(32'hbc3cc487),
	.w3(32'hbc149552),
	.w4(32'h3b3df01b),
	.w5(32'h3c07f311),
	.w6(32'h3c3c229b),
	.w7(32'hba983688),
	.w8(32'hbcb69e10),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e17e4),
	.w1(32'h3abb9fc6),
	.w2(32'h3ceb97cf),
	.w3(32'hbc26bc9c),
	.w4(32'h3c24e7e5),
	.w5(32'h3c71d40c),
	.w6(32'h3bca74cd),
	.w7(32'h3c8c3224),
	.w8(32'hbc2665ce),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7ab22),
	.w1(32'hbb65d412),
	.w2(32'h3b4bf09f),
	.w3(32'hbbf2a7eb),
	.w4(32'h3b5fea94),
	.w5(32'h3ac2c2ba),
	.w6(32'h3c2dc8b5),
	.w7(32'h3ca398b8),
	.w8(32'hbbe96d06),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc981432),
	.w1(32'h3b88d01e),
	.w2(32'h3cbd6b7e),
	.w3(32'hbc9d1515),
	.w4(32'hbaf47cb1),
	.w5(32'h3c25adf1),
	.w6(32'h3ad2f563),
	.w7(32'h3c5e70f1),
	.w8(32'hbcfa649a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2fe21c),
	.w1(32'hba326cec),
	.w2(32'h3dc03d28),
	.w3(32'hbd166dd8),
	.w4(32'hbc778da5),
	.w5(32'h3d2662e9),
	.w6(32'hbb959a8f),
	.w7(32'h3d63303e),
	.w8(32'hbc6faf1e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8e7f9),
	.w1(32'h3ae8518c),
	.w2(32'h3d4ec901),
	.w3(32'hbca62367),
	.w4(32'hbb60788a),
	.w5(32'h3cc064ac),
	.w6(32'h3b29628c),
	.w7(32'h3cf89d2d),
	.w8(32'h3a1533c7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef5723),
	.w1(32'hbbec9997),
	.w2(32'h3bd0be35),
	.w3(32'hbaeafd70),
	.w4(32'hbc3b53ea),
	.w5(32'hbb3ea4d6),
	.w6(32'hbc187844),
	.w7(32'hba019206),
	.w8(32'h3ab0d5a1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9376f92),
	.w1(32'hbb6b4a38),
	.w2(32'hbccc4da9),
	.w3(32'hbc9cdf02),
	.w4(32'hbb245c18),
	.w5(32'h3b8f1241),
	.w6(32'h3bf8bcf4),
	.w7(32'h3ac8b021),
	.w8(32'hbc9906ca),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2f700),
	.w1(32'hb957fba0),
	.w2(32'h3c4e1102),
	.w3(32'hbc8b7322),
	.w4(32'hbb97cea9),
	.w5(32'h3bdebf9a),
	.w6(32'h3b9c15ff),
	.w7(32'h3c8730f8),
	.w8(32'hbbf79d80),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa3757),
	.w1(32'hbcc4e180),
	.w2(32'h3bac0aa6),
	.w3(32'h3be54d52),
	.w4(32'hbb8ba1a6),
	.w5(32'hbc3413ad),
	.w6(32'h3cca1b9c),
	.w7(32'h3ccb5ab0),
	.w8(32'h3b656da7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc845e52),
	.w1(32'hbd0128d6),
	.w2(32'hbd016665),
	.w3(32'h3a19b255),
	.w4(32'h3b77cd73),
	.w5(32'hbb825856),
	.w6(32'h3c21ed54),
	.w7(32'h3c068401),
	.w8(32'hbc65a684),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9eb271),
	.w1(32'hbb9810fb),
	.w2(32'hbb6b8126),
	.w3(32'hbc856b78),
	.w4(32'h3a96bdcd),
	.w5(32'h3c2022b5),
	.w6(32'hbb29e137),
	.w7(32'h3c761cce),
	.w8(32'hbc681eb0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe879e),
	.w1(32'h3c25c96d),
	.w2(32'h3d16411a),
	.w3(32'hbcd0fee5),
	.w4(32'h3adaa2c0),
	.w5(32'h3cbfd1dc),
	.w6(32'h3c0b996b),
	.w7(32'h3cd6a415),
	.w8(32'h3cf40d02),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1b5703),
	.w1(32'h3c358a74),
	.w2(32'hbda8cbd1),
	.w3(32'h3df08735),
	.w4(32'h3c8ab6f8),
	.w5(32'hbd3ed676),
	.w6(32'h3cb697d4),
	.w7(32'hbd1c4b93),
	.w8(32'hba98c384),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ae162),
	.w1(32'h3b2723af),
	.w2(32'h3c26af42),
	.w3(32'hbb860c2d),
	.w4(32'hbb33b411),
	.w5(32'hbb251754),
	.w6(32'h3bb44bfc),
	.w7(32'h3b8cf9dc),
	.w8(32'hbcbe2678),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd21aedb),
	.w1(32'hbc14efea),
	.w2(32'h3c8e2215),
	.w3(32'hbd1a2a12),
	.w4(32'hbc2b0bf0),
	.w5(32'h3c77dec1),
	.w6(32'hbc0a430b),
	.w7(32'h3ca0e794),
	.w8(32'h3ce9aa97),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc75e5b),
	.w1(32'h3c2639f0),
	.w2(32'hbd8ab18a),
	.w3(32'h3d8bb472),
	.w4(32'h3c1116a7),
	.w5(32'hbd0723ec),
	.w6(32'h3acb8880),
	.w7(32'hbd113f61),
	.w8(32'h3cf38c59),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d80fc2d),
	.w1(32'h3b531a70),
	.w2(32'hbd404dce),
	.w3(32'h3d287386),
	.w4(32'hbad31ff4),
	.w5(32'hbcc84087),
	.w6(32'hbc5bfacc),
	.w7(32'hbd14db70),
	.w8(32'h3916f47b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1fcfc),
	.w1(32'hbcc7c637),
	.w2(32'hbe248562),
	.w3(32'hbcc13b01),
	.w4(32'hbd3de599),
	.w5(32'hbd500613),
	.w6(32'hbc0b88bb),
	.w7(32'hbb1d060e),
	.w8(32'hbd9f6c8d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a8036),
	.w1(32'hbc833442),
	.w2(32'hbc2095a2),
	.w3(32'h3ba702f0),
	.w4(32'hbcb800f8),
	.w5(32'hbc822f23),
	.w6(32'hbc2f167e),
	.w7(32'hbbaf8f01),
	.w8(32'hbb5c2d1f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b229a),
	.w1(32'hba88d7c9),
	.w2(32'h3c13ddde),
	.w3(32'hbc347b0b),
	.w4(32'hba985945),
	.w5(32'h3b09db15),
	.w6(32'hba313ac9),
	.w7(32'h3bb73f81),
	.w8(32'hbc8a8341),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60c447),
	.w1(32'h3c46690e),
	.w2(32'h3d070446),
	.w3(32'h3cd3c48b),
	.w4(32'h3c801a53),
	.w5(32'hbbac4943),
	.w6(32'h3c99cb85),
	.w7(32'h3d163709),
	.w8(32'hbc750b05),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdec1d9),
	.w1(32'hbc1ffbd7),
	.w2(32'h3c1a5318),
	.w3(32'hbd0523e9),
	.w4(32'hbc2c76a8),
	.w5(32'h3c9581a9),
	.w6(32'hbc2d2db1),
	.w7(32'h3cc958a0),
	.w8(32'h3bc734b7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb951aa4),
	.w1(32'h3c31efa6),
	.w2(32'h3c2223d2),
	.w3(32'h3c870fc7),
	.w4(32'h3c2c5dc0),
	.w5(32'hbbceed13),
	.w6(32'hbb025719),
	.w7(32'hbc03fedf),
	.w8(32'hbc4b8951),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba993e75),
	.w1(32'hbbc5fe81),
	.w2(32'hbc29e260),
	.w3(32'hbb41516c),
	.w4(32'h3b54be19),
	.w5(32'h3af9292e),
	.w6(32'h3ab6d50a),
	.w7(32'h3c1846f9),
	.w8(32'hbcc2a631),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1fd22c),
	.w1(32'h3bd6c999),
	.w2(32'h3db57f9c),
	.w3(32'hbcf67176),
	.w4(32'hbb83e18f),
	.w5(32'h3d407e0d),
	.w6(32'hba879293),
	.w7(32'h3d590ec7),
	.w8(32'h3ae2fd80),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cedfe),
	.w1(32'hbc22f46f),
	.w2(32'h3ab6ea7c),
	.w3(32'hbc8ac057),
	.w4(32'hbc7e6496),
	.w5(32'hbc1ae7ce),
	.w6(32'h3b96ac1a),
	.w7(32'h3c560e1e),
	.w8(32'hbc6f517b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd46685),
	.w1(32'hb992dc4d),
	.w2(32'h3c9628e2),
	.w3(32'hbcbb7433),
	.w4(32'hbbb9177d),
	.w5(32'h3c998b9b),
	.w6(32'h3bb2948d),
	.w7(32'h3ce4fd44),
	.w8(32'hbc379f4c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68c9a9),
	.w1(32'h3b6a4990),
	.w2(32'h3c947961),
	.w3(32'hbc34ad42),
	.w4(32'h3b7251e1),
	.w5(32'h3c49723c),
	.w6(32'h3bfae111),
	.w7(32'h3c76247e),
	.w8(32'hbc9f53ba),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd41bcaa),
	.w1(32'h3b6866c0),
	.w2(32'h3db2c3a0),
	.w3(32'hbd075876),
	.w4(32'hbbd1ae78),
	.w5(32'h3d289a08),
	.w6(32'h3b93fbae),
	.w7(32'h3d4d1651),
	.w8(32'hbba5c2ff),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1a45),
	.w1(32'h3a729412),
	.w2(32'h3be2e1ba),
	.w3(32'hbbe03bd7),
	.w4(32'hb9b1a81a),
	.w5(32'h3c52a755),
	.w6(32'h3b3a421a),
	.w7(32'h3c805b84),
	.w8(32'h3c86bab6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7219ff),
	.w1(32'h3bfbb6f1),
	.w2(32'hbd280552),
	.w3(32'h3ceeb6b1),
	.w4(32'h3beb7fb5),
	.w5(32'hbcc1843f),
	.w6(32'hbb07527e),
	.w7(32'hbc2d0736),
	.w8(32'h3b75ffbd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9526984),
	.w1(32'hbc1581de),
	.w2(32'hbc646bcd),
	.w3(32'hbbb267b9),
	.w4(32'hbbd80aef),
	.w5(32'hbc88aadf),
	.w6(32'hbaa1e44c),
	.w7(32'hbbeb04dd),
	.w8(32'hbc7c71e5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd8f3),
	.w1(32'hbc52c548),
	.w2(32'hbc728022),
	.w3(32'hbc1dd3e0),
	.w4(32'hbd232cd3),
	.w5(32'hbc868fd2),
	.w6(32'hbced65c0),
	.w7(32'hbc7a3d8b),
	.w8(32'h3b6457a3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bf1ce),
	.w1(32'hbaca6e4a),
	.w2(32'hbc9dab54),
	.w3(32'h3bd63061),
	.w4(32'h3b0b151f),
	.w5(32'hbbcf7b87),
	.w6(32'hbb2ed49a),
	.w7(32'hbb932d1c),
	.w8(32'hba907212),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d199e5b),
	.w1(32'hba34e585),
	.w2(32'hbcbbb7e4),
	.w3(32'h3cdb2db0),
	.w4(32'h3c25525a),
	.w5(32'hbc78867d),
	.w6(32'h3c78b309),
	.w7(32'hbb912bd1),
	.w8(32'hbbb1676b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ccdc5),
	.w1(32'hbc7a3f03),
	.w2(32'hbcda6d66),
	.w3(32'hbb9ee5b9),
	.w4(32'h3aad9090),
	.w5(32'hbc87daa8),
	.w6(32'hbb273c80),
	.w7(32'hbb81f800),
	.w8(32'h3c138608),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bdc3f),
	.w1(32'hbcae0121),
	.w2(32'hbc45f967),
	.w3(32'h3bbb626f),
	.w4(32'h3c732037),
	.w5(32'hba2bdd98),
	.w6(32'h3cc481e2),
	.w7(32'h3cb382dc),
	.w8(32'hbc7273bc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c0dad),
	.w1(32'hbbc5593b),
	.w2(32'hbd221a3f),
	.w3(32'hbb1da0f2),
	.w4(32'hbc7f243e),
	.w5(32'hbcc9360c),
	.w6(32'h3c54090d),
	.w7(32'hbbe0c533),
	.w8(32'hbc63971e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd910a5),
	.w1(32'hbb349dd5),
	.w2(32'h3d14e27b),
	.w3(32'hbcc38486),
	.w4(32'hbcaf5b03),
	.w5(32'h3a9f8247),
	.w6(32'h3bd7e06a),
	.w7(32'h3cbd0ee3),
	.w8(32'h3a14bbaf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1b010),
	.w1(32'h3ac091c1),
	.w2(32'hbc9bc1a7),
	.w3(32'h3c30b2c0),
	.w4(32'h3c971f92),
	.w5(32'hbc1279fa),
	.w6(32'h3ae2d07b),
	.w7(32'hbb94387c),
	.w8(32'h3c0f46de),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d6c1f),
	.w1(32'h3beb88ca),
	.w2(32'hbb09255e),
	.w3(32'hbbdc043a),
	.w4(32'h3bee64a1),
	.w5(32'h3bf296d4),
	.w6(32'hbb57ae70),
	.w7(32'h3ba8f20e),
	.w8(32'h3c7b875a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1d326a),
	.w1(32'hbc223283),
	.w2(32'hbcd4132e),
	.w3(32'h3d0cf73a),
	.w4(32'hb9d0f7c2),
	.w5(32'hbca164c3),
	.w6(32'h3c8b3d2e),
	.w7(32'h3bda327e),
	.w8(32'hbb5f30c9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c680152),
	.w1(32'h3bb1da86),
	.w2(32'hbb869218),
	.w3(32'h3bc8a55b),
	.w4(32'h3abf1333),
	.w5(32'hbc971863),
	.w6(32'hbae6d679),
	.w7(32'hbac1feb9),
	.w8(32'hb94ee62d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d1a3b),
	.w1(32'hbbab7c36),
	.w2(32'hbc0f43f7),
	.w3(32'h3c17049f),
	.w4(32'h3b567a54),
	.w5(32'hbbca576d),
	.w6(32'h3c3dfd23),
	.w7(32'h3b29eb93),
	.w8(32'hbbd4e9d6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f001f),
	.w1(32'h3c0c3566),
	.w2(32'hbbb5c1b1),
	.w3(32'hbcb9e084),
	.w4(32'hbc72230d),
	.w5(32'hb9fb8d2e),
	.w6(32'hbb39682a),
	.w7(32'hbc302676),
	.w8(32'hbbe6d776),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1a4de),
	.w1(32'hbb1e44af),
	.w2(32'hbd81a2cb),
	.w3(32'h3c8f0ea7),
	.w4(32'h39ea4376),
	.w5(32'hbc8eb47f),
	.w6(32'h3c5159d7),
	.w7(32'h3c10e2fe),
	.w8(32'hbc8ca728),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6faa67),
	.w1(32'h3c6dfd43),
	.w2(32'h3c99051e),
	.w3(32'h3c6091d5),
	.w4(32'h3c3c0e16),
	.w5(32'h3b3833e4),
	.w6(32'hbb1510d2),
	.w7(32'h3bb04508),
	.w8(32'hbbd880db),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c9d6b),
	.w1(32'hbc76f500),
	.w2(32'hbc91fde7),
	.w3(32'hbc63f38c),
	.w4(32'hbd2bbd88),
	.w5(32'hbcf1feff),
	.w6(32'hbb866928),
	.w7(32'h3ba2d278),
	.w8(32'h3a1fbda5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac60c6),
	.w1(32'h3b83bd06),
	.w2(32'h3b2982d6),
	.w3(32'h3c0e51f0),
	.w4(32'hbbcb3f6c),
	.w5(32'hbb0a0c69),
	.w6(32'hbbaadcc2),
	.w7(32'h3a3ed302),
	.w8(32'hbb453e0b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fce5f),
	.w1(32'h3b4e68b9),
	.w2(32'h3b69ff0d),
	.w3(32'h3b91e258),
	.w4(32'hbb352b02),
	.w5(32'hbbde7c5c),
	.w6(32'hbbf6cc32),
	.w7(32'hbc0b1e3a),
	.w8(32'h3b652c06),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8563e1),
	.w1(32'hbbf0c613),
	.w2(32'hbc1982dd),
	.w3(32'hbc98d1b9),
	.w4(32'h3bb73e34),
	.w5(32'h3b270213),
	.w6(32'h3c29c698),
	.w7(32'h3c1f8a95),
	.w8(32'hbc38740e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4024bd),
	.w1(32'hbac14b00),
	.w2(32'hbcd28661),
	.w3(32'hbc1b57a1),
	.w4(32'hb8bfdb66),
	.w5(32'hbbbbb963),
	.w6(32'hbba030af),
	.w7(32'hbc470cbf),
	.w8(32'h3c795813),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d32b71d),
	.w1(32'h3bc833b6),
	.w2(32'hbd0fbe2d),
	.w3(32'h3ce47194),
	.w4(32'h3c82f60a),
	.w5(32'hbc8177f6),
	.w6(32'h3ca75e0b),
	.w7(32'h3a35616d),
	.w8(32'hbc1eb631),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2294bd),
	.w1(32'hbc7575eb),
	.w2(32'hbc0c2907),
	.w3(32'hbb2c4dc7),
	.w4(32'hbce7dfe0),
	.w5(32'hbc03e80d),
	.w6(32'hbc8ef82c),
	.w7(32'hbc51ba74),
	.w8(32'h3a8a19f1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b3c2b),
	.w1(32'h3b83e40b),
	.w2(32'hbb152160),
	.w3(32'h3b2802d9),
	.w4(32'hb918ad88),
	.w5(32'hbb2380e9),
	.w6(32'h3ad61336),
	.w7(32'hbaad1b57),
	.w8(32'h3a96788f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd12668),
	.w1(32'hbbb728fb),
	.w2(32'hbc46e8f5),
	.w3(32'hbafe2132),
	.w4(32'hbb8e2e58),
	.w5(32'hbbfd533f),
	.w6(32'hb94cf608),
	.w7(32'hbba6a4d1),
	.w8(32'hbb888e2a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fe6f),
	.w1(32'hb8199e09),
	.w2(32'hbc258a8c),
	.w3(32'hba538515),
	.w4(32'h3ad83297),
	.w5(32'hbb4db119),
	.w6(32'hbc1a9b0f),
	.w7(32'hbc04990e),
	.w8(32'hbcc07226),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd33e6),
	.w1(32'h3c0d5b5c),
	.w2(32'hbc93d09c),
	.w3(32'h3c19f54b),
	.w4(32'h3c225dec),
	.w5(32'hbc638f1a),
	.w6(32'hbb850e94),
	.w7(32'h3cacf69b),
	.w8(32'h3b035c13),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd028b2),
	.w1(32'h3ae0624f),
	.w2(32'hbc327f41),
	.w3(32'h3b0efaa2),
	.w4(32'h3b33db2f),
	.w5(32'hbb86a6aa),
	.w6(32'hbb9c7d1b),
	.w7(32'hbc208069),
	.w8(32'h3c693bd7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db11cf6),
	.w1(32'h3cd09746),
	.w2(32'hbd1f6c8f),
	.w3(32'h3d454cac),
	.w4(32'h3ce0e685),
	.w5(32'h3bbbbf64),
	.w6(32'hbc8e6ec8),
	.w7(32'hbc9284d8),
	.w8(32'hbae36919),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c344d),
	.w1(32'h3af02b01),
	.w2(32'hbb7d865c),
	.w3(32'hb9bc2ec4),
	.w4(32'hb7d53592),
	.w5(32'hba8df98e),
	.w6(32'h3b587524),
	.w7(32'hbb03fca8),
	.w8(32'h3b0338f3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a17c4),
	.w1(32'h3ad60027),
	.w2(32'hbc5db6bf),
	.w3(32'h3bc56462),
	.w4(32'h3a772e74),
	.w5(32'hbbe5e828),
	.w6(32'hbb193114),
	.w7(32'hbc4a199c),
	.w8(32'hba54a4a5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d90f),
	.w1(32'h3b07f0d9),
	.w2(32'hbb8fd454),
	.w3(32'hbbaa8fb4),
	.w4(32'hbb288368),
	.w5(32'hba7c427f),
	.w6(32'hbb02f74c),
	.w7(32'hbbca8d62),
	.w8(32'hbca220bd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9c009),
	.w1(32'hbc3ceca9),
	.w2(32'hbd0ba705),
	.w3(32'hbb868f48),
	.w4(32'hbbcb5847),
	.w5(32'hbcc89fa8),
	.w6(32'hbc031a7f),
	.w7(32'h3c6329b2),
	.w8(32'hbc380ad1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a097d08),
	.w1(32'hbba3dfeb),
	.w2(32'hbc421efc),
	.w3(32'hba00c42a),
	.w4(32'hbba7b65e),
	.w5(32'hbbc7e063),
	.w6(32'hbb6e94eb),
	.w7(32'hbbc4bdcd),
	.w8(32'h3b3bc606),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63059),
	.w1(32'h3b4121e8),
	.w2(32'hbc10f0af),
	.w3(32'h3b8416ab),
	.w4(32'h3b362924),
	.w5(32'hbb7cb2b3),
	.w6(32'h3ba9f1db),
	.w7(32'h39d46603),
	.w8(32'hbabf0530),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25346d),
	.w1(32'hbb15dde5),
	.w2(32'hbc1960e1),
	.w3(32'hb9aa3382),
	.w4(32'hbb259ecb),
	.w5(32'hbb75c50e),
	.w6(32'hba94dcbe),
	.w7(32'hbbcc0ac5),
	.w8(32'h3c6c553d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3daf52e3),
	.w1(32'h3c1022c1),
	.w2(32'hbd2fe68c),
	.w3(32'h3d1ea52b),
	.w4(32'h3c515a9f),
	.w5(32'hbbac43db),
	.w6(32'hbc820621),
	.w7(32'hbcd37963),
	.w8(32'h3b88f209),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d086ec6),
	.w1(32'hbbe4ee57),
	.w2(32'hbd5d4e17),
	.w3(32'h3c85f157),
	.w4(32'h3b95c7aa),
	.w5(32'hbcab0cff),
	.w6(32'hbbd9f9ed),
	.w7(32'hbcc33eb0),
	.w8(32'hbbde0f2b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515d14),
	.w1(32'hbb951a9e),
	.w2(32'hbb9645ad),
	.w3(32'hbb70a263),
	.w4(32'hbbaafd11),
	.w5(32'hbabe04b0),
	.w6(32'hbba605a1),
	.w7(32'h39b3eccc),
	.w8(32'hbc372bd2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc936ebb),
	.w1(32'h3b64db94),
	.w2(32'h3cddb8e6),
	.w3(32'h3cabae9a),
	.w4(32'h3c995c6e),
	.w5(32'hbc1a8adc),
	.w6(32'h390cb63d),
	.w7(32'h3ba6c99f),
	.w8(32'h3acbe79b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6e75),
	.w1(32'hbbbf73b8),
	.w2(32'hbb7fe2df),
	.w3(32'h3bce0ea3),
	.w4(32'h3bdcfa13),
	.w5(32'hba939fd1),
	.w6(32'hbbc68474),
	.w7(32'hbbf36f6a),
	.w8(32'hbc2b9dd6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf35dec),
	.w1(32'h3bb8ed93),
	.w2(32'hbcc953a2),
	.w3(32'h3c51e8a0),
	.w4(32'h3c0c55b3),
	.w5(32'hbc1b370c),
	.w6(32'h3c60d388),
	.w7(32'h3c05f318),
	.w8(32'hbaf38290),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd101a9),
	.w1(32'hbc136d06),
	.w2(32'h3cd76f52),
	.w3(32'hbcfb6f0b),
	.w4(32'hbc9a1237),
	.w5(32'hbc120ec4),
	.w6(32'hbc723971),
	.w7(32'h3cfe3902),
	.w8(32'h3c22f08c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d116784),
	.w1(32'hbb671c96),
	.w2(32'hbceebcf7),
	.w3(32'h3caa20aa),
	.w4(32'h3baa6415),
	.w5(32'hbcd712e9),
	.w6(32'h3c861697),
	.w7(32'hbb563563),
	.w8(32'h3bba20ab),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb91d87),
	.w1(32'h3bbde6a3),
	.w2(32'hbc297400),
	.w3(32'h3cfe31fc),
	.w4(32'h3cacd808),
	.w5(32'hbbb7e591),
	.w6(32'h3c03456d),
	.w7(32'hbb19e730),
	.w8(32'hbafca7dc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd047fb8),
	.w1(32'hbae8d4da),
	.w2(32'h3d4e2489),
	.w3(32'hbcd6dd0a),
	.w4(32'hbcd0bf07),
	.w5(32'h3bc80872),
	.w6(32'h3c58ff61),
	.w7(32'h3d04d251),
	.w8(32'hbb540621),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b998e7c),
	.w1(32'h3b2d791e),
	.w2(32'hbbb27450),
	.w3(32'hbad63ebc),
	.w4(32'hbb3aef08),
	.w5(32'hbb8d5737),
	.w6(32'hbbe155dc),
	.w7(32'hbb27cbaa),
	.w8(32'hbaf7dfcc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fe798),
	.w1(32'hbb611bea),
	.w2(32'h3b3d47be),
	.w3(32'h3a8b1018),
	.w4(32'hbc37a6dc),
	.w5(32'hbbd6226f),
	.w6(32'hba2a8b5a),
	.w7(32'hbbf5e9f3),
	.w8(32'hbba85713),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd4d50),
	.w1(32'h3aebaf4d),
	.w2(32'h3d3f3388),
	.w3(32'hbca9b791),
	.w4(32'hbcc29205),
	.w5(32'h3b3d134a),
	.w6(32'h3c89ecda),
	.w7(32'h3d07932b),
	.w8(32'hbbcda3ac),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd852ad),
	.w1(32'hbb0666b0),
	.w2(32'h3d23b7c2),
	.w3(32'hbc8f3133),
	.w4(32'hbc9f0a05),
	.w5(32'h3bb7589f),
	.w6(32'h3c53ba42),
	.w7(32'h3cd0d5b4),
	.w8(32'hbacf19eb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe396f3),
	.w1(32'hbb11736e),
	.w2(32'hbb23239c),
	.w3(32'hb9a3c774),
	.w4(32'hba646842),
	.w5(32'hbbc88be8),
	.w6(32'hbb766dd5),
	.w7(32'hbc37839e),
	.w8(32'hbc11687a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0954b),
	.w1(32'h3c746f2e),
	.w2(32'h3c9a5a9f),
	.w3(32'hbc1ed494),
	.w4(32'hbbadc235),
	.w5(32'h3bc5295f),
	.w6(32'h3b289004),
	.w7(32'h3c51e09e),
	.w8(32'h3ba70838),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e1845),
	.w1(32'h3a4363f6),
	.w2(32'hbc3e30fa),
	.w3(32'h3c11c777),
	.w4(32'h3b134494),
	.w5(32'hbc044ac1),
	.w6(32'h3b53aad5),
	.w7(32'h38080dd2),
	.w8(32'h3bd8f295),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badd10b),
	.w1(32'hbc352b1a),
	.w2(32'hbc53b7ca),
	.w3(32'hbbdc407c),
	.w4(32'h3cbb88ec),
	.w5(32'h3cd6038d),
	.w6(32'h3c8a9e79),
	.w7(32'hbb00109b),
	.w8(32'hbbd9328d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bbd7e),
	.w1(32'h3b3525b4),
	.w2(32'hbc51bb11),
	.w3(32'h3c8a1d66),
	.w4(32'h3c13a86d),
	.w5(32'hbc85db5b),
	.w6(32'h3c83cc2e),
	.w7(32'hbc459a95),
	.w8(32'hbac1745b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3f840f),
	.w1(32'h3c1e2ad2),
	.w2(32'hbcea8017),
	.w3(32'h3c5f03a7),
	.w4(32'h3c06e492),
	.w5(32'hbc286bff),
	.w6(32'h3c70e0ed),
	.w7(32'h3c1f1712),
	.w8(32'h3a19c328),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d33e0),
	.w1(32'hbb7ac0cc),
	.w2(32'h3cb96305),
	.w3(32'hbacbfc70),
	.w4(32'hbb568e48),
	.w5(32'h3a195377),
	.w6(32'h3c1da471),
	.w7(32'hbb4c59f7),
	.w8(32'h3c52d81d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d52782a),
	.w1(32'h3b8c206d),
	.w2(32'hbce96583),
	.w3(32'h3cc355b6),
	.w4(32'h3c027b80),
	.w5(32'hbae386ea),
	.w6(32'hbca89ecf),
	.w7(32'hbcd17c09),
	.w8(32'hb9b77b33),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf40a9),
	.w1(32'h3b0ad20f),
	.w2(32'hbbc2719c),
	.w3(32'h3a1df80b),
	.w4(32'h3ab011fe),
	.w5(32'hba3e44a1),
	.w6(32'hbb52c9e1),
	.w7(32'hbb81429d),
	.w8(32'h3b081d2b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409160),
	.w1(32'hbc0431f8),
	.w2(32'hbb89ed82),
	.w3(32'hbac06297),
	.w4(32'hbb4be374),
	.w5(32'hbc3bfb3c),
	.w6(32'hbb50c89e),
	.w7(32'hbc503048),
	.w8(32'h3b937965),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf43e15),
	.w1(32'hba40a723),
	.w2(32'hbc41be20),
	.w3(32'h3bbb9107),
	.w4(32'h3b8cda1a),
	.w5(32'hbb5f2221),
	.w6(32'h3aaa223d),
	.w7(32'hbafa251c),
	.w8(32'h3bc0172b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d562c9f),
	.w1(32'h3bd084f0),
	.w2(32'hbd775a1d),
	.w3(32'h3cdc9358),
	.w4(32'h3cc089f3),
	.w5(32'hbc3281e3),
	.w6(32'hbcf0f475),
	.w7(32'hbd3b9ae2),
	.w8(32'hbb1ed5a3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c92d1),
	.w1(32'hbc1c6d7a),
	.w2(32'hbb9094fb),
	.w3(32'h3a32e930),
	.w4(32'hbb7dd787),
	.w5(32'hbb4cf07b),
	.w6(32'hbc399231),
	.w7(32'hbcabb455),
	.w8(32'hbc016177),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87871f),
	.w1(32'hb949d0da),
	.w2(32'h3ca92014),
	.w3(32'hbc5526fc),
	.w4(32'hbc157d30),
	.w5(32'h3b770591),
	.w6(32'h3b156095),
	.w7(32'h3c3b5da2),
	.w8(32'hb9cefd86),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c533a6a),
	.w1(32'h3ac8e605),
	.w2(32'hbc5b3fda),
	.w3(32'h3b4fbb3e),
	.w4(32'hba9804f0),
	.w5(32'hbc02a872),
	.w6(32'hbbfa67f2),
	.w7(32'hbb8ddd60),
	.w8(32'hbc3419f1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc70223),
	.w1(32'h3a9a9804),
	.w2(32'hbb4604d2),
	.w3(32'h3bc1bd79),
	.w4(32'h3aceb5be),
	.w5(32'hbb757bff),
	.w6(32'h3beae0a7),
	.w7(32'h3b29adc8),
	.w8(32'hbbb1d5f6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb041a71),
	.w1(32'hb92574a9),
	.w2(32'hbaff9fcc),
	.w3(32'hbb61bb31),
	.w4(32'hb937e0fc),
	.w5(32'hbb1d6f06),
	.w6(32'hbab4437f),
	.w7(32'hb9398186),
	.w8(32'hbb1b7781),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ff48),
	.w1(32'h3bc78697),
	.w2(32'h3bd4e39a),
	.w3(32'h3a55bc01),
	.w4(32'h3bb6894f),
	.w5(32'h3be510ee),
	.w6(32'hb7561068),
	.w7(32'h3b575d49),
	.w8(32'h3b8d656d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a155b5a),
	.w1(32'hbb8aebe6),
	.w2(32'hbb828a6f),
	.w3(32'hbb008072),
	.w4(32'hbba7f3da),
	.w5(32'hbbe4fadc),
	.w6(32'h3a9f42c4),
	.w7(32'hbbbeb673),
	.w8(32'hbbe98d10),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8153c8),
	.w1(32'hbb43f7b1),
	.w2(32'hbc44febd),
	.w3(32'hbc162e55),
	.w4(32'hbbb6a516),
	.w5(32'hbc2dff28),
	.w6(32'h3ae0dedb),
	.w7(32'h3b34e69d),
	.w8(32'hbb392571),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5399e),
	.w1(32'hbba53a85),
	.w2(32'hbbd30bdf),
	.w3(32'hbc082270),
	.w4(32'hbb14d2bf),
	.w5(32'hbbe5b81b),
	.w6(32'hbb8deb5a),
	.w7(32'h39fd6fa2),
	.w8(32'hbba016be),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf895),
	.w1(32'h3b6da060),
	.w2(32'h3be04f2c),
	.w3(32'hbc02fac2),
	.w4(32'h3bb2111d),
	.w5(32'h3bba2431),
	.w6(32'hbc07e483),
	.w7(32'h39eef406),
	.w8(32'h39b04494),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b71be),
	.w1(32'hb888070c),
	.w2(32'h39fb12e4),
	.w3(32'hb9b85992),
	.w4(32'hba000dd5),
	.w5(32'h3a113597),
	.w6(32'hb8c01bfc),
	.w7(32'hb9e8d50c),
	.w8(32'h3a15000b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e18e0),
	.w1(32'hba189a42),
	.w2(32'hbb0d6c5b),
	.w3(32'h3b254f5f),
	.w4(32'h3a3e6bf9),
	.w5(32'hbb098b86),
	.w6(32'h393ae875),
	.w7(32'hba23208b),
	.w8(32'hbb63178b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec7d2),
	.w1(32'hbb81a996),
	.w2(32'hbbab2177),
	.w3(32'hbb680e3d),
	.w4(32'hbb940dad),
	.w5(32'hbba151cb),
	.w6(32'hbb4632b9),
	.w7(32'hbb48dbb1),
	.w8(32'hbb826165),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923af34),
	.w1(32'h3abfb5ec),
	.w2(32'hb980e3c6),
	.w3(32'hb945f190),
	.w4(32'h3ad3a4bd),
	.w5(32'hb8c07cb5),
	.w6(32'hba0e6e81),
	.w7(32'h3a3022d9),
	.w8(32'hbb1e23e1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21d8a7),
	.w1(32'h3b3ae9ff),
	.w2(32'hbc33f0bb),
	.w3(32'h3a90dc71),
	.w4(32'hba8f3c19),
	.w5(32'hbc1e6fd2),
	.w6(32'h3abadb47),
	.w7(32'hba403ced),
	.w8(32'hbbb04a93),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c5d385),
	.w1(32'h36aa9491),
	.w2(32'h38a1304d),
	.w3(32'h37d7c90b),
	.w4(32'h37cc5cb3),
	.w5(32'h38c5f881),
	.w6(32'h378f23fb),
	.w7(32'h375446ce),
	.w8(32'h38b7212b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa003c9),
	.w1(32'h382e7ba6),
	.w2(32'hbad67fd9),
	.w3(32'h3ab32772),
	.w4(32'h3a8068b9),
	.w5(32'hbac683ed),
	.w6(32'h3b04290d),
	.w7(32'h39f55649),
	.w8(32'h37e4a302),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9274d3),
	.w1(32'h3b60246a),
	.w2(32'h3a0ad9e7),
	.w3(32'h3c43b9eb),
	.w4(32'h3b8d1236),
	.w5(32'h3ae47efd),
	.w6(32'h3c0b07f6),
	.w7(32'h3b632016),
	.w8(32'hb983ebe2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d0018),
	.w1(32'hbbf96cc6),
	.w2(32'hbc1c2610),
	.w3(32'h3ab74406),
	.w4(32'hbb3adbab),
	.w5(32'hbb8c78e0),
	.w6(32'h3b018759),
	.w7(32'hbabb53fa),
	.w8(32'hbb818f98),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc9046),
	.w1(32'hba086d53),
	.w2(32'hb9c6f764),
	.w3(32'hbad47e69),
	.w4(32'h398a85b4),
	.w5(32'h39ba9d0f),
	.w6(32'hba911936),
	.w7(32'hb7e8eaaa),
	.w8(32'h39e3216a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953798),
	.w1(32'hbabeeafb),
	.w2(32'hb9c97c7f),
	.w3(32'hbb0b30cd),
	.w4(32'h3a16d629),
	.w5(32'h39148110),
	.w6(32'hbb25fbd4),
	.w7(32'h35a1a212),
	.w8(32'h38e6b970),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c3186),
	.w1(32'hba79179b),
	.w2(32'hbae019f7),
	.w3(32'hbadbe1b5),
	.w4(32'h39add7a2),
	.w5(32'hbad519d2),
	.w6(32'h3acc1a12),
	.w7(32'h3ac67277),
	.w8(32'hbab05532),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ff683),
	.w1(32'h3bb2b4a3),
	.w2(32'hbab5e099),
	.w3(32'hba38dc52),
	.w4(32'h3b9ec809),
	.w5(32'h3707a904),
	.w6(32'h3a9f5eb2),
	.w7(32'h3bb66054),
	.w8(32'hb998289a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b1de),
	.w1(32'hbbbfbd0e),
	.w2(32'hbc414ca2),
	.w3(32'hbb8a9700),
	.w4(32'hbb6ef799),
	.w5(32'hbc21ffed),
	.w6(32'hbabd3d27),
	.w7(32'hbb75da6d),
	.w8(32'hbba5306f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b387fbf),
	.w1(32'hba38850a),
	.w2(32'hbc1dce3e),
	.w3(32'h3b52e03d),
	.w4(32'hba20b22f),
	.w5(32'hbc131e8c),
	.w6(32'h3b065b9e),
	.w7(32'hba005a54),
	.w8(32'hbc05dc17),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule