module layer_8_featuremap_155(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2f98f),
	.w1(32'h3b9c46b2),
	.w2(32'hbaca7355),
	.w3(32'hba528074),
	.w4(32'hbb7f6a78),
	.w5(32'h3b04fca8),
	.w6(32'h3ba87b37),
	.w7(32'h39234c0a),
	.w8(32'h3bbe6845),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe233d8),
	.w1(32'hbc02bbd9),
	.w2(32'hbb88c074),
	.w3(32'hbb9dfdf3),
	.w4(32'hbc013531),
	.w5(32'hbb11a29c),
	.w6(32'hbb86ad36),
	.w7(32'hbb8b73a1),
	.w8(32'h3ab799f5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b652),
	.w1(32'hbb868c55),
	.w2(32'hb6b64d6d),
	.w3(32'hbbe72aa7),
	.w4(32'h3b5833fb),
	.w5(32'h3c13ee16),
	.w6(32'hbc148f7d),
	.w7(32'hbb403b69),
	.w8(32'h3c64693e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06f96b),
	.w1(32'h3be9ff72),
	.w2(32'hbba1ac48),
	.w3(32'hbaf1576f),
	.w4(32'hbb9cfb66),
	.w5(32'hbb553768),
	.w6(32'h3ab54458),
	.w7(32'hbbe19fce),
	.w8(32'h3aa7046a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb594a7d),
	.w1(32'hbb2bec6f),
	.w2(32'h3b33a3a9),
	.w3(32'hbc1ee4e0),
	.w4(32'hb9bb87e6),
	.w5(32'h3be08ae3),
	.w6(32'hbc00b718),
	.w7(32'h3bcb40aa),
	.w8(32'h3c4a7ce0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8267c6),
	.w1(32'h3c6518e9),
	.w2(32'hbbd38107),
	.w3(32'h3b517f54),
	.w4(32'h382249a3),
	.w5(32'hbbcfd6fc),
	.w6(32'h3c8d32bf),
	.w7(32'hbb822274),
	.w8(32'hbbf6b691),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90f32),
	.w1(32'h39ee2d6f),
	.w2(32'hbaab3e45),
	.w3(32'hba47da57),
	.w4(32'hbc083c3c),
	.w5(32'hbb7486c9),
	.w6(32'hbb9a4051),
	.w7(32'hba143763),
	.w8(32'h3b22b740),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc71b11),
	.w1(32'hbc351211),
	.w2(32'h3b5dd027),
	.w3(32'hbc854342),
	.w4(32'h3b29d7de),
	.w5(32'h3a86fc00),
	.w6(32'hbc4fad0d),
	.w7(32'h3b2657e1),
	.w8(32'hbbbefdcc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba740ab1),
	.w1(32'hb94e9278),
	.w2(32'hbb8449ab),
	.w3(32'hbbd98b04),
	.w4(32'hbb3f4ea3),
	.w5(32'hba5789f6),
	.w6(32'hbc0ed3de),
	.w7(32'hbb9379dc),
	.w8(32'hbb695999),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb21a),
	.w1(32'hbb87ff9a),
	.w2(32'hbbbeb828),
	.w3(32'hbbff1efa),
	.w4(32'hbc220852),
	.w5(32'hbb12612f),
	.w6(32'hbc43ce03),
	.w7(32'hbbc6bd56),
	.w8(32'hbc391eb2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabdae2),
	.w1(32'hbb375e0a),
	.w2(32'hbbbf748b),
	.w3(32'h3a2b2567),
	.w4(32'hbaa685a7),
	.w5(32'h3ae2804b),
	.w6(32'hbb1c7587),
	.w7(32'hbb616937),
	.w8(32'hbaa66cd1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44fc3d),
	.w1(32'hbc1faf89),
	.w2(32'h381be57a),
	.w3(32'h3b957ff5),
	.w4(32'h3b0a54d3),
	.w5(32'h3bb8b35d),
	.w6(32'hb8b9613c),
	.w7(32'h3a222d6c),
	.w8(32'hbb4cf9a4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a352f),
	.w1(32'hbb6d1453),
	.w2(32'hbb49738d),
	.w3(32'hbc027855),
	.w4(32'hbb32572c),
	.w5(32'hbb3a46c3),
	.w6(32'hbb9f5664),
	.w7(32'hbb5cfba8),
	.w8(32'hbb8ecf98),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85b19d),
	.w1(32'hb977b82b),
	.w2(32'h39252496),
	.w3(32'hba61791d),
	.w4(32'hb9fbf7f9),
	.w5(32'hba059f0b),
	.w6(32'hb966c02b),
	.w7(32'hba2973f7),
	.w8(32'hba2d96c9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b48f1),
	.w1(32'hb91b7cd6),
	.w2(32'hb90edbde),
	.w3(32'hb9297508),
	.w4(32'hb96da252),
	.w5(32'hb9657563),
	.w6(32'hb93b2755),
	.w7(32'hb99aba28),
	.w8(32'hb96c0843),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff1519),
	.w1(32'hba20d503),
	.w2(32'hb8ed3298),
	.w3(32'hba13c029),
	.w4(32'hba85bcbf),
	.w5(32'hba25820e),
	.w6(32'hba216633),
	.w7(32'hba961b3a),
	.w8(32'hba382c95),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14604b),
	.w1(32'h3afd95a3),
	.w2(32'h3ae3c288),
	.w3(32'h3a5eb50f),
	.w4(32'h3aa046dd),
	.w5(32'h3b04abaa),
	.w6(32'h3b002fd7),
	.w7(32'h3a1a5b5e),
	.w8(32'h3a58c9f0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff194e),
	.w1(32'hbb9550d3),
	.w2(32'hbb6ee7e8),
	.w3(32'hbc17a618),
	.w4(32'hbb9ff4ca),
	.w5(32'hbb8db990),
	.w6(32'hbc092e85),
	.w7(32'hbbaadcbd),
	.w8(32'hbb970774),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8fe2a),
	.w1(32'hbb605066),
	.w2(32'hbbed96d0),
	.w3(32'hbc33fbaa),
	.w4(32'hb93c3fe4),
	.w5(32'h3aee054e),
	.w6(32'hbb191b2f),
	.w7(32'h3b46f502),
	.w8(32'h3bdf7368),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f337d),
	.w1(32'hbc261606),
	.w2(32'hbc359985),
	.w3(32'hbbbe6d86),
	.w4(32'hbb91f341),
	.w5(32'hbbc1ab6d),
	.w6(32'hbbdedf1f),
	.w7(32'hbb3c6ce6),
	.w8(32'hbc04761b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2af2),
	.w1(32'hbb1cbeca),
	.w2(32'hbb97be41),
	.w3(32'hb7ad32e5),
	.w4(32'hb9c48c0b),
	.w5(32'hbb7639d3),
	.w6(32'hbb4d3f8d),
	.w7(32'hba998847),
	.w8(32'hbb059784),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ec9a6),
	.w1(32'hbbb3a12c),
	.w2(32'hbbc631e0),
	.w3(32'hbc45714f),
	.w4(32'hbbb69e03),
	.w5(32'hbc0732ab),
	.w6(32'hbc21e51a),
	.w7(32'hbbbae154),
	.w8(32'hbbc9a0f2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba462b36),
	.w1(32'hbb9e9af7),
	.w2(32'h3ab3aa27),
	.w3(32'hbb634f9b),
	.w4(32'hba9a20a8),
	.w5(32'h3c0ff5b9),
	.w6(32'h3c0cac61),
	.w7(32'h3c4234d3),
	.w8(32'h3c951cb6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9531a73),
	.w1(32'hb90fe109),
	.w2(32'hba450372),
	.w3(32'h3a86ad86),
	.w4(32'h3aab66de),
	.w5(32'h390751d6),
	.w6(32'h38cb4908),
	.w7(32'h3ac9561f),
	.w8(32'h39872893),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19e612),
	.w1(32'h3ab62e7f),
	.w2(32'h3a30e3b3),
	.w3(32'h3b67d885),
	.w4(32'h3b3075c1),
	.w5(32'h399dc5ef),
	.w6(32'h3b903b80),
	.w7(32'h3ba1c189),
	.w8(32'h3ad24715),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef757a),
	.w1(32'hbb5a4b1f),
	.w2(32'hbb98282e),
	.w3(32'hbb01115b),
	.w4(32'hba2b3e79),
	.w5(32'hba11423a),
	.w6(32'h3a2baae5),
	.w7(32'h3b4afbfb),
	.w8(32'h3b829d6a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac63f6c),
	.w1(32'h3ad60cd3),
	.w2(32'h3ab03b92),
	.w3(32'h3afc23f3),
	.w4(32'h3ae9ef90),
	.w5(32'h3ac4a69c),
	.w6(32'h3b16638d),
	.w7(32'h3afcf00d),
	.w8(32'h3abdaba1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc4d50),
	.w1(32'hbb53ab67),
	.w2(32'hbc3091b7),
	.w3(32'hbca32d0b),
	.w4(32'h3b186f5f),
	.w5(32'hbc5c3842),
	.w6(32'hbc6a7ae2),
	.w7(32'h3cc92f72),
	.w8(32'h3cba762c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2c8a),
	.w1(32'hbb0b3747),
	.w2(32'hbafdaf04),
	.w3(32'hbb6d08d1),
	.w4(32'hbad2f97b),
	.w5(32'hba04c88d),
	.w6(32'hba901ea3),
	.w7(32'h3a8b012d),
	.w8(32'h3aa26cf6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb240c72),
	.w1(32'hbaa17853),
	.w2(32'hb9a65f8b),
	.w3(32'hbad7b6e9),
	.w4(32'hba08f80e),
	.w5(32'hb9cf10ae),
	.w6(32'hbad88b1f),
	.w7(32'hba48c087),
	.w8(32'hba97ccd4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8acc4),
	.w1(32'h3b294ac9),
	.w2(32'h3a2442bc),
	.w3(32'h39ac60e7),
	.w4(32'h3b3b72f4),
	.w5(32'h3ae4d244),
	.w6(32'h3a3d7011),
	.w7(32'h3adb33cd),
	.w8(32'h3a8d5f95),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec145),
	.w1(32'hba0c34db),
	.w2(32'hbb25ffba),
	.w3(32'h385b0e8e),
	.w4(32'h3a502ac4),
	.w5(32'hbaa00b97),
	.w6(32'hba35d0f5),
	.w7(32'h39d8e1ca),
	.w8(32'hbaa69764),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f48fff),
	.w1(32'hb7532c71),
	.w2(32'hb593f862),
	.w3(32'h38ff09fc),
	.w4(32'h385f01ef),
	.w5(32'h36d4821c),
	.w6(32'h39382ffd),
	.w7(32'h38e4211c),
	.w8(32'h388d3912),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3805caa9),
	.w1(32'hb82d7c17),
	.w2(32'h38179f66),
	.w3(32'h380e246c),
	.w4(32'hb884f28f),
	.w5(32'hb7eac595),
	.w6(32'h3885cfc8),
	.w7(32'hb6ec6b83),
	.w8(32'h38299206),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb589e43),
	.w1(32'hba28682b),
	.w2(32'hbb242522),
	.w3(32'hbb203a2e),
	.w4(32'h394ea885),
	.w5(32'hbb18fcfa),
	.w6(32'hbbacaf8a),
	.w7(32'hbb2dd4be),
	.w8(32'hbb92c152),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf1eca),
	.w1(32'hba26edbd),
	.w2(32'hbb162050),
	.w3(32'hbaab82f2),
	.w4(32'h3984fc89),
	.w5(32'h393aff86),
	.w6(32'hba659bd0),
	.w7(32'h3a75b652),
	.w8(32'h3a8c29fb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9112b54),
	.w1(32'hb947b2fe),
	.w2(32'h3989a1f5),
	.w3(32'hb89e7cb7),
	.w4(32'hb94f49bf),
	.w5(32'h3938059a),
	.w6(32'hb85fb8f7),
	.w7(32'h38c615c6),
	.w8(32'h388db4dc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00cf8e),
	.w1(32'hbbb0dea4),
	.w2(32'hbb59c2fd),
	.w3(32'hbbb65d8c),
	.w4(32'hbb3cf680),
	.w5(32'hbb1b8ede),
	.w6(32'hbb89ddac),
	.w7(32'hbb145ba6),
	.w8(32'hbaf5b5e8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915f999),
	.w1(32'hb8c7524f),
	.w2(32'h37e00bec),
	.w3(32'hb8f3e226),
	.w4(32'hb98d5357),
	.w5(32'hb8ec57e4),
	.w6(32'hb9393c11),
	.w7(32'hb998f763),
	.w8(32'hb98ff031),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc792e),
	.w1(32'h39de9133),
	.w2(32'h39cd6e96),
	.w3(32'h3a041788),
	.w4(32'h396266a7),
	.w5(32'h38135e4f),
	.w6(32'h3a296b5b),
	.w7(32'h39df45a7),
	.w8(32'h39d65c54),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb056ad),
	.w1(32'h38061eed),
	.w2(32'hbb8f7bb2),
	.w3(32'hbbe79a14),
	.w4(32'h3b50d3f5),
	.w5(32'hb9dfac24),
	.w6(32'hbbb07086),
	.w7(32'h3b92a73c),
	.w8(32'h39bafd89),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacae300),
	.w1(32'hba82db1a),
	.w2(32'hb9bf2d2b),
	.w3(32'hbae6e5fa),
	.w4(32'h3935ed7f),
	.w5(32'h39d60b5f),
	.w6(32'hbb2ee21a),
	.w7(32'h3992427f),
	.w8(32'h39fe8e71),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0fee5),
	.w1(32'h3a41bd3a),
	.w2(32'h39afa2a1),
	.w3(32'h39e32c13),
	.w4(32'h3a2776dc),
	.w5(32'h39a6c305),
	.w6(32'h39881b76),
	.w7(32'h3a08df1b),
	.w8(32'h389999bb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aadc28),
	.w1(32'h39202d18),
	.w2(32'hba99dad4),
	.w3(32'hba6c3bcc),
	.w4(32'h3a1cb972),
	.w5(32'hb92a8c1b),
	.w6(32'hb8dd8d6c),
	.w7(32'h3aea2f73),
	.w8(32'h3aed7450),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0ffa),
	.w1(32'hbb30fe0a),
	.w2(32'hba839e2b),
	.w3(32'hbbfd9d9c),
	.w4(32'hbb4e2a71),
	.w5(32'hba8c146e),
	.w6(32'hbb24279a),
	.w7(32'h3b39c0ea),
	.w8(32'h3b93a1ee),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e240),
	.w1(32'hb9caac83),
	.w2(32'hba9fa245),
	.w3(32'hbb14a879),
	.w4(32'h3a1b56ab),
	.w5(32'h3a1dea03),
	.w6(32'hbaec62aa),
	.w7(32'h3a9dca00),
	.w8(32'h3a0b06c6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38108e89),
	.w1(32'hb6c0cf97),
	.w2(32'h37948b5b),
	.w3(32'h373e13ad),
	.w4(32'hb80c4fd7),
	.w5(32'hb6a05b42),
	.w6(32'h37d56ed0),
	.w7(32'hb7c2a205),
	.w8(32'h37077ab7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc264c28),
	.w1(32'hbc162cc4),
	.w2(32'hbbbe3488),
	.w3(32'hbc04a0dd),
	.w4(32'hbbb24270),
	.w5(32'hbb3970f4),
	.w6(32'hbb7d6da2),
	.w7(32'hbada43fd),
	.w8(32'h3a719b26),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bdc8f),
	.w1(32'hb9e49b28),
	.w2(32'hba02e5a5),
	.w3(32'hbb41743a),
	.w4(32'hb9aa64a0),
	.w5(32'hb8b5120d),
	.w6(32'hbb381467),
	.w7(32'hb9898e1a),
	.w8(32'hb99a313f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3279a7),
	.w1(32'hbacdfa38),
	.w2(32'hba198f2a),
	.w3(32'hbb73537c),
	.w4(32'hba32ccf8),
	.w5(32'h3aefc485),
	.w6(32'hb9cab113),
	.w7(32'h3b18b8ae),
	.w8(32'h3b33b19f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3de307),
	.w1(32'hbb8c5301),
	.w2(32'hbb92d1da),
	.w3(32'hbbcc9084),
	.w4(32'hba776d37),
	.w5(32'hbb45e820),
	.w6(32'hbb80af2d),
	.w7(32'hba9135c3),
	.w8(32'hbb563299),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb374d1),
	.w1(32'hbab6dcba),
	.w2(32'hbb9d7503),
	.w3(32'hbc8c4b5c),
	.w4(32'hbc4bd027),
	.w5(32'hbc4b66e3),
	.w6(32'hbc2ff871),
	.w7(32'hbb27828f),
	.w8(32'h3a7128a2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3858),
	.w1(32'hbae9adb8),
	.w2(32'hba97d97e),
	.w3(32'hbb37fa1d),
	.w4(32'hbb527f74),
	.w5(32'hba5c4b76),
	.w6(32'h3ad3344e),
	.w7(32'h3ada504d),
	.w8(32'h3aa48982),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbd4c),
	.w1(32'hbb002b5a),
	.w2(32'hbb0a1ab6),
	.w3(32'hbb9cc05d),
	.w4(32'hbac6aaa5),
	.w5(32'h3ae928ae),
	.w6(32'hbb74e166),
	.w7(32'hbad46c8c),
	.w8(32'hba1d934b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9e981),
	.w1(32'hb784269e),
	.w2(32'h37be9b52),
	.w3(32'h38a56339),
	.w4(32'hb838ad6c),
	.w5(32'hb739bd8c),
	.w6(32'h38eb9546),
	.w7(32'hb7c13bdd),
	.w8(32'h379bf910),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bb69),
	.w1(32'hbbbffefa),
	.w2(32'hbb5c31b7),
	.w3(32'hbc008aa5),
	.w4(32'hbb62ffb0),
	.w5(32'h3b18ed9c),
	.w6(32'hba94dcd4),
	.w7(32'h37a663c9),
	.w8(32'h3b7c6600),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bfafc),
	.w1(32'h39dc40c5),
	.w2(32'h39706a72),
	.w3(32'hba904255),
	.w4(32'h3a2f41eb),
	.w5(32'h3a9ed027),
	.w6(32'hba631d36),
	.w7(32'h3a84970b),
	.w8(32'h39edf271),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0fc4),
	.w1(32'h3b3cb42f),
	.w2(32'h3b36fdb5),
	.w3(32'hbb949aff),
	.w4(32'hba9f6266),
	.w5(32'hb8ff8a50),
	.w6(32'hbb32455e),
	.w7(32'h3b7bd7ad),
	.w8(32'h3b5ca8c0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8392ef),
	.w1(32'h3989cd08),
	.w2(32'h39c32530),
	.w3(32'hba8cfdbb),
	.w4(32'hbac1e75d),
	.w5(32'hba15a2ce),
	.w6(32'h3ab7e25c),
	.w7(32'h3b122f81),
	.w8(32'h3b62216c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc49f),
	.w1(32'h39e95b8c),
	.w2(32'h3818aaa7),
	.w3(32'hba7bcec0),
	.w4(32'hb9ef172f),
	.w5(32'hb9a2750f),
	.w6(32'hba018d6f),
	.w7(32'h3aa0b480),
	.w8(32'h3af35213),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa36601),
	.w1(32'h3aa37505),
	.w2(32'h3aeb3a8c),
	.w3(32'h3ad3b499),
	.w4(32'h3a5a2e70),
	.w5(32'h3a7ed577),
	.w6(32'h3ae18794),
	.w7(32'h3ae44578),
	.w8(32'h3a7a706a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09d7f1),
	.w1(32'hb9dc3ac9),
	.w2(32'hb93190f8),
	.w3(32'hb9bb30d6),
	.w4(32'hb9f1dbab),
	.w5(32'hba06088e),
	.w6(32'hb99722e6),
	.w7(32'hb9c9b03c),
	.w8(32'hb9143871),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf63500),
	.w1(32'hbb1e7104),
	.w2(32'hbbad8ee1),
	.w3(32'hbbcc59b9),
	.w4(32'h391c87f7),
	.w5(32'hba736853),
	.w6(32'hbb523d69),
	.w7(32'h3b3bd7b7),
	.w8(32'hb8be8290),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0a938),
	.w1(32'h391d3b78),
	.w2(32'h3802936a),
	.w3(32'hbac732a0),
	.w4(32'hba108884),
	.w5(32'hba0c1ccc),
	.w6(32'hbb47da5f),
	.w7(32'hbb091851),
	.w8(32'hbab8f5f2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988f004),
	.w1(32'h39194c56),
	.w2(32'h3a51b567),
	.w3(32'h3a0c5017),
	.w4(32'h3a0a548d),
	.w5(32'h3a973492),
	.w6(32'h3abb81d4),
	.w7(32'h3aa98037),
	.w8(32'h3a9d4227),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38beeae0),
	.w1(32'h3a6ef9a7),
	.w2(32'h3a6a0cb6),
	.w3(32'hba05e448),
	.w4(32'h3aa9bf49),
	.w5(32'h3aca16fa),
	.w6(32'h3a812511),
	.w7(32'h3b0c5632),
	.w8(32'h3b20d91a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0fa71),
	.w1(32'hbb783441),
	.w2(32'hbb92ff15),
	.w3(32'hbba0875c),
	.w4(32'hbb28165d),
	.w5(32'hbb79f6e7),
	.w6(32'hbbc3a813),
	.w7(32'hbb659764),
	.w8(32'hbb47cd87),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e80a3),
	.w1(32'h3ac26abc),
	.w2(32'h3a62e071),
	.w3(32'h3b197dc3),
	.w4(32'h3b80a048),
	.w5(32'h3b75652c),
	.w6(32'h3b2b9ac6),
	.w7(32'h3b6003de),
	.w8(32'h3aaa1f11),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88cd08),
	.w1(32'h39d2c03b),
	.w2(32'h3ab69032),
	.w3(32'h3a66a9d3),
	.w4(32'h3a26b7a4),
	.w5(32'h3a92b515),
	.w6(32'h3ab97bdd),
	.w7(32'h3a1911df),
	.w8(32'h3a3802de),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a4727),
	.w1(32'h39cc4ed8),
	.w2(32'hbb8905bb),
	.w3(32'hbb5bcd20),
	.w4(32'hb9da8530),
	.w5(32'hb8a68820),
	.w6(32'hba16f78f),
	.w7(32'h3ba90ff0),
	.w8(32'h3c3184ab),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b97f0),
	.w1(32'h3a125bfb),
	.w2(32'h3975b30c),
	.w3(32'h3a26f398),
	.w4(32'h3a20f35a),
	.w5(32'h39d17343),
	.w6(32'h3a365ec2),
	.w7(32'h3a327876),
	.w8(32'h3a0724c7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb7d6c),
	.w1(32'hbbb5db74),
	.w2(32'hbbb49077),
	.w3(32'hbb911fbe),
	.w4(32'hbb4406ad),
	.w5(32'hbb5126d0),
	.w6(32'hbb48c266),
	.w7(32'hbac393f5),
	.w8(32'hbb15561d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cbb6e),
	.w1(32'h3a7c77f4),
	.w2(32'h3a9cf70e),
	.w3(32'h3a01ee44),
	.w4(32'h3a6517c4),
	.w5(32'h3ab709b4),
	.w6(32'h39975b0c),
	.w7(32'h3a0b3e68),
	.w8(32'h3a2ddf6f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c043),
	.w1(32'hbb53625b),
	.w2(32'hbafcfaae),
	.w3(32'hbb9be4be),
	.w4(32'hb9c91a3d),
	.w5(32'h3a5a264e),
	.w6(32'hbb873e15),
	.w7(32'hb856f3c0),
	.w8(32'h3a670f91),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383bd36a),
	.w1(32'h37500554),
	.w2(32'hb79290e4),
	.w3(32'h37f437a5),
	.w4(32'hb750c03a),
	.w5(32'hb66e3d3b),
	.w6(32'h3810090b),
	.w7(32'h3798c539),
	.w8(32'h37b05be1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b31ee),
	.w1(32'h38bb5577),
	.w2(32'h354e35f0),
	.w3(32'h3abaf4c4),
	.w4(32'h3a8a36fa),
	.w5(32'hb9f804cb),
	.w6(32'h3b341015),
	.w7(32'h3b1178f7),
	.w8(32'h38e7f8f2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a10b4),
	.w1(32'hb998702d),
	.w2(32'h3935a91d),
	.w3(32'hb922228a),
	.w4(32'hbb0397f4),
	.w5(32'hb99c81b1),
	.w6(32'hb88815da),
	.w7(32'h39ee8df8),
	.w8(32'hb9f17753),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62fa77),
	.w1(32'hbb4843aa),
	.w2(32'hbbfef8e0),
	.w3(32'hbb9a040d),
	.w4(32'hbb9a12eb),
	.w5(32'hbbcf4754),
	.w6(32'h3b156039),
	.w7(32'hba5c7263),
	.w8(32'h39d82c66),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fe941),
	.w1(32'hbbc30d31),
	.w2(32'hbbc9847e),
	.w3(32'hbbcad8a4),
	.w4(32'hbbbc60c2),
	.w5(32'hbbd0761c),
	.w6(32'hbb86dea7),
	.w7(32'hbba93441),
	.w8(32'hbb860a0e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db8e8),
	.w1(32'hbbea75a6),
	.w2(32'hbc107b03),
	.w3(32'hbc09c15b),
	.w4(32'hbb961b24),
	.w5(32'h3abc1705),
	.w6(32'hbc044a72),
	.w7(32'h3ad7544f),
	.w8(32'hbc23c44f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880ae0),
	.w1(32'hbbaef0e1),
	.w2(32'h3c0d7a94),
	.w3(32'hbbedb70b),
	.w4(32'hb8bb370a),
	.w5(32'h3baa3ff0),
	.w6(32'hbba3f3a9),
	.w7(32'h3b6b16c8),
	.w8(32'h3b9261e1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dfafd),
	.w1(32'h3c284087),
	.w2(32'hbb27325b),
	.w3(32'h3b335fa4),
	.w4(32'hbb738598),
	.w5(32'hbc862b2c),
	.w6(32'h3b417028),
	.w7(32'hbc660c9f),
	.w8(32'h3bc17c94),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2930c9),
	.w1(32'hbc0782a4),
	.w2(32'hbc5639ae),
	.w3(32'hbc11eb19),
	.w4(32'hbc7f7981),
	.w5(32'hbc7f8c13),
	.w6(32'hbbd43eb8),
	.w7(32'hba9024eb),
	.w8(32'hbc41c345),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ae48c),
	.w1(32'hbbd06e65),
	.w2(32'hbc6abab7),
	.w3(32'hbcaf48d0),
	.w4(32'h3ae027e3),
	.w5(32'h398dee81),
	.w6(32'hbcafaabd),
	.w7(32'h3bd4f1a2),
	.w8(32'hbbdcbc2b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3feb76),
	.w1(32'hbc0bf114),
	.w2(32'hbc575fa4),
	.w3(32'hb9f562f5),
	.w4(32'hbbade157),
	.w5(32'h3ada7b3d),
	.w6(32'hbb51bb28),
	.w7(32'h3c9592f0),
	.w8(32'hbc32eb23),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2259dc),
	.w1(32'hbbd32a92),
	.w2(32'h3bc110c7),
	.w3(32'hbc77bdc1),
	.w4(32'hba61d914),
	.w5(32'h3b5669c6),
	.w6(32'h3b97600d),
	.w7(32'h3c23f9a8),
	.w8(32'h3b4af1a1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae75566),
	.w1(32'h3b92c56d),
	.w2(32'hbc370ce8),
	.w3(32'hb9b838c1),
	.w4(32'hbb8237c5),
	.w5(32'hbb308a53),
	.w6(32'hbbad23ed),
	.w7(32'hbb10babd),
	.w8(32'hbb1c405d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc00ba),
	.w1(32'hbb83d846),
	.w2(32'hbc02a1f9),
	.w3(32'hbaeb28e1),
	.w4(32'hbc12e4ac),
	.w5(32'hbc17c1ff),
	.w6(32'h3b222665),
	.w7(32'hbc18e4e2),
	.w8(32'hbc1c681c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0771fe),
	.w1(32'h3a8eb19f),
	.w2(32'hbc5388f9),
	.w3(32'h3b302bb6),
	.w4(32'hbbe1251b),
	.w5(32'hbc2a412a),
	.w6(32'h3a941289),
	.w7(32'hbc130c98),
	.w8(32'hbc380cbd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf91fcb),
	.w1(32'hbbb54487),
	.w2(32'hbc6360e4),
	.w3(32'hbc5a870d),
	.w4(32'hbb0f79c2),
	.w5(32'h3c3d99d7),
	.w6(32'hbb92806d),
	.w7(32'h3cce7625),
	.w8(32'hbd542271),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44ffa6),
	.w1(32'hbc5d1143),
	.w2(32'h3c0b8292),
	.w3(32'hbbffd933),
	.w4(32'hbaf1b05c),
	.w5(32'hbc011090),
	.w6(32'h3c0f5143),
	.w7(32'hbb8c94d2),
	.w8(32'h3c385cc1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abb4d1),
	.w1(32'hbb9a57c7),
	.w2(32'h3ad4dc99),
	.w3(32'h3bdea471),
	.w4(32'h3a3e96cb),
	.w5(32'h3bd9f7f9),
	.w6(32'hbc3fff79),
	.w7(32'h3b94756e),
	.w8(32'hbc1c1b6a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238c63),
	.w1(32'hbac4600f),
	.w2(32'hbbf5fbf3),
	.w3(32'hbc0918d4),
	.w4(32'h38502a6c),
	.w5(32'hba4301f9),
	.w6(32'hbc12dc93),
	.w7(32'h3c30cca3),
	.w8(32'hbc04ff2c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64c56b),
	.w1(32'hbbd52c15),
	.w2(32'hbc24dc7e),
	.w3(32'hbc2321e8),
	.w4(32'hbbbb67b4),
	.w5(32'hbb813d04),
	.w6(32'hbc3c3831),
	.w7(32'hba25b02b),
	.w8(32'hbbda8789),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbab2e),
	.w1(32'h3a3463e7),
	.w2(32'hbbf3cefe),
	.w3(32'h3b5d2d5b),
	.w4(32'hbbb38140),
	.w5(32'hbba1a547),
	.w6(32'hbc458a8c),
	.w7(32'hbbbc6c93),
	.w8(32'hbba8b09f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5aab),
	.w1(32'hbb3eef3d),
	.w2(32'hbbf56dd4),
	.w3(32'hbb3bc037),
	.w4(32'hb9dd0504),
	.w5(32'hbb31574e),
	.w6(32'hbb4b54a9),
	.w7(32'h3c0e8372),
	.w8(32'hbbe6c637),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f18f),
	.w1(32'hbcd84a5e),
	.w2(32'hbc01dd2e),
	.w3(32'hbcc67fa3),
	.w4(32'hbb950a99),
	.w5(32'hbb532bd6),
	.w6(32'hbbc9c0aa),
	.w7(32'h3bbdc751),
	.w8(32'hbc734a34),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936395),
	.w1(32'h3b5ad7a5),
	.w2(32'h3aa5fa58),
	.w3(32'h3b9c9103),
	.w4(32'hbb21fbf6),
	.w5(32'h3b50b9bb),
	.w6(32'hbbf7838d),
	.w7(32'h3c029ee6),
	.w8(32'hbc03b9bb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cb812),
	.w1(32'hbbc36508),
	.w2(32'hbb06d1da),
	.w3(32'hbaf828cf),
	.w4(32'hbabaa933),
	.w5(32'hba293ae4),
	.w6(32'h3c968752),
	.w7(32'hbb93dfa9),
	.w8(32'hbc28f4ec),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820e8f),
	.w1(32'hbb7c41ba),
	.w2(32'h3b4f947f),
	.w3(32'hbbf6136c),
	.w4(32'h3b54b637),
	.w5(32'h3bb173b6),
	.w6(32'hbc5ca302),
	.w7(32'h3a8d125c),
	.w8(32'hbb284192),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53f1c7),
	.w1(32'h3bade0e1),
	.w2(32'h3be3fe3b),
	.w3(32'hbb982b40),
	.w4(32'h3bf7b1e4),
	.w5(32'h3c1364fb),
	.w6(32'hbad40aaf),
	.w7(32'h3c220cc6),
	.w8(32'h3a8e7549),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e837),
	.w1(32'hb899a144),
	.w2(32'hbbffb846),
	.w3(32'hbaad48ac),
	.w4(32'hbae85240),
	.w5(32'hbb9d2294),
	.w6(32'hba283de4),
	.w7(32'hba55457c),
	.w8(32'hbc126745),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a564b13),
	.w1(32'h3ba7fd22),
	.w2(32'hbb8ee649),
	.w3(32'hbacd24a5),
	.w4(32'hbc339af9),
	.w5(32'hbc1216f8),
	.w6(32'h3b20753d),
	.w7(32'h3beb3472),
	.w8(32'hbc1b2dc3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93c4db),
	.w1(32'hbbc8bb72),
	.w2(32'hbbb47ddd),
	.w3(32'hbc008f7e),
	.w4(32'hbbaf0811),
	.w5(32'hbbd06b47),
	.w6(32'hbc5c665a),
	.w7(32'hbb4b64c7),
	.w8(32'hbb06bcc7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb742e01),
	.w1(32'h3a3ead23),
	.w2(32'hbc4da744),
	.w3(32'hbbed7044),
	.w4(32'hbb9f2f28),
	.w5(32'h38bc00ad),
	.w6(32'hbc04514e),
	.w7(32'h3ab3be62),
	.w8(32'hbc97f835),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f40a7),
	.w1(32'hbc7c5c05),
	.w2(32'h3816f40e),
	.w3(32'hbc664383),
	.w4(32'hba4a19f4),
	.w5(32'h3c92748b),
	.w6(32'h3c0b8cbf),
	.w7(32'h3bfacf0e),
	.w8(32'hbb259c49),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca974a),
	.w1(32'hbbe207c8),
	.w2(32'h3be96773),
	.w3(32'hbbaf1906),
	.w4(32'h3c846cde),
	.w5(32'hbc9b31ff),
	.w6(32'h3bbc51bb),
	.w7(32'hbcccbb27),
	.w8(32'h3c9aa0c0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd29c6a5),
	.w1(32'h3ce717c4),
	.w2(32'hbb93527e),
	.w3(32'h3c1408ee),
	.w4(32'hbad0f88f),
	.w5(32'hbb0d0a05),
	.w6(32'hbd265243),
	.w7(32'hbafe1cc6),
	.w8(32'hbb504537),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62b06c),
	.w1(32'h3abf6656),
	.w2(32'h3b652951),
	.w3(32'h38f11247),
	.w4(32'h3b7c3863),
	.w5(32'h3bb6e9d9),
	.w6(32'h3b03b7d9),
	.w7(32'h3b197936),
	.w8(32'h3b7786b2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba383c23),
	.w1(32'hbb8d7ad5),
	.w2(32'h3c0b6280),
	.w3(32'hbb62486f),
	.w4(32'h3be894f4),
	.w5(32'hbc8fbdd7),
	.w6(32'hbbe3daeb),
	.w7(32'hbcfedb9c),
	.w8(32'h3c6be8d4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd19e88),
	.w1(32'h3c921953),
	.w2(32'hbc1cc9ad),
	.w3(32'h3c21c70e),
	.w4(32'h3b6fd336),
	.w5(32'hbad8d824),
	.w6(32'hbce862ad),
	.w7(32'hbbbc5b0e),
	.w8(32'hbc80c847),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b0f63),
	.w1(32'hbb83d84a),
	.w2(32'h3acc1d86),
	.w3(32'hbc511869),
	.w4(32'hb9ea62c7),
	.w5(32'h3c14e72b),
	.w6(32'hbc8971e9),
	.w7(32'h3bf9099b),
	.w8(32'hbc2b5c95),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78d88c),
	.w1(32'h3b7c59dd),
	.w2(32'hba266c2f),
	.w3(32'hbb2ca973),
	.w4(32'hbbae5379),
	.w5(32'hbcb8df92),
	.w6(32'hbbc0d6b0),
	.w7(32'hbced8ebe),
	.w8(32'h3b48b7c0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106523),
	.w1(32'hbc59e933),
	.w2(32'h3b8b82c8),
	.w3(32'hbbb68e5e),
	.w4(32'hb9f1821d),
	.w5(32'hbbe7a270),
	.w6(32'hbc7babe6),
	.w7(32'h3b68fde5),
	.w8(32'h3b8b3409),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21129d),
	.w1(32'hbc59372e),
	.w2(32'hbbd31ea8),
	.w3(32'hbb0614da),
	.w4(32'h3a87f20e),
	.w5(32'h3bbd4593),
	.w6(32'h38d10f3f),
	.w7(32'h3b339934),
	.w8(32'hbc6b1d49),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d8c3),
	.w1(32'h3b55d92f),
	.w2(32'h3b3e2891),
	.w3(32'h3a485dfd),
	.w4(32'h3b027b75),
	.w5(32'h3b41cf32),
	.w6(32'h3bb45c18),
	.w7(32'h3ad7cbae),
	.w8(32'hbb602e9e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bc8a),
	.w1(32'h3b4e7883),
	.w2(32'hbabd278b),
	.w3(32'hbb8e3383),
	.w4(32'h3be21046),
	.w5(32'h3be04080),
	.w6(32'hbc0930f0),
	.w7(32'h3c3b89e3),
	.w8(32'hbbbec230),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ad5ed),
	.w1(32'hb91325c4),
	.w2(32'h38cb20a2),
	.w3(32'hbbe5cbbc),
	.w4(32'h3a680478),
	.w5(32'h3a8b98f0),
	.w6(32'h3c84ad1a),
	.w7(32'h3b2c4ee1),
	.w8(32'h3b86d7ae),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b327b9d),
	.w1(32'h3a3bf12f),
	.w2(32'hbbfdc763),
	.w3(32'h3a88b605),
	.w4(32'hbc000b10),
	.w5(32'hbcad61e5),
	.w6(32'h3b324056),
	.w7(32'hbc7dfc62),
	.w8(32'hbca0a1f0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46ce93),
	.w1(32'hbc3cca58),
	.w2(32'hbb503714),
	.w3(32'hbc9a2223),
	.w4(32'hbc210970),
	.w5(32'hbbfefbb2),
	.w6(32'hbcad560c),
	.w7(32'hbb871789),
	.w8(32'hbc38ddc5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87395f),
	.w1(32'hbc0bedda),
	.w2(32'hbb9bd0c4),
	.w3(32'hbc618d5a),
	.w4(32'hbc0c8204),
	.w5(32'hbb8b5d31),
	.w6(32'hbc7d992d),
	.w7(32'hbbce4d8f),
	.w8(32'hba86e8ee),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b7469),
	.w1(32'hbb9257b1),
	.w2(32'hbb0cde63),
	.w3(32'hbb9302c6),
	.w4(32'h3c4819cd),
	.w5(32'h3c006897),
	.w6(32'hbc3835db),
	.w7(32'h3c10a03f),
	.w8(32'h3b1147a5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a54a),
	.w1(32'h3c7253de),
	.w2(32'h3abc49b4),
	.w3(32'h3b6e8573),
	.w4(32'h3abaf391),
	.w5(32'h3b79a127),
	.w6(32'h3a8f25e4),
	.w7(32'h3b0af74c),
	.w8(32'h3b48a8ef),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c35f6),
	.w1(32'h3bacc685),
	.w2(32'h3c31a8de),
	.w3(32'h3b86e051),
	.w4(32'h3bcca16d),
	.w5(32'hbb8ac845),
	.w6(32'h3b6ced13),
	.w7(32'h3b88dcc4),
	.w8(32'hbc95534c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c157d),
	.w1(32'hbc19f529),
	.w2(32'h3bfbe749),
	.w3(32'hbbe88233),
	.w4(32'hbb1f5176),
	.w5(32'hbb66a4ae),
	.w6(32'h3c3841ec),
	.w7(32'hbc0dbd35),
	.w8(32'h3b946729),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4ca2),
	.w1(32'hbb8b7079),
	.w2(32'hbbd4447f),
	.w3(32'hbc82ca83),
	.w4(32'hbc159c6b),
	.w5(32'hbbc9aa97),
	.w6(32'hbb848cc1),
	.w7(32'hbbfe195f),
	.w8(32'hbc105871),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3132e),
	.w1(32'hbb90e2d7),
	.w2(32'hbc38f5ef),
	.w3(32'hbbb847fd),
	.w4(32'hbbcc4b86),
	.w5(32'hbc2bd617),
	.w6(32'hbbd928a8),
	.w7(32'h39b584ea),
	.w8(32'hbc50d0a0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2808b1),
	.w1(32'hbc3d1306),
	.w2(32'h39571d94),
	.w3(32'hbc629ae3),
	.w4(32'hbb6acf8f),
	.w5(32'hbb5da4f5),
	.w6(32'hbc1d5073),
	.w7(32'h3a26328e),
	.w8(32'hbb94dd70),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule