module layer_10_featuremap_43(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71cc8a),
	.w1(32'hbb588fdc),
	.w2(32'hbc160c77),
	.w3(32'h3bf0ec82),
	.w4(32'h3ae0c5b4),
	.w5(32'hbbbce199),
	.w6(32'h3b874c15),
	.w7(32'h3b91b2ba),
	.w8(32'h3bbcc9ea),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d694),
	.w1(32'h3bccd2a4),
	.w2(32'h3a2702fc),
	.w3(32'hbb3e27de),
	.w4(32'hbb62be52),
	.w5(32'h3c20c324),
	.w6(32'hb9a8e224),
	.w7(32'hbbe0211e),
	.w8(32'h3c054f2f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8b90),
	.w1(32'h3b2bf827),
	.w2(32'hbae30d53),
	.w3(32'h3c52c157),
	.w4(32'h3ac78cdd),
	.w5(32'h3a93e259),
	.w6(32'h3c22d552),
	.w7(32'h3b976efb),
	.w8(32'h3aca7c4e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fcb8e),
	.w1(32'h3c592006),
	.w2(32'h3b84073e),
	.w3(32'h3bd403a4),
	.w4(32'h3bcc6e10),
	.w5(32'h3becc945),
	.w6(32'h3b38b838),
	.w7(32'h3be12681),
	.w8(32'h3bfc0010),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadcec0),
	.w1(32'h3a9a8fd2),
	.w2(32'h3c18c0d3),
	.w3(32'h3c2a18f4),
	.w4(32'h3c3b71e4),
	.w5(32'h3c09b089),
	.w6(32'h3c353461),
	.w7(32'h3bdec966),
	.w8(32'h3ba1557a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49f6af),
	.w1(32'h3b9db381),
	.w2(32'h3abc8f88),
	.w3(32'h3bbfeae1),
	.w4(32'h3c096c4b),
	.w5(32'h3bb83062),
	.w6(32'h3bf69496),
	.w7(32'h3c085ae2),
	.w8(32'h3b55c8a6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97700a),
	.w1(32'hbb5c65e0),
	.w2(32'h3ca36592),
	.w3(32'h3b1f4985),
	.w4(32'h3bba7e28),
	.w5(32'h3c1f54ce),
	.w6(32'h3a81df3a),
	.w7(32'h3ba3a072),
	.w8(32'hbc2db724),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05ba57),
	.w1(32'h3ca2204d),
	.w2(32'hbcb6810e),
	.w3(32'h3ca49463),
	.w4(32'h3c5a3564),
	.w5(32'hbd0245a3),
	.w6(32'h3b4c7757),
	.w7(32'hba983ccb),
	.w8(32'hbcceea10),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ce721),
	.w1(32'hbc8ff2da),
	.w2(32'h3a5b6cca),
	.w3(32'hbd3ed5c4),
	.w4(32'hbce43e3c),
	.w5(32'h3beaea07),
	.w6(32'hbd1ec5da),
	.w7(32'hbcd26c40),
	.w8(32'h3bdc12ea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f652c),
	.w1(32'hba3e7b9d),
	.w2(32'hbb65b220),
	.w3(32'h3bbc2f61),
	.w4(32'h3b6abf17),
	.w5(32'h3c019347),
	.w6(32'h3bcff9cf),
	.w7(32'h3c07d87e),
	.w8(32'h3c62a8d5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1e8b),
	.w1(32'hbbe4ced5),
	.w2(32'hb95d71c1),
	.w3(32'h3babb7d7),
	.w4(32'h3b811f76),
	.w5(32'hba37b797),
	.w6(32'h3c5962f6),
	.w7(32'h3c467631),
	.w8(32'h3b982caa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eae24),
	.w1(32'h3ba39494),
	.w2(32'hbc04c810),
	.w3(32'h3b94f65c),
	.w4(32'hbb86b34d),
	.w5(32'hbbccdb4d),
	.w6(32'h3c27ad41),
	.w7(32'hb952b5cb),
	.w8(32'hbb875acb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc683745),
	.w1(32'hbc3598c7),
	.w2(32'hbc1247e3),
	.w3(32'hbbb7121f),
	.w4(32'hbbca1c0b),
	.w5(32'h3bb23518),
	.w6(32'hb94091dc),
	.w7(32'h39c4bf0f),
	.w8(32'hbb3881d9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b4bb5),
	.w1(32'hbc508fd9),
	.w2(32'hbaa99ead),
	.w3(32'hbbf22975),
	.w4(32'hbb4e8cdd),
	.w5(32'hbc2a56d5),
	.w6(32'hbc22a291),
	.w7(32'hbb8d85c5),
	.w8(32'hbc55218a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88cc02),
	.w1(32'hb9071bb8),
	.w2(32'h3cb0c154),
	.w3(32'hbc892178),
	.w4(32'hbbf23ff3),
	.w5(32'h3cbca742),
	.w6(32'hbcb6d268),
	.w7(32'hbc92b522),
	.w8(32'h3c02f114),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d052f9b),
	.w1(32'h3c69e8aa),
	.w2(32'hbbcb8baf),
	.w3(32'h3d25ef26),
	.w4(32'h3ccd2f46),
	.w5(32'h3b532956),
	.w6(32'h3cea4550),
	.w7(32'h3ce9cc65),
	.w8(32'h3c1655b2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122620),
	.w1(32'hbbd914a6),
	.w2(32'hbbf1434f),
	.w3(32'h3b1c0861),
	.w4(32'h3ac749c2),
	.w5(32'hbbef0660),
	.w6(32'h3c2d7a5f),
	.w7(32'h3c1710f2),
	.w8(32'hbbd9775d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81438f),
	.w1(32'hbab2f616),
	.w2(32'hbb482563),
	.w3(32'hbc1d1663),
	.w4(32'hbbab6298),
	.w5(32'hbb2fddac),
	.w6(32'hbc41e446),
	.w7(32'hbbed832c),
	.w8(32'hbb98346f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9419ea),
	.w1(32'hbbcb8980),
	.w2(32'hbb062640),
	.w3(32'hbc1b21bf),
	.w4(32'hbb2d2ba0),
	.w5(32'hbb785fe1),
	.w6(32'h3b001485),
	.w7(32'hbb64bb3d),
	.w8(32'h3a8ab2c9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5d60),
	.w1(32'hbb867758),
	.w2(32'h3b842a09),
	.w3(32'hbb5df0cb),
	.w4(32'h398fb954),
	.w5(32'h39e28efd),
	.w6(32'hbb8f8090),
	.w7(32'hbb8feb1c),
	.w8(32'hbbb8fe5b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9cf2),
	.w1(32'hbbce1fcc),
	.w2(32'h3a139bea),
	.w3(32'hbc211d5e),
	.w4(32'h3ad5d4e7),
	.w5(32'h3b8ff924),
	.w6(32'hbbd5ceab),
	.w7(32'h3b4de87c),
	.w8(32'hbb3c11ad),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab068),
	.w1(32'h3a9e21c5),
	.w2(32'h3bb6c5f4),
	.w3(32'h3b18d566),
	.w4(32'h3b040803),
	.w5(32'h3b059c3e),
	.w6(32'h38dc6c67),
	.w7(32'h3a441855),
	.w8(32'hbb94d485),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac4371),
	.w1(32'h3b937f60),
	.w2(32'h3bf320f6),
	.w3(32'hbab39f81),
	.w4(32'h3b3aa112),
	.w5(32'h3b331909),
	.w6(32'hbbe9f9a3),
	.w7(32'hb7c9eb56),
	.w8(32'hbab57bd9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91c6c9),
	.w1(32'h3c267894),
	.w2(32'hbb2322db),
	.w3(32'h3a867f51),
	.w4(32'h3b94257c),
	.w5(32'h3bb25ce4),
	.w6(32'hbc0b0538),
	.w7(32'hbb47e336),
	.w8(32'hbb0ea113),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122600),
	.w1(32'hbc0ead59),
	.w2(32'h3a10caad),
	.w3(32'hbb349c5b),
	.w4(32'hb9992a60),
	.w5(32'hbc5fbc10),
	.w6(32'hbb07ca27),
	.w7(32'hbb6a84ae),
	.w8(32'hbbbab45e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed2ee0),
	.w1(32'h3a5481a9),
	.w2(32'hba4c4b52),
	.w3(32'hbc74eb94),
	.w4(32'hbb158aa5),
	.w5(32'hbb0006a2),
	.w6(32'hbca84bcf),
	.w7(32'hbbbcb5c1),
	.w8(32'h3bcccd0e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98035ee),
	.w1(32'hbab7ecce),
	.w2(32'h3ac76d3b),
	.w3(32'h3bfacc8d),
	.w4(32'h3b6c21ae),
	.w5(32'h3a00de49),
	.w6(32'h3bee98cf),
	.w7(32'h399d06c6),
	.w8(32'h39ed9459),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aea47),
	.w1(32'h39ab60e0),
	.w2(32'h3a80380f),
	.w3(32'h3b63052a),
	.w4(32'h3ac90494),
	.w5(32'h3ba603f7),
	.w6(32'h38bd9d35),
	.w7(32'h3acb74b2),
	.w8(32'hbbe792d5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c69dc),
	.w1(32'h3c0c97a5),
	.w2(32'hbb586f3a),
	.w3(32'hb982a576),
	.w4(32'hbb33c67c),
	.w5(32'hbc3c710d),
	.w6(32'h3ae37d87),
	.w7(32'h3bc338c9),
	.w8(32'hbbccbfc8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb16696),
	.w1(32'hbc097582),
	.w2(32'h3b21531b),
	.w3(32'hbbeccfe6),
	.w4(32'h3bed8fcf),
	.w5(32'h3a76df77),
	.w6(32'hbbea0d01),
	.w7(32'hbc17e1a4),
	.w8(32'hba8849c1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7036e8),
	.w1(32'hbab31a01),
	.w2(32'h3bb88278),
	.w3(32'hb9c3b392),
	.w4(32'hbaecc711),
	.w5(32'hbc99125e),
	.w6(32'hbb66f6ba),
	.w7(32'h3a7eea12),
	.w8(32'hbb82273c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca2234),
	.w1(32'hbc23e549),
	.w2(32'hbadf2f39),
	.w3(32'hba919c74),
	.w4(32'hbbdc2fa5),
	.w5(32'hbb7c712f),
	.w6(32'hbc2c1f6a),
	.w7(32'hbb90ee27),
	.w8(32'hbbcb25e2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fde7eb),
	.w1(32'hbbf0e591),
	.w2(32'h3a039366),
	.w3(32'hbbdf45b0),
	.w4(32'hbb24994f),
	.w5(32'hbb273919),
	.w6(32'hbbc7ee90),
	.w7(32'hbc0fc55e),
	.w8(32'hba1b0603),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dfe2d),
	.w1(32'hbaa2bdb2),
	.w2(32'h3c47d450),
	.w3(32'hbb433a8f),
	.w4(32'h3b2a672f),
	.w5(32'hbc625da1),
	.w6(32'hba8bac0f),
	.w7(32'h3addac82),
	.w8(32'h3bcca994),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf786ad),
	.w1(32'hbc0f6ce4),
	.w2(32'hbb91684f),
	.w3(32'hbc992628),
	.w4(32'h3c8cf150),
	.w5(32'hbb0ac766),
	.w6(32'h3cd3aeca),
	.w7(32'hbc13a0d1),
	.w8(32'hbb4900d6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d98a),
	.w1(32'hb8ea859a),
	.w2(32'h3c99dc3e),
	.w3(32'hbba08c0b),
	.w4(32'hbb4667fa),
	.w5(32'hbc9f0002),
	.w6(32'hbb62d9f0),
	.w7(32'hbbf37a0d),
	.w8(32'h3bd04d50),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5cf1),
	.w1(32'hbcde09fe),
	.w2(32'h3a92bbd1),
	.w3(32'hbc98fb31),
	.w4(32'h3d55de1c),
	.w5(32'h3b43c940),
	.w6(32'h3d509b92),
	.w7(32'hbba5a588),
	.w8(32'h39adccb1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbef137),
	.w1(32'hba069ebd),
	.w2(32'hbc19a821),
	.w3(32'hb7b8b998),
	.w4(32'h3b27c0a4),
	.w5(32'h3c96caa4),
	.w6(32'hbae2b76c),
	.w7(32'h3981a002),
	.w8(32'hbbc28f73),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1b9fb),
	.w1(32'h3c93ee9b),
	.w2(32'hbc06212c),
	.w3(32'h3c292fe4),
	.w4(32'hbc69a97f),
	.w5(32'hbc04c3f1),
	.w6(32'hbc7c9be3),
	.w7(32'hbac70034),
	.w8(32'h3a033342),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a0a31),
	.w1(32'h3acb2ba4),
	.w2(32'hbb8f40d1),
	.w3(32'h3aea5933),
	.w4(32'h3b489f4b),
	.w5(32'hba15c035),
	.w6(32'hbc670efc),
	.w7(32'h3baedd1c),
	.w8(32'hbbb36dc8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ea1b),
	.w1(32'hba92d142),
	.w2(32'h3bb83678),
	.w3(32'hbbdcc6d3),
	.w4(32'hbbfef0c1),
	.w5(32'h3c501028),
	.w6(32'hbb780379),
	.w7(32'h382077b1),
	.w8(32'hbaad8322),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1813db),
	.w1(32'h3b46c864),
	.w2(32'h3b4d5d72),
	.w3(32'hbbb61afa),
	.w4(32'hbbc7a6c6),
	.w5(32'h3b135a93),
	.w6(32'h3b894279),
	.w7(32'h3c338aac),
	.w8(32'hbb3b2133),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397c56),
	.w1(32'h3b4e4687),
	.w2(32'hb683551b),
	.w3(32'hbbdef2bc),
	.w4(32'hbb03159e),
	.w5(32'h3b29874f),
	.w6(32'hb9e339bf),
	.w7(32'h3c0a2812),
	.w8(32'h38ee4bbe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6423f),
	.w1(32'h3a9ed44c),
	.w2(32'hbbdab9c3),
	.w3(32'h3a9c60c5),
	.w4(32'h38aa5db3),
	.w5(32'hbc0f3cd2),
	.w6(32'h3aa9e484),
	.w7(32'hbb6da569),
	.w8(32'h3b448f77),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dac4f),
	.w1(32'h3bd0e921),
	.w2(32'hbbf1309c),
	.w3(32'h3b9b7770),
	.w4(32'h3993555e),
	.w5(32'h3d22c425),
	.w6(32'hba960904),
	.w7(32'hbbf00483),
	.w8(32'h3bf9f19d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce71541),
	.w1(32'h3cc57e39),
	.w2(32'h3bd5b006),
	.w3(32'h3d01309e),
	.w4(32'hbb8dac35),
	.w5(32'h3c22132c),
	.w6(32'h3c71ed9a),
	.w7(32'h3ce963da),
	.w8(32'h3b86110d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36b293),
	.w1(32'h3beda77c),
	.w2(32'h3bbc1ae6),
	.w3(32'h3bf47daf),
	.w4(32'h3b25f332),
	.w5(32'hbb67b6e2),
	.w6(32'h3be2d2e6),
	.w7(32'h3c97b4ff),
	.w8(32'hbba9a048),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fe581),
	.w1(32'hbb2ae911),
	.w2(32'hbb406214),
	.w3(32'hbbfefe3e),
	.w4(32'h3998e9a6),
	.w5(32'hb8158e71),
	.w6(32'h3c52614b),
	.w7(32'hbbd2371d),
	.w8(32'hbb691611),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abff573),
	.w1(32'hbabcc01e),
	.w2(32'hbb37135c),
	.w3(32'hba9c3407),
	.w4(32'hbbac271f),
	.w5(32'hbc1be401),
	.w6(32'h399215dc),
	.w7(32'hbb640d7b),
	.w8(32'hbc14c68d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a0df0),
	.w1(32'hba8e3154),
	.w2(32'hbbdde7c3),
	.w3(32'hba236af4),
	.w4(32'hbbde3b6a),
	.w5(32'hbc850f51),
	.w6(32'hbc9992e6),
	.w7(32'hbae8ce1e),
	.w8(32'h3c89af60),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2943e),
	.w1(32'h3cb33de0),
	.w2(32'hbc116ac5),
	.w3(32'h3bd90fce),
	.w4(32'h3ab03575),
	.w5(32'hb855d514),
	.w6(32'h3bdf0d5c),
	.w7(32'hbc8f5923),
	.w8(32'h3bdaed9c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d11ab),
	.w1(32'h3ced3034),
	.w2(32'hbbf5a761),
	.w3(32'h3cc90b24),
	.w4(32'hbcb6abf8),
	.w5(32'hbc9c6c57),
	.w6(32'hbcbeab42),
	.w7(32'hbb53f65e),
	.w8(32'h3c0cc597),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a1b14),
	.w1(32'h3c516ea8),
	.w2(32'h3b074f18),
	.w3(32'h3b50e16c),
	.w4(32'h3b2cf27d),
	.w5(32'hbb344877),
	.w6(32'h3b0d8e46),
	.w7(32'hbb9c2197),
	.w8(32'h3b7aefa0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc217898),
	.w1(32'h3b20d0a6),
	.w2(32'hbc6765dd),
	.w3(32'h3c1e5333),
	.w4(32'hbadcae3d),
	.w5(32'h3bddf403),
	.w6(32'hbc144ea0),
	.w7(32'hbc06f970),
	.w8(32'h3c66ad83),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc462410),
	.w1(32'h3c0ee101),
	.w2(32'h3cb6572c),
	.w3(32'h3c8e43ae),
	.w4(32'hbc5e9ce0),
	.w5(32'h3bd5a2da),
	.w6(32'hbc83cf52),
	.w7(32'hbc16f55e),
	.w8(32'h3bc89bbd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f0504),
	.w1(32'hbc73e8b2),
	.w2(32'h3b424f25),
	.w3(32'hbc8305fd),
	.w4(32'h3d15f74c),
	.w5(32'h3b397115),
	.w6(32'h3ca67a5c),
	.w7(32'hbc1fb3b6),
	.w8(32'hbbb97f7c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23652d),
	.w1(32'hba4d84a0),
	.w2(32'h3b789488),
	.w3(32'hbc5c29c4),
	.w4(32'h3b959b71),
	.w5(32'h3b2686a2),
	.w6(32'h393adb4f),
	.w7(32'hbaabc984),
	.w8(32'h3b6c277f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e51f),
	.w1(32'h39009dba),
	.w2(32'hbb082b25),
	.w3(32'h3b150614),
	.w4(32'hb9f8f143),
	.w5(32'hbbbdcfbc),
	.w6(32'h39b66333),
	.w7(32'hbb608dc7),
	.w8(32'hbb2f6af0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe871a2),
	.w1(32'h3b1daba1),
	.w2(32'h3bdbbfd2),
	.w3(32'hbab1cae2),
	.w4(32'h3bf41b1e),
	.w5(32'hbb95e310),
	.w6(32'h3a82756c),
	.w7(32'h3b7dabb5),
	.w8(32'h3b7d5e7b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96b995),
	.w1(32'h3a96b5a8),
	.w2(32'hbb2f9618),
	.w3(32'h3b8fec3e),
	.w4(32'h3ab2f0ad),
	.w5(32'h3b574a73),
	.w6(32'h3a278220),
	.w7(32'hb6427252),
	.w8(32'hbc4bc775),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37045fc8),
	.w1(32'h3c071013),
	.w2(32'hbb459b20),
	.w3(32'hb87be1c7),
	.w4(32'hbc2a01db),
	.w5(32'h3bb447dc),
	.w6(32'hbbab4890),
	.w7(32'h3b4771d7),
	.w8(32'hbc45a382),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf46288),
	.w1(32'hbc31ee11),
	.w2(32'hbbc356f4),
	.w3(32'hbc4420c5),
	.w4(32'hbc4fa3f0),
	.w5(32'hbc245c1e),
	.w6(32'hbbb95442),
	.w7(32'h3c17d0df),
	.w8(32'hbb2242e5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6699cc),
	.w1(32'hbb2cbe42),
	.w2(32'h3b0e241e),
	.w3(32'hbbacce43),
	.w4(32'hbc223e52),
	.w5(32'hbb20ca8c),
	.w6(32'hbc04ec4c),
	.w7(32'hba8eb3fe),
	.w8(32'hba5ac72f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01faba),
	.w1(32'hbb4cb146),
	.w2(32'h3be30941),
	.w3(32'h3c0e3f26),
	.w4(32'h3b9c61da),
	.w5(32'hbcadbb64),
	.w6(32'hbb8a1737),
	.w7(32'hbc13aa0f),
	.w8(32'h3bbe4630),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabff76),
	.w1(32'hbc6a5a2c),
	.w2(32'h3acdf8be),
	.w3(32'hbc8848c1),
	.w4(32'h3ba83746),
	.w5(32'h3b77a503),
	.w6(32'hbc4639b0),
	.w7(32'hbc93db1c),
	.w8(32'h3b28bf83),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b79d7),
	.w1(32'h3a61efea),
	.w2(32'h3bcb3b36),
	.w3(32'h3b52d709),
	.w4(32'h398c5cf4),
	.w5(32'h3b65fd82),
	.w6(32'h3b29ead3),
	.w7(32'hba53d2be),
	.w8(32'hbb18fd8f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad83332),
	.w1(32'h3b74e7af),
	.w2(32'hbb57f411),
	.w3(32'h38a0056d),
	.w4(32'hb993e4cd),
	.w5(32'hbc2a9984),
	.w6(32'hbba878c0),
	.w7(32'hbaca1c9b),
	.w8(32'hbc98b05b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3900a6),
	.w1(32'hbb90adbb),
	.w2(32'hbc0adb8f),
	.w3(32'hbcbcd47f),
	.w4(32'hbce7f8b5),
	.w5(32'hbcb3a471),
	.w6(32'hbc866bca),
	.w7(32'hbc530c80),
	.w8(32'h3c2eacbd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e3e21),
	.w1(32'h3ae187ff),
	.w2(32'h3b5f84c4),
	.w3(32'h3c090aff),
	.w4(32'h3c80b2d1),
	.w5(32'h3a1c501e),
	.w6(32'h3be4aa9b),
	.w7(32'hbc8a9b05),
	.w8(32'h390f6b94),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214a27),
	.w1(32'h3a9fef38),
	.w2(32'hbb01f6e6),
	.w3(32'hbb079cbd),
	.w4(32'hbae2df87),
	.w5(32'h3aac21de),
	.w6(32'hba8c6888),
	.w7(32'h3ae5c546),
	.w8(32'h3bfd3284),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eab84),
	.w1(32'hbb0d10e5),
	.w2(32'hba3d0832),
	.w3(32'h3ace4e73),
	.w4(32'hbb3861e3),
	.w5(32'h3a475321),
	.w6(32'hbb902634),
	.w7(32'h3b1aee40),
	.w8(32'hba8584b2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac98a),
	.w1(32'hbb995843),
	.w2(32'h3b03e2a6),
	.w3(32'hbaea46e0),
	.w4(32'h3b83733a),
	.w5(32'h3c76bdce),
	.w6(32'h3b8d61d3),
	.w7(32'hb9438fc7),
	.w8(32'h3bf07ef9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d3551),
	.w1(32'h3af75cf5),
	.w2(32'hbc51c780),
	.w3(32'h3aecf637),
	.w4(32'h3aca3e20),
	.w5(32'hbc6125fb),
	.w6(32'h3bbdc01f),
	.w7(32'h3c3c8f3f),
	.w8(32'h3c0490b0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82b061),
	.w1(32'h3aa9cbd1),
	.w2(32'hba8996f1),
	.w3(32'h3c5adbd2),
	.w4(32'h3c03c1bb),
	.w5(32'h3a944d1b),
	.w6(32'h3ba01570),
	.w7(32'hbc8b154d),
	.w8(32'hb830ca7a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d749ef),
	.w1(32'h3ae5962c),
	.w2(32'hbc5e2bee),
	.w3(32'hbb057a72),
	.w4(32'hbb062f24),
	.w5(32'hbc41162f),
	.w6(32'hbadb66af),
	.w7(32'h3b06a7a4),
	.w8(32'hbc4cec7b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d36ad),
	.w1(32'hbbab8c1d),
	.w2(32'hbb16875a),
	.w3(32'hbc47c857),
	.w4(32'hbc5d4962),
	.w5(32'hbc047d77),
	.w6(32'hbc00de8c),
	.w7(32'hba803eb2),
	.w8(32'h3cc5e484),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a83c8),
	.w1(32'h3bd14955),
	.w2(32'hbc1415f5),
	.w3(32'h3c978bea),
	.w4(32'h3cb0600a),
	.w5(32'hbc6eab1e),
	.w6(32'hbb6084ea),
	.w7(32'hbc886738),
	.w8(32'h3c77c2e7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3fe8a),
	.w1(32'h3b690c2b),
	.w2(32'h3be19176),
	.w3(32'h3cbe8cec),
	.w4(32'h3ca4d7bd),
	.w5(32'h39c0d3ca),
	.w6(32'hbb78e24a),
	.w7(32'hbcb38f48),
	.w8(32'hbc05739b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71d866),
	.w1(32'hbb741d68),
	.w2(32'h3b39dcdc),
	.w3(32'hbbcd3dac),
	.w4(32'hbbe6adda),
	.w5(32'hba74d04a),
	.w6(32'h3b91aaa1),
	.w7(32'hbbd591a6),
	.w8(32'h3a87ce46),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868e8f),
	.w1(32'h39cacb4e),
	.w2(32'hbaa8c8ea),
	.w3(32'hbb30bfa5),
	.w4(32'hbac7e798),
	.w5(32'hbaa82e05),
	.w6(32'hba916431),
	.w7(32'h3ab2f86b),
	.w8(32'hbb1c245b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824459),
	.w1(32'h3a8881ef),
	.w2(32'hba8008d9),
	.w3(32'h3a37af96),
	.w4(32'h3b786c03),
	.w5(32'hba9c8bbf),
	.w6(32'h388c7f76),
	.w7(32'h3721e629),
	.w8(32'hbb51f133),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc39e7),
	.w1(32'hbaebd4b0),
	.w2(32'hbc107b5a),
	.w3(32'hba818464),
	.w4(32'hba33d076),
	.w5(32'hbb541f66),
	.w6(32'hbaed2668),
	.w7(32'h3adc4408),
	.w8(32'h3be9539e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bba7),
	.w1(32'hb98a2d4c),
	.w2(32'h3af1bff7),
	.w3(32'h3a9bd2ac),
	.w4(32'hbc3a5cd4),
	.w5(32'h3c6f68dd),
	.w6(32'h3a1076de),
	.w7(32'hba51f476),
	.w8(32'hbc18a852),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48436),
	.w1(32'hbba33d71),
	.w2(32'hbb552916),
	.w3(32'hbc8e68af),
	.w4(32'hbc29dba6),
	.w5(32'hb9254f95),
	.w6(32'hba733543),
	.w7(32'h3bae3630),
	.w8(32'h3ae1b5c1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d7e9),
	.w1(32'hbb6f69a1),
	.w2(32'hbc19f966),
	.w3(32'h3b0de718),
	.w4(32'h3b632798),
	.w5(32'h3937f51d),
	.w6(32'hba33e268),
	.w7(32'h3ae20dc0),
	.w8(32'h3b9afb4e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a682),
	.w1(32'h3b9f8d52),
	.w2(32'h3b4facaa),
	.w3(32'h3c0251f9),
	.w4(32'hbcacbe5a),
	.w5(32'h3b926a89),
	.w6(32'hbcb36a40),
	.w7(32'hbc41d42a),
	.w8(32'h3b34c5cc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10cfd0),
	.w1(32'h3b2ebea9),
	.w2(32'hba34cf58),
	.w3(32'hbae3fba9),
	.w4(32'h3b1cabd9),
	.w5(32'hbb106db8),
	.w6(32'hbb3c2313),
	.w7(32'h3b034020),
	.w8(32'hba25fb4c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6a760),
	.w1(32'h3aaf801a),
	.w2(32'hbadd2505),
	.w3(32'hb9cc44ae),
	.w4(32'hbbba057f),
	.w5(32'hbcba9c85),
	.w6(32'hbb7dffe1),
	.w7(32'hbb8357a2),
	.w8(32'h3c915539),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc18909),
	.w1(32'h3c85ac2b),
	.w2(32'h3bf8b4b2),
	.w3(32'h3ba0a3c1),
	.w4(32'h3bd407d6),
	.w5(32'h3bb434d4),
	.w6(32'h3c09743a),
	.w7(32'hbc76ca5a),
	.w8(32'hbb899ad1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96abc4),
	.w1(32'h3b072971),
	.w2(32'h3b3cdc8f),
	.w3(32'hbbb53e77),
	.w4(32'h3adb832c),
	.w5(32'hbbc71d9c),
	.w6(32'hbbf95b4e),
	.w7(32'h3c111787),
	.w8(32'hba33db3e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb416e),
	.w1(32'hbaf2b3ae),
	.w2(32'hbae45172),
	.w3(32'hbbd1328f),
	.w4(32'hbbce8db6),
	.w5(32'h3a9db2c4),
	.w6(32'hba08ee9d),
	.w7(32'h3b7189f5),
	.w8(32'hbc2aa273),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad421d7),
	.w1(32'hbc28959f),
	.w2(32'hbb0c8c53),
	.w3(32'hbb759d61),
	.w4(32'hba8a5273),
	.w5(32'h3a145a81),
	.w6(32'hb9e32d9d),
	.w7(32'h3ad8945b),
	.w8(32'h3a666837),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d512c),
	.w1(32'h3a694a1c),
	.w2(32'hba63742b),
	.w3(32'h3b21a80f),
	.w4(32'h3aa36623),
	.w5(32'hbaab0431),
	.w6(32'h35143cc6),
	.w7(32'hbafbedda),
	.w8(32'h3ab8f78a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af66e0b),
	.w1(32'hbb0dc871),
	.w2(32'hbbf6c81c),
	.w3(32'h3a0e83ca),
	.w4(32'hbb3a615c),
	.w5(32'hbc8f7f28),
	.w6(32'h3b0fa33d),
	.w7(32'h39f68ccd),
	.w8(32'h3c0c9000),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca05c3f),
	.w1(32'h3c05ba4b),
	.w2(32'hbbf8be65),
	.w3(32'h3c767292),
	.w4(32'h3bea7392),
	.w5(32'h3afc072d),
	.w6(32'h3b9cb864),
	.w7(32'hbc771456),
	.w8(32'hbb0a4006),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83c7ed),
	.w1(32'h3bebb802),
	.w2(32'hbba8aa04),
	.w3(32'h3cd6f7ae),
	.w4(32'hbc0aac27),
	.w5(32'hbadc9fe3),
	.w6(32'hbcda10b7),
	.w7(32'hbaf67f9a),
	.w8(32'hbc12cd03),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb960e69),
	.w1(32'h3ae10c55),
	.w2(32'hbb8f7e4b),
	.w3(32'hbc4059d1),
	.w4(32'hbb083c89),
	.w5(32'hbbdd922b),
	.w6(32'hbb4dff1f),
	.w7(32'hbba0f774),
	.w8(32'hbbdb520e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb195d3),
	.w1(32'hbbc6935f),
	.w2(32'hbc484c51),
	.w3(32'hbc110976),
	.w4(32'hbc4cae69),
	.w5(32'hbca0cb6b),
	.w6(32'h3a9297b2),
	.w7(32'h3afc671b),
	.w8(32'h3b9cf3a3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb29d56),
	.w1(32'hba1e50bf),
	.w2(32'h3a89b114),
	.w3(32'hbab2b9bf),
	.w4(32'h3b822c1e),
	.w5(32'h3ba79b01),
	.w6(32'h3aa9fcfb),
	.w7(32'hbc1f53a8),
	.w8(32'hbaea8e1c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b3c74),
	.w1(32'h3aa0d488),
	.w2(32'h3b676a5b),
	.w3(32'h3b9ff393),
	.w4(32'h3ab0a77d),
	.w5(32'hbc050098),
	.w6(32'h3b1d396a),
	.w7(32'h3b78b7e8),
	.w8(32'hbc765921),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f1c0f),
	.w1(32'hbbdc0253),
	.w2(32'h3bc44c4b),
	.w3(32'hbcb70c4c),
	.w4(32'hbca2652b),
	.w5(32'hbc7669b1),
	.w6(32'hbc9e8093),
	.w7(32'hbbb135d9),
	.w8(32'hbc2e502d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc443209),
	.w1(32'hbcd48716),
	.w2(32'h3c35ddf4),
	.w3(32'hbc6db773),
	.w4(32'hbb43ee9a),
	.w5(32'hbbf5fe7c),
	.w6(32'hbcbc1d0d),
	.w7(32'hbcb71064),
	.w8(32'hbbb68af5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0245b),
	.w1(32'hbbd11ad8),
	.w2(32'h3b19f9a5),
	.w3(32'hbbe0fdae),
	.w4(32'hbae0fa87),
	.w5(32'h3ad09fb8),
	.w6(32'hbac63bbb),
	.w7(32'h3b51a551),
	.w8(32'h3bcaf8ea),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2b42),
	.w1(32'h3bc34b90),
	.w2(32'h3bdc18f4),
	.w3(32'h3bd54a41),
	.w4(32'hbbc15f38),
	.w5(32'hbb849563),
	.w6(32'hbc1d521f),
	.w7(32'hbc20457a),
	.w8(32'h3a0a149d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc881c),
	.w1(32'h3b46ced1),
	.w2(32'hbb1eb19a),
	.w3(32'h3b1c9507),
	.w4(32'h3b700dcd),
	.w5(32'hbb14ac12),
	.w6(32'h3b46c119),
	.w7(32'h3b8f1dd1),
	.w8(32'h3b9722cc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe7759),
	.w1(32'h3b5b6a8b),
	.w2(32'h3b5dbea4),
	.w3(32'h3addbc60),
	.w4(32'h3c303a73),
	.w5(32'h3b54a4c4),
	.w6(32'h3ab279cb),
	.w7(32'hbb366d3c),
	.w8(32'hba276157),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266c7e),
	.w1(32'h3b14f5f7),
	.w2(32'h3afb60e2),
	.w3(32'hbb039d13),
	.w4(32'h3b31b77f),
	.w5(32'h39e6d0f0),
	.w6(32'h3ac561a0),
	.w7(32'hbb55251e),
	.w8(32'hbb324a92),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be35676),
	.w1(32'h3aaa8dd4),
	.w2(32'hbb2176ad),
	.w3(32'h3a04f4b7),
	.w4(32'h3a7571e5),
	.w5(32'h3ba2ea75),
	.w6(32'h3b831114),
	.w7(32'h3b8a9b1f),
	.w8(32'hbb41579c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32dfa2),
	.w1(32'h3a49d119),
	.w2(32'h3baa9280),
	.w3(32'hbbe4ce91),
	.w4(32'h3bfa4f19),
	.w5(32'hbbb88795),
	.w6(32'h3b266b63),
	.w7(32'h3c444555),
	.w8(32'hbb64057a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5f816),
	.w1(32'hbbece339),
	.w2(32'h3b3fb602),
	.w3(32'hbc03055a),
	.w4(32'hbae42b2e),
	.w5(32'hbc0cd24a),
	.w6(32'hbbbbfb58),
	.w7(32'hbc47590a),
	.w8(32'hbc022941),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f31e1f),
	.w1(32'hbbd1711e),
	.w2(32'h3acde7b2),
	.w3(32'hbc387040),
	.w4(32'hbbd8be52),
	.w5(32'hb9aade6d),
	.w6(32'hbb9f20da),
	.w7(32'h3c075622),
	.w8(32'hbb3424a2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1949ac),
	.w1(32'h3b35cefc),
	.w2(32'h3c763cd4),
	.w3(32'hbbd75154),
	.w4(32'hbb732759),
	.w5(32'hbb7a7a95),
	.w6(32'h3b006068),
	.w7(32'h3bcac3ea),
	.w8(32'hbaf202a1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97e4d8),
	.w1(32'hbb7ee7f8),
	.w2(32'h3b89ae75),
	.w3(32'hbc6178fa),
	.w4(32'h3cbc4ad3),
	.w5(32'h3ba98f1a),
	.w6(32'h3cfa3670),
	.w7(32'hba46f33d),
	.w8(32'hbbf770a6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc55d),
	.w1(32'hbb0ffa18),
	.w2(32'h3c6041c2),
	.w3(32'hbc5d4d4c),
	.w4(32'hbb474115),
	.w5(32'hbc30afd0),
	.w6(32'hbc11ead3),
	.w7(32'h3b8727e6),
	.w8(32'h3a966505),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484a92),
	.w1(32'hbc6c062a),
	.w2(32'h3b4976f3),
	.w3(32'hbc8ff67c),
	.w4(32'h3cef3db6),
	.w5(32'hb9875f60),
	.w6(32'h3cadee68),
	.w7(32'h3bf81ff6),
	.w8(32'hbb9c2687),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e89cb),
	.w1(32'h3ba3f0f6),
	.w2(32'h3a85cd7f),
	.w3(32'h3b4d0064),
	.w4(32'h3ac3f193),
	.w5(32'hbad1a079),
	.w6(32'hbac79ef9),
	.w7(32'h3b202f90),
	.w8(32'h3b200cfc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba928c4),
	.w1(32'hbb6edca0),
	.w2(32'h3bd6da46),
	.w3(32'hb9fe9bd4),
	.w4(32'h39a214c6),
	.w5(32'hb959bc7f),
	.w6(32'h3b9572ac),
	.w7(32'h3bd27af5),
	.w8(32'h37c87ea5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25436f),
	.w1(32'h3b661da8),
	.w2(32'hbc36a997),
	.w3(32'h3b177aab),
	.w4(32'hbad23ec3),
	.w5(32'hbc8222c4),
	.w6(32'hbb73f8e8),
	.w7(32'hbad60a9d),
	.w8(32'h3bae960e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17cf2c),
	.w1(32'hbb54874e),
	.w2(32'h3b19a9fc),
	.w3(32'hbb9311d9),
	.w4(32'hbaee2733),
	.w5(32'hbc31ea4e),
	.w6(32'hbc439f50),
	.w7(32'hbc84e754),
	.w8(32'hbc4f20f3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ab97),
	.w1(32'hbc9278d7),
	.w2(32'hbc00481b),
	.w3(32'hbc96df69),
	.w4(32'hbc5591cb),
	.w5(32'hbc305fbf),
	.w6(32'hbd08b56f),
	.w7(32'hbc42532a),
	.w8(32'hbb64a70f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5221b2),
	.w1(32'hbadd5a7a),
	.w2(32'hbb3809fa),
	.w3(32'hbc0f5eb6),
	.w4(32'hbc2da2fb),
	.w5(32'hba8f93e8),
	.w6(32'hbbde0603),
	.w7(32'hbaba4468),
	.w8(32'hbb8d421c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae42cd5),
	.w1(32'hbb240db9),
	.w2(32'hbaa23705),
	.w3(32'hbaab05c1),
	.w4(32'hbb9b36bf),
	.w5(32'hbb9900a9),
	.w6(32'hbbd70aba),
	.w7(32'hbbc4f376),
	.w8(32'hbb4e2fc0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb172690),
	.w1(32'hb9d7895d),
	.w2(32'hbab127a9),
	.w3(32'hbb974a4c),
	.w4(32'hbba094f1),
	.w5(32'hb929a1d6),
	.w6(32'hbb05b379),
	.w7(32'hbadcb77e),
	.w8(32'h3b057f89),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718ad5),
	.w1(32'hbbd3bc6a),
	.w2(32'h3bfff6e7),
	.w3(32'h3ac07f52),
	.w4(32'h3b17b076),
	.w5(32'h3af07282),
	.w6(32'h3c682bfa),
	.w7(32'hb8065b41),
	.w8(32'hbb82469f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d46bc),
	.w1(32'hba5b3885),
	.w2(32'hbb4da005),
	.w3(32'hbb4ceabe),
	.w4(32'hbb43741f),
	.w5(32'hbc9885e1),
	.w6(32'hbb974e3d),
	.w7(32'h3b87b13d),
	.w8(32'hbc2b0c74),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2c50b),
	.w1(32'h3abe48fc),
	.w2(32'h3b8e08e5),
	.w3(32'h3b4fb2e2),
	.w4(32'h3b3cf2f8),
	.w5(32'h3c08b275),
	.w6(32'hbadfd354),
	.w7(32'hbbb0c49e),
	.w8(32'hbc27959a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1525),
	.w1(32'hbbc5fd7e),
	.w2(32'h3b9cb109),
	.w3(32'hbcd3809c),
	.w4(32'hbb6f883b),
	.w5(32'hba1dfef1),
	.w6(32'hbc2e07e9),
	.w7(32'hbb9e49ae),
	.w8(32'hbc68d057),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecd276),
	.w1(32'h3b45f92e),
	.w2(32'hbc1c0295),
	.w3(32'hbc959b94),
	.w4(32'hbbb4cc96),
	.w5(32'h3c051b66),
	.w6(32'hbc010177),
	.w7(32'h3c0cf287),
	.w8(32'hbbecb975),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960ed2),
	.w1(32'hbbadbf5e),
	.w2(32'hba7c625b),
	.w3(32'hbb61ddbb),
	.w4(32'h3ac682d1),
	.w5(32'hbc2dc005),
	.w6(32'h3a976493),
	.w7(32'h3c23deba),
	.w8(32'hbc1b1162),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca703e),
	.w1(32'h3bbc7dc8),
	.w2(32'h3c40071b),
	.w3(32'hbbe99608),
	.w4(32'h3b799891),
	.w5(32'h3c20e6f6),
	.w6(32'hbc4f1672),
	.w7(32'hbc5feead),
	.w8(32'hbc761e34),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd8790),
	.w1(32'hbc336ec7),
	.w2(32'h3b930091),
	.w3(32'hbcf652e1),
	.w4(32'hbc0e9993),
	.w5(32'hba24f9f8),
	.w6(32'h3bb0fd1a),
	.w7(32'h3be55d63),
	.w8(32'hbae4752d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacd0c),
	.w1(32'h3af6ad93),
	.w2(32'hbc5e84b1),
	.w3(32'hbc4bbd1a),
	.w4(32'hbbab1274),
	.w5(32'h3cf21ee0),
	.w6(32'hba0213eb),
	.w7(32'h3bd33229),
	.w8(32'h3bdae38a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfac1a0),
	.w1(32'h3d0fb84e),
	.w2(32'h3c3617e5),
	.w3(32'h3d2b5a6d),
	.w4(32'hbc9462f0),
	.w5(32'h3b96c26b),
	.w6(32'hbc930577),
	.w7(32'h3c465527),
	.w8(32'h3c03da97),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ab5aa),
	.w1(32'h3ad9f6de),
	.w2(32'hbb8b160b),
	.w3(32'h3a63ce82),
	.w4(32'hbc45f432),
	.w5(32'hba92c190),
	.w6(32'hb98d6843),
	.w7(32'h3c6c3612),
	.w8(32'h39b10bd4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3744e8),
	.w1(32'h3b09d0d5),
	.w2(32'h3b7fbdef),
	.w3(32'hb93b3b44),
	.w4(32'hbb8ef963),
	.w5(32'hbc5d8305),
	.w6(32'hbb319994),
	.w7(32'hba433c00),
	.w8(32'h3c445cab),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a9a02),
	.w1(32'hbb4be601),
	.w2(32'h3bf1be20),
	.w3(32'h3bf1e2b8),
	.w4(32'h3bc7d452),
	.w5(32'h3b96b22f),
	.w6(32'h3b1c97f4),
	.w7(32'hbbdc5f38),
	.w8(32'hb88ee3f7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a9f0),
	.w1(32'h39f74fca),
	.w2(32'h3b4aa339),
	.w3(32'h3b3422d9),
	.w4(32'h3bad5db1),
	.w5(32'h3bb5c87d),
	.w6(32'h3bf93f7c),
	.w7(32'h3b992860),
	.w8(32'h3b4ad667),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8c86c),
	.w1(32'h3a596ac6),
	.w2(32'hbae5bab4),
	.w3(32'hbb3e1a32),
	.w4(32'h3c32f699),
	.w5(32'hbb66477d),
	.w6(32'h3bb92bb9),
	.w7(32'h3c4230e7),
	.w8(32'hbb178f16),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadefd05),
	.w1(32'hbae337e3),
	.w2(32'h3bf19e26),
	.w3(32'hbb10640d),
	.w4(32'h362e5ae6),
	.w5(32'h3a1553cc),
	.w6(32'hba906064),
	.w7(32'h3aaf8fd8),
	.w8(32'hbb4dc365),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351f56),
	.w1(32'h3b3a3342),
	.w2(32'hba23a6af),
	.w3(32'hbc020dc3),
	.w4(32'hbc3b902d),
	.w5(32'hba80dc34),
	.w6(32'hbbd2ec1c),
	.w7(32'h3b46d956),
	.w8(32'h39d7874a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0869c8),
	.w1(32'hba21656b),
	.w2(32'hbb1075fb),
	.w3(32'hb966e56d),
	.w4(32'h3a58db38),
	.w5(32'h3b39ddb7),
	.w6(32'h3b8a6ea5),
	.w7(32'h3ad724ab),
	.w8(32'h3bcee921),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910bf84),
	.w1(32'hb8408f1e),
	.w2(32'hbc39a683),
	.w3(32'h3af025e5),
	.w4(32'hbaa78717),
	.w5(32'h3ccbb15d),
	.w6(32'h3b338960),
	.w7(32'hbb7137d2),
	.w8(32'h3bc92b06),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978f1d),
	.w1(32'h3ccb1ad4),
	.w2(32'h39469a2f),
	.w3(32'h3cca244f),
	.w4(32'hbc6498d1),
	.w5(32'hbb56ff10),
	.w6(32'hbbdca141),
	.w7(32'h3c32caee),
	.w8(32'hba41c99a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab17397),
	.w1(32'h382d839e),
	.w2(32'hbae5a884),
	.w3(32'h3899f62d),
	.w4(32'h3b054e72),
	.w5(32'hbb188e64),
	.w6(32'h3b2b37e1),
	.w7(32'h3b10c3e8),
	.w8(32'hbb38f654),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c6daa),
	.w1(32'hbb6dfdba),
	.w2(32'h3af205ba),
	.w3(32'hbb214e75),
	.w4(32'hbafc9902),
	.w5(32'hbc0c5778),
	.w6(32'hba4e3c09),
	.w7(32'h39fac288),
	.w8(32'hbc2204b3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fa405),
	.w1(32'hbc11cded),
	.w2(32'h3b9de4d9),
	.w3(32'hbc3fb764),
	.w4(32'hba4e79a9),
	.w5(32'h3ad05949),
	.w6(32'hbb9d89b8),
	.w7(32'h3ac0feb3),
	.w8(32'h3b48fc6d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926606),
	.w1(32'h3b847133),
	.w2(32'h3b477645),
	.w3(32'hbabea6e5),
	.w4(32'h3ad8cbdc),
	.w5(32'hbaeba709),
	.w6(32'hbaaee400),
	.w7(32'h3b320df9),
	.w8(32'hba32145d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9efa39),
	.w1(32'hbc325fc0),
	.w2(32'h3a0f048a),
	.w3(32'hbc30404b),
	.w4(32'hbbe04270),
	.w5(32'hbac7ddc7),
	.w6(32'h3b667339),
	.w7(32'hbb59b80d),
	.w8(32'h3ab58f0f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890701),
	.w1(32'h3b731b1f),
	.w2(32'hbc389316),
	.w3(32'h3b649b08),
	.w4(32'hbbb37e09),
	.w5(32'hbc3d2849),
	.w6(32'hbc2f1925),
	.w7(32'hbc1f6cbc),
	.w8(32'hbc15a1d3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85190),
	.w1(32'hbc2710b6),
	.w2(32'hbacf5315),
	.w3(32'hbca13c58),
	.w4(32'hbc41321f),
	.w5(32'h3a35da12),
	.w6(32'h3a232538),
	.w7(32'hbae182c4),
	.w8(32'hbc17f227),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73b4a7),
	.w1(32'hb98e8be3),
	.w2(32'hbb240d5c),
	.w3(32'hbbe5471f),
	.w4(32'hbc6e6cf2),
	.w5(32'hbb30a7fe),
	.w6(32'hbbca4206),
	.w7(32'h3a8c81d6),
	.w8(32'hba7332d5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e07a),
	.w1(32'hbb6ed68e),
	.w2(32'hbb8c0759),
	.w3(32'hbb89a285),
	.w4(32'hbaf0ef5c),
	.w5(32'hbb30a09f),
	.w6(32'hbb64fed0),
	.w7(32'hbad1e925),
	.w8(32'h3beca204),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad8e09),
	.w1(32'h3be38ada),
	.w2(32'h3c48f926),
	.w3(32'h3b8994ba),
	.w4(32'h3b12da5a),
	.w5(32'hbb8db8cb),
	.w6(32'hbb63b13a),
	.w7(32'hbb03fc35),
	.w8(32'hbaa12738),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9037),
	.w1(32'hbbeb1326),
	.w2(32'h3c0574e7),
	.w3(32'hbade6477),
	.w4(32'h3c31469f),
	.w5(32'hbc54bfc7),
	.w6(32'h3c9aae4f),
	.w7(32'h3bb73d56),
	.w8(32'h3ce64e9a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d457c),
	.w1(32'h3c93b10f),
	.w2(32'hba918326),
	.w3(32'h3d31f8b9),
	.w4(32'h3d0d95a2),
	.w5(32'hb8034788),
	.w6(32'h3bf280b9),
	.w7(32'hbc38b71a),
	.w8(32'h3b05896f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813fbb),
	.w1(32'hbbc2299a),
	.w2(32'h3b37e365),
	.w3(32'hbc47aee8),
	.w4(32'hbbdf65f4),
	.w5(32'h3b6f06a1),
	.w6(32'hbb0e7db8),
	.w7(32'hbb148c58),
	.w8(32'h3b49ab4f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3b3b1),
	.w1(32'hbb0ee870),
	.w2(32'h393d06e5),
	.w3(32'h3b5d84b2),
	.w4(32'hbb558ebc),
	.w5(32'h398993ac),
	.w6(32'h3b172211),
	.w7(32'h3b03e0f0),
	.w8(32'hbaa86e24),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9386c7),
	.w1(32'hbaa0dd0d),
	.w2(32'hbbf6e144),
	.w3(32'h3b82687e),
	.w4(32'h3b5bd8ce),
	.w5(32'hbc4587b0),
	.w6(32'h3b09cc41),
	.w7(32'h3aa184fb),
	.w8(32'h3c5f9605),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd037c54),
	.w1(32'hbca47b2c),
	.w2(32'hba978d5e),
	.w3(32'hbd383a75),
	.w4(32'hbd112c7a),
	.w5(32'h3aa8077d),
	.w6(32'hbbd9e912),
	.w7(32'h3aac9d18),
	.w8(32'hbab5ae94),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147113),
	.w1(32'h3a957105),
	.w2(32'h3b637aa4),
	.w3(32'h39452b87),
	.w4(32'hb90c57c4),
	.w5(32'h3b732f3b),
	.w6(32'hba61bc44),
	.w7(32'h3a91dba9),
	.w8(32'h3a0c7983),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31bdca),
	.w1(32'h3b303d5f),
	.w2(32'hbbb09bc9),
	.w3(32'h3bee30be),
	.w4(32'h3badf173),
	.w5(32'hbc5ac18d),
	.w6(32'h3ade59b2),
	.w7(32'h3ba1a6d5),
	.w8(32'h3c13fb99),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9cd38),
	.w1(32'hbc5cfe53),
	.w2(32'h3b5667c7),
	.w3(32'hbd16508d),
	.w4(32'hbcc0983c),
	.w5(32'hbb4e9911),
	.w6(32'hbc0b1848),
	.w7(32'h3b418edc),
	.w8(32'hb9bb4f71),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0b1b),
	.w1(32'hbb6aa999),
	.w2(32'h3b70c64b),
	.w3(32'h3a8c4d69),
	.w4(32'hbaf71687),
	.w5(32'h3bf552b7),
	.w6(32'h385d69cd),
	.w7(32'h3b6081a6),
	.w8(32'hbc4dafcf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc584e5),
	.w1(32'h3c621f7f),
	.w2(32'h3a0a05ba),
	.w3(32'h3d150da4),
	.w4(32'h3cd64595),
	.w5(32'h3b7a8470),
	.w6(32'h3bec3cdf),
	.w7(32'hb9c5b5de),
	.w8(32'hbb96876a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb076d3c),
	.w1(32'hbb34aea6),
	.w2(32'hbb98f7c2),
	.w3(32'h3b6f1086),
	.w4(32'h3b178fb3),
	.w5(32'hbb9a1f50),
	.w6(32'h3927165d),
	.w7(32'hbad5bf44),
	.w8(32'h3befbec7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123d06),
	.w1(32'h3b7c997b),
	.w2(32'hba438964),
	.w3(32'hbc223bf9),
	.w4(32'hba070be6),
	.w5(32'hbb9282ff),
	.w6(32'h3bdf1c17),
	.w7(32'h3c964f40),
	.w8(32'hbbd52829),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3818df),
	.w1(32'h3b8b8a18),
	.w2(32'hbb0f55fe),
	.w3(32'hbbdc5164),
	.w4(32'hbb012cb1),
	.w5(32'hbbd4f658),
	.w6(32'hbbb63391),
	.w7(32'hbbabe00d),
	.w8(32'hbc21132d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dd0f9),
	.w1(32'hbab380ac),
	.w2(32'h3b277a66),
	.w3(32'hbbf552ee),
	.w4(32'hba540d2c),
	.w5(32'hbae7fb0a),
	.w6(32'hbb265ec8),
	.w7(32'hbc11e3da),
	.w8(32'h3b9bd096),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b503efb),
	.w1(32'hb9ac5b2f),
	.w2(32'h39a7637b),
	.w3(32'h3a5f646b),
	.w4(32'hbb745894),
	.w5(32'hbb3bf6e9),
	.w6(32'hbb0ad7d1),
	.w7(32'hb97e1f7f),
	.w8(32'hbc1d704c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3eba0),
	.w1(32'h3b09e98d),
	.w2(32'hba31f026),
	.w3(32'h3a065281),
	.w4(32'h3b587085),
	.w5(32'hbb965d79),
	.w6(32'hbb269a7f),
	.w7(32'hbb56fe05),
	.w8(32'h3a965c53),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847ecfd),
	.w1(32'h3a2285cd),
	.w2(32'hbc8db962),
	.w3(32'hbb8174a5),
	.w4(32'hbb14435c),
	.w5(32'hbb69d897),
	.w6(32'hbb2d6740),
	.w7(32'hbac822f6),
	.w8(32'hbc1eafe1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30757e),
	.w1(32'hbca8e31c),
	.w2(32'hba2462a5),
	.w3(32'h3a72807d),
	.w4(32'hbbfb1a09),
	.w5(32'h3a847c31),
	.w6(32'hbbe02084),
	.w7(32'hbc767dd2),
	.w8(32'h3b112e2f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78cecd6),
	.w1(32'hbb55a437),
	.w2(32'hba2564f0),
	.w3(32'hbbcfe4e8),
	.w4(32'h38e6890b),
	.w5(32'hbb58fb73),
	.w6(32'hbacae173),
	.w7(32'hbaf9d891),
	.w8(32'hbb5911df),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872200),
	.w1(32'hbbc89d0a),
	.w2(32'hbb20aa3d),
	.w3(32'hba4d06db),
	.w4(32'hb98743af),
	.w5(32'hbb5ba562),
	.w6(32'hbba0d867),
	.w7(32'hbb8b5aed),
	.w8(32'hbb81ffa4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafde131),
	.w1(32'h3b41b899),
	.w2(32'h3b1ab3f4),
	.w3(32'h3b146f8a),
	.w4(32'h3b6a7522),
	.w5(32'h3931896e),
	.w6(32'hb9652f4f),
	.w7(32'h3b45b215),
	.w8(32'h3b101e99),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11e068),
	.w1(32'h3c160a2f),
	.w2(32'hbb1b610d),
	.w3(32'hbb8bfb89),
	.w4(32'hba0efdce),
	.w5(32'h3c07173e),
	.w6(32'hbb805090),
	.w7(32'hbb24ea37),
	.w8(32'hbcd9fc16),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0bb985),
	.w1(32'h3c973e96),
	.w2(32'hba0a1214),
	.w3(32'h3d5e3047),
	.w4(32'h3d242403),
	.w5(32'hbb2f4832),
	.w6(32'h3bc6ccca),
	.w7(32'hbb95f359),
	.w8(32'hbb152207),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e6ec2),
	.w1(32'h3ac4d0ab),
	.w2(32'h3acd90bb),
	.w3(32'h3b9078d2),
	.w4(32'h3a4534f9),
	.w5(32'h3bfd6473),
	.w6(32'hbb3dbcb1),
	.w7(32'h3afee920),
	.w8(32'h3b142b12),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90aca),
	.w1(32'hbb1ffe57),
	.w2(32'h3b2ea18d),
	.w3(32'h3b244d13),
	.w4(32'hb9f79200),
	.w5(32'hbbc71759),
	.w6(32'hb9db7f81),
	.w7(32'hbb033c1a),
	.w8(32'hbbe8f95f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63f8910),
	.w1(32'h3aeaa9b1),
	.w2(32'hba23e751),
	.w3(32'h39b1e30b),
	.w4(32'hbba7a0da),
	.w5(32'h3af2ae68),
	.w6(32'hbb15760e),
	.w7(32'hbb8a8085),
	.w8(32'h3b8057ac),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad41523),
	.w1(32'hbb8cc6d1),
	.w2(32'h3acff446),
	.w3(32'h388e97ef),
	.w4(32'h3a5bb721),
	.w5(32'hbb3ca56f),
	.w6(32'hb845a2a6),
	.w7(32'hbb0c9c5f),
	.w8(32'hbb92a971),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a757),
	.w1(32'h3ba4c51e),
	.w2(32'hbb66e5a6),
	.w3(32'h39c3030c),
	.w4(32'hbad0f202),
	.w5(32'hbbf3f289),
	.w6(32'hbb9ee7c7),
	.w7(32'hbbd34405),
	.w8(32'hbb8dc3ac),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac76b56),
	.w1(32'hbad0e997),
	.w2(32'h3b401477),
	.w3(32'hbc09394d),
	.w4(32'hbc22eea2),
	.w5(32'h3b3aba4a),
	.w6(32'hbb818dad),
	.w7(32'hbc0cee0b),
	.w8(32'hbaf3b544),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f078c),
	.w1(32'h3aa6e088),
	.w2(32'h3ae8e696),
	.w3(32'hbb10bde5),
	.w4(32'h3a3bd532),
	.w5(32'hbb1f1f6f),
	.w6(32'hbaea5585),
	.w7(32'h3a587cb1),
	.w8(32'hbbdcaba2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b104b8b),
	.w1(32'h3b8b55f3),
	.w2(32'hbb846d06),
	.w3(32'h3b2a7c97),
	.w4(32'h3b1810a2),
	.w5(32'hbb9e36ff),
	.w6(32'hbb0df8b0),
	.w7(32'hbbbce37e),
	.w8(32'hbbbfe021),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf5f3e),
	.w1(32'h3bba0d61),
	.w2(32'h39a409c8),
	.w3(32'hbb4e6b20),
	.w4(32'h3bb1312d),
	.w5(32'h3b0b241a),
	.w6(32'hbb0047b9),
	.w7(32'h3b191ce5),
	.w8(32'h3b8d2fa5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0379b),
	.w1(32'h3ac18c30),
	.w2(32'h3b59a926),
	.w3(32'hbb84694d),
	.w4(32'hbb3018ca),
	.w5(32'h39015c6f),
	.w6(32'hbbe6aa0c),
	.w7(32'hbc2b3858),
	.w8(32'hba1c791a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac021ad),
	.w1(32'h3b327cf7),
	.w2(32'h3a83d006),
	.w3(32'h3ba54fa7),
	.w4(32'h3b97c9aa),
	.w5(32'h3b49a747),
	.w6(32'h3b0011de),
	.w7(32'h3bad474e),
	.w8(32'h3bb4e867),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0c27e),
	.w1(32'hbb0c4498),
	.w2(32'h3abf4063),
	.w3(32'hb9b43790),
	.w4(32'hbba143fd),
	.w5(32'h3b3b331f),
	.w6(32'h3ad4d105),
	.w7(32'hbaeda720),
	.w8(32'hba95d1f0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c360a),
	.w1(32'h3b9db72b),
	.w2(32'hbaedc7fe),
	.w3(32'h3b0085be),
	.w4(32'h3bc6811c),
	.w5(32'h3ae3335b),
	.w6(32'h3a590f6d),
	.w7(32'h3b8f5855),
	.w8(32'h3b3ce90b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9201cc),
	.w1(32'h3aef33d3),
	.w2(32'hbad2f6d0),
	.w3(32'hbb292563),
	.w4(32'h3ad23f50),
	.w5(32'h3bde6f25),
	.w6(32'h3ac2074f),
	.w7(32'h3b54704a),
	.w8(32'h3ac300d8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9760ef),
	.w1(32'h3b064f38),
	.w2(32'hba3b1604),
	.w3(32'h3c2329c8),
	.w4(32'h3ba17d2e),
	.w5(32'h3b76815d),
	.w6(32'h3b0776f1),
	.w7(32'hbab17f12),
	.w8(32'hbc00df78),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa892ba),
	.w1(32'hba1b0416),
	.w2(32'h3bbd2bd9),
	.w3(32'hbaa112b5),
	.w4(32'hba0b19f6),
	.w5(32'h3b6b25f3),
	.w6(32'hbb638a3f),
	.w7(32'hbb8d043f),
	.w8(32'h3ba2eb80),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becf2d9),
	.w1(32'h3b50eac9),
	.w2(32'hbc2ca51d),
	.w3(32'h3bd65b02),
	.w4(32'h3ba918b2),
	.w5(32'hbc076c04),
	.w6(32'h3b9c9e1a),
	.w7(32'h3b991a69),
	.w8(32'h3ca66264),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b6801),
	.w1(32'hbd02d35e),
	.w2(32'h3ada9e26),
	.w3(32'hbd42c77f),
	.w4(32'hbd1f01e9),
	.w5(32'h3a150ab7),
	.w6(32'hbba7b80f),
	.w7(32'hba66292f),
	.w8(32'h39f85c40),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e83e),
	.w1(32'hbb216ada),
	.w2(32'h3b4d36ac),
	.w3(32'h3ae77548),
	.w4(32'hbaf1ec98),
	.w5(32'h3b34ba6b),
	.w6(32'hb99532d9),
	.w7(32'h3ae03182),
	.w8(32'h3b18eeed),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282554),
	.w1(32'hbb564031),
	.w2(32'h3aaeb2b8),
	.w3(32'h3add8338),
	.w4(32'hbb8140ba),
	.w5(32'hbb277d62),
	.w6(32'hbb3c2852),
	.w7(32'hbbbc4792),
	.w8(32'hba96029d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8c94),
	.w1(32'h3ab8105f),
	.w2(32'h3baf5922),
	.w3(32'hbae34ad5),
	.w4(32'hbb77548c),
	.w5(32'h3b176713),
	.w6(32'hbaf943a2),
	.w7(32'hbb17fdc7),
	.w8(32'hb9e947da),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fe46c),
	.w1(32'h3b9d84f3),
	.w2(32'h3984788e),
	.w3(32'h3ba48830),
	.w4(32'h3b1d7832),
	.w5(32'hb9dd20ef),
	.w6(32'h3b5f15dd),
	.w7(32'hba1e892c),
	.w8(32'hba6a5e70),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806f79),
	.w1(32'h3af64238),
	.w2(32'hbb4e8f20),
	.w3(32'hb9c74869),
	.w4(32'h3b0b627c),
	.w5(32'hba67dacd),
	.w6(32'hbb88f1f2),
	.w7(32'hbb521d64),
	.w8(32'hbbc23360),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b3007),
	.w1(32'hbb4efc39),
	.w2(32'h3ad209cc),
	.w3(32'h3a62b1e7),
	.w4(32'hb8d3c594),
	.w5(32'hbbef9109),
	.w6(32'hbaefd87e),
	.w7(32'hba8ff5a4),
	.w8(32'hbc36633f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accdd14),
	.w1(32'h3b255b2a),
	.w2(32'hbc8cf175),
	.w3(32'hbb65484f),
	.w4(32'h39d7ba91),
	.w5(32'hba8e2860),
	.w6(32'hbc00b96e),
	.w7(32'hba3b1693),
	.w8(32'hbca41f79),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef0296),
	.w1(32'hbc06ba33),
	.w2(32'hbac45169),
	.w3(32'h3cd66154),
	.w4(32'h3c512877),
	.w5(32'hbb814538),
	.w6(32'h3a88ff71),
	.w7(32'hbc1fedbb),
	.w8(32'hbb9ff837),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d94a),
	.w1(32'h3b8849e5),
	.w2(32'h3a040eac),
	.w3(32'hb9fc11d2),
	.w4(32'h39c84342),
	.w5(32'h3b256747),
	.w6(32'hbbd0bf0e),
	.w7(32'hbb6d49fb),
	.w8(32'hbb1693c1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8899d),
	.w1(32'h3a6b320a),
	.w2(32'h3a87efe0),
	.w3(32'h3b521afb),
	.w4(32'hbb626a2b),
	.w5(32'h3b3f68f0),
	.w6(32'hbb43f46c),
	.w7(32'h3a000bce),
	.w8(32'hbb622e30),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b097d12),
	.w1(32'h3affd666),
	.w2(32'hbb5a195c),
	.w3(32'h3ba8106a),
	.w4(32'h3b7815cc),
	.w5(32'hbb7fea42),
	.w6(32'hbb055bcc),
	.w7(32'h3a903f1e),
	.w8(32'hbb4c07b8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4387de),
	.w1(32'h3b8e1e01),
	.w2(32'hbb0274d0),
	.w3(32'hbbb34754),
	.w4(32'hb965c975),
	.w5(32'hbbc3b60e),
	.w6(32'hbc2b9eba),
	.w7(32'hbb8e153f),
	.w8(32'h3b620c65),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec891),
	.w1(32'hbc0c07e4),
	.w2(32'hbb933774),
	.w3(32'hbca6d0a2),
	.w4(32'hbc8447a3),
	.w5(32'hbbcf7886),
	.w6(32'hbb8937f9),
	.w7(32'hbb21ac41),
	.w8(32'hbbda75d6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a32fc),
	.w1(32'hbb8bd311),
	.w2(32'hbce79531),
	.w3(32'hbba77da1),
	.w4(32'hbbdda967),
	.w5(32'hbcd0322b),
	.w6(32'hbbcdbff6),
	.w7(32'hbb77c946),
	.w8(32'h3bc90913),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd85bddd),
	.w1(32'hbd676e8e),
	.w2(32'hbb4a5024),
	.w3(32'hbda6a1cd),
	.w4(32'hbd8c4774),
	.w5(32'hba7faf67),
	.w6(32'hbceb421d),
	.w7(32'hbca5c785),
	.w8(32'hba6b3c06),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea82a4),
	.w1(32'h39e74c74),
	.w2(32'hbbac9712),
	.w3(32'hbaaeeccf),
	.w4(32'h3af71182),
	.w5(32'h3aa8a1d3),
	.w6(32'hbb555552),
	.w7(32'hb9e1e8d3),
	.w8(32'hbaab9c60),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22abbf),
	.w1(32'hbaf7cb15),
	.w2(32'hbb56a362),
	.w3(32'h3ab507f9),
	.w4(32'h3b118963),
	.w5(32'h3a78a066),
	.w6(32'hbbdeaecc),
	.w7(32'hbb622fe5),
	.w8(32'h3b0db7db),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9463f4),
	.w1(32'hbac1cf2f),
	.w2(32'h396952bb),
	.w3(32'hbba3b75f),
	.w4(32'h3b20e1ba),
	.w5(32'h3b316675),
	.w6(32'h3aaf3a89),
	.w7(32'h3b58ba40),
	.w8(32'hbb9a6278),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0ec7),
	.w1(32'h3bc18ec8),
	.w2(32'h39b61b9e),
	.w3(32'hbb835e1c),
	.w4(32'hb8cf8fee),
	.w5(32'hbb2d6ab6),
	.w6(32'hbbd89e7e),
	.w7(32'h3af884b3),
	.w8(32'hbb2afdfd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbb755),
	.w1(32'h3b1d0b8d),
	.w2(32'h3a6d39f7),
	.w3(32'hb9a7b990),
	.w4(32'hba4659e1),
	.w5(32'hbb2cb5c8),
	.w6(32'hbaf8024a),
	.w7(32'hbb7aed9e),
	.w8(32'h3bb22a11),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168cfc),
	.w1(32'hbb0b3d3f),
	.w2(32'hbb0b0b03),
	.w3(32'hbbc755da),
	.w4(32'hbba7a2c4),
	.w5(32'h3b900343),
	.w6(32'h3b1b44a3),
	.w7(32'h3b50990f),
	.w8(32'h3b9699a9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada0ebf),
	.w1(32'hbad1465f),
	.w2(32'hb9b85b23),
	.w3(32'hba839a20),
	.w4(32'hb92a9032),
	.w5(32'h3b266d6a),
	.w6(32'h38a20e56),
	.w7(32'hbacef29b),
	.w8(32'hbbf3caf7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4d2a2),
	.w1(32'hb9961e74),
	.w2(32'h3c767a45),
	.w3(32'h37b47d81),
	.w4(32'hb87acb62),
	.w5(32'h3c28742e),
	.w6(32'hbc0c804c),
	.w7(32'hbbaa3dad),
	.w8(32'h3c2bc08d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cc4a1),
	.w1(32'h3c6eac26),
	.w2(32'hbba2e9c4),
	.w3(32'h3c7c733e),
	.w4(32'h3c8bf6ba),
	.w5(32'h3b5a852d),
	.w6(32'h3c85f983),
	.w7(32'h3c84a101),
	.w8(32'hba05e441),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69d824),
	.w1(32'hbc2b7723),
	.w2(32'h3c1ef955),
	.w3(32'h3ba93f50),
	.w4(32'hbb882e6c),
	.w5(32'h3b820710),
	.w6(32'h3b7a4972),
	.w7(32'hbbd5eb9e),
	.w8(32'h3b9b8f70),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a6133),
	.w1(32'h3c4cda46),
	.w2(32'h3ac7ebe6),
	.w3(32'h3bc0c3de),
	.w4(32'h3bc3dca8),
	.w5(32'h3b64166a),
	.w6(32'h3bbdbbb3),
	.w7(32'h3be0798b),
	.w8(32'h3c96f3de),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b95f1),
	.w1(32'hbbe145e2),
	.w2(32'hbaebeef0),
	.w3(32'hbc6284d9),
	.w4(32'hbc3812b1),
	.w5(32'h39d06297),
	.w6(32'h3bfb6c6a),
	.w7(32'h3bd74e12),
	.w8(32'hbac71469),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8a14),
	.w1(32'hbb8fc4bc),
	.w2(32'h3c042dd9),
	.w3(32'hbb79c598),
	.w4(32'hba93f141),
	.w5(32'hb8396a4e),
	.w6(32'h3a3a7629),
	.w7(32'hbbdd1a59),
	.w8(32'h3bc46fff),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af41dcf),
	.w1(32'h3b7c0b74),
	.w2(32'h3b5204ea),
	.w3(32'hbb79c28f),
	.w4(32'h3b8a42c0),
	.w5(32'hb8ea55aa),
	.w6(32'hbb007d41),
	.w7(32'h3bb4ad66),
	.w8(32'hbb4958f2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb400c65),
	.w1(32'h3b29e77c),
	.w2(32'hbb55df40),
	.w3(32'hbb2e3ddc),
	.w4(32'h38428a3e),
	.w5(32'hba67953a),
	.w6(32'hbbda0068),
	.w7(32'hbae2b2ee),
	.w8(32'hbac247e8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3ed5),
	.w1(32'hb932447c),
	.w2(32'hbb9ad0e3),
	.w3(32'hba253871),
	.w4(32'hba0d3376),
	.w5(32'hba18ae4c),
	.w6(32'h3b63385e),
	.w7(32'hba4d21ef),
	.w8(32'hbb449ce6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe3c02),
	.w1(32'h3aa2be49),
	.w2(32'hbbd6b515),
	.w3(32'h3b07c5e7),
	.w4(32'h3ab550b3),
	.w5(32'hbc01028e),
	.w6(32'hba24fcb2),
	.w7(32'hbbb8197e),
	.w8(32'hbc13661c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5b36),
	.w1(32'hbae61d46),
	.w2(32'hb847a0bb),
	.w3(32'hbc08b841),
	.w4(32'hbbaaf616),
	.w5(32'hb8f66717),
	.w6(32'hbb95388e),
	.w7(32'hbad95bc1),
	.w8(32'hbab3fada),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0531c1),
	.w1(32'h3a8c4ee2),
	.w2(32'h3ab84f71),
	.w3(32'hbb55b95b),
	.w4(32'h3aca31aa),
	.w5(32'hbb93f157),
	.w6(32'hbb6cb316),
	.w7(32'h3a6192b2),
	.w8(32'hbb2831fb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a243cce),
	.w1(32'hb9e3c0fc),
	.w2(32'hbb7ffad8),
	.w3(32'hbb2d3730),
	.w4(32'hb95dacaf),
	.w5(32'hbba91649),
	.w6(32'hbaf325a2),
	.w7(32'h3a819f04),
	.w8(32'hbc01fdd5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3116d),
	.w1(32'hbb7548d4),
	.w2(32'hba2da1a1),
	.w3(32'h3b15a501),
	.w4(32'hb9511089),
	.w5(32'hbb12c54b),
	.w6(32'hbb394314),
	.w7(32'hbbaa1486),
	.w8(32'hbb3023dc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f44a3d),
	.w1(32'h3bd27d97),
	.w2(32'h3aa2256d),
	.w3(32'hba250bb6),
	.w4(32'h3bc532d6),
	.w5(32'hbb4e3445),
	.w6(32'hbb3e327a),
	.w7(32'hb9adfe38),
	.w8(32'hbb00fef1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef35d6),
	.w1(32'hba9bd6ca),
	.w2(32'h39aa83f4),
	.w3(32'hba4c2601),
	.w4(32'hbacb27d1),
	.w5(32'hbb075200),
	.w6(32'hbb809d48),
	.w7(32'hba57d698),
	.w8(32'hbbec377a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4286f3),
	.w1(32'h3b6e17fd),
	.w2(32'h3bd7ced8),
	.w3(32'hbabb262f),
	.w4(32'hbb361eee),
	.w5(32'h3b079b00),
	.w6(32'hbbd0a7ea),
	.w7(32'hbbb2e935),
	.w8(32'hbac5a6bd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c370102),
	.w1(32'h3c000837),
	.w2(32'hbb47e6b8),
	.w3(32'h3bb63d9b),
	.w4(32'h3b840d22),
	.w5(32'hbc1e6d0a),
	.w6(32'hbae748bf),
	.w7(32'hba60b803),
	.w8(32'hbc07e211),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df482),
	.w1(32'h3a9d1017),
	.w2(32'hbb8c3fda),
	.w3(32'hbb427589),
	.w4(32'hbbb40a0e),
	.w5(32'hba9bbb87),
	.w6(32'hbc07fc25),
	.w7(32'hbbfe1d43),
	.w8(32'hba9e33d9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c00f7),
	.w1(32'h3b9998a1),
	.w2(32'h3b04934a),
	.w3(32'hba94abfa),
	.w4(32'hb8d896f3),
	.w5(32'hbb5268c9),
	.w6(32'h3aba4503),
	.w7(32'h3a9e65ce),
	.w8(32'hbacb84c2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34600),
	.w1(32'h3bd5af33),
	.w2(32'hbb23e7f7),
	.w3(32'h3ad136f0),
	.w4(32'h3b0f742a),
	.w5(32'hb9ab8c29),
	.w6(32'h3aa400d2),
	.w7(32'hbb468879),
	.w8(32'h38654c2b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0d8c0),
	.w1(32'h399893db),
	.w2(32'h3b507f5e),
	.w3(32'hbb5a2803),
	.w4(32'hba353eb7),
	.w5(32'hbb9a4bb1),
	.w6(32'hbb3ddff5),
	.w7(32'hbb323666),
	.w8(32'hbb92e912),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbedf10),
	.w1(32'h3b6f8567),
	.w2(32'h3b0d803c),
	.w3(32'h3be65991),
	.w4(32'h3ad9934c),
	.w5(32'hbb3e8911),
	.w6(32'hbb541351),
	.w7(32'h3ad21f04),
	.w8(32'hbb9f588b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74e052),
	.w1(32'h3b0a8e9b),
	.w2(32'hbb810355),
	.w3(32'h3b7baf5b),
	.w4(32'h3aba4365),
	.w5(32'hbb99ec5d),
	.w6(32'h3b0e49a1),
	.w7(32'h3a2b2ad5),
	.w8(32'hbb474c41),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16ebd1),
	.w1(32'h39ab498d),
	.w2(32'hbace1102),
	.w3(32'hbb270598),
	.w4(32'h3b24f4e2),
	.w5(32'h3b2d7d07),
	.w6(32'hbbf543f4),
	.w7(32'hbb62e3bc),
	.w8(32'h3bbeb3fc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9169a15),
	.w1(32'hbb589e13),
	.w2(32'hbb7f7421),
	.w3(32'h3b805626),
	.w4(32'h3b0c09e8),
	.w5(32'hbc0b4152),
	.w6(32'h3b627ef6),
	.w7(32'h3b903d5d),
	.w8(32'hbbfbbd99),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ede9),
	.w1(32'hbbaa86c2),
	.w2(32'hb9c7c6ff),
	.w3(32'hbc20c11d),
	.w4(32'hbc0af889),
	.w5(32'hbb4e8645),
	.w6(32'hbc0a902d),
	.w7(32'hbbeb753e),
	.w8(32'hb92ce227),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc61723),
	.w1(32'h3bbacdc1),
	.w2(32'hbb58be0b),
	.w3(32'hba7a202b),
	.w4(32'h3b594dba),
	.w5(32'hbb8c4992),
	.w6(32'hbaa38691),
	.w7(32'hbb8f996d),
	.w8(32'hbb23901d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaffc79),
	.w1(32'hbbaac6f1),
	.w2(32'hbb5014dd),
	.w3(32'hbbcada3f),
	.w4(32'hbb939283),
	.w5(32'hbb82f2af),
	.w6(32'hbc02925c),
	.w7(32'hbc00d711),
	.w8(32'hb9f13261),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6091),
	.w1(32'hbb40b77b),
	.w2(32'h3baf6e96),
	.w3(32'hbbc9e419),
	.w4(32'hbaa76b3c),
	.w5(32'hbb0cd116),
	.w6(32'hba4206d9),
	.w7(32'hbadaa34d),
	.w8(32'hbac7ff47),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d653),
	.w1(32'h3b715bc6),
	.w2(32'h39fd88b3),
	.w3(32'h3ae328a4),
	.w4(32'hbb7eca96),
	.w5(32'hbaefccb9),
	.w6(32'hba55ebd4),
	.w7(32'hba6b2630),
	.w8(32'h3a41203c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1660),
	.w1(32'hb9a7bf18),
	.w2(32'h3be1d221),
	.w3(32'hbb384ca5),
	.w4(32'hbb3e7e31),
	.w5(32'h3c06372f),
	.w6(32'h3a4366e6),
	.w7(32'h3a53294b),
	.w8(32'h3b160499),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c390dca),
	.w1(32'h3c5dbed3),
	.w2(32'h3a3c69ff),
	.w3(32'h3c77fa71),
	.w4(32'h3c8b0b81),
	.w5(32'hbb16abd5),
	.w6(32'h3c33aae7),
	.w7(32'h3c3cd1cc),
	.w8(32'h3bb0ee93),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9206e9),
	.w1(32'h3b151ec2),
	.w2(32'hbbaa12b0),
	.w3(32'hbc306ba1),
	.w4(32'hbba81ee8),
	.w5(32'h3b0965de),
	.w6(32'h39987015),
	.w7(32'h3badd3e5),
	.w8(32'hbb2b85fe),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322483),
	.w1(32'h3b8becd1),
	.w2(32'hba768670),
	.w3(32'hbbe2357f),
	.w4(32'h3b9c3715),
	.w5(32'hb999ca34),
	.w6(32'hbc38c1ee),
	.w7(32'hbb3b3b0f),
	.w8(32'hbb481502),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae8360),
	.w1(32'hbb895fea),
	.w2(32'h3b2d0b9d),
	.w3(32'hbb227b92),
	.w4(32'hbb6451a4),
	.w5(32'hbb0335ba),
	.w6(32'hbb512ffb),
	.w7(32'hbb5a5527),
	.w8(32'h3a0c6743),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23d2f7),
	.w1(32'h3b53c5f7),
	.w2(32'hbb4851b5),
	.w3(32'h38fa99e5),
	.w4(32'hbb559105),
	.w5(32'h3b2641ab),
	.w6(32'hbaece718),
	.w7(32'hbb0aca8e),
	.w8(32'h3b4d761a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42611a),
	.w1(32'h3bd34f75),
	.w2(32'hbb532ce3),
	.w3(32'hba7b94d0),
	.w4(32'h3b44260f),
	.w5(32'hbb6a4028),
	.w6(32'hbab6015b),
	.w7(32'h3b03166c),
	.w8(32'hbb2a0581),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56eca9),
	.w1(32'hb9c73523),
	.w2(32'h3956e171),
	.w3(32'h3a88cfb2),
	.w4(32'h3b04cfbf),
	.w5(32'hbbdd033d),
	.w6(32'hba766531),
	.w7(32'hbac749b1),
	.w8(32'hbba570b5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule