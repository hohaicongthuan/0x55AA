module layer_10_featuremap_27(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8d20),
	.w1(32'h3c942966),
	.w2(32'hbc819897),
	.w3(32'hbcc63a68),
	.w4(32'h3c45d97f),
	.w5(32'h3baaa1dc),
	.w6(32'hbcad1280),
	.w7(32'h3b2dcff2),
	.w8(32'h3c51e0dc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3c316),
	.w1(32'hbc2a9983),
	.w2(32'hba50399b),
	.w3(32'hbc61d087),
	.w4(32'hbb3b2f2a),
	.w5(32'hbc4b30b7),
	.w6(32'hbc0a6396),
	.w7(32'hbc4880fc),
	.w8(32'hbc5c58be),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cb187),
	.w1(32'hbcb048bf),
	.w2(32'hbb5a2a92),
	.w3(32'h3d01ecfe),
	.w4(32'hbbf68f7a),
	.w5(32'hbb9aafeb),
	.w6(32'h3c8613c5),
	.w7(32'h3c83e948),
	.w8(32'h3a3018b2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a942cf3),
	.w1(32'h3bbeda6b),
	.w2(32'h3b42ae2c),
	.w3(32'h39df8924),
	.w4(32'hbb4153c5),
	.w5(32'h3c1f52e0),
	.w6(32'hbb83bc31),
	.w7(32'h3bb85534),
	.w8(32'hbb206b29),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d36e4),
	.w1(32'hbb267b3b),
	.w2(32'hbb028e2b),
	.w3(32'h3bf8c00c),
	.w4(32'hbc3cba73),
	.w5(32'h3afed3b3),
	.w6(32'h3bd12777),
	.w7(32'hbbeff354),
	.w8(32'hb9ad48b5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0949d1),
	.w1(32'h3c2519de),
	.w2(32'hb7787879),
	.w3(32'h3c47ba6e),
	.w4(32'h3cd8a5da),
	.w5(32'hbb86b701),
	.w6(32'hbb8bf41e),
	.w7(32'h3cc2e025),
	.w8(32'hbb904b96),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd93ab),
	.w1(32'h3bd9673d),
	.w2(32'h3be49e86),
	.w3(32'h3bd1dbfe),
	.w4(32'h3c1351f8),
	.w5(32'h3bc01fbc),
	.w6(32'h396cdc55),
	.w7(32'h3b9c89d3),
	.w8(32'h3aa15cef),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca65677),
	.w1(32'h3c0de12e),
	.w2(32'hbbada41d),
	.w3(32'h3ccac709),
	.w4(32'h3c409fb9),
	.w5(32'h3c047105),
	.w6(32'h3cc9c8cb),
	.w7(32'h3b126a18),
	.w8(32'h3c48dfe5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc88f),
	.w1(32'h3bb0145c),
	.w2(32'hbbfba503),
	.w3(32'hbcbb3d8a),
	.w4(32'hbb9d4528),
	.w5(32'hbc23834c),
	.w6(32'hbc5c62df),
	.w7(32'hbc6b7755),
	.w8(32'hbc16fa1c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c9b85),
	.w1(32'hbbf4062e),
	.w2(32'h3bbdc005),
	.w3(32'hbbb8c8b6),
	.w4(32'hbc27377c),
	.w5(32'h3bf5888d),
	.w6(32'h3aaff303),
	.w7(32'hbb6894be),
	.w8(32'h3c077756),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cdeb3),
	.w1(32'hbb77734f),
	.w2(32'h3bee9dee),
	.w3(32'h3bc13fd0),
	.w4(32'hbbd9300c),
	.w5(32'hbc034ac9),
	.w6(32'h3c06bc30),
	.w7(32'hbad1f5fe),
	.w8(32'hbbbbee47),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a92d9),
	.w1(32'hba2f4da9),
	.w2(32'h3bc2cdf5),
	.w3(32'hbbc7eded),
	.w4(32'hbc26b05e),
	.w5(32'h3bc0a203),
	.w6(32'hbba665a0),
	.w7(32'hbc04d211),
	.w8(32'h399b9af4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e2eaf),
	.w1(32'hbc18a9eb),
	.w2(32'h392a4c7b),
	.w3(32'h3ac2de7b),
	.w4(32'hbc290cde),
	.w5(32'h3a8f019d),
	.w6(32'h3c161ad7),
	.w7(32'hbb872e09),
	.w8(32'h39e24bdc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a320ad4),
	.w1(32'hb9908736),
	.w2(32'hbba9bc10),
	.w3(32'hbb5cdbe5),
	.w4(32'hbb5509ca),
	.w5(32'h3b90f763),
	.w6(32'hbbad44f7),
	.w7(32'hbc1639a8),
	.w8(32'hbb6f3f32),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07363),
	.w1(32'hbc5a8236),
	.w2(32'hbc58ed8a),
	.w3(32'h3c0c1c29),
	.w4(32'h3ac73927),
	.w5(32'hbc1696ef),
	.w6(32'h3c2447b3),
	.w7(32'hbada9ed5),
	.w8(32'hbc139b0f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394098),
	.w1(32'h3c0bd430),
	.w2(32'h3bc8f556),
	.w3(32'h3c815df2),
	.w4(32'h3c4bfb92),
	.w5(32'h3c01287c),
	.w6(32'h3c5c0f27),
	.w7(32'h3c3eddbf),
	.w8(32'h3c204a6d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f3fb6),
	.w1(32'hbbe38fe2),
	.w2(32'h3b9791a7),
	.w3(32'h3badd7e3),
	.w4(32'hbc12eac5),
	.w5(32'hba641c22),
	.w6(32'h3c04eb4d),
	.w7(32'hbb94904a),
	.w8(32'hbb412e10),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d62f0),
	.w1(32'h3c8beadc),
	.w2(32'h3b0edfc7),
	.w3(32'h3c9bc6f5),
	.w4(32'h3c838b9f),
	.w5(32'h3c087892),
	.w6(32'h3c6b9360),
	.w7(32'h3c13f688),
	.w8(32'hba99a012),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b361a80),
	.w1(32'hba7b6602),
	.w2(32'h3ca40220),
	.w3(32'hba8dea5b),
	.w4(32'h38ba4c4b),
	.w5(32'h3d2516a1),
	.w6(32'h3bd96ead),
	.w7(32'hbbcde9be),
	.w8(32'h3c8dad70),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72bf8),
	.w1(32'hbc5e9bab),
	.w2(32'hbb21b304),
	.w3(32'h3b40b9f7),
	.w4(32'hbc422f94),
	.w5(32'hbb491d02),
	.w6(32'h3cb1f4f3),
	.w7(32'hbc2ea279),
	.w8(32'hbbee902f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00320a),
	.w1(32'h3bb742a1),
	.w2(32'h3bae0c1e),
	.w3(32'h3afd8a64),
	.w4(32'h3c255fb8),
	.w5(32'h3bf891cd),
	.w6(32'hbb15d3fa),
	.w7(32'h3bfc3cbd),
	.w8(32'h3ba15aa3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6ba1f),
	.w1(32'h3b9fbc29),
	.w2(32'h3a351f3e),
	.w3(32'hbc6bfb9e),
	.w4(32'hbb1de8b7),
	.w5(32'h3c56f97a),
	.w6(32'hbb1a0536),
	.w7(32'hbc059a56),
	.w8(32'h3c8323d2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9efde7),
	.w1(32'h3b52fe21),
	.w2(32'h3bb69ed7),
	.w3(32'h3c67930e),
	.w4(32'hbbe546cd),
	.w5(32'h3c11c17e),
	.w6(32'h3c273981),
	.w7(32'hbb62b61a),
	.w8(32'h3c55fcab),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5828),
	.w1(32'hbc5df76d),
	.w2(32'h3b0441cc),
	.w3(32'h3c508b0d),
	.w4(32'hbc438ab8),
	.w5(32'h3b2db22c),
	.w6(32'h3c9f0310),
	.w7(32'hbb1bc4ec),
	.w8(32'h3b7866ee),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad83484),
	.w1(32'hbc3f3bd1),
	.w2(32'hbb15e671),
	.w3(32'h3c0bee0c),
	.w4(32'hbbccf736),
	.w5(32'h3c0fc125),
	.w6(32'h3c81688c),
	.w7(32'h3a915784),
	.w8(32'h3cec53f0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6487d5),
	.w1(32'hbc59dd39),
	.w2(32'h3bb4c1f6),
	.w3(32'hbc152533),
	.w4(32'hbc8d192f),
	.w5(32'h3b925cb6),
	.w6(32'h3b98e55c),
	.w7(32'hbca2f953),
	.w8(32'hbb6cca1d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31b8d2),
	.w1(32'hbbd53ae8),
	.w2(32'h3a02bf83),
	.w3(32'h3bff72d4),
	.w4(32'h3b09c81a),
	.w5(32'hb8c5d10d),
	.w6(32'h3bd498f1),
	.w7(32'hbb687a00),
	.w8(32'h3a5125ee),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc299b),
	.w1(32'hbb73b3b5),
	.w2(32'h39125440),
	.w3(32'h3b3cf9d8),
	.w4(32'h3a910d2e),
	.w5(32'h3b06237e),
	.w6(32'hbb6fb79f),
	.w7(32'hbb979b9b),
	.w8(32'hbc366156),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb899396),
	.w1(32'hba0ec48f),
	.w2(32'h3c22ad8f),
	.w3(32'hbbce0898),
	.w4(32'h3a6bb8d7),
	.w5(32'h3bb3fd4b),
	.w6(32'hbb131590),
	.w7(32'h3acbde19),
	.w8(32'hbc061c9e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9346e8),
	.w1(32'hbd1d24fb),
	.w2(32'hbb834738),
	.w3(32'h3d1e9728),
	.w4(32'hbd1d11ee),
	.w5(32'h3c2042c9),
	.w6(32'h3c56c301),
	.w7(32'hbcf0fda8),
	.w8(32'h3c3c4e5b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba694fa7),
	.w1(32'hbb454a7e),
	.w2(32'h3c0bc876),
	.w3(32'hbaaa51d4),
	.w4(32'hbb4ee6f7),
	.w5(32'hba99bdfd),
	.w6(32'hba57c5be),
	.w7(32'hba7683d3),
	.w8(32'hbc0e4bfc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c305971),
	.w1(32'hbbab236b),
	.w2(32'h3ae7ec92),
	.w3(32'h3c5fb51c),
	.w4(32'h3b2689d7),
	.w5(32'h3a7e7653),
	.w6(32'hbb259434),
	.w7(32'h3b92da96),
	.w8(32'hbc423f14),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8cf2a),
	.w1(32'hbc0a91ba),
	.w2(32'h3b9c9d91),
	.w3(32'h3c506019),
	.w4(32'hbc2dec46),
	.w5(32'h3b273002),
	.w6(32'h3c477b7c),
	.w7(32'hbb951292),
	.w8(32'h3b7f377d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9064f7),
	.w1(32'h3937b71c),
	.w2(32'h3b78f812),
	.w3(32'h3aee4136),
	.w4(32'hbb1a2141),
	.w5(32'h3bd1b664),
	.w6(32'h3b0942a0),
	.w7(32'h3a53e3db),
	.w8(32'h3c5c1c05),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada95b),
	.w1(32'hbc832998),
	.w2(32'hb983fa96),
	.w3(32'h3bc35cfe),
	.w4(32'hbc2d62fd),
	.w5(32'hb9814d35),
	.w6(32'h3bdd4e09),
	.w7(32'hbc41bf26),
	.w8(32'hbb590c8f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d484),
	.w1(32'h3aac6b4d),
	.w2(32'h3c9dbb00),
	.w3(32'h3aafe1ff),
	.w4(32'h3ae868b8),
	.w5(32'h3c9554c0),
	.w6(32'hba8218cc),
	.w7(32'hbae13a89),
	.w8(32'hbbe5dc5f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48f86e),
	.w1(32'hbd067922),
	.w2(32'h3bbff5b1),
	.w3(32'h3cfb42cd),
	.w4(32'hbd543816),
	.w5(32'hbbbcb56f),
	.w6(32'h3d277fc9),
	.w7(32'hbcd6d10b),
	.w8(32'h3a1484ae),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c18e03),
	.w1(32'hbcbd1799),
	.w2(32'hbc224e72),
	.w3(32'h3c09c571),
	.w4(32'hbc790cd8),
	.w5(32'h3a32d43e),
	.w6(32'h3c854e40),
	.w7(32'hba60c75e),
	.w8(32'h3c38c9be),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896f056),
	.w1(32'hbc432b49),
	.w2(32'hbafce772),
	.w3(32'h39383f3e),
	.w4(32'h3ac77d75),
	.w5(32'h3bed48ac),
	.w6(32'h3b927d03),
	.w7(32'h3c4b9f6a),
	.w8(32'h3c940a17),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baffc95),
	.w1(32'hbc0b50b6),
	.w2(32'hbb0b0da0),
	.w3(32'h3afe940b),
	.w4(32'hbc80c9fd),
	.w5(32'hbb9ed2b1),
	.w6(32'h3c00a58e),
	.w7(32'hbc803977),
	.w8(32'hbb2627b7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cf33a),
	.w1(32'hb72b3404),
	.w2(32'hbb85d621),
	.w3(32'hba5f326d),
	.w4(32'hbaa05376),
	.w5(32'h3c5bb092),
	.w6(32'hbc05722d),
	.w7(32'hbb48d9f0),
	.w8(32'h3bb5855a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8e29),
	.w1(32'h3bc5c751),
	.w2(32'hbc47ca0b),
	.w3(32'h3c028c43),
	.w4(32'h3c3563c9),
	.w5(32'hbc2ad02c),
	.w6(32'h3bf30bf3),
	.w7(32'h3c215ec6),
	.w8(32'hbb17f9cc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a5bd5),
	.w1(32'hbbc4224d),
	.w2(32'hbb6b2638),
	.w3(32'h3c4c8728),
	.w4(32'hbc5c995c),
	.w5(32'hbb5db699),
	.w6(32'h3c14ef64),
	.w7(32'hbb9e913d),
	.w8(32'hbbb7a409),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ddfb8),
	.w1(32'hbbaa26b6),
	.w2(32'hba4c3466),
	.w3(32'h3c396799),
	.w4(32'hbb48f365),
	.w5(32'h3c71a520),
	.w6(32'h3c598003),
	.w7(32'hbb31626f),
	.w8(32'h3ce4d911),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8892e),
	.w1(32'h3b7a59c5),
	.w2(32'hbb9dac6c),
	.w3(32'h3aacf142),
	.w4(32'h3bd1b285),
	.w5(32'h3c08f3c4),
	.w6(32'hbc1d6b14),
	.w7(32'hbca97e4d),
	.w8(32'hbbc78f4c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addc067),
	.w1(32'hbb405cde),
	.w2(32'hbc3d083d),
	.w3(32'h3c6d0b70),
	.w4(32'h3b81a912),
	.w5(32'h3aecfa0b),
	.w6(32'h3b598cec),
	.w7(32'hbc48ae6c),
	.w8(32'h3bb19334),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03d21b),
	.w1(32'h3c035c05),
	.w2(32'h3b9d79fe),
	.w3(32'h3c8eeec8),
	.w4(32'h3b1cccfe),
	.w5(32'h3abaec3d),
	.w6(32'h3d15cb64),
	.w7(32'hbbabd538),
	.w8(32'h3be94217),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67ac78),
	.w1(32'hbb3d6507),
	.w2(32'hb907d9ae),
	.w3(32'h3be47403),
	.w4(32'hbb42a950),
	.w5(32'h3b9faa1d),
	.w6(32'h3c9e5673),
	.w7(32'h3aff3c13),
	.w8(32'hbabb5e7d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c852f),
	.w1(32'hbb2f2e51),
	.w2(32'h3b43f5f5),
	.w3(32'hb81814b7),
	.w4(32'hba1a05bd),
	.w5(32'hbc5d61ba),
	.w6(32'hb9cf6b1e),
	.w7(32'hbb65561d),
	.w8(32'hbca66b8b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40092),
	.w1(32'h3b690115),
	.w2(32'h3c3d6e8d),
	.w3(32'hbbf8f848),
	.w4(32'h3cd75c29),
	.w5(32'h3cdea0c5),
	.w6(32'hbbc8f4c6),
	.w7(32'h3cb4380c),
	.w8(32'h3c34fbe8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c158),
	.w1(32'hbb5e0d3d),
	.w2(32'h3af5fbc1),
	.w3(32'hbc11a9bf),
	.w4(32'h3b7b4c29),
	.w5(32'h3c1cb5ac),
	.w6(32'hba06751e),
	.w7(32'hbb232c6c),
	.w8(32'h3c1a2661),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9cf3),
	.w1(32'h3c414a3a),
	.w2(32'h3be17e68),
	.w3(32'hbbb47e5d),
	.w4(32'h3bde8bc9),
	.w5(32'h3c9e6c99),
	.w6(32'hbc2ddd0b),
	.w7(32'h3980500f),
	.w8(32'h3c843102),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6cdf),
	.w1(32'h3c0630c6),
	.w2(32'h3bc03b12),
	.w3(32'hbc21a0d8),
	.w4(32'h3bd2ff8c),
	.w5(32'h3b2e046b),
	.w6(32'hbacdfbc8),
	.w7(32'h3c1e7f83),
	.w8(32'hbb5e9492),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48ed27),
	.w1(32'h3bb26236),
	.w2(32'h3d0a2e8b),
	.w3(32'h3baba0d4),
	.w4(32'h3a67dd84),
	.w5(32'h3cc0b306),
	.w6(32'hba614a8f),
	.w7(32'h3bedd42a),
	.w8(32'h3bae3a4f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb25019),
	.w1(32'hbcd1b8a5),
	.w2(32'h3b43e183),
	.w3(32'h3cc57150),
	.w4(32'hbcbc8043),
	.w5(32'h3c45b5c4),
	.w6(32'h3bbf1658),
	.w7(32'hbb6f80b1),
	.w8(32'hb90024d3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d112),
	.w1(32'hbc340cc0),
	.w2(32'hbc15da58),
	.w3(32'h3c095f3d),
	.w4(32'hbbc1a1ba),
	.w5(32'hbb525ff5),
	.w6(32'h3ba3323f),
	.w7(32'h3bb13677),
	.w8(32'h3b17de69),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2578db),
	.w1(32'hbc698184),
	.w2(32'h3a225e49),
	.w3(32'h3be1be92),
	.w4(32'hbc4ce00b),
	.w5(32'hbad8bf12),
	.w6(32'hbbf24034),
	.w7(32'hbca734e2),
	.w8(32'h3ab01314),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85de37),
	.w1(32'h3be8603a),
	.w2(32'h3a5f2ddf),
	.w3(32'hba451016),
	.w4(32'h3bd5c4e7),
	.w5(32'hbac518ed),
	.w6(32'hbb90d063),
	.w7(32'hba05d306),
	.w8(32'hbbe26da6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e2801),
	.w1(32'hba9bf2df),
	.w2(32'h3b7a19d5),
	.w3(32'hbb694568),
	.w4(32'hbb93a5b9),
	.w5(32'h3abd6ed1),
	.w6(32'hbbff9406),
	.w7(32'hbbd77ab7),
	.w8(32'hbc078174),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab32512),
	.w1(32'hba82d8dc),
	.w2(32'h3bb1df21),
	.w3(32'hba1ba5ce),
	.w4(32'h3b85f107),
	.w5(32'hbb3e76d9),
	.w6(32'hbc10f97d),
	.w7(32'h3b555ce1),
	.w8(32'hbc785afb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0019),
	.w1(32'h397f5be3),
	.w2(32'hbc801a94),
	.w3(32'h3a96eaa1),
	.w4(32'h3b986f83),
	.w5(32'hbc78fd4a),
	.w6(32'h3b971391),
	.w7(32'h3c2900d7),
	.w8(32'h3b18979b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c596fc1),
	.w1(32'h3addf089),
	.w2(32'hbc26e726),
	.w3(32'h3c9c8454),
	.w4(32'hbc0420cb),
	.w5(32'hbc425eee),
	.w6(32'h3c3d0f6e),
	.w7(32'hba93ce76),
	.w8(32'hbc914d84),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1e9f6),
	.w1(32'hbbca4ea6),
	.w2(32'h3b01a3f1),
	.w3(32'h3b9a593b),
	.w4(32'hbba4aa23),
	.w5(32'h3c278bc1),
	.w6(32'h3aa622dd),
	.w7(32'h3b8be472),
	.w8(32'h39361994),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90f8ea),
	.w1(32'h3b0c22a8),
	.w2(32'h3c354064),
	.w3(32'h3a1929a6),
	.w4(32'hbab6bdce),
	.w5(32'h3c1cf97b),
	.w6(32'hbb6f3815),
	.w7(32'hbb646ba5),
	.w8(32'hbad0a77e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6968f),
	.w1(32'hbb92d984),
	.w2(32'hb89100d1),
	.w3(32'h3bbd2246),
	.w4(32'hbad12ed9),
	.w5(32'h3a868ef0),
	.w6(32'hbbaa1d8b),
	.w7(32'h3b346ba4),
	.w8(32'h3aa8c8e5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba555b92),
	.w1(32'h3a9984f0),
	.w2(32'hbad1e204),
	.w3(32'hbb388cb9),
	.w4(32'hb93e0503),
	.w5(32'hba83a7bc),
	.w6(32'hbb64ac4e),
	.w7(32'hbb42e22f),
	.w8(32'h39227372),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89718b),
	.w1(32'h3c4e0bfa),
	.w2(32'h3c697be4),
	.w3(32'h3c71a25b),
	.w4(32'h3b56509c),
	.w5(32'h3c944250),
	.w6(32'h3c0f757e),
	.w7(32'hbaaa8f8e),
	.w8(32'hba15d198),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897675),
	.w1(32'h3c0bd48f),
	.w2(32'hba4b7bb3),
	.w3(32'h3c4823aa),
	.w4(32'h3c6d467f),
	.w5(32'h3c93c9ff),
	.w6(32'h3ccdffbb),
	.w7(32'h3ab99fda),
	.w8(32'h3cbc4585),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa24e4),
	.w1(32'hba7a7901),
	.w2(32'h3c0d9e49),
	.w3(32'h3bc8c001),
	.w4(32'h3b3816ee),
	.w5(32'h3c53d1b3),
	.w6(32'h3c90d2a5),
	.w7(32'h3bea9431),
	.w8(32'h3c22c19f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362efe),
	.w1(32'hbca44b3e),
	.w2(32'hbbc00ee4),
	.w3(32'h3c2ed2c7),
	.w4(32'hbc2a1ca9),
	.w5(32'h3b5c85ea),
	.w6(32'h3cb89b45),
	.w7(32'h3b88bb5e),
	.w8(32'h3cb50c6f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3e8a6),
	.w1(32'h3b574c89),
	.w2(32'hbbfea8a9),
	.w3(32'hbb23241e),
	.w4(32'h3b10b5a2),
	.w5(32'hbb8042e4),
	.w6(32'hbb1f5921),
	.w7(32'h3b160455),
	.w8(32'hba9bb20b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe74c),
	.w1(32'h3ad701d4),
	.w2(32'hbc689bd4),
	.w3(32'h3b085107),
	.w4(32'hb904cddb),
	.w5(32'hbbd65c4f),
	.w6(32'h3ae3d2d3),
	.w7(32'hbc27e614),
	.w8(32'h3aa10d23),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69bf0c),
	.w1(32'h3c952503),
	.w2(32'hba6c95bc),
	.w3(32'h3b7823cf),
	.w4(32'h3bbe7b8f),
	.w5(32'h3a376fa0),
	.w6(32'h3ca12932),
	.w7(32'hbc368450),
	.w8(32'h3b95acaa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e65f),
	.w1(32'hbc7453f0),
	.w2(32'hbb7e75eb),
	.w3(32'hbb8a9a1d),
	.w4(32'hba91f7bf),
	.w5(32'hba2a0517),
	.w6(32'hbc7426f7),
	.w7(32'h3bd97133),
	.w8(32'hbb646a07),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba341699),
	.w1(32'hbb6d700d),
	.w2(32'h3b41af91),
	.w3(32'h3a324486),
	.w4(32'hbafbabfa),
	.w5(32'hbb9fe69e),
	.w6(32'hba704419),
	.w7(32'hbb84ef23),
	.w8(32'hbb639e4d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11248f),
	.w1(32'h3c5835cb),
	.w2(32'h3ca91184),
	.w3(32'h3ad66757),
	.w4(32'h3c16502e),
	.w5(32'h3c91e26e),
	.w6(32'h3b7eb8e8),
	.w7(32'h3b1bde11),
	.w8(32'h3c2089d6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed790),
	.w1(32'hbb8f6fdd),
	.w2(32'h3c8a96c8),
	.w3(32'h3b1640bc),
	.w4(32'h3c2008dc),
	.w5(32'h3c756613),
	.w6(32'hb88c0e6a),
	.w7(32'h3c2e5f6c),
	.w8(32'h3c3e6401),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5d1c),
	.w1(32'hbcc5b087),
	.w2(32'hbc307ae3),
	.w3(32'hba7c5ef3),
	.w4(32'hbc389840),
	.w5(32'hbb69a5c9),
	.w6(32'hbc8b15be),
	.w7(32'hb9efb816),
	.w8(32'h3b856bc2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60b79),
	.w1(32'h3c25353b),
	.w2(32'h3bba6e2a),
	.w3(32'h3c1029b6),
	.w4(32'hbbb9d969),
	.w5(32'h3ae76a60),
	.w6(32'h3c9fc30f),
	.w7(32'hbc2c83ef),
	.w8(32'h3b8f7772),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3d516),
	.w1(32'h3b9fb7fa),
	.w2(32'h3b16ba35),
	.w3(32'h3b324015),
	.w4(32'h3b13c1e0),
	.w5(32'h3bbace9a),
	.w6(32'h3b160af7),
	.w7(32'h3ac576a2),
	.w8(32'hba5c2379),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dbb0c),
	.w1(32'h39f40e7b),
	.w2(32'h39aff6ab),
	.w3(32'hbb248d5e),
	.w4(32'hba4d10b0),
	.w5(32'h3b061515),
	.w6(32'h3c0b9cc2),
	.w7(32'hbb5885b8),
	.w8(32'h3afe67eb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e5075),
	.w1(32'hbb160281),
	.w2(32'h3c91d3f9),
	.w3(32'hba8a455e),
	.w4(32'hbb9813f9),
	.w5(32'h3c57c5ce),
	.w6(32'hba9f4c99),
	.w7(32'hbbb1a230),
	.w8(32'hbc12c44f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc906844),
	.w1(32'hbbb1845e),
	.w2(32'hbbeed65d),
	.w3(32'h3ba22d26),
	.w4(32'hbbe75064),
	.w5(32'hbbaaaf55),
	.w6(32'h3d05a7ce),
	.w7(32'h3bd5acb2),
	.w8(32'hbc2aa5a6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc048aa6),
	.w1(32'h3b46338a),
	.w2(32'hbc67347b),
	.w3(32'h370740c8),
	.w4(32'hb953b596),
	.w5(32'hbc21b848),
	.w6(32'h3b84f540),
	.w7(32'h3b81b69a),
	.w8(32'hb8931d34),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88355d),
	.w1(32'h3c5d93f3),
	.w2(32'hbc747928),
	.w3(32'h3c3e3ec4),
	.w4(32'h3bac04ff),
	.w5(32'h3baaf8d6),
	.w6(32'h3c80802d),
	.w7(32'hbbc348ac),
	.w8(32'h3ca279b0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1575d3),
	.w1(32'h3c2ea26a),
	.w2(32'hba9da546),
	.w3(32'hbc3a981e),
	.w4(32'h3c6241f6),
	.w5(32'h395e0d72),
	.w6(32'hbc6e6aa0),
	.w7(32'h3bcb46dc),
	.w8(32'hbab2c6d8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf32bd8),
	.w1(32'h3b31c1e8),
	.w2(32'hb9f7d218),
	.w3(32'h3c3b0fbc),
	.w4(32'hb883fb47),
	.w5(32'h3ac53de8),
	.w6(32'h3c2bb074),
	.w7(32'hbb510558),
	.w8(32'h3bd46e3c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff6c6d),
	.w1(32'hba9d5cd8),
	.w2(32'h3b838fc4),
	.w3(32'h39d5aa3a),
	.w4(32'h3aca6ae4),
	.w5(32'h3cc21275),
	.w6(32'hb9ce4e2c),
	.w7(32'hba5734ad),
	.w8(32'h3cc94db5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f3a1),
	.w1(32'h3bbe5a32),
	.w2(32'hbbd1563c),
	.w3(32'hbc0bf626),
	.w4(32'h3c3c548f),
	.w5(32'h3bd58845),
	.w6(32'h3b1aa918),
	.w7(32'h3b8cc1be),
	.w8(32'h3c08e2bf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c550c0d),
	.w1(32'hba231ae6),
	.w2(32'h3c047850),
	.w3(32'h3cd9845a),
	.w4(32'h3baaafd3),
	.w5(32'h3baf3e40),
	.w6(32'h3cc4ffb2),
	.w7(32'h3c06b069),
	.w8(32'hbb66d6da),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90e3da),
	.w1(32'hbc3aa91a),
	.w2(32'h3ba53bba),
	.w3(32'h3a855509),
	.w4(32'hbbb3a815),
	.w5(32'h3c1baace),
	.w6(32'hbbedc596),
	.w7(32'hbb84334a),
	.w8(32'hba8449ed),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb533b2),
	.w1(32'h3c93e7d0),
	.w2(32'h3c056d9d),
	.w3(32'h3c808bbb),
	.w4(32'h3c4ea1c5),
	.w5(32'h3b1a0f3c),
	.w6(32'h3b4bb928),
	.w7(32'h3c342b4b),
	.w8(32'hba205698),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade32df),
	.w1(32'hbc2d68ec),
	.w2(32'h39987d52),
	.w3(32'h3b2f056e),
	.w4(32'hbb856e52),
	.w5(32'h3b17b5e7),
	.w6(32'h3ba85c00),
	.w7(32'h3b7e88dd),
	.w8(32'h3bb945d2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0930d2),
	.w1(32'h3a5f6085),
	.w2(32'h3c8b598d),
	.w3(32'h3c040d5a),
	.w4(32'hbb0db251),
	.w5(32'h3c426eb8),
	.w6(32'h3c504e3b),
	.w7(32'h3b31440b),
	.w8(32'h3baf2737),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83d112),
	.w1(32'h3bd01dbf),
	.w2(32'h3bed27a1),
	.w3(32'hbb3138d1),
	.w4(32'h3b8ba0e4),
	.w5(32'hbb1d4f38),
	.w6(32'hb9b42cac),
	.w7(32'h3b01926a),
	.w8(32'hbc0c088c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552b01),
	.w1(32'h3be69664),
	.w2(32'hbaa9f514),
	.w3(32'hbb2eaa5a),
	.w4(32'h3ce65a46),
	.w5(32'h3c5665c2),
	.w6(32'hbc4f78e7),
	.w7(32'h3cb893fc),
	.w8(32'h3bf53a3e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0845ec),
	.w1(32'hbbafe09c),
	.w2(32'hbc4f464c),
	.w3(32'hbb861788),
	.w4(32'hbb87cb4c),
	.w5(32'hbc917b0d),
	.w6(32'h3b5cacd5),
	.w7(32'h3988a8b9),
	.w8(32'hbbc5578d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc579c),
	.w1(32'hbc0f159e),
	.w2(32'h3ca4ab7d),
	.w3(32'h3d159960),
	.w4(32'hbc0b1436),
	.w5(32'h3cc5acc1),
	.w6(32'h3cfe21ef),
	.w7(32'h3bfb6700),
	.w8(32'h3c50c200),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c156),
	.w1(32'hbc405e4c),
	.w2(32'h3c4ded60),
	.w3(32'hbb5bdbf8),
	.w4(32'hbb3e3bc5),
	.w5(32'h3c5e79db),
	.w6(32'hba40c99a),
	.w7(32'h3c2ebed0),
	.w8(32'h3c18f9f4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceefe9a),
	.w1(32'h3b5ce5d6),
	.w2(32'hbae6268e),
	.w3(32'h3cadfe10),
	.w4(32'hbbbde1ca),
	.w5(32'hbc64a313),
	.w6(32'h3c3a0436),
	.w7(32'hbbd86fdb),
	.w8(32'hbb8930ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464ff2),
	.w1(32'hbc8f93d0),
	.w2(32'h3c007fc6),
	.w3(32'h3c9a010d),
	.w4(32'hbbe2b2f9),
	.w5(32'h3c090964),
	.w6(32'h3b9fdedf),
	.w7(32'h3c6734c9),
	.w8(32'h3c0311ad),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a25d3),
	.w1(32'hbcc67ae0),
	.w2(32'hbb293f94),
	.w3(32'h3c504c83),
	.w4(32'h3b0ea08a),
	.w5(32'h3c2bc95d),
	.w6(32'hbb54ce1e),
	.w7(32'h3b47f1ec),
	.w8(32'h3c82cbdf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad2c3b),
	.w1(32'h3c6a116c),
	.w2(32'h3c0eac32),
	.w3(32'h3c864982),
	.w4(32'h3c06bc5b),
	.w5(32'h3c1ecffa),
	.w6(32'h3c0529e1),
	.w7(32'h3925da87),
	.w8(32'h3acd8053),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7fe0e),
	.w1(32'h3ad6035b),
	.w2(32'hbb337efa),
	.w3(32'hbb43f765),
	.w4(32'h3acf5c0b),
	.w5(32'h3bf9fd26),
	.w6(32'hbb5b6ef7),
	.w7(32'hba9de5e8),
	.w8(32'h3cb6fbdb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cedf461),
	.w1(32'h3cc4f2af),
	.w2(32'h3be33e8e),
	.w3(32'h3c9bf082),
	.w4(32'h3bf2a6fe),
	.w5(32'h3c134ef2),
	.w6(32'h3c216b99),
	.w7(32'hbc51b173),
	.w8(32'h3bf1f067),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe4618),
	.w1(32'hbbb81272),
	.w2(32'h39499d6a),
	.w3(32'hbc12c23b),
	.w4(32'hbb65b25e),
	.w5(32'h3bcefe33),
	.w6(32'hbbc69d39),
	.w7(32'hbc0b983a),
	.w8(32'h3c455fe2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8931b9b),
	.w1(32'h3b674b28),
	.w2(32'hbc4ca15c),
	.w3(32'hbb61f1c7),
	.w4(32'h3af32fdc),
	.w5(32'hbc43d685),
	.w6(32'hbb6e409b),
	.w7(32'hbbd630ab),
	.w8(32'hbada5310),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e556),
	.w1(32'h3c00659e),
	.w2(32'hbc3ece01),
	.w3(32'h3c31da4b),
	.w4(32'hb8c71b63),
	.w5(32'hbbc131fe),
	.w6(32'h3bd6c4b9),
	.w7(32'h3aa267b9),
	.w8(32'h3afe8278),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c454b91),
	.w1(32'hbc990be0),
	.w2(32'h3b1ddc03),
	.w3(32'h3c0f069f),
	.w4(32'hbc88fc29),
	.w5(32'h3b0bdc9e),
	.w6(32'h3c6642a3),
	.w7(32'hbca40560),
	.w8(32'hbbfeafb7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14aaf7),
	.w1(32'hbca06643),
	.w2(32'hbc01f7f9),
	.w3(32'h3c985ae5),
	.w4(32'hbbebdb1e),
	.w5(32'hbbbbd0e2),
	.w6(32'h3bfecbe7),
	.w7(32'h3bc09744),
	.w8(32'h3bdc742d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5d0bc),
	.w1(32'hbbdae3c2),
	.w2(32'hbbf8e2fc),
	.w3(32'h3c39fe2c),
	.w4(32'hbc18c3e4),
	.w5(32'h3c1ffbc5),
	.w6(32'hbb064721),
	.w7(32'hbbc7a4f9),
	.w8(32'h3c92868b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ab11),
	.w1(32'h3bd76499),
	.w2(32'h3bf4a174),
	.w3(32'hbb9ea443),
	.w4(32'hbaf3b115),
	.w5(32'h3b995a4e),
	.w6(32'h3be37e7d),
	.w7(32'hbc2528ef),
	.w8(32'hbb495e54),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96102e),
	.w1(32'hbc6f28dd),
	.w2(32'hbbe3e669),
	.w3(32'h3c395b0a),
	.w4(32'hbbf2dfc5),
	.w5(32'hbc875c1a),
	.w6(32'h3cf007bb),
	.w7(32'hb9b16ebf),
	.w8(32'hbc819637),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb52c6c),
	.w1(32'h3b8db8d2),
	.w2(32'h3bcb005d),
	.w3(32'h3cabd842),
	.w4(32'hbbc7183a),
	.w5(32'h3bbfa58e),
	.w6(32'h3c203056),
	.w7(32'hbac557c2),
	.w8(32'h3c121d35),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6bc21),
	.w1(32'hbc825da8),
	.w2(32'hba5f2684),
	.w3(32'h3c6d50c1),
	.w4(32'hbbff5263),
	.w5(32'hbaf149db),
	.w6(32'h3bbde77a),
	.w7(32'h3b463cfa),
	.w8(32'hbab0734a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28c5b9),
	.w1(32'hbb836e09),
	.w2(32'h3a1b5b02),
	.w3(32'hbb1b6f3e),
	.w4(32'hbb72ea2f),
	.w5(32'hbabdcdd9),
	.w6(32'hba99cc9c),
	.w7(32'h3af3e725),
	.w8(32'h3b611217),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93663d),
	.w1(32'h39a126fc),
	.w2(32'h3a48030f),
	.w3(32'hba2b657d),
	.w4(32'hbba930be),
	.w5(32'hba3949f2),
	.w6(32'h3b6489c9),
	.w7(32'h3ac5c24f),
	.w8(32'hbaedd289),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3657e),
	.w1(32'h3abbc825),
	.w2(32'h3c9dadf0),
	.w3(32'h3a08f0e6),
	.w4(32'hbafc48d5),
	.w5(32'h3c9d1700),
	.w6(32'hba3a0f76),
	.w7(32'h3af1bf27),
	.w8(32'h3ba2ef30),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcb773),
	.w1(32'hbc237bd3),
	.w2(32'h3bff4e3c),
	.w3(32'hbc113c42),
	.w4(32'hbba4f7ca),
	.w5(32'hbb33a30d),
	.w6(32'hbc73cdd6),
	.w7(32'h39eb03e0),
	.w8(32'hbc736fa0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079348),
	.w1(32'hbb9c1202),
	.w2(32'hbb095407),
	.w3(32'h3bc7c5ea),
	.w4(32'hbc134417),
	.w5(32'hbc178c60),
	.w6(32'hbbb187a5),
	.w7(32'h3c09ea50),
	.w8(32'h3a980fd8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0b53b),
	.w1(32'hb9ced8e1),
	.w2(32'h3a8eb0cd),
	.w3(32'hbb8a6743),
	.w4(32'hb9c4cf1b),
	.w5(32'hba6b2d3b),
	.w6(32'hbae24733),
	.w7(32'h3c51dbfe),
	.w8(32'hbaa7b1c3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2db95),
	.w1(32'h3a54ea14),
	.w2(32'h39083a05),
	.w3(32'h3b63cae5),
	.w4(32'h3aeace04),
	.w5(32'hbb01e4fe),
	.w6(32'hbaefdfc7),
	.w7(32'hbb1879c4),
	.w8(32'hbb88275b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c1191),
	.w1(32'hbba9ad7c),
	.w2(32'h3c21d52b),
	.w3(32'hbaadce0a),
	.w4(32'hbbcc7023),
	.w5(32'h3c078fd9),
	.w6(32'h3b0ecf1e),
	.w7(32'hbb7f01f2),
	.w8(32'hbb17cdba),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21d8b4),
	.w1(32'h3ac9d17e),
	.w2(32'h3b3f116c),
	.w3(32'h3ba6c23f),
	.w4(32'hbb9e919f),
	.w5(32'h3af1a6f1),
	.w6(32'h3c68db38),
	.w7(32'hbc1f1249),
	.w8(32'hba387ee7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a24e3),
	.w1(32'h3b7347fc),
	.w2(32'h3c03f134),
	.w3(32'hb9dcabc2),
	.w4(32'h3b2e3029),
	.w5(32'h3c852e08),
	.w6(32'hbab0d108),
	.w7(32'h3a078034),
	.w8(32'h3c89f935),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92097d),
	.w1(32'h3c05fa8d),
	.w2(32'hbbe97110),
	.w3(32'hbca907ac),
	.w4(32'h3bcd4d8b),
	.w5(32'h3c080fd1),
	.w6(32'hbb6de278),
	.w7(32'hbbbe8110),
	.w8(32'h3c567d05),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74ca7e),
	.w1(32'h3c9df020),
	.w2(32'hbc039657),
	.w3(32'hbbd936e8),
	.w4(32'h3b14e042),
	.w5(32'h3be79666),
	.w6(32'h3c947f5d),
	.w7(32'hbc97221d),
	.w8(32'h3b639c57),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe697a1),
	.w1(32'h3cb74bfe),
	.w2(32'h39f3d9d9),
	.w3(32'hbac72680),
	.w4(32'h3c4f5095),
	.w5(32'h3c5e3c0e),
	.w6(32'h3b993c73),
	.w7(32'hbc07a7df),
	.w8(32'h3b58d658),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ff24b),
	.w1(32'hbad14e5e),
	.w2(32'hbc1b8c46),
	.w3(32'h3c76028a),
	.w4(32'hbcacec72),
	.w5(32'hbaa001c1),
	.w6(32'h3c8ecb4b),
	.w7(32'hbc56fc5b),
	.w8(32'hbb3794bf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6920),
	.w1(32'h3ca23707),
	.w2(32'h3b0bc927),
	.w3(32'h3b03193c),
	.w4(32'h3d247dc2),
	.w5(32'h3b29f5c2),
	.w6(32'h3b30772c),
	.w7(32'h3d24c6f1),
	.w8(32'hbc51e684),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ec012),
	.w1(32'hbbcbfbaa),
	.w2(32'hbb0e02d6),
	.w3(32'h3bfa8d93),
	.w4(32'h3c05dffc),
	.w5(32'hbc5b98d1),
	.w6(32'h3a820862),
	.w7(32'h3bdea1da),
	.w8(32'hbb18c048),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ea7b),
	.w1(32'hbb2d6d4e),
	.w2(32'h3c3be456),
	.w3(32'h3bea4bea),
	.w4(32'hbb3f15ca),
	.w5(32'h3b9e4fbd),
	.w6(32'hb8c69a6c),
	.w7(32'h3b3bc51a),
	.w8(32'hbbfe03b1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff0729),
	.w1(32'h3b2d559e),
	.w2(32'hbc3bf187),
	.w3(32'h3b552e89),
	.w4(32'h3bb670bf),
	.w5(32'hbb142175),
	.w6(32'hbc0ed621),
	.w7(32'h3c27d28a),
	.w8(32'h3cac6f86),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf02132),
	.w1(32'hbb88861f),
	.w2(32'h3b4974de),
	.w3(32'h3bee88ee),
	.w4(32'h3b946e3e),
	.w5(32'h3b1299d7),
	.w6(32'hbc8b784c),
	.w7(32'hbbdc20e7),
	.w8(32'hb95a75c5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06c6cd),
	.w1(32'h3b886944),
	.w2(32'h3c8f9b7e),
	.w3(32'h3bfa1a89),
	.w4(32'h3b5836b9),
	.w5(32'h3c8b1f9a),
	.w6(32'h3c001522),
	.w7(32'hbad4393e),
	.w8(32'hbb043efe),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b440e95),
	.w1(32'hbb54cac4),
	.w2(32'hbc07b96e),
	.w3(32'h3a605202),
	.w4(32'hbbace6f3),
	.w5(32'hbbb61d96),
	.w6(32'hbb14fe34),
	.w7(32'hbabdafc5),
	.w8(32'h3bddc989),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73b49b),
	.w1(32'h3b8b88bb),
	.w2(32'h3c5b1e94),
	.w3(32'h3c176e64),
	.w4(32'hbbb8de9f),
	.w5(32'h3b2dd30e),
	.w6(32'h3ba4e3cb),
	.w7(32'hba8b5e38),
	.w8(32'hbaf91330),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e015),
	.w1(32'h3b407683),
	.w2(32'h3bc2504a),
	.w3(32'h3c7fbb6e),
	.w4(32'h3c25b8c3),
	.w5(32'h3c1d7929),
	.w6(32'h3a96be9a),
	.w7(32'h3bbf3155),
	.w8(32'h3b2c3b33),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ebf3),
	.w1(32'hbb3f8c8a),
	.w2(32'hbb56ad31),
	.w3(32'h3b8c3314),
	.w4(32'hbafb81cf),
	.w5(32'hbc2e4c69),
	.w6(32'h3c187f3f),
	.w7(32'h3b76c4be),
	.w8(32'hbb748747),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99c9dd),
	.w1(32'h3b1103cd),
	.w2(32'h3bfb7c20),
	.w3(32'h3c20301a),
	.w4(32'hba86b739),
	.w5(32'h3b9fd5d4),
	.w6(32'h3bec41cf),
	.w7(32'hbb0e99bd),
	.w8(32'h3b43e0d5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb8f89),
	.w1(32'hbaf8ee8d),
	.w2(32'hbb0845bb),
	.w3(32'h3821bed2),
	.w4(32'hbafc00a8),
	.w5(32'h3bbb42b4),
	.w6(32'hb939ccac),
	.w7(32'h39fb8f48),
	.w8(32'h3b069cb7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bf8e4),
	.w1(32'hbc3c1dc8),
	.w2(32'h3c0a2fdd),
	.w3(32'h3bd54645),
	.w4(32'h3b54f814),
	.w5(32'h3bf589d3),
	.w6(32'h3bc32204),
	.w7(32'h3b325a53),
	.w8(32'h3b9e5de5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33570f),
	.w1(32'hbb9818fd),
	.w2(32'hbae0a92b),
	.w3(32'h3c374847),
	.w4(32'h3c6fea21),
	.w5(32'hbb5413d3),
	.w6(32'hb9bdeef8),
	.w7(32'h3ca1ae8a),
	.w8(32'h39c55914),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72e8d1a),
	.w1(32'h39afa68a),
	.w2(32'hba373d52),
	.w3(32'hba5c2ff1),
	.w4(32'hba5f5020),
	.w5(32'hbab37b73),
	.w6(32'hbb17deff),
	.w7(32'h3ab222f9),
	.w8(32'h38a2efcc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5063eb),
	.w1(32'hba8e33a6),
	.w2(32'h3b1c818b),
	.w3(32'hbb750711),
	.w4(32'hbb441e91),
	.w5(32'h3a1fe527),
	.w6(32'hba80458f),
	.w7(32'hbab50044),
	.w8(32'h3aeabf4a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6529c),
	.w1(32'hbaa601fd),
	.w2(32'h3b5cf9fd),
	.w3(32'h3ae8412e),
	.w4(32'h3ad7434f),
	.w5(32'h3b6092cc),
	.w6(32'h3b2af836),
	.w7(32'hbaf66b70),
	.w8(32'hba03a200),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc0f56),
	.w1(32'hbbb57a2c),
	.w2(32'hbc5d424b),
	.w3(32'h3bad70a1),
	.w4(32'hbb7f433f),
	.w5(32'hbc024806),
	.w6(32'h3c1b165d),
	.w7(32'hbb44523b),
	.w8(32'h3bf1ca2f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c832174),
	.w1(32'hbc0a7c63),
	.w2(32'h3ae51026),
	.w3(32'h3c678a0f),
	.w4(32'hbbd4746e),
	.w5(32'h3bb3cc9c),
	.w6(32'h3c659d00),
	.w7(32'hbb2ee2ba),
	.w8(32'h3bf9f47c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69ed0),
	.w1(32'h3ab95cac),
	.w2(32'hbc539f02),
	.w3(32'hbb9c3cdd),
	.w4(32'h3b64f229),
	.w5(32'hbc7302b0),
	.w6(32'hbaef54e3),
	.w7(32'h3b20ad00),
	.w8(32'hbb9afd10),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c853f04),
	.w1(32'hbaab3e68),
	.w2(32'h3b2eb820),
	.w3(32'h3ccd05bc),
	.w4(32'hbbff1db3),
	.w5(32'hbb53c0ec),
	.w6(32'h3cb970e6),
	.w7(32'h3b876619),
	.w8(32'hbb18a143),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260af8),
	.w1(32'hbc061f4a),
	.w2(32'hba836cc1),
	.w3(32'h3b9e098a),
	.w4(32'hbc62e519),
	.w5(32'hbb80350d),
	.w6(32'h3beb83f3),
	.w7(32'hbb5f3701),
	.w8(32'h3aa17bdf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2883ec),
	.w1(32'h3b3da0f5),
	.w2(32'h3c1c29e6),
	.w3(32'h3b726312),
	.w4(32'hbb185d38),
	.w5(32'h3c714d7d),
	.w6(32'hbaca0513),
	.w7(32'hbb51c398),
	.w8(32'h3adc41e4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cdf52),
	.w1(32'hbb2e1c4f),
	.w2(32'hbbfb5dbc),
	.w3(32'h3b982c94),
	.w4(32'h3b71e574),
	.w5(32'hbb5a13c3),
	.w6(32'h3c056f33),
	.w7(32'h3adc66af),
	.w8(32'h3bbc41a6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44df4e),
	.w1(32'h39d898dd),
	.w2(32'h3c20ee27),
	.w3(32'hbc14c46f),
	.w4(32'h3ca5b973),
	.w5(32'h3c3f162a),
	.w6(32'hbc362270),
	.w7(32'h3bffad95),
	.w8(32'h3c1f7ef6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7caca),
	.w1(32'hbb9b1c5c),
	.w2(32'h38d9b2fd),
	.w3(32'hbc5d0c43),
	.w4(32'hb9fccd23),
	.w5(32'h3a8044b1),
	.w6(32'hbbb436c4),
	.w7(32'h3b9be67c),
	.w8(32'h390633fc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af3f6a),
	.w1(32'hbbe3275f),
	.w2(32'hbb36a144),
	.w3(32'h3b8dbf6b),
	.w4(32'hbb04c849),
	.w5(32'h3a875956),
	.w6(32'h3bc20615),
	.w7(32'hba110766),
	.w8(32'h3b994fc6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf5871),
	.w1(32'hbb3d5d54),
	.w2(32'h3c1d551b),
	.w3(32'h3b50d642),
	.w4(32'h3b7eb35b),
	.w5(32'h3ab34570),
	.w6(32'h3b97bc9b),
	.w7(32'hb997b395),
	.w8(32'h38c8163c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a303b5d),
	.w1(32'hbc828a2f),
	.w2(32'hbafd960e),
	.w3(32'h3c19ca32),
	.w4(32'h3b0f0d80),
	.w5(32'hbae0fc92),
	.w6(32'h3bc3b5f6),
	.w7(32'h3bd0c5ec),
	.w8(32'h3a9db23d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f512bf),
	.w1(32'h39d6d583),
	.w2(32'hbb87e276),
	.w3(32'h392cabb1),
	.w4(32'hba21d270),
	.w5(32'h3a8420f4),
	.w6(32'h3ac225a8),
	.w7(32'h3b04a1c9),
	.w8(32'h3b564764),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc163de),
	.w1(32'h3a94dc74),
	.w2(32'h3b5fdd40),
	.w3(32'h3afafae0),
	.w4(32'h3b7f3b2b),
	.w5(32'hbb966c4d),
	.w6(32'h3bc6b681),
	.w7(32'h3ae26baa),
	.w8(32'hbb102541),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c4b1f),
	.w1(32'h3b2b6734),
	.w2(32'h3afd893d),
	.w3(32'h3c05b74c),
	.w4(32'h3a264a0e),
	.w5(32'hbb3209db),
	.w6(32'h3c08ca2f),
	.w7(32'h3b092382),
	.w8(32'hba78efd0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81683a),
	.w1(32'hb8e7eba0),
	.w2(32'h3b8ae94b),
	.w3(32'hbbd55a9d),
	.w4(32'hbb101569),
	.w5(32'h3a9fdeaa),
	.w6(32'hbb391a3a),
	.w7(32'h3ab79e12),
	.w8(32'hbb71ffd8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ff44b),
	.w1(32'h39a95356),
	.w2(32'hbb6553b6),
	.w3(32'h3c00c3f3),
	.w4(32'hbbff6814),
	.w5(32'h3ae58300),
	.w6(32'hb902f7d2),
	.w7(32'hbbd573f0),
	.w8(32'h3af73043),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ccc87),
	.w1(32'hbb37e272),
	.w2(32'h3b3f6af6),
	.w3(32'hbabfb246),
	.w4(32'hbb1b4103),
	.w5(32'h3a59a2c2),
	.w6(32'hbb0b5a8e),
	.w7(32'hbb5c0ade),
	.w8(32'h3c130faa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeedf4b),
	.w1(32'hbbccf745),
	.w2(32'hb9f243da),
	.w3(32'hbc275b9b),
	.w4(32'hbca99b65),
	.w5(32'hbb352a01),
	.w6(32'hba35c9c1),
	.w7(32'h3bcf30b6),
	.w8(32'hba580266),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9e42),
	.w1(32'h3a0b13f6),
	.w2(32'hbb5943b7),
	.w3(32'hbbb1c8e4),
	.w4(32'hbaee1801),
	.w5(32'h3ac10eab),
	.w6(32'hbb76a1ba),
	.w7(32'h3aed115d),
	.w8(32'hb927f274),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb019df5),
	.w1(32'h3aaa6d0d),
	.w2(32'h3a918721),
	.w3(32'hbb73383a),
	.w4(32'hbbcbf99e),
	.w5(32'hbaedb7d4),
	.w6(32'h3b9676e0),
	.w7(32'hbb65666e),
	.w8(32'hbb88a810),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef545),
	.w1(32'hbc450447),
	.w2(32'hbac7ad99),
	.w3(32'h3c1505b7),
	.w4(32'h3bab6d0f),
	.w5(32'h3b0533b2),
	.w6(32'h3b81802a),
	.w7(32'h3b815707),
	.w8(32'h3ba68b2d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39933b),
	.w1(32'hbc114372),
	.w2(32'hbb77d24b),
	.w3(32'h3c45d81e),
	.w4(32'hba497cb8),
	.w5(32'h3b5a27c6),
	.w6(32'h3c578b5a),
	.w7(32'hb931ccd1),
	.w8(32'h3aca5eeb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd39745),
	.w1(32'hbb80e659),
	.w2(32'h3c1ff753),
	.w3(32'hbc6203aa),
	.w4(32'hbc32b102),
	.w5(32'h3ba8c947),
	.w6(32'hbbabf4d6),
	.w7(32'hbbdfd14a),
	.w8(32'hbc25cb5a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b587a),
	.w1(32'hbbca70de),
	.w2(32'hbb4ac398),
	.w3(32'h3b0de8d0),
	.w4(32'hbab74103),
	.w5(32'h3b8c34dc),
	.w6(32'hbb52a612),
	.w7(32'hbc1d5459),
	.w8(32'h3b05761a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22dae7),
	.w1(32'hbb7434bf),
	.w2(32'h3b202fe4),
	.w3(32'h3bb0b0c5),
	.w4(32'hba755599),
	.w5(32'hbaac5489),
	.w6(32'hbaa1e25e),
	.w7(32'hbb7c1332),
	.w8(32'hbba88e21),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c327400),
	.w1(32'hbc16b2ed),
	.w2(32'h3c3f9b09),
	.w3(32'h3c89bb73),
	.w4(32'h3c3f983a),
	.w5(32'h3c1f1920),
	.w6(32'h3ca211d2),
	.w7(32'h3c6c7a3b),
	.w8(32'hbb0f0824),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6d5a),
	.w1(32'hbbb51878),
	.w2(32'hbb8ed787),
	.w3(32'h3c301dc3),
	.w4(32'h3c31624f),
	.w5(32'h3b484c4d),
	.w6(32'h3c3996d8),
	.w7(32'h3b01bc83),
	.w8(32'h3b97fd91),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3faf8b),
	.w1(32'h3b9920b4),
	.w2(32'hbba9e461),
	.w3(32'h3bb85999),
	.w4(32'hba070e5d),
	.w5(32'hbb02672a),
	.w6(32'h3c33c7bc),
	.w7(32'h3a85d442),
	.w8(32'h3bb5d9c0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f47ff),
	.w1(32'hba982243),
	.w2(32'hbae367b3),
	.w3(32'hbba09ad3),
	.w4(32'h39fc310a),
	.w5(32'h3a09bf5c),
	.w6(32'h3c0cdbba),
	.w7(32'h3c0c2991),
	.w8(32'hbb6f6933),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdadfcc),
	.w1(32'h3b062561),
	.w2(32'h3bd1c51e),
	.w3(32'h3c09e15f),
	.w4(32'h3abc50d6),
	.w5(32'hbb82dd87),
	.w6(32'h3b21973a),
	.w7(32'hbb7329e4),
	.w8(32'hba8919ee),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b957),
	.w1(32'h3b530a39),
	.w2(32'h3baafa77),
	.w3(32'hbb292c10),
	.w4(32'h3b9dbd31),
	.w5(32'h3a5eddf9),
	.w6(32'hbbecd816),
	.w7(32'hbc5593d1),
	.w8(32'hbc767f0e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c264b3c),
	.w1(32'h3ad21681),
	.w2(32'h3be75139),
	.w3(32'hbb9ad2b3),
	.w4(32'hbc5ffea7),
	.w5(32'h3c109354),
	.w6(32'hbc8c6aab),
	.w7(32'hbb5bb0b3),
	.w8(32'h3b75a51e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be32c5d),
	.w1(32'hbb244abe),
	.w2(32'h3bbc6257),
	.w3(32'h3bb30b30),
	.w4(32'h3bcb5eef),
	.w5(32'hbaceb506),
	.w6(32'h3b993cb3),
	.w7(32'h3b96c2ce),
	.w8(32'hbc1b8fd0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a512),
	.w1(32'h3acbfd0f),
	.w2(32'h3ba53a4c),
	.w3(32'h3a5075f1),
	.w4(32'hbc0e190c),
	.w5(32'h3b8d043e),
	.w6(32'hbc67b31a),
	.w7(32'hbabcdaef),
	.w8(32'hba880525),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57c0c6),
	.w1(32'h3b58ab5d),
	.w2(32'hbc067227),
	.w3(32'h3b7b26b8),
	.w4(32'h3bd8703f),
	.w5(32'hbb8020ab),
	.w6(32'hb707cfe7),
	.w7(32'hb899f7a0),
	.w8(32'h39f3b7d3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf3fb4),
	.w1(32'hbb8db2ef),
	.w2(32'h3a58e6e5),
	.w3(32'hbc5bd07a),
	.w4(32'hbaeead8b),
	.w5(32'hbba80cfd),
	.w6(32'h3be70761),
	.w7(32'h3c205c3d),
	.w8(32'h3bb48d3e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3219d6),
	.w1(32'hbb8b9e14),
	.w2(32'hba15016e),
	.w3(32'hbb8b4b6b),
	.w4(32'hbc31b3e7),
	.w5(32'hba8cd107),
	.w6(32'h3bd8498a),
	.w7(32'h3b448f7a),
	.w8(32'hbbaecf40),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab0fb),
	.w1(32'h3acb60f2),
	.w2(32'h3c00afdc),
	.w3(32'h3ca869ac),
	.w4(32'h3c144dff),
	.w5(32'h3c53b336),
	.w6(32'h3acf0a15),
	.w7(32'h3c3733ee),
	.w8(32'h3bb7b1cb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ad7f9),
	.w1(32'h3bd23cde),
	.w2(32'h3b4a1ccb),
	.w3(32'h3c2071f9),
	.w4(32'h3c33304c),
	.w5(32'hba952d7d),
	.w6(32'hb9666cb4),
	.w7(32'h3b94baa1),
	.w8(32'hbb4ae9ea),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfa358),
	.w1(32'h3a880422),
	.w2(32'hbb26d512),
	.w3(32'h3a7a58ee),
	.w4(32'h3bbe1a4d),
	.w5(32'hbbe3e459),
	.w6(32'h3b2119bf),
	.w7(32'h3c0df4bb),
	.w8(32'hbb20e94f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4add1e),
	.w1(32'h3b7dd4c6),
	.w2(32'h3bb2370a),
	.w3(32'h3bff3644),
	.w4(32'hba00b623),
	.w5(32'h3c7e9486),
	.w6(32'h3c556415),
	.w7(32'hbb5422f9),
	.w8(32'h3c28a982),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7705d4),
	.w1(32'hbc009278),
	.w2(32'h3bb045f0),
	.w3(32'h3c689c16),
	.w4(32'hbba65ac9),
	.w5(32'h3bbcebf6),
	.w6(32'h3c6f830e),
	.w7(32'hbc2425a4),
	.w8(32'hbaafa7d4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde6fc8),
	.w1(32'hbad5267b),
	.w2(32'h3be534a8),
	.w3(32'h3bac8399),
	.w4(32'h3bd29458),
	.w5(32'hbc393327),
	.w6(32'hba5b7613),
	.w7(32'hbb1909ff),
	.w8(32'hbc5a440d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca25a2b),
	.w1(32'h3c67240b),
	.w2(32'hba04c378),
	.w3(32'hbbb9d0fb),
	.w4(32'h3c9437bf),
	.w5(32'h3a270ab3),
	.w6(32'hbcc72e0a),
	.w7(32'hbc6c8eda),
	.w8(32'h3a788f3f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c049),
	.w1(32'hbb8d3f6a),
	.w2(32'hbc029040),
	.w3(32'hbae75251),
	.w4(32'hbaf4f7bb),
	.w5(32'hbb66c812),
	.w6(32'hb85b4f80),
	.w7(32'h3a11b4e4),
	.w8(32'h3c90c623),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a59fd),
	.w1(32'hbbb73d8d),
	.w2(32'hba19448a),
	.w3(32'hbc5114e6),
	.w4(32'hbba0e624),
	.w5(32'hba9010cd),
	.w6(32'h3cd3b0e1),
	.w7(32'h3cbe00c0),
	.w8(32'h393cca30),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b50b6),
	.w1(32'hbbb67006),
	.w2(32'h3b7d8bfd),
	.w3(32'hb978348f),
	.w4(32'hb9c0f36a),
	.w5(32'h3b8fed95),
	.w6(32'h3a70410c),
	.w7(32'h3b8746ac),
	.w8(32'h3a57f04a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8865f),
	.w1(32'hbac9b85a),
	.w2(32'h3c1d9f49),
	.w3(32'h3bcd7cf8),
	.w4(32'hba6d58d4),
	.w5(32'h3c4d7ccc),
	.w6(32'h3bad332a),
	.w7(32'h3b7ab729),
	.w8(32'h3c4a9236),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c270190),
	.w1(32'hbc1bcc40),
	.w2(32'hba49f9c5),
	.w3(32'h3c22c98a),
	.w4(32'hbc89c2eb),
	.w5(32'hbb81cd8d),
	.w6(32'h3bc9785c),
	.w7(32'hbba98510),
	.w8(32'hbabb6464),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbd6d6),
	.w1(32'hbc0d734b),
	.w2(32'hbb07da62),
	.w3(32'hbc0bb491),
	.w4(32'hbb25fa73),
	.w5(32'hbae41bd1),
	.w6(32'hbbe68edb),
	.w7(32'h3b916edf),
	.w8(32'hbb1a7b3e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e51f8),
	.w1(32'hbbaadce8),
	.w2(32'hbab60e43),
	.w3(32'h3ae76935),
	.w4(32'hbbd59882),
	.w5(32'h3b311744),
	.w6(32'h3b3a1e12),
	.w7(32'hbba5f70f),
	.w8(32'h3b822a4e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfe813),
	.w1(32'hbae66170),
	.w2(32'hba86541f),
	.w3(32'h3b882c33),
	.w4(32'hb9f716b9),
	.w5(32'h3a8cb972),
	.w6(32'h3ba88ee6),
	.w7(32'hbb389d6c),
	.w8(32'h3ba124fb),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43634),
	.w1(32'hba796483),
	.w2(32'hbb2444e9),
	.w3(32'h3ab61dec),
	.w4(32'h3b4000d6),
	.w5(32'h3be445ab),
	.w6(32'hba69ff76),
	.w7(32'h3b24c1c6),
	.w8(32'h3c197fc8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56c2f3),
	.w1(32'h3b866370),
	.w2(32'h3bdada9f),
	.w3(32'h3bcc8a2e),
	.w4(32'hbb8a5c96),
	.w5(32'h3bd22af0),
	.w6(32'h3c3f2b58),
	.w7(32'hbb5b1f93),
	.w8(32'h3befe426),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c29f1),
	.w1(32'hbbe9e926),
	.w2(32'hbb27cfbd),
	.w3(32'h3c5d13ca),
	.w4(32'h3c7f3732),
	.w5(32'hbb272472),
	.w6(32'h3cb33e96),
	.w7(32'h3cb84c02),
	.w8(32'hbbde18fc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd89c),
	.w1(32'hbbba5fa8),
	.w2(32'h3b0010aa),
	.w3(32'h3a96214d),
	.w4(32'hbbfa0968),
	.w5(32'h3b823a38),
	.w6(32'hbb098d09),
	.w7(32'hbbb4c3bb),
	.w8(32'h3bf0a4a9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92b5ba),
	.w1(32'hbb397432),
	.w2(32'hbc4cb559),
	.w3(32'h3beee30e),
	.w4(32'hbbba6dd8),
	.w5(32'hbc04ebdb),
	.w6(32'h3c4bee31),
	.w7(32'h3ae09537),
	.w8(32'hba304340),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc814bc),
	.w1(32'hbc491466),
	.w2(32'hbc4a1463),
	.w3(32'h39bf438b),
	.w4(32'hbb077b5b),
	.w5(32'hbbcb5060),
	.w6(32'h3c40d02d),
	.w7(32'h3c89a153),
	.w8(32'h3c39d310),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d7ab7),
	.w1(32'hbb4142ef),
	.w2(32'hbbaf0832),
	.w3(32'h3a2459ec),
	.w4(32'h3bfdcf3e),
	.w5(32'hbbcaa866),
	.w6(32'h3c72cbfb),
	.w7(32'h3c8059d5),
	.w8(32'hbb891286),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff0f07),
	.w1(32'hbbb14c08),
	.w2(32'hba4dcdc1),
	.w3(32'h3b973589),
	.w4(32'hbb41e58f),
	.w5(32'h3c136633),
	.w6(32'h3c4099fc),
	.w7(32'hbbba3319),
	.w8(32'h3bfe4402),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afab5d4),
	.w1(32'h3a06c3a5),
	.w2(32'hb998b948),
	.w3(32'h3bfc781a),
	.w4(32'h3b6a1918),
	.w5(32'h3aaf4dae),
	.w6(32'h3bc652a4),
	.w7(32'h399710d6),
	.w8(32'hb9751f0a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb497f01),
	.w1(32'hbc23a40f),
	.w2(32'h3b6ad124),
	.w3(32'h3b9af716),
	.w4(32'hbbb3891d),
	.w5(32'h3b3aee43),
	.w6(32'h3c265794),
	.w7(32'hb9ced662),
	.w8(32'h3bdc3b5b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ac388),
	.w1(32'h3a91dbe4),
	.w2(32'h3c382808),
	.w3(32'h3b08d75a),
	.w4(32'h3a92c270),
	.w5(32'h3c6cecf4),
	.w6(32'h3ba79710),
	.w7(32'h3baf2357),
	.w8(32'h3c872741),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ee8a6),
	.w1(32'h3bce268b),
	.w2(32'h3aa4634f),
	.w3(32'h3c0abc71),
	.w4(32'hbb4b1452),
	.w5(32'h3b1b8a05),
	.w6(32'h3bbcdfb8),
	.w7(32'hbb0b05f2),
	.w8(32'h3c3ed5d8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c035036),
	.w1(32'hba84c7a4),
	.w2(32'hbc43a62f),
	.w3(32'h3c323404),
	.w4(32'h3bd15324),
	.w5(32'hbb87d408),
	.w6(32'h3c7f00d2),
	.w7(32'h3bcd26e2),
	.w8(32'h3bafe80a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a745163),
	.w1(32'h3b30403a),
	.w2(32'h3c35ab84),
	.w3(32'h3c01fc8c),
	.w4(32'h3b136378),
	.w5(32'h3ca9d208),
	.w6(32'h3c772aab),
	.w7(32'hb9d5970a),
	.w8(32'h3c0b0ab3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb2444),
	.w1(32'hbc0466e5),
	.w2(32'h3b413906),
	.w3(32'hbb976472),
	.w4(32'hbbfb3ecc),
	.w5(32'h3bb96836),
	.w6(32'h3c0d8ece),
	.w7(32'hbb92eca3),
	.w8(32'h3c0823b5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36a3c6),
	.w1(32'h3b66388b),
	.w2(32'h3ad4769a),
	.w3(32'h3c71f694),
	.w4(32'h3c0d1106),
	.w5(32'h3c0c1d2a),
	.w6(32'h3ba4d263),
	.w7(32'h3a4912dc),
	.w8(32'hbbf77a34),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163b22),
	.w1(32'hbafb0226),
	.w2(32'h3c53faed),
	.w3(32'hba89d295),
	.w4(32'hbaa11a72),
	.w5(32'h3bda213a),
	.w6(32'hba586d53),
	.w7(32'hbab3e496),
	.w8(32'hbc558094),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1c1cd),
	.w1(32'h35ee132c),
	.w2(32'hba0d4daf),
	.w3(32'hbbdd04fa),
	.w4(32'hbbf18854),
	.w5(32'hbbef77ca),
	.w6(32'hbc7049a3),
	.w7(32'hbb29affa),
	.w8(32'hbbacf9c8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d9e5),
	.w1(32'h3b6079e7),
	.w2(32'h3acd85a0),
	.w3(32'h39e7a65b),
	.w4(32'hbc62d37f),
	.w5(32'hb9de313c),
	.w6(32'h3ae69a52),
	.w7(32'hbbc39090),
	.w8(32'hbb82155d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf74f7b),
	.w1(32'hb9dcc2f9),
	.w2(32'h3b9e9213),
	.w3(32'h3bcac93d),
	.w4(32'h3a90efb3),
	.w5(32'h3b92af15),
	.w6(32'h3bcd4e80),
	.w7(32'h3b1bd0cc),
	.w8(32'h3b4a9b6e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75d504),
	.w1(32'h3bf23791),
	.w2(32'h3992ba49),
	.w3(32'h3c40ad51),
	.w4(32'h3c1fa5d6),
	.w5(32'hb97cbb13),
	.w6(32'h3c077a98),
	.w7(32'hba808b4e),
	.w8(32'hbb518604),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf591d9),
	.w1(32'hbc0e0c35),
	.w2(32'hbbc0406d),
	.w3(32'h3b532a7d),
	.w4(32'hbb0c6cfd),
	.w5(32'h3b29a2bf),
	.w6(32'h3b71787a),
	.w7(32'h3a5e6786),
	.w8(32'h3ba73a25),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc3db0),
	.w1(32'hbbc8bb86),
	.w2(32'h393312b1),
	.w3(32'h3c101c23),
	.w4(32'hbae117a4),
	.w5(32'hbbdf8db4),
	.w6(32'h3c1df5a3),
	.w7(32'hb9c66412),
	.w8(32'h39b57433),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b731f2c),
	.w1(32'h3b38b1df),
	.w2(32'h398cb7da),
	.w3(32'hbc311b66),
	.w4(32'hbc0450ed),
	.w5(32'h3bc3f70f),
	.w6(32'hbc118d58),
	.w7(32'hbb329798),
	.w8(32'h3b8f3426),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f21dc),
	.w1(32'h3bc8e9c1),
	.w2(32'h3b9dd8ac),
	.w3(32'h3c5bb23b),
	.w4(32'h3c097749),
	.w5(32'h394d0a3f),
	.w6(32'h3b3f0408),
	.w7(32'hbc029106),
	.w8(32'hbb2450f4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb666cff6),
	.w1(32'hba1bd623),
	.w2(32'h3b2accba),
	.w3(32'hbbd9764d),
	.w4(32'hbab9a8af),
	.w5(32'hbc239af6),
	.w6(32'hbc010658),
	.w7(32'h3b658ac8),
	.w8(32'hbc2a5f20),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f89c7),
	.w1(32'h3c381319),
	.w2(32'hbb3c5f02),
	.w3(32'hbb2be622),
	.w4(32'h3c69549f),
	.w5(32'hbbbda8d8),
	.w6(32'hbc603666),
	.w7(32'hbb9bdebf),
	.w8(32'hbb81c424),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3be420),
	.w1(32'hbb8361d3),
	.w2(32'h3b41a822),
	.w3(32'hbb6c3416),
	.w4(32'hbb14dc96),
	.w5(32'h3b654783),
	.w6(32'hbabbe39e),
	.w7(32'hbaf8a9a3),
	.w8(32'h398f550c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be75fc7),
	.w1(32'h3b306f34),
	.w2(32'h3ae1c62e),
	.w3(32'h3c0d98f4),
	.w4(32'h3b8dc244),
	.w5(32'h3cbfcd18),
	.w6(32'h3bf6bc41),
	.w7(32'h3c14f438),
	.w8(32'h3c668aa1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc62b),
	.w1(32'hbbf4a5dd),
	.w2(32'hbbe1f9b8),
	.w3(32'h3ca58552),
	.w4(32'h3b67e334),
	.w5(32'h3c9d1e0d),
	.w6(32'h3cb71060),
	.w7(32'h3b42b67b),
	.w8(32'h3c969da6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5517fd),
	.w1(32'hbc414c42),
	.w2(32'h3adbead8),
	.w3(32'h3c6dca87),
	.w4(32'h3b033a6c),
	.w5(32'h3bc0b229),
	.w6(32'h3cd63989),
	.w7(32'h3c8b66ce),
	.w8(32'hba9733a3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb07710),
	.w1(32'h3b0fc8da),
	.w2(32'h3a985a60),
	.w3(32'h3cbf8a19),
	.w4(32'h3be0ab38),
	.w5(32'h3bdcc894),
	.w6(32'h3c817fd3),
	.w7(32'h3b93a5c4),
	.w8(32'hbb66867c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc04b2f),
	.w1(32'h3bb7027a),
	.w2(32'h3bf117c5),
	.w3(32'h3c18ccdd),
	.w4(32'h3b8db5f6),
	.w5(32'h3baff746),
	.w6(32'h3b61b5c6),
	.w7(32'h3b264d54),
	.w8(32'h3ba47d30),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb875d39),
	.w1(32'h398b4949),
	.w2(32'h3b9a6c6c),
	.w3(32'hbc0de205),
	.w4(32'hbbec75ef),
	.w5(32'h3a954537),
	.w6(32'hbab6de26),
	.w7(32'hbc0b086c),
	.w8(32'h3af7ab80),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe25f),
	.w1(32'h3a83ebf1),
	.w2(32'h3bb21522),
	.w3(32'hbadc8513),
	.w4(32'h3b0b19b9),
	.w5(32'h3bc36403),
	.w6(32'hba5f1557),
	.w7(32'h3bc029e4),
	.w8(32'h3ba37f8b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2084ec),
	.w1(32'hb939837d),
	.w2(32'hbbb17131),
	.w3(32'h3a42ee37),
	.w4(32'h3b5742c0),
	.w5(32'hbbc36ab9),
	.w6(32'h3b078749),
	.w7(32'h3baed397),
	.w8(32'h3b77837b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0386ff),
	.w1(32'hbaed84c0),
	.w2(32'hbbf51252),
	.w3(32'h3b3e4961),
	.w4(32'h3b402e8e),
	.w5(32'hbbd67d41),
	.w6(32'h3bdbc6e3),
	.w7(32'h3b97b701),
	.w8(32'hbb4d0d71),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784c86),
	.w1(32'h3c3fd491),
	.w2(32'h3ae23f1b),
	.w3(32'hbba23230),
	.w4(32'h3be23bb3),
	.w5(32'hbbdb38f8),
	.w6(32'hbc14a506),
	.w7(32'hbb5fe781),
	.w8(32'hbaa98aef),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9022),
	.w1(32'h3c24fd64),
	.w2(32'h3c71c4ad),
	.w3(32'hbb61c0ca),
	.w4(32'hb7c699f3),
	.w5(32'hbc48df95),
	.w6(32'hbb931a2b),
	.w7(32'h3abe07e4),
	.w8(32'hbc840ad5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82bc06),
	.w1(32'h3b2d26dc),
	.w2(32'h3979c3e2),
	.w3(32'h3b940aeb),
	.w4(32'h3b82955e),
	.w5(32'h3c6801a7),
	.w6(32'hbc942bc3),
	.w7(32'hbc7b4a9c),
	.w8(32'h3bedd477),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6ed5b),
	.w1(32'h39dce8e6),
	.w2(32'h3c6d86de),
	.w3(32'h3c38a508),
	.w4(32'hbbbb70fa),
	.w5(32'h3c1d2245),
	.w6(32'h3b3c1450),
	.w7(32'hbb730a05),
	.w8(32'h3adbc48f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b0aed),
	.w1(32'h3c58d140),
	.w2(32'h3b79abbf),
	.w3(32'h3c9648c8),
	.w4(32'h3a8bd80d),
	.w5(32'hbac3f6a5),
	.w6(32'h3bcf4dba),
	.w7(32'hbb9c47a9),
	.w8(32'hbc0d1c69),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3800fd),
	.w1(32'h3a882670),
	.w2(32'h3bda611a),
	.w3(32'h3c35e964),
	.w4(32'h3c3467e8),
	.w5(32'hbb1f58c4),
	.w6(32'hbae08986),
	.w7(32'hbbe6717a),
	.w8(32'hbc089c9a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8184cd1),
	.w1(32'hba996351),
	.w2(32'h391107c1),
	.w3(32'hbbfa8f9c),
	.w4(32'hbbb817e9),
	.w5(32'h39369e61),
	.w6(32'hbbfc38d9),
	.w7(32'hbbce3679),
	.w8(32'h39d361a2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e4eac),
	.w1(32'h3a978a78),
	.w2(32'h3b406cc5),
	.w3(32'h3af333f9),
	.w4(32'h3a988833),
	.w5(32'hbb1b5b98),
	.w6(32'h3a8919a6),
	.w7(32'hbabedd05),
	.w8(32'hbb12846c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b976ec0),
	.w1(32'hbb53c01b),
	.w2(32'hb9c2f833),
	.w3(32'h3b1c1f3a),
	.w4(32'h3b872765),
	.w5(32'hb92c2631),
	.w6(32'h3a24f620),
	.w7(32'h39c1ae6f),
	.w8(32'h39cdc6a0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce86f4),
	.w1(32'h3b0f328f),
	.w2(32'hbbae6394),
	.w3(32'hb93e6540),
	.w4(32'h3b082e7f),
	.w5(32'hbbe3d80a),
	.w6(32'h3a2ab575),
	.w7(32'h3a6be078),
	.w8(32'h37048e59),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba471fe),
	.w1(32'h3b540041),
	.w2(32'h3b3a003c),
	.w3(32'h3ba579a4),
	.w4(32'hbbbfa933),
	.w5(32'h3c94abee),
	.w6(32'h3c9b08d6),
	.w7(32'h3c13cda1),
	.w8(32'h3cc5889c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3df150),
	.w1(32'hbc1331f4),
	.w2(32'h3c0e792d),
	.w3(32'h3bd0f207),
	.w4(32'hbb3c718d),
	.w5(32'hbc236e52),
	.w6(32'h3ccc90d9),
	.w7(32'h3c7cf48a),
	.w8(32'hbc760781),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80e0e6),
	.w1(32'h3c3b9c46),
	.w2(32'h3b7a96b6),
	.w3(32'hba8d5160),
	.w4(32'h3c17d85d),
	.w5(32'h3b608d11),
	.w6(32'hbcb22330),
	.w7(32'hbc6b4963),
	.w8(32'h3b260981),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b96f),
	.w1(32'h3b030c07),
	.w2(32'h3b139ff1),
	.w3(32'h3bd235b1),
	.w4(32'h3b9329ac),
	.w5(32'h3adb8a00),
	.w6(32'h3b5e2bf8),
	.w7(32'h39d50f1a),
	.w8(32'h3b13bca0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd9a60),
	.w1(32'hba6ae746),
	.w2(32'hbc021bfc),
	.w3(32'hbb17b9c6),
	.w4(32'hbb8763d6),
	.w5(32'hbb892fac),
	.w6(32'h392fa37d),
	.w7(32'hb9cad439),
	.w8(32'hbacb114d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae14295),
	.w1(32'hbae09655),
	.w2(32'h3ad00a33),
	.w3(32'h3b8632ac),
	.w4(32'h3b9ecb36),
	.w5(32'h3a1fc1f7),
	.w6(32'hbb038003),
	.w7(32'hbb73c52d),
	.w8(32'hbb644a52),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f67d4),
	.w1(32'h3b6e1ff5),
	.w2(32'h3b3bf7fe),
	.w3(32'hb93c8b86),
	.w4(32'h3a0e3cda),
	.w5(32'h3b862cb4),
	.w6(32'hbba50e21),
	.w7(32'hbb3d2bec),
	.w8(32'hbb5d1f92),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caecaad),
	.w1(32'h3bc95962),
	.w2(32'h3ca7790c),
	.w3(32'h3c805dea),
	.w4(32'hbb81e683),
	.w5(32'h3c8c0f07),
	.w6(32'h3c039d37),
	.w7(32'hbb9cb658),
	.w8(32'h3be4353a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a114194),
	.w1(32'h398d57a3),
	.w2(32'h3c18cd28),
	.w3(32'h3c21ea74),
	.w4(32'hbc4d13b7),
	.w5(32'h3ca5af3a),
	.w6(32'h3bd62782),
	.w7(32'h3b143517),
	.w8(32'h3c55da3b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf436ad),
	.w1(32'hbbe38d5f),
	.w2(32'hbc3aa5b1),
	.w3(32'h3c2b369b),
	.w4(32'hbc14a6d1),
	.w5(32'h3b406fed),
	.w6(32'h3c98aeaa),
	.w7(32'h3af8b7d1),
	.w8(32'h3b80e39f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule