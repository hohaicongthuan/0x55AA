module layer_10_featuremap_442(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b27eb),
	.w1(32'h3b14bdcb),
	.w2(32'hbb06d3c7),
	.w3(32'h3acc5ade),
	.w4(32'hba9a6f62),
	.w5(32'hbb13068a),
	.w6(32'hb95272a2),
	.w7(32'hbadfd663),
	.w8(32'hba2c83c7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad02cf),
	.w1(32'hbb80a96b),
	.w2(32'hbbe3d999),
	.w3(32'hbc855049),
	.w4(32'h3b0cf99b),
	.w5(32'hb9c400e2),
	.w6(32'hbc63bf01),
	.w7(32'hbbaccecf),
	.w8(32'hbbd65ea7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29ab40),
	.w1(32'h3b951bac),
	.w2(32'hbaf89b6b),
	.w3(32'hbb4e59e6),
	.w4(32'h3b106c7f),
	.w5(32'hbb3cddac),
	.w6(32'hbbaba9ed),
	.w7(32'h38c09a3a),
	.w8(32'hba64faa8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4419fc),
	.w1(32'h3ad72eeb),
	.w2(32'h3bc53595),
	.w3(32'h3b76b0d9),
	.w4(32'h3a713853),
	.w5(32'h3a7eb6ee),
	.w6(32'h3acd95e8),
	.w7(32'h3bfe2412),
	.w8(32'hbb2cef9b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd35f),
	.w1(32'hbb049cc9),
	.w2(32'hb9ad88e4),
	.w3(32'h3b026303),
	.w4(32'hbaf1d19f),
	.w5(32'h39312dd7),
	.w6(32'h3b0db570),
	.w7(32'h3b4ca68c),
	.w8(32'h3ac05da7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fa0b2),
	.w1(32'h3b6b3a39),
	.w2(32'h39e4161e),
	.w3(32'h3aafbe68),
	.w4(32'hbb03ea96),
	.w5(32'h3bf6ec70),
	.w6(32'h3ab93977),
	.w7(32'hba8ba24f),
	.w8(32'h3c85ad05),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c276dbe),
	.w1(32'hbc3be420),
	.w2(32'hbc9d1820),
	.w3(32'h3bbeb3c8),
	.w4(32'hbc23dfad),
	.w5(32'hbcb3e6bc),
	.w6(32'h3ad9104b),
	.w7(32'hbb12f587),
	.w8(32'hbc653ba9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ad46),
	.w1(32'hbc2f3269),
	.w2(32'hbc450c2e),
	.w3(32'hbc8b0de3),
	.w4(32'hbb2f5224),
	.w5(32'h3b181254),
	.w6(32'hbc12175e),
	.w7(32'hbc84e10a),
	.w8(32'hbba725b6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb848359),
	.w1(32'h3b645877),
	.w2(32'h3bc847db),
	.w3(32'h3b1973b9),
	.w4(32'h3b4864be),
	.w5(32'h3b20b62b),
	.w6(32'hba11c3da),
	.w7(32'h3b9bd16a),
	.w8(32'h39f866e7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510117),
	.w1(32'hbb766854),
	.w2(32'hbd09ac1d),
	.w3(32'hbb4ce8dc),
	.w4(32'h3bfa22bd),
	.w5(32'hbca09288),
	.w6(32'hbc497a86),
	.w7(32'h3bb2f86f),
	.w8(32'hbc8417dd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e6cf),
	.w1(32'hbb416b77),
	.w2(32'hbbd11d23),
	.w3(32'hba2c86ed),
	.w4(32'hba905775),
	.w5(32'hbb32b540),
	.w6(32'h3b465fab),
	.w7(32'h3b5b6b77),
	.w8(32'hbb0c43c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2abaa),
	.w1(32'h3c0a2f8e),
	.w2(32'hbc89d224),
	.w3(32'hbc2d3d4c),
	.w4(32'h3b573f9a),
	.w5(32'hbcc8ff82),
	.w6(32'hbbf5e14f),
	.w7(32'h3bb81c48),
	.w8(32'hbcba1ffa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030287),
	.w1(32'h3b0e621c),
	.w2(32'hbcf26430),
	.w3(32'h3b816d91),
	.w4(32'h3c092eda),
	.w5(32'hbc811d98),
	.w6(32'h3aa408e2),
	.w7(32'h3c5a895a),
	.w8(32'hbc5f4db5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2078fe),
	.w1(32'hbb8419af),
	.w2(32'hbc31fcc0),
	.w3(32'hbb89c9ae),
	.w4(32'hbb3890a4),
	.w5(32'hbc0e7b37),
	.w6(32'hbc0fbc49),
	.w7(32'hbbb3103e),
	.w8(32'hbba4691f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178179),
	.w1(32'hbaa7544d),
	.w2(32'hbc1f5691),
	.w3(32'hbbebc3ed),
	.w4(32'h3bc4f4d8),
	.w5(32'h3a323182),
	.w6(32'hbc6235e7),
	.w7(32'h3a816b84),
	.w8(32'hbc02c425),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f9a98),
	.w1(32'hbc12b425),
	.w2(32'hbcea86e3),
	.w3(32'hbbfe2a2d),
	.w4(32'h3b232dbe),
	.w5(32'hbc49010e),
	.w6(32'hbc4b68ff),
	.w7(32'hbb17ed5a),
	.w8(32'hbcacec3a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f29aa),
	.w1(32'h3a5f2013),
	.w2(32'h3b8cf1ba),
	.w3(32'hbb826747),
	.w4(32'hbb006199),
	.w5(32'hbb299a8f),
	.w6(32'hbb7f5d2d),
	.w7(32'hbab1f315),
	.w8(32'hbb439933),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b923e),
	.w1(32'hbbf93024),
	.w2(32'hbceb5e01),
	.w3(32'hbc7a9bd1),
	.w4(32'hbb0b3ff6),
	.w5(32'hbccce4ed),
	.w6(32'hbc6f06d9),
	.w7(32'hbba9f741),
	.w8(32'hbcb9e36c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870d90),
	.w1(32'hbb3dbe01),
	.w2(32'hbc7ddfaa),
	.w3(32'h3b0c562b),
	.w4(32'hbbb2596a),
	.w5(32'hbc5b446d),
	.w6(32'hbaccf187),
	.w7(32'hbabd7583),
	.w8(32'hbc14b66e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf41460),
	.w1(32'h3b4b5107),
	.w2(32'h398b875e),
	.w3(32'hba3566a0),
	.w4(32'hb86a8c7b),
	.w5(32'hbb7d1e8c),
	.w6(32'h3a345b14),
	.w7(32'h3b9d5c4d),
	.w8(32'h3af6c6f2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d4eb),
	.w1(32'hbac1c444),
	.w2(32'hbb9cf120),
	.w3(32'hbb3206d5),
	.w4(32'hbb96c0a9),
	.w5(32'h3a841660),
	.w6(32'hbb9d889c),
	.w7(32'h3a1930d8),
	.w8(32'h3ba56a6d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6013),
	.w1(32'h3c115732),
	.w2(32'h3b28d231),
	.w3(32'h3badd9a6),
	.w4(32'h3c03364a),
	.w5(32'h3c6e528e),
	.w6(32'hbb8f79b7),
	.w7(32'h3b91e121),
	.w8(32'h3b9607b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd52f19e),
	.w1(32'hbc6b74a4),
	.w2(32'hbd02ccb4),
	.w3(32'hbcf1924e),
	.w4(32'h3b2999ed),
	.w5(32'hbce0202f),
	.w6(32'hbd3cd627),
	.w7(32'hbc76e08e),
	.w8(32'hbd4fd594),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb12c90),
	.w1(32'h3b8632d0),
	.w2(32'hbcde7a4b),
	.w3(32'hbc17de21),
	.w4(32'h3c4e566d),
	.w5(32'hbc6dffb7),
	.w6(32'hbc75f0dd),
	.w7(32'h3c1e585e),
	.w8(32'hbc8a96d5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd019c41),
	.w1(32'h3af4120e),
	.w2(32'hbb781b8c),
	.w3(32'hbcb252e6),
	.w4(32'h3cad3d9d),
	.w5(32'h3c3267ba),
	.w6(32'hbd078387),
	.w7(32'h3becca7c),
	.w8(32'hbbd84cc7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911207d),
	.w1(32'h3ad57397),
	.w2(32'h3bd393e1),
	.w3(32'h3c5b8120),
	.w4(32'h3b201358),
	.w5(32'h3c46de4f),
	.w6(32'h3c4a4835),
	.w7(32'hba0b6191),
	.w8(32'h3b3673ad),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be371a6),
	.w1(32'h3b9eb83e),
	.w2(32'h3b90f73b),
	.w3(32'h3c35a43c),
	.w4(32'h39e55c1a),
	.w5(32'h3c82f174),
	.w6(32'h3b656706),
	.w7(32'hbb9a5228),
	.w8(32'h3ab7889e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3c9dc),
	.w1(32'hbb867b54),
	.w2(32'h3aa8d023),
	.w3(32'h3af3e290),
	.w4(32'h39da2d47),
	.w5(32'h3b441202),
	.w6(32'hbc43500f),
	.w7(32'hbb794707),
	.w8(32'h3b5183be),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad012e),
	.w1(32'h3ba63a5a),
	.w2(32'h3a849381),
	.w3(32'hb98c689e),
	.w4(32'h3b42cd9f),
	.w5(32'hb9857cfa),
	.w6(32'hb92e8fe5),
	.w7(32'hbb059ab8),
	.w8(32'hbb69c7ec),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf601a),
	.w1(32'h3bcc9bdb),
	.w2(32'hbb3ec751),
	.w3(32'hbb0ee3ee),
	.w4(32'h3c219808),
	.w5(32'h3b54909b),
	.w6(32'hbc1cfcae),
	.w7(32'h3c00cb1c),
	.w8(32'h3bc769e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273a4a),
	.w1(32'hba0258ec),
	.w2(32'hba556851),
	.w3(32'hb92dd75e),
	.w4(32'h39d4c171),
	.w5(32'hbb7648e7),
	.w6(32'h39caca8e),
	.w7(32'hb98aefc0),
	.w8(32'hbb885771),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba354da2),
	.w1(32'h3a53e1b5),
	.w2(32'hbaf55f1b),
	.w3(32'hbab932a9),
	.w4(32'h3b2243b7),
	.w5(32'hbb09fcde),
	.w6(32'hba1de3b8),
	.w7(32'h3b65b6c6),
	.w8(32'hba2e40e6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd4b3),
	.w1(32'hbb56dd80),
	.w2(32'hbc898eb6),
	.w3(32'h3a7553d1),
	.w4(32'h3b9e7654),
	.w5(32'hbc3c0a05),
	.w6(32'hbba85fae),
	.w7(32'h3b3313b2),
	.w8(32'hbbe743b4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc882204),
	.w1(32'hbb1966f4),
	.w2(32'hba907452),
	.w3(32'hbc2e1c0c),
	.w4(32'h3a9b7c6b),
	.w5(32'hbb9e11d0),
	.w6(32'hbc1e5e7e),
	.w7(32'h39993503),
	.w8(32'hbbd89113),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca78bc),
	.w1(32'h3b99d34e),
	.w2(32'h382674db),
	.w3(32'hbb0ed6b9),
	.w4(32'h3a6a5ff9),
	.w5(32'hbb872727),
	.w6(32'hbb736791),
	.w7(32'hbb2ddeeb),
	.w8(32'h39db7083),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db72a),
	.w1(32'hbad78776),
	.w2(32'hbc13ad20),
	.w3(32'h3ba62216),
	.w4(32'h3a195890),
	.w5(32'hbbac9485),
	.w6(32'h3b542cb9),
	.w7(32'hbafb72e3),
	.w8(32'hbc092c60),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd33fa7),
	.w1(32'hba3269be),
	.w2(32'hbcf7e104),
	.w3(32'hbc984dbe),
	.w4(32'h3c1a82bd),
	.w5(32'hbc4378b6),
	.w6(32'hbc3f8b26),
	.w7(32'h3c9729b9),
	.w8(32'hbca74473),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7d5cdb),
	.w1(32'h3c1fe5e8),
	.w2(32'h3c289590),
	.w3(32'hbd25adbd),
	.w4(32'h3c8c9549),
	.w5(32'h3c9c58b2),
	.w6(32'hbd853b5c),
	.w7(32'hbbbb3f3f),
	.w8(32'hbb20a819),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2251f0),
	.w1(32'h3aeba267),
	.w2(32'hbb3b8b6b),
	.w3(32'hbd092512),
	.w4(32'h3bbba177),
	.w5(32'hbbbebfe5),
	.w6(32'hbd50645b),
	.w7(32'hbc6f6f24),
	.w8(32'hbcb49391),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc362a3c),
	.w1(32'h3aebfce5),
	.w2(32'h3b1aacb2),
	.w3(32'hbc1cb16f),
	.w4(32'h3ba36609),
	.w5(32'h3c0758b9),
	.w6(32'hbc52e950),
	.w7(32'h3a47ad8a),
	.w8(32'hba0ce0a7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9029a),
	.w1(32'hbb59c733),
	.w2(32'hbba39387),
	.w3(32'h3b507d60),
	.w4(32'hbb1fd0cd),
	.w5(32'hbad2945f),
	.w6(32'h3a083b81),
	.w7(32'h3a65cd78),
	.w8(32'hb9e37120),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb84f28),
	.w1(32'hbb04dec7),
	.w2(32'hb9a326f8),
	.w3(32'hbb891788),
	.w4(32'hbb279b3c),
	.w5(32'h3b05a94e),
	.w6(32'hba58276e),
	.w7(32'h39592877),
	.w8(32'hb89a56b8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5eed9a),
	.w1(32'hba2f5cd6),
	.w2(32'hbb91ed52),
	.w3(32'hbc7da246),
	.w4(32'hbae27519),
	.w5(32'hbbb406b1),
	.w6(32'hbc66c4b4),
	.w7(32'hb80d3582),
	.w8(32'hbc0e9fbc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6704a),
	.w1(32'hbc3f4814),
	.w2(32'hbd118380),
	.w3(32'hbba5a53a),
	.w4(32'h3a6d17d4),
	.w5(32'hbc999a1d),
	.w6(32'hbc70f3ab),
	.w7(32'hbc1310e4),
	.w8(32'hbcd36892),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcaf7e),
	.w1(32'hbb08314c),
	.w2(32'hbcc48f6c),
	.w3(32'hbc09916b),
	.w4(32'h3c50c0ff),
	.w5(32'hbb9896d8),
	.w6(32'hbc5b9d19),
	.w7(32'h3c160811),
	.w8(32'hbc463b7b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccaefc0),
	.w1(32'hbb5f7a37),
	.w2(32'hbd02f06a),
	.w3(32'hbac59b6b),
	.w4(32'h3c8a0cf8),
	.w5(32'hbc121192),
	.w6(32'hbc87f559),
	.w7(32'h3c08d034),
	.w8(32'hbc892428),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc11821),
	.w1(32'hb980e229),
	.w2(32'hbc6ebaa2),
	.w3(32'hbc9f7ed2),
	.w4(32'h3bc477b2),
	.w5(32'hbb7f7fbb),
	.w6(32'hbcd61feb),
	.w7(32'hbc04e130),
	.w8(32'hbc9fe6db),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba265f21),
	.w1(32'hbbbd0518),
	.w2(32'hbcb4ec34),
	.w3(32'hbb9d85a4),
	.w4(32'hbafa414d),
	.w5(32'hbc834fe3),
	.w6(32'hbc22fc21),
	.w7(32'hbc01d98f),
	.w8(32'hbca26867),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c8582),
	.w1(32'h3b4bad6d),
	.w2(32'h3b55fe8b),
	.w3(32'hbb67fb97),
	.w4(32'hb706fd4a),
	.w5(32'hb98acfc1),
	.w6(32'hba8bac78),
	.w7(32'hbb20803a),
	.w8(32'h3b44ca0e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0acff6),
	.w1(32'h3b98ecf2),
	.w2(32'h3b909cfa),
	.w3(32'h38f8a924),
	.w4(32'h3ac7bef2),
	.w5(32'h3b6728e8),
	.w6(32'h389cec61),
	.w7(32'hb9d175b3),
	.w8(32'h3b2c68b3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb348d0),
	.w1(32'h3a99b6dc),
	.w2(32'hbb1e093a),
	.w3(32'h3b21c638),
	.w4(32'hbae086f2),
	.w5(32'hba15e13e),
	.w6(32'hb9e599ab),
	.w7(32'hbbb1fa37),
	.w8(32'h3ae2bfa7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab36c),
	.w1(32'hbad8f352),
	.w2(32'hbc8d313f),
	.w3(32'hbb418405),
	.w4(32'h3bdccb52),
	.w5(32'hbba044d3),
	.w6(32'hbc0156b4),
	.w7(32'h3b68a69c),
	.w8(32'hba1bf190),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c3565),
	.w1(32'h3a36de07),
	.w2(32'hbc145e46),
	.w3(32'hbbe499ff),
	.w4(32'h3aa9e0c2),
	.w5(32'hbbdbf816),
	.w6(32'hbbabc426),
	.w7(32'h3aed2eb2),
	.w8(32'hbb124683),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc268b17),
	.w1(32'hbc1591d0),
	.w2(32'hbd0d7ac5),
	.w3(32'hbb9bec70),
	.w4(32'hb898b154),
	.w5(32'hbca1a652),
	.w6(32'hbbee1e05),
	.w7(32'hba5a44ec),
	.w8(32'hbc59a632),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb973ba2d),
	.w1(32'hbb3ed3c5),
	.w2(32'h3b02cbed),
	.w3(32'h3a0c2d90),
	.w4(32'hbb96456d),
	.w5(32'h3a88d852),
	.w6(32'hbba7cbff),
	.w7(32'hbbfbbb9d),
	.w8(32'hbbb61332),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c040ee4),
	.w1(32'h3a9f2297),
	.w2(32'h373eb8b2),
	.w3(32'h3c4a231a),
	.w4(32'h3b26e18b),
	.w5(32'h3a135423),
	.w6(32'h3c09cc16),
	.w7(32'h3a989632),
	.w8(32'h3b020e41),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978ab18),
	.w1(32'hbb0ad186),
	.w2(32'hbb43d9cb),
	.w3(32'hb99bc2a2),
	.w4(32'hbb9ba68b),
	.w5(32'hbab5ce47),
	.w6(32'hba8042ae),
	.w7(32'hbae3e5f8),
	.w8(32'h3adca488),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13f546),
	.w1(32'h36ca8e94),
	.w2(32'h3bbf3d92),
	.w3(32'hb9c58ca3),
	.w4(32'h3a1a145a),
	.w5(32'h3b3ed342),
	.w6(32'hbabcd943),
	.w7(32'h3bdbffd5),
	.w8(32'h3b8678a0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9adb4),
	.w1(32'h3b2bb579),
	.w2(32'h3a941e69),
	.w3(32'hbb7c6ecd),
	.w4(32'h3b947045),
	.w5(32'h3b90ce30),
	.w6(32'hbbf814af),
	.w7(32'h3a39ad73),
	.w8(32'hbb367a95),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aebe3),
	.w1(32'h3babc532),
	.w2(32'h3b546644),
	.w3(32'hbacbbbec),
	.w4(32'h3bba068c),
	.w5(32'h3c2431d7),
	.w6(32'h3999cbe1),
	.w7(32'hbb45d6e4),
	.w8(32'hbaa902c6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ce11),
	.w1(32'hbafccc4d),
	.w2(32'hbc1d4ed0),
	.w3(32'h3c02a272),
	.w4(32'hbb38cb68),
	.w5(32'hbb0af4f0),
	.w6(32'hbb908cf0),
	.w7(32'hbc373012),
	.w8(32'hbc3359a1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94fe7),
	.w1(32'hbbbe9a04),
	.w2(32'hbc25a951),
	.w3(32'hbbbf371f),
	.w4(32'hbae8253d),
	.w5(32'hbbcf7ad2),
	.w6(32'hbc0ffa0b),
	.w7(32'hbad66a95),
	.w8(32'hbc0f840e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e24c),
	.w1(32'hbb7112bb),
	.w2(32'hbad15678),
	.w3(32'h3b996cf8),
	.w4(32'hbbd21e11),
	.w5(32'hbb6dba6a),
	.w6(32'h3b907427),
	.w7(32'hbb220207),
	.w8(32'hba731b80),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd406c5),
	.w1(32'hbae33a6a),
	.w2(32'hba7202d5),
	.w3(32'hb9f6bd6b),
	.w4(32'hbaf5dc0e),
	.w5(32'hbbac1ae4),
	.w6(32'h3b695a93),
	.w7(32'hbb1cb956),
	.w8(32'hbad1c787),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb203874),
	.w1(32'h39a6fb08),
	.w2(32'h391fa61e),
	.w3(32'hbb8924f4),
	.w4(32'hbacb0447),
	.w5(32'hbb886344),
	.w6(32'hbb870e07),
	.w7(32'h3a3c8680),
	.w8(32'h3a3a13e4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9a05),
	.w1(32'hbb27626b),
	.w2(32'hb9b10767),
	.w3(32'h3ac866bc),
	.w4(32'hba3b916f),
	.w5(32'h3a691438),
	.w6(32'h3b00f822),
	.w7(32'h3ac21a5f),
	.w8(32'h3b7de11c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0dc56),
	.w1(32'hbc1ba6f9),
	.w2(32'hbcaef8c5),
	.w3(32'hbb8fa247),
	.w4(32'hbbeef6df),
	.w5(32'hbc451cbe),
	.w6(32'hbb0a6cb6),
	.w7(32'hbc0e5858),
	.w8(32'hbc26e503),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcb2e9),
	.w1(32'h3ac28394),
	.w2(32'hbce2b343),
	.w3(32'hba9de345),
	.w4(32'h3c7fd9e4),
	.w5(32'hbc7013f8),
	.w6(32'hbcdbef3f),
	.w7(32'hbb599938),
	.w8(32'hbd04906c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca30f8c),
	.w1(32'hbb858fc6),
	.w2(32'hbcbf128d),
	.w3(32'hbc0bd064),
	.w4(32'h3c141cdb),
	.w5(32'hbc7fe439),
	.w6(32'hbd0ad322),
	.w7(32'hbc5d2233),
	.w8(32'hbcee9dab),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1485b0),
	.w1(32'h3cb5085b),
	.w2(32'hbc497933),
	.w3(32'hbc587c28),
	.w4(32'h3d4746e3),
	.w5(32'h3cb9c900),
	.w6(32'hbd215954),
	.w7(32'h3cebbd00),
	.w8(32'hbbd70a5d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996fe9),
	.w1(32'hba18127c),
	.w2(32'hbab38f07),
	.w3(32'h3a5290bf),
	.w4(32'hbb0d284e),
	.w5(32'hbacf106c),
	.w6(32'h3adc5ed6),
	.w7(32'hbaf2b9fc),
	.w8(32'hbb147849),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85a6136),
	.w1(32'h393fe79a),
	.w2(32'h39ee6110),
	.w3(32'hba2818fa),
	.w4(32'hba5d7730),
	.w5(32'hb8cb2f91),
	.w6(32'hb96fc47c),
	.w7(32'h3a93ad22),
	.w8(32'h3ac7bdbf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45c67f),
	.w1(32'h395e4545),
	.w2(32'h3a807878),
	.w3(32'h39db25e7),
	.w4(32'h38eda722),
	.w5(32'h3abb1a49),
	.w6(32'h3a4bfbc6),
	.w7(32'h3a92a6a9),
	.w8(32'h3aa15ab0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb80b3),
	.w1(32'h3b59b371),
	.w2(32'hbb210424),
	.w3(32'h3a880040),
	.w4(32'h3b006db3),
	.w5(32'hbb129453),
	.w6(32'h39dd852e),
	.w7(32'h399727ba),
	.w8(32'hbb309cbf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398253fa),
	.w1(32'hba6e8491),
	.w2(32'hba02effd),
	.w3(32'h3a4ee455),
	.w4(32'hbb06008e),
	.w5(32'hbb1327b5),
	.w6(32'hb87e26c3),
	.w7(32'hbac2e5d9),
	.w8(32'hba4f0837),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2120),
	.w1(32'hbb060bcb),
	.w2(32'hbc07d03a),
	.w3(32'hbb490bf3),
	.w4(32'hbacb0aca),
	.w5(32'hbbbcb52d),
	.w6(32'hbb5d178e),
	.w7(32'h38381527),
	.w8(32'hbb4637ac),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6062fb),
	.w1(32'hb82b24ee),
	.w2(32'hbc425ff3),
	.w3(32'hbbd956d4),
	.w4(32'h3bb3d3b7),
	.w5(32'hbafd8edf),
	.w6(32'hbc543140),
	.w7(32'hbad3c598),
	.w8(32'hbc7d8807),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc892710),
	.w1(32'hbb37ae78),
	.w2(32'hbc58a2ef),
	.w3(32'hbbda6290),
	.w4(32'h3c268e4e),
	.w5(32'h3b8adec1),
	.w6(32'hbc289f74),
	.w7(32'h3c0166c6),
	.w8(32'hbb1e5af3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4e35),
	.w1(32'hbb47d406),
	.w2(32'hbc85a45b),
	.w3(32'hbae5fc07),
	.w4(32'h3b7eda46),
	.w5(32'hbc048ce8),
	.w6(32'hbbb58af4),
	.w7(32'h3ad4ef51),
	.w8(32'hbc1cf2d5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e3c9b),
	.w1(32'h3afbc690),
	.w2(32'hbc1783c6),
	.w3(32'h3a8dd86e),
	.w4(32'h3aeb58bb),
	.w5(32'hbbcaae32),
	.w6(32'hba0bea35),
	.w7(32'h3b945d12),
	.w8(32'hbb3e9579),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd32f4),
	.w1(32'hba983610),
	.w2(32'hbc2b952d),
	.w3(32'hbaeac69c),
	.w4(32'h3bc75dd0),
	.w5(32'hbb977d03),
	.w6(32'hbbb0e1d4),
	.w7(32'h3b83dfc8),
	.w8(32'hbb59051b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfddd3),
	.w1(32'hb96558f5),
	.w2(32'hbc6a426d),
	.w3(32'h3b0b9b14),
	.w4(32'hbacaccde),
	.w5(32'hbc4c8fbf),
	.w6(32'hb8edcd4e),
	.w7(32'h3a7cb254),
	.w8(32'hbc125702),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1b848),
	.w1(32'hba4f4968),
	.w2(32'hb9ac370e),
	.w3(32'h39d28f55),
	.w4(32'hb99e711c),
	.w5(32'hb9e5f2c9),
	.w6(32'h39c311fc),
	.w7(32'h39965554),
	.w8(32'h3a66954a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399890a8),
	.w1(32'h3a02bb68),
	.w2(32'h39459587),
	.w3(32'h39d76b44),
	.w4(32'h39f72ae6),
	.w5(32'hb8bad48c),
	.w6(32'h3a61105c),
	.w7(32'hb875d835),
	.w8(32'hba1dfbdb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87acae),
	.w1(32'hb91a489e),
	.w2(32'h39fade81),
	.w3(32'h382921ef),
	.w4(32'hba8300a4),
	.w5(32'h3a74be25),
	.w6(32'h3ab5adc8),
	.w7(32'hb9c51fff),
	.w8(32'hb8016280),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a34c4),
	.w1(32'h3ac7c464),
	.w2(32'h3b1beadb),
	.w3(32'hbaad204e),
	.w4(32'h3b100a8e),
	.w5(32'h3aeffe5a),
	.w6(32'hba7ee999),
	.w7(32'h38ecb99a),
	.w8(32'h3ac5f3f9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd765c2),
	.w1(32'hbbbe1d72),
	.w2(32'hbafa9322),
	.w3(32'hbcaa8d45),
	.w4(32'h3a0b867e),
	.w5(32'h3bdba8ea),
	.w6(32'hbcce4dbd),
	.w7(32'h3939cf46),
	.w8(32'hb9c2228e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d96269),
	.w1(32'h3b420029),
	.w2(32'hb83ab8a7),
	.w3(32'h39f55713),
	.w4(32'h3bac88a0),
	.w5(32'h3b328205),
	.w6(32'hbb39f485),
	.w7(32'h3b1ae682),
	.w8(32'hb9ab557b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9000ec),
	.w1(32'hbbfeea92),
	.w2(32'hbc83e2d4),
	.w3(32'hbbc80e96),
	.w4(32'h39b7af0c),
	.w5(32'hbc0551ae),
	.w6(32'hbc45a3b7),
	.w7(32'hbb21a11a),
	.w8(32'hbc606a3f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8f7c2),
	.w1(32'hbc1cb94a),
	.w2(32'hbc9528a5),
	.w3(32'hbccd14d8),
	.w4(32'hbbfd47ab),
	.w5(32'hbc7d101f),
	.w6(32'hbceeece2),
	.w7(32'hbc4d0ba3),
	.w8(32'hbca3ab6a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9e03),
	.w1(32'h3b4e2dd4),
	.w2(32'h3aec1e68),
	.w3(32'hbc10eaef),
	.w4(32'h3a836793),
	.w5(32'h3b2d6bfd),
	.w6(32'hbc9d5858),
	.w7(32'hba284833),
	.w8(32'hbbb9cf9d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc184038),
	.w1(32'hbaf343d4),
	.w2(32'hbc9329af),
	.w3(32'hbbcc9902),
	.w4(32'h3bfcd6ec),
	.w5(32'hbbdec28d),
	.w6(32'hbc0566d9),
	.w7(32'h3bed8e0a),
	.w8(32'hbc12b072),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b52e9),
	.w1(32'h3c61a551),
	.w2(32'h3af850f7),
	.w3(32'h3b37d9aa),
	.w4(32'h3c7b16d2),
	.w5(32'h3ba6f498),
	.w6(32'hbb545dd6),
	.w7(32'h3c709406),
	.w8(32'h3bf83dbe),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6be69),
	.w1(32'hbc1eeb85),
	.w2(32'hbcbc52bf),
	.w3(32'hbc41190e),
	.w4(32'h3a95e0e2),
	.w5(32'hbc124c04),
	.w6(32'hbc9ced9a),
	.w7(32'hbb1da73f),
	.w8(32'hbc8259a4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83b895),
	.w1(32'hbbccb286),
	.w2(32'hbc4b29ff),
	.w3(32'hbc4e088f),
	.w4(32'hbac76fbe),
	.w5(32'hbb220a85),
	.w6(32'hbc6abbb8),
	.w7(32'hbb0c0aa7),
	.w8(32'hbbe1c08a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc87b4f),
	.w1(32'h3b6d25be),
	.w2(32'h3b9e4f62),
	.w3(32'hbc771213),
	.w4(32'h3c1a3b0e),
	.w5(32'h3c0b02dd),
	.w6(32'hbcb0d801),
	.w7(32'h3bb0dab3),
	.w8(32'h3bc1b9b3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34803),
	.w1(32'hb9e553af),
	.w2(32'h3a2752b0),
	.w3(32'h39e5fffb),
	.w4(32'hbab1b502),
	.w5(32'hba094c26),
	.w6(32'h3a3ea875),
	.w7(32'hb9c1870a),
	.w8(32'h3a055408),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6be4af),
	.w1(32'hbba3a42a),
	.w2(32'hbcd5ccca),
	.w3(32'hbbca1b77),
	.w4(32'h3bf1b1b2),
	.w5(32'hbc18ff63),
	.w6(32'hbc6a0875),
	.w7(32'hbabfb833),
	.w8(32'hbc8b30ce),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233ff0),
	.w1(32'hba36d624),
	.w2(32'hbc934332),
	.w3(32'hbba0af4f),
	.w4(32'h3b9486a0),
	.w5(32'hbc301032),
	.w6(32'hbc1119b4),
	.w7(32'h3b0898c7),
	.w8(32'hbc34dae3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7616e9),
	.w1(32'h3ad1e2dc),
	.w2(32'hbccadc05),
	.w3(32'hbb1a69da),
	.w4(32'h3ca6596d),
	.w5(32'hbaef4adc),
	.w6(32'hbb9138ee),
	.w7(32'h3c6b6f84),
	.w8(32'hbc7ab9c5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8b5b6f),
	.w1(32'h3b848c83),
	.w2(32'h3c86de9a),
	.w3(32'hbd3ced74),
	.w4(32'h3cb96304),
	.w5(32'h3cb66383),
	.w6(32'hbd6dda2b),
	.w7(32'h3aa053c5),
	.w8(32'hbb12d256),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc933fef),
	.w1(32'h3abe2d49),
	.w2(32'hbc9f652d),
	.w3(32'hbb337ce8),
	.w4(32'h3c647a9a),
	.w5(32'hbac0c16c),
	.w6(32'hbc6f046e),
	.w7(32'h3c02a87c),
	.w8(32'hbbdd3eb8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e3a80),
	.w1(32'hbbc10210),
	.w2(32'hbc94fb4c),
	.w3(32'hbc54ad4b),
	.w4(32'hba1cd325),
	.w5(32'hbc4e6f12),
	.w6(32'hbb69db9e),
	.w7(32'h3bdb781b),
	.w8(32'hbc328d25),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc84d),
	.w1(32'h3a83c2dd),
	.w2(32'h3aa1329f),
	.w3(32'h391fb6a7),
	.w4(32'h399671a6),
	.w5(32'h3afea1ed),
	.w6(32'h3ad653eb),
	.w7(32'h3a9951e2),
	.w8(32'h3b29b2d4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf942e0),
	.w1(32'hbc55c439),
	.w2(32'hbcd6641a),
	.w3(32'hbca6dad5),
	.w4(32'h3b574543),
	.w5(32'hbc1b84dc),
	.w6(32'hbc61784c),
	.w7(32'h3c095f5d),
	.w8(32'hbba5b5aa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b688f),
	.w1(32'h3c02841a),
	.w2(32'hbbb4cd47),
	.w3(32'h3a1e8586),
	.w4(32'h3c02d291),
	.w5(32'hbbbb1e0d),
	.w6(32'hba0845f1),
	.w7(32'h3c259176),
	.w8(32'hbb831e3a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39901fc8),
	.w1(32'h3a9edac0),
	.w2(32'hba4c556e),
	.w3(32'h3980db57),
	.w4(32'h3a8053de),
	.w5(32'hb90cf7c2),
	.w6(32'h39df9ddf),
	.w7(32'h39e008a5),
	.w8(32'h39545d8e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7e530),
	.w1(32'hbb8e4570),
	.w2(32'hbb67e1e4),
	.w3(32'hbb421597),
	.w4(32'hba897e51),
	.w5(32'hbaea961b),
	.w6(32'hbba71184),
	.w7(32'hbaf72709),
	.w8(32'hbb5a14cf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15752c),
	.w1(32'hbb6d0e05),
	.w2(32'hbc795595),
	.w3(32'hbb4cf058),
	.w4(32'h3adfadf0),
	.w5(32'hbbcdddb1),
	.w6(32'hbbf71a45),
	.w7(32'hbb594c81),
	.w8(32'hbc613550),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6b2f),
	.w1(32'h3b2a5d9d),
	.w2(32'hbbfe11cb),
	.w3(32'hba1a1d6e),
	.w4(32'h3c1cb385),
	.w5(32'h3b6ffa3f),
	.w6(32'hbc0e3444),
	.w7(32'h3bb3fead),
	.w8(32'hb904fdf4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82d10d),
	.w1(32'hbae429b7),
	.w2(32'h3aaa0bdf),
	.w3(32'hbc7200d2),
	.w4(32'h39878bcc),
	.w5(32'h3b346b08),
	.w6(32'hbcb0be0d),
	.w7(32'hbbe11fd4),
	.w8(32'hbbaa7ff2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66da67),
	.w1(32'hbacfe403),
	.w2(32'hbc26289d),
	.w3(32'hbbf13669),
	.w4(32'h3ba7bf25),
	.w5(32'h3a7a5c70),
	.w6(32'hbc327f6c),
	.w7(32'h39c27a63),
	.w8(32'hbbbd94e1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30747b),
	.w1(32'h3bbd0cdb),
	.w2(32'h39992d22),
	.w3(32'hbb4edd67),
	.w4(32'h3c06a24f),
	.w5(32'h3b1982eb),
	.w6(32'hbc36b1b7),
	.w7(32'h3a943676),
	.w8(32'hbc168fa3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803801),
	.w1(32'hbbdb43f7),
	.w2(32'hbc9185e7),
	.w3(32'hbb6f98a6),
	.w4(32'h39da0519),
	.w5(32'hbc2a94b9),
	.w6(32'hbb169921),
	.w7(32'hba2c1aac),
	.w8(32'hbc364169),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5aa80),
	.w1(32'h3aed68ac),
	.w2(32'hbbf60f36),
	.w3(32'hba416cab),
	.w4(32'h3be3b9dc),
	.w5(32'hbad8a746),
	.w6(32'hbbf42a87),
	.w7(32'h3ba1bcfc),
	.w8(32'hbb7f97af),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a4dba),
	.w1(32'h3adfe7f8),
	.w2(32'h3a9ed1d6),
	.w3(32'hbaa8655a),
	.w4(32'h3aadfe90),
	.w5(32'h3a23cb81),
	.w6(32'hbaa137ea),
	.w7(32'h3abc7d8f),
	.w8(32'h3813b49b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad396e4),
	.w1(32'hbaa2869a),
	.w2(32'h381aa2eb),
	.w3(32'hba1c54c6),
	.w4(32'hba20d529),
	.w5(32'hb8bbd985),
	.w6(32'hba24fd8f),
	.w7(32'hbad93e77),
	.w8(32'hba77b752),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b4d6),
	.w1(32'h3ac2ed50),
	.w2(32'h39d580d2),
	.w3(32'hb9812fcb),
	.w4(32'h3a60049d),
	.w5(32'h3a1569d8),
	.w6(32'h38741ee3),
	.w7(32'h3b56611c),
	.w8(32'h3b277910),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a897bb9),
	.w1(32'h39d7ca20),
	.w2(32'h3ac956ca),
	.w3(32'h3a2cf12b),
	.w4(32'hb89e3d9f),
	.w5(32'h3ad2784c),
	.w6(32'hb9772965),
	.w7(32'h3a2a0e49),
	.w8(32'h3a8b7c08),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fccd2),
	.w1(32'h3a9bdc9c),
	.w2(32'hbc227dc3),
	.w3(32'hba3db910),
	.w4(32'h3c2373c8),
	.w5(32'hbaa9ef9a),
	.w6(32'hbbfa0907),
	.w7(32'h3bd9b5dc),
	.w8(32'hbbb1aee3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03461b),
	.w1(32'h3a274e5b),
	.w2(32'h3909cf73),
	.w3(32'hbb15361c),
	.w4(32'h3b23115b),
	.w5(32'h3a47e004),
	.w6(32'hbabc81f6),
	.w7(32'h3b1dd31a),
	.w8(32'h384c84a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319c47),
	.w1(32'hba3ac64e),
	.w2(32'hbc0ffc32),
	.w3(32'hb9ab5bc6),
	.w4(32'hbab8eb1c),
	.w5(32'hbba0a60f),
	.w6(32'h3acc4990),
	.w7(32'hbad75988),
	.w8(32'hbbd8cfc0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc3edb),
	.w1(32'hbb9e07f1),
	.w2(32'h3a2793a8),
	.w3(32'hbc9f8107),
	.w4(32'h3b1ee62d),
	.w5(32'h3bc300be),
	.w6(32'hbcee3ab9),
	.w7(32'hbb9a03ed),
	.w8(32'hbb8794b3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59e17),
	.w1(32'hb9c8ec5d),
	.w2(32'hba301c10),
	.w3(32'h3a1c5e64),
	.w4(32'h36f6c03b),
	.w5(32'hb8c68877),
	.w6(32'h3ae93a48),
	.w7(32'hb8fbec70),
	.w8(32'h39982381),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a28d),
	.w1(32'h3a8a5709),
	.w2(32'hba51b3f4),
	.w3(32'h3a8bd158),
	.w4(32'h3a8a2049),
	.w5(32'h3a49ef5d),
	.w6(32'h38b2d2a3),
	.w7(32'h3ab47077),
	.w8(32'h3901e78f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958d0eb),
	.w1(32'h39b7fedb),
	.w2(32'hb99fec05),
	.w3(32'hbaa968d0),
	.w4(32'hba8b63b9),
	.w5(32'hbac5e235),
	.w6(32'hb8fd1590),
	.w7(32'hb8d6191b),
	.w8(32'h3a19229a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4c7f2),
	.w1(32'hbb848f82),
	.w2(32'hbb1cc5a3),
	.w3(32'hbb9f3b08),
	.w4(32'hbb9973b1),
	.w5(32'hba955786),
	.w6(32'hbbb1a38b),
	.w7(32'hbbc88bd3),
	.w8(32'hbbbc596d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbb39f),
	.w1(32'hbc1c7c28),
	.w2(32'hbc8706cf),
	.w3(32'h3c15203e),
	.w4(32'hbace48d2),
	.w5(32'hbc80f430),
	.w6(32'hba1ba547),
	.w7(32'hbc4840fb),
	.w8(32'hbca313cd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89dc94),
	.w1(32'hbbb66d5e),
	.w2(32'hbcaeb5a6),
	.w3(32'hb9e7ae73),
	.w4(32'h3b29c42b),
	.w5(32'hbc432f2a),
	.w6(32'hbb360d07),
	.w7(32'hb9c81dde),
	.w8(32'hbc42e218),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c5b80),
	.w1(32'hba9ec0f0),
	.w2(32'hbb10571f),
	.w3(32'hb992b70c),
	.w4(32'hba42b76b),
	.w5(32'h3a7dcb55),
	.w6(32'h39f433c7),
	.w7(32'h393b728a),
	.w8(32'hb8929ab0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8596),
	.w1(32'h3a183721),
	.w2(32'hbb9d07de),
	.w3(32'hbb1fc0b3),
	.w4(32'h3b43a42c),
	.w5(32'hbaa91936),
	.w6(32'hbbecf86f),
	.w7(32'hbb21dc02),
	.w8(32'hbbbc65e3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a402),
	.w1(32'h395d65f0),
	.w2(32'hbb806fa8),
	.w3(32'hbbae86f0),
	.w4(32'h3acf69f5),
	.w5(32'hbb3b952a),
	.w6(32'hbc091a1b),
	.w7(32'h3b4c6dab),
	.w8(32'hbb3195f2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba184cc),
	.w1(32'hba9f53eb),
	.w2(32'hbc172b08),
	.w3(32'h39b9aadd),
	.w4(32'h3b832e0b),
	.w5(32'hbb13e00b),
	.w6(32'hbbae94b2),
	.w7(32'h39d6a33e),
	.w8(32'hbba960f2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7847c4),
	.w1(32'hbc1d9d02),
	.w2(32'hbc8e0a8b),
	.w3(32'hbc14966f),
	.w4(32'h3b0bbc9e),
	.w5(32'hbb9b49a9),
	.w6(32'hbc1eaabb),
	.w7(32'hba91f3b5),
	.w8(32'hbbdb9d5c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b844),
	.w1(32'hbb5f568d),
	.w2(32'hbcbdd3f1),
	.w3(32'hbb17efcb),
	.w4(32'h3a50232b),
	.w5(32'hbc8b40c5),
	.w6(32'hbb3d480c),
	.w7(32'h3a9b30d5),
	.w8(32'hbc7db24e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc821ca9),
	.w1(32'hb918c8a0),
	.w2(32'hbb6da302),
	.w3(32'hbc0c88d1),
	.w4(32'h3bc86d5e),
	.w5(32'h3b72cd83),
	.w6(32'hbc7750df),
	.w7(32'h3b2de8b9),
	.w8(32'hbb300fce),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc544247),
	.w1(32'hbbc4d0b2),
	.w2(32'hbc602c15),
	.w3(32'hbb876232),
	.w4(32'h3abb8987),
	.w5(32'hbb882f03),
	.w6(32'hbb946eed),
	.w7(32'hba6a31b2),
	.w8(32'hbc16b650),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86afef),
	.w1(32'hbc02c534),
	.w2(32'hbcb7d760),
	.w3(32'hbc1de6f5),
	.w4(32'hba068d11),
	.w5(32'hbc74a191),
	.w6(32'hbc229773),
	.w7(32'h39e8a68a),
	.w8(32'hbc55693c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98e5c4),
	.w1(32'hb8e98275),
	.w2(32'h3a619e8a),
	.w3(32'hbc05cb59),
	.w4(32'h3bce7221),
	.w5(32'h3bfa6693),
	.w6(32'hbc7fe842),
	.w7(32'h3abbe8fa),
	.w8(32'hba4ae495),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f4f9),
	.w1(32'hbadbe46e),
	.w2(32'hbc413c1d),
	.w3(32'hbb9b8188),
	.w4(32'h3b23c228),
	.w5(32'hbbd05779),
	.w6(32'hbbc2c686),
	.w7(32'hba35e2a5),
	.w8(32'hbc2ffd42),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4f8da),
	.w1(32'h3926e0b2),
	.w2(32'hbb9c3eff),
	.w3(32'h3ab89b19),
	.w4(32'h3b32964f),
	.w5(32'hba846c2d),
	.w6(32'hbac652d8),
	.w7(32'h3ac97ce4),
	.w8(32'hbb2fe9d3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5d27d),
	.w1(32'h3c0efa31),
	.w2(32'h3c51a92a),
	.w3(32'hbcad932e),
	.w4(32'h3c07465e),
	.w5(32'h3c737e2d),
	.w6(32'hbcd2d01e),
	.w7(32'h3a8c30b7),
	.w8(32'h3bd9be34),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc729998),
	.w1(32'hbb8b1310),
	.w2(32'h3a803a6c),
	.w3(32'hbc3384a4),
	.w4(32'hbb0fc68a),
	.w5(32'h3b79607f),
	.w6(32'hbc726566),
	.w7(32'hbb98b22f),
	.w8(32'hbb807dd9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e021d0),
	.w1(32'hb9c5be8a),
	.w2(32'hb9c4a698),
	.w3(32'hba79b8cc),
	.w4(32'hba94fd69),
	.w5(32'hb9d71083),
	.w6(32'h3a0ab2a0),
	.w7(32'hb9fad62e),
	.w8(32'hba1695e5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643b9a),
	.w1(32'h3a8ee374),
	.w2(32'h3a8e147f),
	.w3(32'hba34282c),
	.w4(32'h3a3637b6),
	.w5(32'h3a43df2a),
	.w6(32'h397c00a5),
	.w7(32'h3b0143d1),
	.w8(32'h3aaf97f0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718b83),
	.w1(32'hbb01891e),
	.w2(32'hbb178af5),
	.w3(32'hbb84df93),
	.w4(32'h3ae26d5c),
	.w5(32'h3ae080e8),
	.w6(32'hbb3a7cc9),
	.w7(32'h3a7f75f3),
	.w8(32'h3b0d2f88),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca473d),
	.w1(32'hbb541d74),
	.w2(32'h3a7d28dd),
	.w3(32'hbc6e0386),
	.w4(32'h3b9f3829),
	.w5(32'h3c05939f),
	.w6(32'hbc9f812d),
	.w7(32'h3a1f6ce8),
	.w8(32'hbb3ea236),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffc6cc),
	.w1(32'h3b0e17dc),
	.w2(32'hbc8a4c1e),
	.w3(32'h3ac8a8b8),
	.w4(32'h3c538bd3),
	.w5(32'hbb95d975),
	.w6(32'hba235a04),
	.w7(32'h3c0677c2),
	.w8(32'hbc09bedd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89894ef),
	.w1(32'h3800db1a),
	.w2(32'hba153950),
	.w3(32'h3a8f0b33),
	.w4(32'hb9ceea55),
	.w5(32'hb9b23304),
	.w6(32'h3a8257d2),
	.w7(32'h395a6768),
	.w8(32'h3a450e21),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf72108),
	.w1(32'hbbc15614),
	.w2(32'hbcae08be),
	.w3(32'hba9dd457),
	.w4(32'h3b9066da),
	.w5(32'hbc5554d3),
	.w6(32'hbbb193c6),
	.w7(32'h3aacd618),
	.w8(32'hbc4abddf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068a86),
	.w1(32'hbb1e2416),
	.w2(32'hbc0d2ecd),
	.w3(32'hbb9cc4dc),
	.w4(32'h3aec0e45),
	.w5(32'hbb33d080),
	.w6(32'hbbd5d35c),
	.w7(32'h3a853b77),
	.w8(32'hbb86b633),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be881),
	.w1(32'hbb0808c7),
	.w2(32'hbc98425b),
	.w3(32'hbba30808),
	.w4(32'h3a2bca88),
	.w5(32'hbc1e2446),
	.w6(32'h3ae9d74b),
	.w7(32'h3b9e46f8),
	.w8(32'hbc11d80d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050feb),
	.w1(32'h3be03d13),
	.w2(32'hbc0c7001),
	.w3(32'h39543c1c),
	.w4(32'h3c83f7e2),
	.w5(32'h3af37e08),
	.w6(32'hbc40c645),
	.w7(32'h3c57cd5b),
	.w8(32'h3abcdc68),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cfea8),
	.w1(32'hbb88f071),
	.w2(32'hbb24a7cd),
	.w3(32'hbc5f574f),
	.w4(32'hbbb2d49e),
	.w5(32'hbb9a233c),
	.w6(32'hbc8324cf),
	.w7(32'hbbcd85f6),
	.w8(32'hbbde4541),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54f301),
	.w1(32'hb9076c08),
	.w2(32'h3aa5bd5c),
	.w3(32'h3b32e03d),
	.w4(32'hba38c5c2),
	.w5(32'h39aacd03),
	.w6(32'h3acefc69),
	.w7(32'hba60fd0a),
	.w8(32'h398b0d88),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b0161),
	.w1(32'h3b66e0d0),
	.w2(32'h3ae4375e),
	.w3(32'hbba90976),
	.w4(32'h3c09ff91),
	.w5(32'h3bce2a5f),
	.w6(32'hbc653c58),
	.w7(32'h3a8aef51),
	.w8(32'hbb392397),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd041cca),
	.w1(32'hbbecc025),
	.w2(32'hbbaca8d2),
	.w3(32'hbcc5f12c),
	.w4(32'hbbfabcf4),
	.w5(32'hbbcfd357),
	.w6(32'hbcef3d60),
	.w7(32'hbc1bfe32),
	.w8(32'hbc75927f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8282ba),
	.w1(32'h3c031864),
	.w2(32'h3acafa01),
	.w3(32'hbb0ed3ef),
	.w4(32'h3c214c20),
	.w5(32'h3b87a15f),
	.w6(32'hbc2acd3b),
	.w7(32'h3b9a11a8),
	.w8(32'hb9ec10cb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a9579),
	.w1(32'hb9378f89),
	.w2(32'hbb4e6255),
	.w3(32'hb9975213),
	.w4(32'hbb6cdf03),
	.w5(32'hbb6ffda4),
	.w6(32'hba5cf548),
	.w7(32'hbaab76f9),
	.w8(32'hbb8f0b51),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4ddf6),
	.w1(32'hbb2f75dc),
	.w2(32'hbaf2c71d),
	.w3(32'hbaa11df3),
	.w4(32'hbabdd73c),
	.w5(32'hbace70b4),
	.w6(32'hbadc0049),
	.w7(32'hbaada2c1),
	.w8(32'hbb275d88),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670bab),
	.w1(32'hbbbec402),
	.w2(32'hbc472470),
	.w3(32'hbc0fc8bd),
	.w4(32'h397aad6d),
	.w5(32'hbbf8e24b),
	.w6(32'hbc36e6ef),
	.w7(32'hbb77b663),
	.w8(32'hbc2e200a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60e91),
	.w1(32'h3a7cf3c6),
	.w2(32'hbac38241),
	.w3(32'h3afc3d85),
	.w4(32'h3a1e9f54),
	.w5(32'hb9e0d2f2),
	.w6(32'h3addf46d),
	.w7(32'h3b3ed1c5),
	.w8(32'h3ad8cb6a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed3986),
	.w1(32'h3b040de5),
	.w2(32'hbb94262d),
	.w3(32'hb98df0bf),
	.w4(32'h3bdd88af),
	.w5(32'h3a23cb33),
	.w6(32'hbbb50dca),
	.w7(32'h3bb08a14),
	.w8(32'h3ae1910d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a14cf),
	.w1(32'h3ac23907),
	.w2(32'hb9abb79f),
	.w3(32'h3ae9cc14),
	.w4(32'h3af7fcc0),
	.w5(32'h3a13e444),
	.w6(32'h3b1587bc),
	.w7(32'h3b0833e5),
	.w8(32'h3aa6f5a8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0548e9),
	.w1(32'h3c1a654f),
	.w2(32'hbc35cf61),
	.w3(32'h3c113421),
	.w4(32'h3c190c1c),
	.w5(32'hbbee8815),
	.w6(32'h3a92808c),
	.w7(32'h3ba93940),
	.w8(32'hbc02b3ec),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4dadd),
	.w1(32'h3a2682d4),
	.w2(32'h3a615f82),
	.w3(32'h3a89c147),
	.w4(32'h39097b2a),
	.w5(32'h3a5c7b4e),
	.w6(32'h3b0a4263),
	.w7(32'h394256df),
	.w8(32'hba11e88c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993d274),
	.w1(32'h395f9063),
	.w2(32'h3abcc4a3),
	.w3(32'hb9b29df8),
	.w4(32'h37aa1b59),
	.w5(32'h3ac1e46b),
	.w6(32'hba238425),
	.w7(32'h37acf001),
	.w8(32'hb9087401),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f179c),
	.w1(32'hbb0aa371),
	.w2(32'hbb06b7fb),
	.w3(32'hbc44b9f7),
	.w4(32'h3b2372a8),
	.w5(32'h3af33bf9),
	.w6(32'hbc8f4992),
	.w7(32'hbb79cf67),
	.w8(32'hbbc981cb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1d89e),
	.w1(32'hbaa71f25),
	.w2(32'hbc809519),
	.w3(32'hbc30914d),
	.w4(32'h38e2a49a),
	.w5(32'hbcc128fd),
	.w6(32'hbc96ecab),
	.w7(32'hbb05d922),
	.w8(32'hbcd33b03),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f8f54),
	.w1(32'h3b8db00e),
	.w2(32'hb9eaf200),
	.w3(32'hba31d3fb),
	.w4(32'h3b61ee3f),
	.w5(32'hbaad8ee0),
	.w6(32'hbb9853d7),
	.w7(32'h3ae29d74),
	.w8(32'hbb409481),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40f08e),
	.w1(32'h3a8aac05),
	.w2(32'hbc48798b),
	.w3(32'hbb6a4658),
	.w4(32'h3c18656d),
	.w5(32'hbb875a14),
	.w6(32'hbbd364c2),
	.w7(32'h3bd0b507),
	.w8(32'hbbf19512),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b9e43),
	.w1(32'hb8062108),
	.w2(32'hbb63ef78),
	.w3(32'hbb88bed4),
	.w4(32'hba3b7a8c),
	.w5(32'hbb12415e),
	.w6(32'hbb4bd210),
	.w7(32'h3a996481),
	.w8(32'h3a4c95b5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c6ed7),
	.w1(32'h3ab14884),
	.w2(32'hbcf3123e),
	.w3(32'hbba92af0),
	.w4(32'h3c49a627),
	.w5(32'hbc5ad485),
	.w6(32'hbc3390e4),
	.w7(32'h3ba13752),
	.w8(32'hbcaa89c5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc725a9a),
	.w1(32'hbaba46fd),
	.w2(32'hbc9f792b),
	.w3(32'hbc13f722),
	.w4(32'h3bc6f534),
	.w5(32'hbbcbd56e),
	.w6(32'hbc71dcae),
	.w7(32'h3afb4945),
	.w8(32'hbc516c89),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d36fa),
	.w1(32'hbbb546bc),
	.w2(32'hbce14df6),
	.w3(32'h3998f339),
	.w4(32'h3a571479),
	.w5(32'hbca2ee5d),
	.w6(32'hbb3d0ea0),
	.w7(32'hba145df5),
	.w8(32'hbc93c4d4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cdd70),
	.w1(32'hb9de6d7b),
	.w2(32'h39b28b35),
	.w3(32'hbab97a87),
	.w4(32'h381181ce),
	.w5(32'h3add4fd3),
	.w6(32'hbb15a593),
	.w7(32'h39e836a8),
	.w8(32'h39e03a84),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ca76),
	.w1(32'hbbd561f8),
	.w2(32'hbc304a21),
	.w3(32'hbb5d8f75),
	.w4(32'hbb519bf7),
	.w5(32'hbbdad85f),
	.w6(32'hbb0966b9),
	.w7(32'hba6cafee),
	.w8(32'hbbcaacca),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef363f),
	.w1(32'h39e9fb2e),
	.w2(32'h3a8350b7),
	.w3(32'hb9e91853),
	.w4(32'h3ac3d7a0),
	.w5(32'h3a840854),
	.w6(32'hb87d541c),
	.w7(32'h3aab62f6),
	.w8(32'h3a9d5cfa),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1e51c),
	.w1(32'h3b4a8655),
	.w2(32'hbbbc8637),
	.w3(32'h3b9bead3),
	.w4(32'h3b772e64),
	.w5(32'hbae668e0),
	.w6(32'h3a7eb4eb),
	.w7(32'h3ae1dcbb),
	.w8(32'hbba082c7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a873b),
	.w1(32'h3a36f17a),
	.w2(32'h3887ce0d),
	.w3(32'hbb683f83),
	.w4(32'hba843e9b),
	.w5(32'h39c0b8f4),
	.w6(32'hbb8e80fc),
	.w7(32'hba905214),
	.w8(32'hbb20d879),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03922),
	.w1(32'h3a59f588),
	.w2(32'hbc470117),
	.w3(32'hbba6fcc1),
	.w4(32'h3bc8a5ac),
	.w5(32'hbb6d50ef),
	.w6(32'hbbf27a5a),
	.w7(32'h3b510516),
	.w8(32'hbbe21bc9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d082b5),
	.w1(32'h3a87f83b),
	.w2(32'hb8023596),
	.w3(32'h3a238a46),
	.w4(32'h39e6cbb1),
	.w5(32'h388c8781),
	.w6(32'h3ac09051),
	.w7(32'h3a357dd7),
	.w8(32'h39082daa),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39675775),
	.w1(32'hb8ffcf84),
	.w2(32'hba49e723),
	.w3(32'h3a58fa99),
	.w4(32'h39abbcbb),
	.w5(32'h39aeb5cf),
	.w6(32'h3a1f9515),
	.w7(32'h3ab0867f),
	.w8(32'hba3271c1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f00fb),
	.w1(32'h3ab71273),
	.w2(32'h3a2e9c06),
	.w3(32'hbb3adf17),
	.w4(32'h3bacc041),
	.w5(32'h3baf6f17),
	.w6(32'hbbb58641),
	.w7(32'h3a97ea2d),
	.w8(32'h39dd9402),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d584b),
	.w1(32'hbbdcbb45),
	.w2(32'hbc7e727c),
	.w3(32'hbc0de155),
	.w4(32'hbb8a7562),
	.w5(32'hbc3c465b),
	.w6(32'hbc6e2636),
	.w7(32'hbc1a4ee2),
	.w8(32'hbc873785),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb08177),
	.w1(32'h3b9ae29b),
	.w2(32'hbb7040fc),
	.w3(32'hbbe3a78d),
	.w4(32'h3ae5f9d1),
	.w5(32'hba0a4377),
	.w6(32'hbb3f3924),
	.w7(32'h3bda3381),
	.w8(32'hbb0a20ed),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9f5a),
	.w1(32'h393bcdad),
	.w2(32'hbae7b944),
	.w3(32'hbb27d352),
	.w4(32'h3a6ddbd9),
	.w5(32'hbace1ff7),
	.w6(32'hbb400f0a),
	.w7(32'h3a00fdef),
	.w8(32'hbb1a652e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeed157),
	.w1(32'hbbb47346),
	.w2(32'hbd2c4f2d),
	.w3(32'h3bb5c90a),
	.w4(32'h3bbb6070),
	.w5(32'hbcb12c67),
	.w6(32'h3c22e02a),
	.w7(32'h3b8195ec),
	.w8(32'hbcc45548),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1efe89),
	.w1(32'hbc200c57),
	.w2(32'hbc6732d6),
	.w3(32'hbd03da9d),
	.w4(32'hb9fab67e),
	.w5(32'hba26a29c),
	.w6(32'hbd08128b),
	.w7(32'hbb0f1652),
	.w8(32'hbbbf5af3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c6a16),
	.w1(32'h3a129186),
	.w2(32'hbabe0691),
	.w3(32'h3b0ad286),
	.w4(32'hb98abf63),
	.w5(32'hbb4acb43),
	.w6(32'h3a9da160),
	.w7(32'h39eb5273),
	.w8(32'hbb4ebded),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9209d7),
	.w1(32'hba1822a0),
	.w2(32'hba78db02),
	.w3(32'hba329db7),
	.w4(32'hb9f88d0a),
	.w5(32'hba963363),
	.w6(32'hb98c586a),
	.w7(32'hb9e68b39),
	.w8(32'hbac4e6a3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3366c7),
	.w1(32'h3aadf74b),
	.w2(32'h3a97d5f9),
	.w3(32'hba9cae51),
	.w4(32'h3a2515e8),
	.w5(32'hb99b8259),
	.w6(32'hbb11edde),
	.w7(32'h39741188),
	.w8(32'hba5cdfb1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ad4a7),
	.w1(32'h3a705fc6),
	.w2(32'h38cdd288),
	.w3(32'h3860ce6b),
	.w4(32'h3a669801),
	.w5(32'hb9128ffb),
	.w6(32'h38edfc78),
	.w7(32'h3aac29a2),
	.w8(32'h3a54a491),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac428a),
	.w1(32'hbaecfdf7),
	.w2(32'hbbaec58c),
	.w3(32'hbaa13904),
	.w4(32'hbb2c7957),
	.w5(32'hbba4fea7),
	.w6(32'hbb69a70f),
	.w7(32'hbb73ca7d),
	.w8(32'hbba77e4a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8298b6),
	.w1(32'hbba3a74f),
	.w2(32'hbc4d2169),
	.w3(32'hbbf26fc3),
	.w4(32'h3b54e216),
	.w5(32'hbbb930be),
	.w6(32'hbc485a40),
	.w7(32'h3a23bea6),
	.w8(32'hbc46c7f2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc903f7b),
	.w1(32'hba329132),
	.w2(32'hbc6dbe61),
	.w3(32'hbbbc6b45),
	.w4(32'h3c390d34),
	.w5(32'h3b84236c),
	.w6(32'hbc46b421),
	.w7(32'h3be4296f),
	.w8(32'hbabb7204),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d774f),
	.w1(32'h3b2f3302),
	.w2(32'hba0c95d8),
	.w3(32'hbb191bf5),
	.w4(32'h3b41680a),
	.w5(32'h3adb49ac),
	.w6(32'hbb946c4e),
	.w7(32'h37b4df4c),
	.w8(32'hbb27c0e1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0088),
	.w1(32'hbb631fc7),
	.w2(32'hbcb47f3a),
	.w3(32'hbb34abd5),
	.w4(32'h3c0f4199),
	.w5(32'hbc05aa93),
	.w6(32'hbc157645),
	.w7(32'h3b6f54ee),
	.w8(32'hbc69c431),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70a397),
	.w1(32'hbb50056b),
	.w2(32'hbbf494e4),
	.w3(32'h3a03a73b),
	.w4(32'hba7cbbb4),
	.w5(32'hbb9ba8fd),
	.w6(32'hba9d1a95),
	.w7(32'hbb2c4f09),
	.w8(32'hbbc66061),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94510c),
	.w1(32'hbad85dde),
	.w2(32'hbb14c2a8),
	.w3(32'hbadca952),
	.w4(32'hbb82823e),
	.w5(32'hbb327962),
	.w6(32'hba80e5f2),
	.w7(32'h3929e454),
	.w8(32'h3a920c16),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5afb87),
	.w1(32'hbb5e7632),
	.w2(32'h3aff409e),
	.w3(32'hbb23df5d),
	.w4(32'hbb45e91e),
	.w5(32'h3b18c536),
	.w6(32'hba110354),
	.w7(32'hba6a21a0),
	.w8(32'h3abca063),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b7807),
	.w1(32'h3a4a09e7),
	.w2(32'h3ad65d11),
	.w3(32'h3b3c1855),
	.w4(32'hb82f0b87),
	.w5(32'hb98fc4ea),
	.w6(32'h3b48c51a),
	.w7(32'h38c34774),
	.w8(32'h3a3c5186),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20b106),
	.w1(32'h3b72641a),
	.w2(32'hb9b278ca),
	.w3(32'hbb5ea44a),
	.w4(32'h3c12f168),
	.w5(32'h3ba0ac9e),
	.w6(32'hbc0cc81b),
	.w7(32'h3aadaee4),
	.w8(32'hba5e4565),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd33dae),
	.w1(32'h3b3860b1),
	.w2(32'hbaef11b0),
	.w3(32'hbc84bd9b),
	.w4(32'h3c02fd40),
	.w5(32'h3b0d79c8),
	.w6(32'hbcff5ee1),
	.w7(32'hbb4b2334),
	.w8(32'hbc3f41c8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97cc14),
	.w1(32'hb92548c1),
	.w2(32'hbc32e7d2),
	.w3(32'hbc2b98f0),
	.w4(32'h3bf0d558),
	.w5(32'hbb345c01),
	.w6(32'hbc8c463b),
	.w7(32'hba970748),
	.w8(32'hbc2fe612),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32ac8),
	.w1(32'hbb3a2f0d),
	.w2(32'hbb34fb47),
	.w3(32'hbbc92940),
	.w4(32'hbae7c376),
	.w5(32'hba18bca9),
	.w6(32'hbc12037b),
	.w7(32'hbb90ab83),
	.w8(32'hbbc9296d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbf0e3),
	.w1(32'hbb1d70a3),
	.w2(32'hbc0c3a5c),
	.w3(32'hbc78cf1a),
	.w4(32'h3c3259a4),
	.w5(32'h3b80f91d),
	.w6(32'hbcbeaa5e),
	.w7(32'hb9e24885),
	.w8(32'hbc013201),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57241b),
	.w1(32'hb5c1ae74),
	.w2(32'hbc4805f4),
	.w3(32'hbabf180a),
	.w4(32'h3b75660c),
	.w5(32'hbbdfa306),
	.w6(32'hbb9c2001),
	.w7(32'h3adab4d3),
	.w8(32'hbbaf479d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134877),
	.w1(32'h3c099d21),
	.w2(32'hbc8f5cf3),
	.w3(32'hba75c792),
	.w4(32'h3c95ff7f),
	.w5(32'hba3f986a),
	.w6(32'hbb6357dd),
	.w7(32'h3c8c4a8e),
	.w8(32'hbbe97c0d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803832),
	.w1(32'hb9aa74ee),
	.w2(32'h39b9103b),
	.w3(32'h3b6f02f1),
	.w4(32'h382ce89f),
	.w5(32'h39c7d0ce),
	.w6(32'h3b83c45e),
	.w7(32'h39994f68),
	.w8(32'h3a0cd430),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bca8d),
	.w1(32'hb9a02461),
	.w2(32'h39df5d5b),
	.w3(32'hb897cfb4),
	.w4(32'hba87824b),
	.w5(32'hba5bc0bf),
	.w6(32'hb9d289ed),
	.w7(32'h395d4a1a),
	.w8(32'h3a3fc3da),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8293e0),
	.w1(32'h3b26d494),
	.w2(32'hbc5bb37f),
	.w3(32'hb9ef43a8),
	.w4(32'h3c4d00d5),
	.w5(32'hbbc94c0b),
	.w6(32'hbc832110),
	.w7(32'hb9e32709),
	.w8(32'hbca7b58b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80525f),
	.w1(32'hb94d00dd),
	.w2(32'hbcc52b23),
	.w3(32'hbba6bfdb),
	.w4(32'h3c014d50),
	.w5(32'hbc9ba388),
	.w6(32'hbc57ee94),
	.w7(32'h3b1cbe37),
	.w8(32'hbca6c71f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0be66),
	.w1(32'hba50734d),
	.w2(32'hbc589a2e),
	.w3(32'hbbbe2727),
	.w4(32'h3c3ab2a7),
	.w5(32'hbb98532a),
	.w6(32'hbc815173),
	.w7(32'h3aebf522),
	.w8(32'hbc50c570),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf314a),
	.w1(32'hbb719f87),
	.w2(32'hbb3d1b93),
	.w3(32'hbc082358),
	.w4(32'hbc0180bc),
	.w5(32'hbb51e0b3),
	.w6(32'h38810b41),
	.w7(32'h3a9f523f),
	.w8(32'hbade1f0b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97dc2f),
	.w1(32'hbae945c6),
	.w2(32'hba9e9dae),
	.w3(32'h3a01eb2d),
	.w4(32'hbb04ad2f),
	.w5(32'hba9c9116),
	.w6(32'hba39a812),
	.w7(32'hba23d2d7),
	.w8(32'h3a7372cc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b06a7),
	.w1(32'hbaa48c62),
	.w2(32'h3a4cfcde),
	.w3(32'hbb61fe64),
	.w4(32'hb8b00948),
	.w5(32'h3a559321),
	.w6(32'hbac4e5d1),
	.w7(32'hbb1a64c9),
	.w8(32'hbb06ad13),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35c8e),
	.w1(32'h3c2fe07e),
	.w2(32'hbc538eaf),
	.w3(32'hbba73db7),
	.w4(32'h3b44c03a),
	.w5(32'hbc63b86c),
	.w6(32'hbbb4b621),
	.w7(32'h3bbee2d2),
	.w8(32'hbc24eb86),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31d104),
	.w1(32'hbbcdfede),
	.w2(32'hbcc8110d),
	.w3(32'hbb547c73),
	.w4(32'h3b8a3d9d),
	.w5(32'hbc44b070),
	.w6(32'hbb9d9bd3),
	.w7(32'h3a722254),
	.w8(32'hbc8a5855),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc35b9),
	.w1(32'hbb5a2e4c),
	.w2(32'hbbbabb5d),
	.w3(32'hbbb51f5f),
	.w4(32'hbb6bfd75),
	.w5(32'hbbb6d808),
	.w6(32'hbb87d158),
	.w7(32'hbb6c15e2),
	.w8(32'hbc233380),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc560f7f),
	.w1(32'h3bfc99d3),
	.w2(32'h3bcf54bc),
	.w3(32'hbc18a102),
	.w4(32'h3c0fd7d0),
	.w5(32'h3bda8ebb),
	.w6(32'hbc9a2280),
	.w7(32'h3b0ab0cc),
	.w8(32'hba3d43e6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c54bc),
	.w1(32'hba42d702),
	.w2(32'hbc0545f3),
	.w3(32'hbc0f1719),
	.w4(32'h3c28b050),
	.w5(32'h3b6a4a7c),
	.w6(32'hbc802da2),
	.w7(32'h3adb26f9),
	.w8(32'hbba997b5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94c0d1),
	.w1(32'h3a4ec0ed),
	.w2(32'h3ac53462),
	.w3(32'h3a30d4b0),
	.w4(32'hba08cba8),
	.w5(32'h3822f94c),
	.w6(32'h3abedc56),
	.w7(32'hbb652845),
	.w8(32'hb9d4b5b3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad7a25),
	.w1(32'h39eb8610),
	.w2(32'hba9d8574),
	.w3(32'hb9a42366),
	.w4(32'hbacb704c),
	.w5(32'hbb13213f),
	.w6(32'h39e70ae8),
	.w7(32'hb91a9ed5),
	.w8(32'h39ff2d7d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a5810),
	.w1(32'hba07322c),
	.w2(32'hba989337),
	.w3(32'h3ae266ea),
	.w4(32'hbb5d7577),
	.w5(32'hbb9510e2),
	.w6(32'h3b032252),
	.w7(32'hbb2f693b),
	.w8(32'hb9b507a0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0fe2),
	.w1(32'h3a17bb68),
	.w2(32'hb9a31bdd),
	.w3(32'hbb0934c3),
	.w4(32'h3b07d9d6),
	.w5(32'h3a2fc73a),
	.w6(32'h39c6394f),
	.w7(32'h3ac3d1d6),
	.w8(32'h39929e81),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b6aa7),
	.w1(32'hbb6206e2),
	.w2(32'hbba6b05d),
	.w3(32'hb9018dba),
	.w4(32'hbb9be4e3),
	.w5(32'hbb8b0295),
	.w6(32'hbab3b215),
	.w7(32'hbb6a484c),
	.w8(32'hbb7d9730),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62ce06),
	.w1(32'hbb6a6eae),
	.w2(32'hbc86ad81),
	.w3(32'hbad73e3f),
	.w4(32'h3c1023a0),
	.w5(32'hbc30f69f),
	.w6(32'hbc1aebcb),
	.w7(32'hbac294ee),
	.w8(32'hbca3548a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85dd54),
	.w1(32'hbb6746d4),
	.w2(32'hbbd91e9b),
	.w3(32'hbc5c9df5),
	.w4(32'h3a4f267a),
	.w5(32'hbaa4715b),
	.w6(32'hbc83bfd0),
	.w7(32'hbb8c5d24),
	.w8(32'hbbf9bdc6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39335955),
	.w1(32'hb96a9a2d),
	.w2(32'h39b9f8ae),
	.w3(32'h39f6fa5d),
	.w4(32'hbb07c86c),
	.w5(32'h38c79a69),
	.w6(32'h3a93e096),
	.w7(32'hbad046f2),
	.w8(32'hb950bff8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd46f70),
	.w1(32'h3be484dc),
	.w2(32'hbc97f38f),
	.w3(32'hbb211ca6),
	.w4(32'h3b9b2260),
	.w5(32'hbc6f371c),
	.w6(32'h3b43ddce),
	.w7(32'h3c00c0e1),
	.w8(32'hbc542750),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a45d),
	.w1(32'hbaba5206),
	.w2(32'hbc1b0682),
	.w3(32'hb9e50056),
	.w4(32'h3b006c2c),
	.w5(32'hbb5d1253),
	.w6(32'h39593d68),
	.w7(32'h3a9d1436),
	.w8(32'hbb9b0608),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc074e),
	.w1(32'hba88d640),
	.w2(32'hba111a52),
	.w3(32'hba5f606e),
	.w4(32'hbafed108),
	.w5(32'hbb01660f),
	.w6(32'hb953af79),
	.w7(32'hbaa2aa27),
	.w8(32'hbaee3182),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1502),
	.w1(32'h3b3bcd32),
	.w2(32'hbb9fc3e5),
	.w3(32'h39080581),
	.w4(32'h3b54f845),
	.w5(32'hbb86f99b),
	.w6(32'hbab68f5a),
	.w7(32'h3a3c6e8f),
	.w8(32'hbbafcaaf),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ce0a2),
	.w1(32'h3aaefd31),
	.w2(32'h3a829029),
	.w3(32'hb944cebd),
	.w4(32'h3ae00c28),
	.w5(32'h3a4e93dc),
	.w6(32'hb83210f3),
	.w7(32'h3aceb41c),
	.w8(32'h3ac1dbad),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3820e6f7),
	.w1(32'hbac13a0e),
	.w2(32'h3acb5f40),
	.w3(32'h3a31067b),
	.w4(32'hbac2a12c),
	.w5(32'h3a3ebf13),
	.w6(32'hb870d437),
	.w7(32'hba5f05bc),
	.w8(32'hba953dc6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0c0fc),
	.w1(32'hba99fc5a),
	.w2(32'hba5d9f9d),
	.w3(32'h397ccbc4),
	.w4(32'hbab23002),
	.w5(32'h3a87794b),
	.w6(32'hba52d545),
	.w7(32'h3ad7d378),
	.w8(32'h3b08f176),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eabfa),
	.w1(32'hba6467c2),
	.w2(32'hbaac1e65),
	.w3(32'h3aacf15b),
	.w4(32'hbad1ccde),
	.w5(32'h3a2e9962),
	.w6(32'h3a8582a7),
	.w7(32'h3a826138),
	.w8(32'h3a2b9461),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7f13),
	.w1(32'h3ab1619b),
	.w2(32'hbb7436c3),
	.w3(32'hbbb46505),
	.w4(32'hba515fb5),
	.w5(32'h37bd7596),
	.w6(32'hbc15024c),
	.w7(32'hba89933a),
	.w8(32'hbadee227),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b504e),
	.w1(32'hbc0d1e48),
	.w2(32'hbd034f5f),
	.w3(32'hba8ba323),
	.w4(32'hbb3099d9),
	.w5(32'hbcaea9f3),
	.w6(32'hbb50d1c3),
	.w7(32'h38b7e1bc),
	.w8(32'hbc8669ec),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc62fe2),
	.w1(32'hbb887013),
	.w2(32'hbc695065),
	.w3(32'hba7e5793),
	.w4(32'h3b8a0068),
	.w5(32'hbc0996f3),
	.w6(32'hb9e585c4),
	.w7(32'h3b8b9b06),
	.w8(32'hbba306e7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3ee1),
	.w1(32'hbb732159),
	.w2(32'hbc91afda),
	.w3(32'hbaff625a),
	.w4(32'hbac12853),
	.w5(32'hbc82df90),
	.w6(32'hbad73107),
	.w7(32'h396e755b),
	.w8(32'hbc295fa5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca9b18),
	.w1(32'h38de0c90),
	.w2(32'h3abacae4),
	.w3(32'hb8161cb9),
	.w4(32'h3a2e00cd),
	.w5(32'h3b1b5e74),
	.w6(32'h3aaebc37),
	.w7(32'hb9a373da),
	.w8(32'h3a698926),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52e38d),
	.w1(32'hba25b14f),
	.w2(32'h3a1d28e4),
	.w3(32'h3ab8a50c),
	.w4(32'hba858c6a),
	.w5(32'h3ab1becc),
	.w6(32'h3a5c9b75),
	.w7(32'hbaa69ffc),
	.w8(32'h389cf3b4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae513b5),
	.w1(32'hbaa94e50),
	.w2(32'h39753288),
	.w3(32'h3a9d0ff6),
	.w4(32'hba3bd886),
	.w5(32'h3b02d52d),
	.w6(32'h39aded02),
	.w7(32'hba1656a4),
	.w8(32'h3a08972f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8a46e),
	.w1(32'h3a91c661),
	.w2(32'h3a2ee31a),
	.w3(32'h3a79eb68),
	.w4(32'h3ad293b5),
	.w5(32'h3aeec596),
	.w6(32'h39bf0225),
	.w7(32'h3b21a3bc),
	.w8(32'h3b1dcc63),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6985c6),
	.w1(32'hbc149a3c),
	.w2(32'hbc75127a),
	.w3(32'hbb820704),
	.w4(32'h3a2a6564),
	.w5(32'hbb9273c7),
	.w6(32'hbba5593f),
	.w7(32'hbaf38eb0),
	.w8(32'hbc30ed2a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd02d4),
	.w1(32'hba24b330),
	.w2(32'hb838744f),
	.w3(32'hba87c76b),
	.w4(32'hbb17c7a8),
	.w5(32'h3a050aad),
	.w6(32'hb992ee8f),
	.w7(32'hbadcbce7),
	.w8(32'h39fb222a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7f040),
	.w1(32'h3b966c4c),
	.w2(32'h3aa0b1e0),
	.w3(32'hbaa04184),
	.w4(32'h3b0d08cc),
	.w5(32'hb9f7ff53),
	.w6(32'hbbf93f12),
	.w7(32'hbad4a31d),
	.w8(32'hbb897c47),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53c7e9),
	.w1(32'hbab7a156),
	.w2(32'hbb7b2069),
	.w3(32'hbb6f684f),
	.w4(32'hbac7f1c3),
	.w5(32'hbad3430f),
	.w6(32'hbb86086f),
	.w7(32'h38be616c),
	.w8(32'hb9fbd8f7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81cb22),
	.w1(32'hba278249),
	.w2(32'h38eecec7),
	.w3(32'hbab8f3c3),
	.w4(32'hba4c6420),
	.w5(32'hba95c051),
	.w6(32'hbaf1e838),
	.w7(32'hba32dd4e),
	.w8(32'h3896b9eb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19cc9d),
	.w1(32'h3b4620c0),
	.w2(32'hbaa5a992),
	.w3(32'hba11cfe9),
	.w4(32'h3b5c16e5),
	.w5(32'hb9193416),
	.w6(32'hba8b34be),
	.w7(32'h3ab9caa7),
	.w8(32'hbb32869b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c98b7),
	.w1(32'hbac554ea),
	.w2(32'hb95e0b77),
	.w3(32'hba875f8b),
	.w4(32'hbae5d7da),
	.w5(32'h3ac069e7),
	.w6(32'hba8417d9),
	.w7(32'h3afd0eda),
	.w8(32'h3ae53c01),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c9bc),
	.w1(32'hbc354856),
	.w2(32'hbce0ba4a),
	.w3(32'hbbdd69be),
	.w4(32'hbb16945a),
	.w5(32'hbc4cd697),
	.w6(32'hbbb316b4),
	.w7(32'hba1b80a1),
	.w8(32'hbc2eae65),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b93eb),
	.w1(32'h3ab9c916),
	.w2(32'h3ab832e3),
	.w3(32'h379f9d11),
	.w4(32'hb9ff574e),
	.w5(32'hbb191066),
	.w6(32'h3ad208c0),
	.w7(32'hbb1697f4),
	.w8(32'hbbb7ece8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2238d),
	.w1(32'h39b29934),
	.w2(32'hb9b56251),
	.w3(32'hbc54cd2d),
	.w4(32'h3bb3fe20),
	.w5(32'h3b969187),
	.w6(32'hbcdf3341),
	.w7(32'hbbf14ecd),
	.w8(32'hbb93a304),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule