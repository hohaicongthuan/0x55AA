module layer_10_featuremap_462(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9833083),
	.w1(32'hb7a982b9),
	.w2(32'h394a137a),
	.w3(32'h398c2d7c),
	.w4(32'h38df7fd3),
	.w5(32'h3976058b),
	.w6(32'hb890b1e4),
	.w7(32'h393adbf4),
	.w8(32'h38e35a43),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab7169),
	.w1(32'h3a8452c5),
	.w2(32'hba97127d),
	.w3(32'hbadcd700),
	.w4(32'h3b1cc97f),
	.w5(32'h3adc21c6),
	.w6(32'hbb23f936),
	.w7(32'hbac4619b),
	.w8(32'hbbae062f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f425ba),
	.w1(32'h3a279dfd),
	.w2(32'hb7cfa0df),
	.w3(32'h388cf485),
	.w4(32'h3a089b28),
	.w5(32'hb942d670),
	.w6(32'h3927e6de),
	.w7(32'h3a16a1a3),
	.w8(32'hb90a832d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68b243),
	.w1(32'hb90b6783),
	.w2(32'h3b2046d1),
	.w3(32'hbb091934),
	.w4(32'hbb300b0c),
	.w5(32'hbb702f1a),
	.w6(32'hbb1e8da8),
	.w7(32'hbb0c3c34),
	.w8(32'hb9b64131),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8551d52),
	.w1(32'hb832e926),
	.w2(32'hb998a461),
	.w3(32'hb8c97063),
	.w4(32'h3905a171),
	.w5(32'hb8520c42),
	.w6(32'hb972b667),
	.w7(32'hb8a81aaf),
	.w8(32'h391fc3eb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952647a),
	.w1(32'h3943fbe6),
	.w2(32'h36e55080),
	.w3(32'hb954c364),
	.w4(32'h370d3c5a),
	.w5(32'h388f1476),
	.w6(32'hb8b50dbf),
	.w7(32'hb9fa8174),
	.w8(32'hb9992a2a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb797b),
	.w1(32'hbb996ad9),
	.w2(32'h3b96767d),
	.w3(32'hbc111fad),
	.w4(32'hbc295c7d),
	.w5(32'h399c6fb9),
	.w6(32'hbb9979e3),
	.w7(32'hbb74ef11),
	.w8(32'hbb006b15),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd053fbc),
	.w1(32'hbc9653f0),
	.w2(32'hbb76143c),
	.w3(32'hbd179b4c),
	.w4(32'hbcc8db3f),
	.w5(32'hbc20217e),
	.w6(32'hbcdd8bd3),
	.w7(32'hbc491da6),
	.w8(32'h3c229cb8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979885e),
	.w1(32'hb98e2927),
	.w2(32'hba16a95a),
	.w3(32'h39ef42da),
	.w4(32'hb9a79a04),
	.w5(32'hb9e07fa4),
	.w6(32'h39db7de3),
	.w7(32'hb9a88ff9),
	.w8(32'hb959d86a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2e77),
	.w1(32'h3bc87ee2),
	.w2(32'h3c1e57cd),
	.w3(32'hbbfe27b8),
	.w4(32'h3ad9c727),
	.w5(32'h3b66af9a),
	.w6(32'hbc356f01),
	.w7(32'h3ba710f8),
	.w8(32'h3c1beddc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c3f8e),
	.w1(32'hb9e90e2d),
	.w2(32'hba344e17),
	.w3(32'h39b082d9),
	.w4(32'h3823862c),
	.w5(32'hb9b67db0),
	.w6(32'h391fcca8),
	.w7(32'h38d094b8),
	.w8(32'h38b5064e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a51e1),
	.w1(32'hbbbdca48),
	.w2(32'h3be9db22),
	.w3(32'hbc3e25f6),
	.w4(32'hbbd8c7fc),
	.w5(32'h3ac7a12b),
	.w6(32'hbc00ab8d),
	.w7(32'h3a7a4b09),
	.w8(32'h3b5efd8e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a0575),
	.w1(32'hba0bc6a2),
	.w2(32'h3bbbfed5),
	.w3(32'hbc46f9f0),
	.w4(32'hbb7d81fc),
	.w5(32'h3a0d2491),
	.w6(32'hbbf5f9d2),
	.w7(32'h3bac000e),
	.w8(32'h3c02e236),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80a106),
	.w1(32'hb880b7b6),
	.w2(32'hbbc3e218),
	.w3(32'h3ad231ee),
	.w4(32'h3b00116e),
	.w5(32'hbb4e7dd4),
	.w6(32'h3b667571),
	.w7(32'h3a618e23),
	.w8(32'hbad47a79),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1a97),
	.w1(32'h3b164f5a),
	.w2(32'h3aaaa7e0),
	.w3(32'hba26b8c0),
	.w4(32'h3b9f5966),
	.w5(32'h3bb121a9),
	.w6(32'hbaad24a8),
	.w7(32'hbabaeafe),
	.w8(32'hbb890d4e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4596d9),
	.w1(32'hbb2d8ca9),
	.w2(32'h3c646fff),
	.w3(32'hbc362aa5),
	.w4(32'h3b3478ee),
	.w5(32'h3c6144e9),
	.w6(32'hbc374486),
	.w7(32'h3b97c085),
	.w8(32'h3b879277),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c811b6),
	.w1(32'hb819ea8f),
	.w2(32'h391d9de1),
	.w3(32'h3a50f75f),
	.w4(32'hb92eb211),
	.w5(32'hb9fa9cae),
	.w6(32'h3a27e921),
	.w7(32'hb9167203),
	.w8(32'hba2da757),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3a326),
	.w1(32'hbc1a639d),
	.w2(32'h3c57eab0),
	.w3(32'hbcf889d5),
	.w4(32'hbca0ff2b),
	.w5(32'hbc694f18),
	.w6(32'hbc0ad137),
	.w7(32'h3c3dabae),
	.w8(32'h3ca9a750),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc304b16),
	.w1(32'hbab7eb51),
	.w2(32'h3c0fded7),
	.w3(32'hbc434c35),
	.w4(32'hbbe9e9f7),
	.w5(32'hbb058c97),
	.w6(32'hbb918e19),
	.w7(32'h3b9846bd),
	.w8(32'h3c2fd7cc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01d903),
	.w1(32'hb9bc4738),
	.w2(32'hba01c474),
	.w3(32'h3679fe55),
	.w4(32'h399d908d),
	.w5(32'hb8bef014),
	.w6(32'hb9c12279),
	.w7(32'h399e2553),
	.w8(32'hb9b53a81),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883b672),
	.w1(32'hb94cf70c),
	.w2(32'hb9cc39b9),
	.w3(32'h39837bcd),
	.w4(32'hba366fe6),
	.w5(32'hb9a98dc8),
	.w6(32'hb7d0050a),
	.w7(32'hb962806f),
	.w8(32'h394b5199),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c177923),
	.w1(32'h3b3d916e),
	.w2(32'hb959841e),
	.w3(32'h3bb8b1f7),
	.w4(32'h3a1b9b4f),
	.w5(32'hbb2b88ef),
	.w6(32'h3b63402b),
	.w7(32'hba8273e5),
	.w8(32'hbb9ee79d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfbf773),
	.w1(32'hbc8544f6),
	.w2(32'h3c8ca2d2),
	.w3(32'hbca2bede),
	.w4(32'hbc4c9d96),
	.w5(32'h3b305b7c),
	.w6(32'hbcf33eab),
	.w7(32'h3c180d25),
	.w8(32'h3c10b308),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bc319),
	.w1(32'h3bfb80be),
	.w2(32'h3ba0c01d),
	.w3(32'hbb85f7d5),
	.w4(32'h3b32348b),
	.w5(32'h3b4098ed),
	.w6(32'hbb8ddc16),
	.w7(32'h3bf73c7f),
	.w8(32'h3b916124),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca5b08),
	.w1(32'h3c937b88),
	.w2(32'h3c36917c),
	.w3(32'h3b3071c7),
	.w4(32'h3b5a8ca1),
	.w5(32'h3c0a556d),
	.w6(32'h3b83b97b),
	.w7(32'h3bd5b7a2),
	.w8(32'hbaa33184),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89fdf08),
	.w1(32'hb9602274),
	.w2(32'hb98ad0ce),
	.w3(32'hba7e4e8b),
	.w4(32'hba133b92),
	.w5(32'hb9aec023),
	.w6(32'hb9dd1b67),
	.w7(32'hb9b04f1d),
	.w8(32'hba0913a5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3721f8f9),
	.w1(32'hb8e04879),
	.w2(32'hb84d64e9),
	.w3(32'hb8cb50c9),
	.w4(32'hb70f226e),
	.w5(32'h3900b92a),
	.w6(32'hb9251337),
	.w7(32'h3735f68f),
	.w8(32'h39b237bc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf24d5b),
	.w1(32'hbc973d33),
	.w2(32'hbc2fabde),
	.w3(32'h3c1123dd),
	.w4(32'hbd2994be),
	.w5(32'hbc6a4a3b),
	.w6(32'h3cb2fce1),
	.w7(32'hbd009446),
	.w8(32'hbbeea231),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b517c),
	.w1(32'h3a014dc0),
	.w2(32'hba96c45f),
	.w3(32'h39e2511a),
	.w4(32'h3a18db6d),
	.w5(32'hba35f55f),
	.w6(32'hb9130aba),
	.w7(32'hba01c3b8),
	.w8(32'hbabbaae6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3386c7),
	.w1(32'h3c0bb03f),
	.w2(32'h393874ec),
	.w3(32'h3cbba562),
	.w4(32'hbc26877d),
	.w5(32'hbc4dab23),
	.w6(32'h3cbe49aa),
	.w7(32'hbbfd3633),
	.w8(32'hbc92fef1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39483f4c),
	.w1(32'h3a128f11),
	.w2(32'h3a877172),
	.w3(32'h39ec7058),
	.w4(32'h3a0403c9),
	.w5(32'h3a9d9348),
	.w6(32'h39535588),
	.w7(32'h389db18e),
	.w8(32'h38be2c20),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3d3b7),
	.w1(32'h39327b6b),
	.w2(32'h35fd6f19),
	.w3(32'h3a3e792e),
	.w4(32'hb6c5683b),
	.w5(32'hb878e799),
	.w6(32'h39561972),
	.w7(32'h398797e5),
	.w8(32'h389356de),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe32d),
	.w1(32'h3a187628),
	.w2(32'h3b6e2461),
	.w3(32'hbba6798f),
	.w4(32'hbb056ef6),
	.w5(32'hbadddf97),
	.w6(32'hbb23d3c8),
	.w7(32'h3b3524e9),
	.w8(32'h3b91af19),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92efff),
	.w1(32'h3b5e6ba6),
	.w2(32'hba9ee3ba),
	.w3(32'h3ad144b1),
	.w4(32'h3b685088),
	.w5(32'h3a30529a),
	.w6(32'h3b09b344),
	.w7(32'h3b2cd623),
	.w8(32'hbafb6a5a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac1fd1),
	.w1(32'h3a6390f6),
	.w2(32'h3a337fb9),
	.w3(32'h395f8282),
	.w4(32'hb94f1974),
	.w5(32'hb9e60a0b),
	.w6(32'hbac8a132),
	.w7(32'hb8c1f68c),
	.w8(32'h3ace604b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0ef32),
	.w1(32'hbbf037f2),
	.w2(32'h39ec9058),
	.w3(32'hbc175a36),
	.w4(32'hbc7f2c39),
	.w5(32'hbbecd555),
	.w6(32'hbb7515b1),
	.w7(32'h3a26adf4),
	.w8(32'h3bc617d8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd24a814),
	.w1(32'hbc44cdf4),
	.w2(32'hbc8dacaf),
	.w3(32'hbc3ca40c),
	.w4(32'hbc27e694),
	.w5(32'h3c93702e),
	.w6(32'hbc1f287d),
	.w7(32'h3c3e7c4e),
	.w8(32'h3c9042be),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10360c),
	.w1(32'h3c2228d5),
	.w2(32'hbc0f637b),
	.w3(32'h3c7f2764),
	.w4(32'hb962a819),
	.w5(32'hbba0051b),
	.w6(32'h3bfaf641),
	.w7(32'hbcaa9bdd),
	.w8(32'hbd02a0ae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d55434d),
	.w1(32'h3b939f4d),
	.w2(32'hbc1cf9bf),
	.w3(32'h3d12a148),
	.w4(32'hbbd38635),
	.w5(32'hbcbdc24b),
	.w6(32'h3d0b9d35),
	.w7(32'hbc3adc38),
	.w8(32'hbd0535b7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b559270),
	.w1(32'h3ab44180),
	.w2(32'hb9fc96dd),
	.w3(32'hbaa9aa6a),
	.w4(32'hba8f9245),
	.w5(32'hba81b062),
	.w6(32'hbaa8f94b),
	.w7(32'hbb633eb1),
	.w8(32'hbbbac426),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c5c85),
	.w1(32'hb9f75e40),
	.w2(32'hb9c5ab17),
	.w3(32'h36821832),
	.w4(32'hb9dddb55),
	.w5(32'hb9ab9193),
	.w6(32'hb843f0cf),
	.w7(32'hba58651c),
	.w8(32'hba22b277),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09e6d0),
	.w1(32'h3a4037b6),
	.w2(32'h39127f49),
	.w3(32'h3a357950),
	.w4(32'h39e6570e),
	.w5(32'h3996f5da),
	.w6(32'h398c2870),
	.w7(32'h388a3ba7),
	.w8(32'hb6beef8e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba490f07),
	.w1(32'hb99b71e1),
	.w2(32'hbafeeda6),
	.w3(32'hb9c07b63),
	.w4(32'hb90a2223),
	.w5(32'hbad6204e),
	.w6(32'hba5b9ada),
	.w7(32'h385bd805),
	.w8(32'hba9eebc3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77a861),
	.w1(32'hbb4dd86f),
	.w2(32'h3c179419),
	.w3(32'hbcafef3c),
	.w4(32'hbbd40516),
	.w5(32'h3b8c1129),
	.w6(32'hbc83bd15),
	.w7(32'h3bde7015),
	.w8(32'h3c9646f9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f3785),
	.w1(32'h3c40df05),
	.w2(32'h3c0c646b),
	.w3(32'h3aebc43b),
	.w4(32'h3bb220d8),
	.w5(32'h3be4b404),
	.w6(32'h3ba4b088),
	.w7(32'h3bbb3887),
	.w8(32'h3a0bbf96),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57cc9),
	.w1(32'h3c6ba6c1),
	.w2(32'h3c69a8bd),
	.w3(32'hbba578d3),
	.w4(32'h3b1c2c30),
	.w5(32'h3c4aaa3f),
	.w6(32'h3ad0af33),
	.w7(32'h3c88d81d),
	.w8(32'h3c5c2a64),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5aa71),
	.w1(32'h3bf1e837),
	.w2(32'h3c15f07e),
	.w3(32'hbb3e4c40),
	.w4(32'h3abcdd45),
	.w5(32'h3b55eceb),
	.w6(32'hbac63621),
	.w7(32'h3b08341a),
	.w8(32'h3bb2d124),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd22962),
	.w1(32'hbc3a70cc),
	.w2(32'h3be22c67),
	.w3(32'hbce1385d),
	.w4(32'hbcb28adb),
	.w5(32'hbc9c5bb5),
	.w6(32'hbc1bcf46),
	.w7(32'h3b58b436),
	.w8(32'h3c6d49f2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8550a15),
	.w1(32'hb89fee9f),
	.w2(32'h396c1581),
	.w3(32'h3773f856),
	.w4(32'hb8a2bc77),
	.w5(32'h390d6a36),
	.w6(32'h39802575),
	.w7(32'h39c830a0),
	.w8(32'h39c242ba),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070919),
	.w1(32'h3a42e669),
	.w2(32'h3a4a5cd7),
	.w3(32'hb99d142c),
	.w4(32'hb99ac674),
	.w5(32'h3989f2c9),
	.w6(32'h39c26d1e),
	.w7(32'hb8da87a3),
	.w8(32'hb8eee099),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d198ae),
	.w1(32'h3770340b),
	.w2(32'hb9dd9e2d),
	.w3(32'h39ebc9e4),
	.w4(32'hb9dc8f12),
	.w5(32'hb9c094ee),
	.w6(32'h3a734fd5),
	.w7(32'hb9d92eed),
	.w8(32'hb9819b4d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5730f),
	.w1(32'h3aaa2dd4),
	.w2(32'h3b8052bc),
	.w3(32'hbbda95eb),
	.w4(32'hbabdf384),
	.w5(32'h3ac68487),
	.w6(32'hb7dd3a2c),
	.w7(32'h3b992385),
	.w8(32'h3b1f4e97),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83320e),
	.w1(32'hb9a7ea2a),
	.w2(32'h3b32d970),
	.w3(32'hbb1aea70),
	.w4(32'hbb196958),
	.w5(32'hb81cb9a8),
	.w6(32'hbac7c287),
	.w7(32'h3a903d84),
	.w8(32'h3b807291),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc53e66),
	.w1(32'hbbbe7bd6),
	.w2(32'h3c44137d),
	.w3(32'hbcb720ff),
	.w4(32'hbc7c8498),
	.w5(32'hbc011480),
	.w6(32'hbc1612c8),
	.w7(32'h3bb637fb),
	.w8(32'h3c9fb407),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab45071),
	.w1(32'h383eae8b),
	.w2(32'h3ada429f),
	.w3(32'hbbc4a974),
	.w4(32'hbb87a3ab),
	.w5(32'hbb19d330),
	.w6(32'h3b884598),
	.w7(32'h3b81624e),
	.w8(32'h3bc0a3a0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c7915),
	.w1(32'hb71c822a),
	.w2(32'hb9864977),
	.w3(32'h3732f1f8),
	.w4(32'h3971808c),
	.w5(32'h39aa000c),
	.w6(32'hb8d96d75),
	.w7(32'hb8b0d9cc),
	.w8(32'h398ab398),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37401193),
	.w1(32'h39b10e05),
	.w2(32'h398d6c08),
	.w3(32'h396b2bf9),
	.w4(32'h39eac956),
	.w5(32'h3a0919e7),
	.w6(32'h3a426511),
	.w7(32'hb97341e9),
	.w8(32'hb6b8f93a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad0fc),
	.w1(32'h3a940097),
	.w2(32'h3a9e2d43),
	.w3(32'h3a2a7eb8),
	.w4(32'hba6cc6da),
	.w5(32'hba89458b),
	.w6(32'h3a77cf07),
	.w7(32'hb80fd5cf),
	.w8(32'hba0702f1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf70e),
	.w1(32'h38ed6bfa),
	.w2(32'h388237bf),
	.w3(32'h348dcdcc),
	.w4(32'hba3c01bd),
	.w5(32'hba8c8ee2),
	.w6(32'hb9dfae38),
	.w7(32'hbaae1057),
	.w8(32'hbadb5b35),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39661635),
	.w1(32'hb9ca208f),
	.w2(32'h3addea1f),
	.w3(32'h39df712e),
	.w4(32'hbab1cec0),
	.w5(32'hbac3993b),
	.w6(32'h3aa74e27),
	.w7(32'h3ab87c94),
	.w8(32'h3ab78088),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe67846),
	.w1(32'hbb1e693e),
	.w2(32'h3bab085c),
	.w3(32'hbc1a2be8),
	.w4(32'hbbd01284),
	.w5(32'hbb5c3cd3),
	.w6(32'hbb622c81),
	.w7(32'h3bac2ffb),
	.w8(32'h3c109f6d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf045f8),
	.w1(32'hbb86d602),
	.w2(32'h3c65017f),
	.w3(32'hbc1cbe6c),
	.w4(32'hbc522967),
	.w5(32'h3b466899),
	.w6(32'hbad802a7),
	.w7(32'h3b234bff),
	.w8(32'h3c02d2b6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38330049),
	.w1(32'h39acd025),
	.w2(32'hb9a3e260),
	.w3(32'hb6b9c7ce),
	.w4(32'h39aba9ff),
	.w5(32'hb9f69fe7),
	.w6(32'h392f671e),
	.w7(32'h39b1889f),
	.w8(32'hb9804979),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b26729),
	.w1(32'hb9aea92f),
	.w2(32'hb898c372),
	.w3(32'hb89af6bf),
	.w4(32'hb99120cb),
	.w5(32'h39a8dd43),
	.w6(32'h38660cc5),
	.w7(32'hb974a5ad),
	.w8(32'hb98a7a43),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dca26),
	.w1(32'h3a1bd893),
	.w2(32'h39da86bd),
	.w3(32'h39393951),
	.w4(32'h3a40bb47),
	.w5(32'h39e80bbd),
	.w6(32'h3869b7d3),
	.w7(32'h3a70b4c8),
	.w8(32'h3a329227),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c8dae),
	.w1(32'h398f0e34),
	.w2(32'h38d8d35c),
	.w3(32'h3a3dca2e),
	.w4(32'h3a1c5b7d),
	.w5(32'h3a252753),
	.w6(32'h3a83866f),
	.w7(32'h39fe6d8d),
	.w8(32'h39307cd0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc02e48),
	.w1(32'hbb05026c),
	.w2(32'h3c69c54c),
	.w3(32'hbc847291),
	.w4(32'hbc13d6b5),
	.w5(32'h3b12a57f),
	.w6(32'hbcc9f8d9),
	.w7(32'hbc02b9ab),
	.w8(32'h3c490aa2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7d4d),
	.w1(32'h3c594874),
	.w2(32'h3c660dab),
	.w3(32'hbcabd336),
	.w4(32'hbc659309),
	.w5(32'hbbda31f8),
	.w6(32'h3b7109a8),
	.w7(32'h3cdc15ff),
	.w8(32'h3ce1dfa2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0085c7),
	.w1(32'h3b6d984b),
	.w2(32'h3bd34c68),
	.w3(32'hbcaaedc1),
	.w4(32'hbc459674),
	.w5(32'hbbd8147a),
	.w6(32'hbc1457e3),
	.w7(32'h3c9fc0da),
	.w8(32'h3c924061),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c18f0),
	.w1(32'h3cd6d0b4),
	.w2(32'h3b8a04cc),
	.w3(32'h3c04261d),
	.w4(32'h3bfef219),
	.w5(32'h3bc62ea8),
	.w6(32'h3bc658c0),
	.w7(32'hbac86799),
	.w8(32'hbc8507f5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26891),
	.w1(32'h3bcc7773),
	.w2(32'h3c68ffa0),
	.w3(32'h3bbdfc4b),
	.w4(32'h3ba6f125),
	.w5(32'h3aec9fb4),
	.w6(32'hbae80c0c),
	.w7(32'hbbdbc9a0),
	.w8(32'hbc8b9386),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39875f),
	.w1(32'hbaf56a5e),
	.w2(32'hbbc6c0f0),
	.w3(32'hbc39ca55),
	.w4(32'h39bea935),
	.w5(32'hbc1eb9bc),
	.w6(32'hbc92e033),
	.w7(32'h3c205d98),
	.w8(32'h3aba3689),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370981fa),
	.w1(32'h3bb87b22),
	.w2(32'h3b596705),
	.w3(32'hbb9c60b5),
	.w4(32'h3bc33caf),
	.w5(32'h3a96219b),
	.w6(32'h3a37e981),
	.w7(32'h3b52107e),
	.w8(32'h3bc7c4da),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd3441),
	.w1(32'hbb9ef071),
	.w2(32'h3bafeda2),
	.w3(32'h3b9b9a9c),
	.w4(32'h388ac094),
	.w5(32'h3bce4533),
	.w6(32'h3b734627),
	.w7(32'h3b327a14),
	.w8(32'h3b6299c6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d37c),
	.w1(32'h3a83539e),
	.w2(32'h3b75d549),
	.w3(32'hbc00200c),
	.w4(32'h3ae0b898),
	.w5(32'h3bc030c2),
	.w6(32'hbc65731a),
	.w7(32'h39f8a2c1),
	.w8(32'h3ba991a6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6adb9f),
	.w1(32'hbbc525fa),
	.w2(32'h3c8d268f),
	.w3(32'hba1c140f),
	.w4(32'hbb4f2931),
	.w5(32'h3c7d8b06),
	.w6(32'hbc252ee0),
	.w7(32'hbc33438c),
	.w8(32'hbba866d5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda4b0c),
	.w1(32'hbc16c4f2),
	.w2(32'hbb95a081),
	.w3(32'hbb93b4fa),
	.w4(32'hbc93ce32),
	.w5(32'hbca1af88),
	.w6(32'hbbf42e9d),
	.w7(32'hbb2361d2),
	.w8(32'h3b16d30b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4782a4),
	.w1(32'h3c18ef6c),
	.w2(32'hbbf055ec),
	.w3(32'h3be55287),
	.w4(32'h3c8dbe6d),
	.w5(32'hbc08c137),
	.w6(32'h3bec1336),
	.w7(32'h3c20cd4e),
	.w8(32'h3bb0b489),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d97f8),
	.w1(32'h3b98f946),
	.w2(32'h370e2926),
	.w3(32'hbcdfabf3),
	.w4(32'h3bfdc762),
	.w5(32'h3b8e29ef),
	.w6(32'hbc55d252),
	.w7(32'h3be76b63),
	.w8(32'h3b63c95e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc329f9),
	.w1(32'hbbd1a856),
	.w2(32'h3b889576),
	.w3(32'hbcced2ff),
	.w4(32'hbb1f1181),
	.w5(32'hba2a709b),
	.w6(32'hbcf744dc),
	.w7(32'hbb8d8783),
	.w8(32'h3b0b646f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb9515),
	.w1(32'h3bac5165),
	.w2(32'h3b0e3e26),
	.w3(32'h3bb4fa03),
	.w4(32'h3b2ddfe4),
	.w5(32'h3c956ea0),
	.w6(32'h3af2af95),
	.w7(32'hbb27cc87),
	.w8(32'h3baf55ff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b8b3),
	.w1(32'hbb740a46),
	.w2(32'h39ecd141),
	.w3(32'hbb3294eb),
	.w4(32'hbc2d1daf),
	.w5(32'hbc3c1815),
	.w6(32'h3ae16be1),
	.w7(32'hbb736322),
	.w8(32'h3b4dd6f4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe9bc8),
	.w1(32'hbc1e18aa),
	.w2(32'hbbd2e64a),
	.w3(32'h3a8b4078),
	.w4(32'hbbc7dee5),
	.w5(32'h3bea9aac),
	.w6(32'h3bc83d33),
	.w7(32'h3b97ce73),
	.w8(32'h3c490cfc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7639eb),
	.w1(32'h3bbf4413),
	.w2(32'h3b9948aa),
	.w3(32'h3bf9e33c),
	.w4(32'h3c479019),
	.w5(32'h3bdbd6a3),
	.w6(32'h3b9f8a70),
	.w7(32'h3a665370),
	.w8(32'hbb6be413),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e4511),
	.w1(32'hb9fc9361),
	.w2(32'hbb3fa411),
	.w3(32'hbb219ec5),
	.w4(32'hbb4a1064),
	.w5(32'hbc22f9a7),
	.w6(32'h3b8df4b4),
	.w7(32'hbaff41d3),
	.w8(32'h3a86033c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b553190),
	.w1(32'h3c4f470e),
	.w2(32'h3bc61215),
	.w3(32'hbbc8263f),
	.w4(32'h3c004f24),
	.w5(32'hbbbfa60f),
	.w6(32'h3b7abfdc),
	.w7(32'hb9d46cdc),
	.w8(32'hbc214224),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17fd2c),
	.w1(32'h3b992548),
	.w2(32'hbbd09505),
	.w3(32'hbc2b53a0),
	.w4(32'h3bd45877),
	.w5(32'h3c23378e),
	.w6(32'hbbfe09bd),
	.w7(32'hbb455bbe),
	.w8(32'h3c022116),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9dd82),
	.w1(32'h3c8bd7b6),
	.w2(32'h3bd71744),
	.w3(32'hbc19e5c9),
	.w4(32'h3c4598fe),
	.w5(32'h3c1fc624),
	.w6(32'hbaffbeec),
	.w7(32'h3c550f48),
	.w8(32'h3cb6a476),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2055f),
	.w1(32'h3c36d339),
	.w2(32'h3c255f8d),
	.w3(32'h3b7e2f18),
	.w4(32'hbad9bc2a),
	.w5(32'h3bc31065),
	.w6(32'h3c22c13c),
	.w7(32'h3920cdd3),
	.w8(32'hba8cce3f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30f884),
	.w1(32'hb9ca368a),
	.w2(32'h39a91775),
	.w3(32'hbc2d296b),
	.w4(32'hbb0d7150),
	.w5(32'hbccc6538),
	.w6(32'hbc19e391),
	.w7(32'h3c818cd2),
	.w8(32'h3c1f8fcc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dc30a),
	.w1(32'h3b832b5c),
	.w2(32'hbc256868),
	.w3(32'hbb87cb72),
	.w4(32'hba165aaa),
	.w5(32'hbcbb75bf),
	.w6(32'h3a0dfe8e),
	.w7(32'hbc5c24a0),
	.w8(32'hbccc795f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1040c9),
	.w1(32'hbc4272e0),
	.w2(32'h3c89b755),
	.w3(32'hbc388a62),
	.w4(32'hbbd7d8bd),
	.w5(32'h3ca0d01d),
	.w6(32'hbcc9421d),
	.w7(32'hbc3277a8),
	.w8(32'h3c4b77cf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2860ba),
	.w1(32'h3c1a1c13),
	.w2(32'h3c33e8d7),
	.w3(32'h39b7aeb4),
	.w4(32'h3ab77000),
	.w5(32'h3c1d2a58),
	.w6(32'hbc4a3d57),
	.w7(32'hbbf1d438),
	.w8(32'hbc49d85a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca3d4),
	.w1(32'h3c2722d2),
	.w2(32'h3d067874),
	.w3(32'hbc2e6fd3),
	.w4(32'h3a9e8531),
	.w5(32'h3cab3bc6),
	.w6(32'hbc39f135),
	.w7(32'hbbcb5e72),
	.w8(32'hbb3e941d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befd4c8),
	.w1(32'h3bd947bd),
	.w2(32'h3c234c5d),
	.w3(32'h3aa5f0b3),
	.w4(32'h3b3698b9),
	.w5(32'h3bcd6202),
	.w6(32'hbc9b892c),
	.w7(32'hbb49ac87),
	.w8(32'h3b077be2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5514b4),
	.w1(32'h3ba9bfa1),
	.w2(32'hba1b1b12),
	.w3(32'h3a84e956),
	.w4(32'hbaed3b31),
	.w5(32'hbc6f377a),
	.w6(32'h3b3ae959),
	.w7(32'hbca047c5),
	.w8(32'hbca8383f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ea52),
	.w1(32'hbc181b39),
	.w2(32'hbbb57d8f),
	.w3(32'h3c064c14),
	.w4(32'hbc20ebff),
	.w5(32'hbbb78041),
	.w6(32'hbb18d069),
	.w7(32'hb99a3051),
	.w8(32'h3b64d3ba),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73cb1d),
	.w1(32'h3810cce2),
	.w2(32'h3c3e6a24),
	.w3(32'hbc58570c),
	.w4(32'hb9b2a49d),
	.w5(32'hbbd4ca6e),
	.w6(32'hbadd8aca),
	.w7(32'h3c7d5485),
	.w8(32'h3c87f52b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1fd0),
	.w1(32'h3b029749),
	.w2(32'h3c98c262),
	.w3(32'h3b01b979),
	.w4(32'hbb937d13),
	.w5(32'hbc3ca25e),
	.w6(32'hbc191dd9),
	.w7(32'hbbae2ab9),
	.w8(32'h3aa4f812),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68b3a4),
	.w1(32'hbca2f256),
	.w2(32'hbbcb12b3),
	.w3(32'hbcac6eab),
	.w4(32'hbca7363c),
	.w5(32'h3befe898),
	.w6(32'hbc6fc61e),
	.w7(32'h3c89615e),
	.w8(32'h3d237566),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8bb5),
	.w1(32'hbbcf9a7c),
	.w2(32'hbc4ee7b1),
	.w3(32'hbc6e3c6a),
	.w4(32'hbc09d6fc),
	.w5(32'hbcba2250),
	.w6(32'hbc801ae9),
	.w7(32'hbceed406),
	.w8(32'hbd48f8af),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43ec25),
	.w1(32'h3c5f76ad),
	.w2(32'h3c5db7d3),
	.w3(32'hbc0364e8),
	.w4(32'hbae197d9),
	.w5(32'h3c69f1b8),
	.w6(32'hbbb94bfd),
	.w7(32'h3b43a489),
	.w8(32'h3a97b5d4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95076a),
	.w1(32'hbad1c4d3),
	.w2(32'hbbc56bd2),
	.w3(32'h3bc1dee0),
	.w4(32'hbada4a10),
	.w5(32'hbc65096a),
	.w6(32'hbc292acb),
	.w7(32'h39ec91e6),
	.w8(32'h3c9e26de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc738eca),
	.w1(32'h3a070104),
	.w2(32'hbc35de12),
	.w3(32'hbba1a7b9),
	.w4(32'h3c1392ca),
	.w5(32'hbc6e18db),
	.w6(32'hbbd6f3c8),
	.w7(32'hbb6b5bc6),
	.w8(32'hbb4c30e1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5167bc),
	.w1(32'hbc1ba79a),
	.w2(32'hbc89987c),
	.w3(32'hbd6f93ec),
	.w4(32'hbc089338),
	.w5(32'h3bf1296d),
	.w6(32'hbd1c58c1),
	.w7(32'h3ba53354),
	.w8(32'h3c24dcec),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d88dd),
	.w1(32'hbbeb0b27),
	.w2(32'hbbbf4c59),
	.w3(32'hbc0dca79),
	.w4(32'hbbdbf52f),
	.w5(32'hbc047aaa),
	.w6(32'hbbd43a5c),
	.w7(32'h3c343c2a),
	.w8(32'h3c3af651),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51c4c9),
	.w1(32'h3b1b6f9b),
	.w2(32'h3be753a6),
	.w3(32'h3c767a2f),
	.w4(32'h3bd6aec7),
	.w5(32'h3c72af6e),
	.w6(32'h3c9d5380),
	.w7(32'h3bb2afb0),
	.w8(32'h3b6434a9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd5472),
	.w1(32'hbb9707c8),
	.w2(32'hbb6af4a7),
	.w3(32'hbc68f587),
	.w4(32'h3b31c2a8),
	.w5(32'h3c0f83d6),
	.w6(32'hbc82e03e),
	.w7(32'hbbd474c3),
	.w8(32'h3a9ea833),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d73ff),
	.w1(32'hbb518fdc),
	.w2(32'hba5f76f1),
	.w3(32'hbc28cb1a),
	.w4(32'hbbe5c765),
	.w5(32'hbafe72ac),
	.w6(32'hbc7055dc),
	.w7(32'h3c14b90a),
	.w8(32'h3c0db911),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a8c8),
	.w1(32'h3bccff1f),
	.w2(32'h3be4dd07),
	.w3(32'h393299d1),
	.w4(32'h3a0499d0),
	.w5(32'hbbc7b65d),
	.w6(32'h3b9d9e79),
	.w7(32'h3a83f026),
	.w8(32'hbc302afe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021fe1),
	.w1(32'h3c84907a),
	.w2(32'h3c9055ad),
	.w3(32'h3b86514a),
	.w4(32'h3c481b0a),
	.w5(32'hbbfd09e0),
	.w6(32'h3b14bfce),
	.w7(32'hbc027069),
	.w8(32'hbc830a91),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8abf9),
	.w1(32'hb925ab04),
	.w2(32'h3b845621),
	.w3(32'hbb956d08),
	.w4(32'hbb5a3316),
	.w5(32'hbb674066),
	.w6(32'hbc20b677),
	.w7(32'hba7bf663),
	.w8(32'hbab24e18),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbecd5d),
	.w1(32'h3bc3155e),
	.w2(32'h3cc89cb6),
	.w3(32'hbc6020b5),
	.w4(32'hbcb158d2),
	.w5(32'h3b96f99a),
	.w6(32'hbbcbfd2b),
	.w7(32'h3c36dfea),
	.w8(32'h3d4a1e07),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad885b8),
	.w1(32'hbc4c131e),
	.w2(32'h3ca08ddc),
	.w3(32'h3c6f69d5),
	.w4(32'h3bc10c37),
	.w5(32'h3d5a9eda),
	.w6(32'h3c757dfa),
	.w7(32'hbc0302ee),
	.w8(32'h3c1021b3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134e03),
	.w1(32'h3bd6f845),
	.w2(32'h3b10713a),
	.w3(32'hbc49368f),
	.w4(32'h3a572a91),
	.w5(32'hbab496e3),
	.w6(32'hbcaa9a8d),
	.w7(32'h3c1c12ea),
	.w8(32'h3b6e91c3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20ddb7),
	.w1(32'hbb96384a),
	.w2(32'h3b60be40),
	.w3(32'hbc846ae0),
	.w4(32'hbc22f6b5),
	.w5(32'h3bd247cc),
	.w6(32'hbc1d5902),
	.w7(32'h39ec05e3),
	.w8(32'h3c1ca413),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb96d95),
	.w1(32'hbb72e3cc),
	.w2(32'h3bef0206),
	.w3(32'h3c11d4be),
	.w4(32'hbb9ccdeb),
	.w5(32'h3b089e40),
	.w6(32'h3bbdd85d),
	.w7(32'h3b9ce94b),
	.w8(32'h3879eb7d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c321bcb),
	.w1(32'h3c514c42),
	.w2(32'h3ce1a4a3),
	.w3(32'h3cbf9651),
	.w4(32'h3c002973),
	.w5(32'h3bde1760),
	.w6(32'h3c37667b),
	.w7(32'hbc80f166),
	.w8(32'hbd05f173),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befd50b),
	.w1(32'hbc5984d4),
	.w2(32'hbc775deb),
	.w3(32'hbc94d912),
	.w4(32'hbc2927b3),
	.w5(32'hbc5c3be4),
	.w6(32'hbd03501b),
	.w7(32'hbbf8172d),
	.w8(32'h39992a8c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba292),
	.w1(32'hbbc1c69b),
	.w2(32'hbb2d5785),
	.w3(32'hbbeca840),
	.w4(32'hbcb48336),
	.w5(32'hbc45f94b),
	.w6(32'h3b3947ef),
	.w7(32'hbc097584),
	.w8(32'h3b97a507),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3fd14),
	.w1(32'h3b3ce315),
	.w2(32'hba5289a3),
	.w3(32'h3cb79692),
	.w4(32'h3af1070f),
	.w5(32'h3bc1f229),
	.w6(32'h3c70060f),
	.w7(32'hbb375a9b),
	.w8(32'hbb9947c6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3645),
	.w1(32'hbc5988b1),
	.w2(32'h39c4549b),
	.w3(32'hbbd16578),
	.w4(32'hbc727caa),
	.w5(32'h3aa3d8f2),
	.w6(32'hbc2885f6),
	.w7(32'hbb711482),
	.w8(32'h3ba0a30e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd18a),
	.w1(32'h3b77fda7),
	.w2(32'h3abc7c7e),
	.w3(32'h3be3d521),
	.w4(32'hbb888643),
	.w5(32'h3c368941),
	.w6(32'h3c9d7496),
	.w7(32'hbc1184e9),
	.w8(32'h3badaea9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae428),
	.w1(32'hbc102a86),
	.w2(32'hb995a7ce),
	.w3(32'h3c808ab1),
	.w4(32'hbc8a8340),
	.w5(32'h3b82f807),
	.w6(32'h3bb0e953),
	.w7(32'hbc3d1363),
	.w8(32'h3b092184),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa37ab),
	.w1(32'hbbd14359),
	.w2(32'h3c3cc869),
	.w3(32'h3c9fe24f),
	.w4(32'h3bc48208),
	.w5(32'h3c6bfa43),
	.w6(32'h3c3b9966),
	.w7(32'h3a5a1688),
	.w8(32'hbaa3adfc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525dc2),
	.w1(32'hbb8aedf1),
	.w2(32'h3c6741f5),
	.w3(32'h3a528515),
	.w4(32'h3bc210eb),
	.w5(32'h3cb367f5),
	.w6(32'hba224ce3),
	.w7(32'hbbc16331),
	.w8(32'h3b909dc7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf48933),
	.w1(32'hbbcf7d13),
	.w2(32'h3b867a98),
	.w3(32'hba8d162b),
	.w4(32'hbbb39c13),
	.w5(32'hbc14e504),
	.w6(32'hba278dfd),
	.w7(32'hbc0b5506),
	.w8(32'hbc0bd071),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32557a),
	.w1(32'hbbcc0c1c),
	.w2(32'h3cd53634),
	.w3(32'hbcce36c7),
	.w4(32'hbd0073c1),
	.w5(32'hbc9f23e5),
	.w6(32'hbc585ee4),
	.w7(32'h3b00ae39),
	.w8(32'h3c6f69ac),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd19d17),
	.w1(32'hbae21154),
	.w2(32'h3c122665),
	.w3(32'hbc04ccb3),
	.w4(32'hbc0a0310),
	.w5(32'hbbb08823),
	.w6(32'hbc5086d0),
	.w7(32'h3b4226c3),
	.w8(32'h3c835b4b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ee2d5),
	.w1(32'hbbe4c1c0),
	.w2(32'hbb8608af),
	.w3(32'hbc743966),
	.w4(32'hbbe17746),
	.w5(32'hbbb6b80c),
	.w6(32'hbba23c1b),
	.w7(32'hbb5a11c8),
	.w8(32'h3a5af759),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f5586),
	.w1(32'hbb68fd15),
	.w2(32'hbc21ea12),
	.w3(32'hbbeb2450),
	.w4(32'hbb5f8d52),
	.w5(32'hbc413adc),
	.w6(32'hbb1efcc9),
	.w7(32'h3b04bab1),
	.w8(32'hbcb0c48a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01be43),
	.w1(32'hbb735002),
	.w2(32'h3c516aa3),
	.w3(32'hbae714cf),
	.w4(32'h3c162f21),
	.w5(32'h3d13b78f),
	.w6(32'hbbf6299d),
	.w7(32'h3a9a3000),
	.w8(32'h3c496943),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060656),
	.w1(32'hbad379d3),
	.w2(32'h3ba505e3),
	.w3(32'h3b51bc3e),
	.w4(32'h3ae7a378),
	.w5(32'h3c04a6fd),
	.w6(32'h3b8f389d),
	.w7(32'h3c07de66),
	.w8(32'h3c01e337),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68c7ae),
	.w1(32'hba2eb3a5),
	.w2(32'h3a86b922),
	.w3(32'h3b095560),
	.w4(32'hbbb0e412),
	.w5(32'h3b1b4e17),
	.w6(32'hbb22c6a3),
	.w7(32'hbb9b1c6e),
	.w8(32'hbbac2b97),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a2a43),
	.w1(32'hbc3310ac),
	.w2(32'h3bd1bca8),
	.w3(32'hbc6c585f),
	.w4(32'hbc549852),
	.w5(32'hbc5c8226),
	.w6(32'hbc30a53c),
	.w7(32'hbb8c22d6),
	.w8(32'h3c6ca795),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69f558),
	.w1(32'h3b9b5907),
	.w2(32'h3bdb225e),
	.w3(32'h3b78717a),
	.w4(32'h3b8197f6),
	.w5(32'h3be7c3fc),
	.w6(32'h3b93c50b),
	.w7(32'hbc1926c7),
	.w8(32'hbcaa1139),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1661fd),
	.w1(32'hbc048b6b),
	.w2(32'h3c29854e),
	.w3(32'hbc1a8abb),
	.w4(32'h3c3beb91),
	.w5(32'h3cbb845d),
	.w6(32'hbc18270f),
	.w7(32'h3b54e04f),
	.w8(32'h3c97e5f2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5fe28),
	.w1(32'hbba20077),
	.w2(32'h3c893f6c),
	.w3(32'hbd0b4c60),
	.w4(32'hbca5b228),
	.w5(32'hbc4f25cb),
	.w6(32'hbc899403),
	.w7(32'hbc3243c9),
	.w8(32'hbaf2c0a6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67a16e),
	.w1(32'h3b58e4d5),
	.w2(32'hbb7b712f),
	.w3(32'hbca57d38),
	.w4(32'hbb3ac222),
	.w5(32'hbad8dca3),
	.w6(32'hbbba2786),
	.w7(32'h3c1f0919),
	.w8(32'h3c7dde79),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e56ff),
	.w1(32'hbba6628d),
	.w2(32'h3b618d4d),
	.w3(32'hbb92b9e1),
	.w4(32'hbc9464ce),
	.w5(32'hbc172527),
	.w6(32'hbb7da6dc),
	.w7(32'hbc11be06),
	.w8(32'hba0577d6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054a3f),
	.w1(32'h3c3abc8a),
	.w2(32'h3b6d3620),
	.w3(32'h3c43ff3a),
	.w4(32'h3c29c9f9),
	.w5(32'hbb4b9ba1),
	.w6(32'h3c19aa13),
	.w7(32'h3b79aae0),
	.w8(32'hbc0e3019),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5625a5),
	.w1(32'h3b97eba9),
	.w2(32'h3c275788),
	.w3(32'h3c6f71a6),
	.w4(32'hbc9a3c3f),
	.w5(32'hbca686fc),
	.w6(32'h3c9da39d),
	.w7(32'hbc93fa7e),
	.w8(32'hbc841931),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d11d),
	.w1(32'hbc2a9d0b),
	.w2(32'h3a8b8c87),
	.w3(32'hbbaa9daf),
	.w4(32'hbc4fe547),
	.w5(32'h3b37f8d1),
	.w6(32'h3a90f486),
	.w7(32'hbbf2d0e6),
	.w8(32'h3bbdd336),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ce60),
	.w1(32'h3c2ca91c),
	.w2(32'h3b674f1a),
	.w3(32'h3bb6c218),
	.w4(32'h3c15d516),
	.w5(32'h3b562c02),
	.w6(32'h3bf482c5),
	.w7(32'h3b44bc84),
	.w8(32'h3aff3154),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947350),
	.w1(32'h3bd95230),
	.w2(32'h3c313679),
	.w3(32'hbbb2f76c),
	.w4(32'h3c169b10),
	.w5(32'h3c67d90d),
	.w6(32'hbb02ede0),
	.w7(32'h3aaea311),
	.w8(32'h3bc00e95),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874503),
	.w1(32'h3bf37aba),
	.w2(32'h3babfab6),
	.w3(32'h3c021d8f),
	.w4(32'h3c58b9ff),
	.w5(32'hbb9aba4f),
	.w6(32'h3c1dc20a),
	.w7(32'h3c6eb9f3),
	.w8(32'hbb92250d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc8e52),
	.w1(32'hbbfb69c4),
	.w2(32'hba9b3316),
	.w3(32'hbd0385a2),
	.w4(32'hbc5bef28),
	.w5(32'h3a938c80),
	.w6(32'hbcbd8b4a),
	.w7(32'hbc946b4a),
	.w8(32'hbc02817a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9aa37),
	.w1(32'hb70a1a04),
	.w2(32'h37168e7e),
	.w3(32'hbc5869c7),
	.w4(32'h3c3ec3e3),
	.w5(32'hbb365682),
	.w6(32'hbb74a399),
	.w7(32'h3ca507c5),
	.w8(32'h3cb5f080),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b5c62),
	.w1(32'hbb2b875e),
	.w2(32'hbaa23bbd),
	.w3(32'hba5e6eef),
	.w4(32'h3ac50bb7),
	.w5(32'hbb83b2bb),
	.w6(32'hbb586b8e),
	.w7(32'h3a74c3af),
	.w8(32'hbc15d199),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e97b),
	.w1(32'h3aec4bf5),
	.w2(32'hbb6fdbb1),
	.w3(32'hbc6d59b5),
	.w4(32'h3c645e81),
	.w5(32'hb9251dbd),
	.w6(32'hbc8ecb7d),
	.w7(32'h3b60a567),
	.w8(32'hbb01970e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3575fd),
	.w1(32'h3b8f30a0),
	.w2(32'h3c16b4c7),
	.w3(32'h3a502d3a),
	.w4(32'h3b6482d6),
	.w5(32'h3c0d51ab),
	.w6(32'hbbde6c3e),
	.w7(32'h3b10f36f),
	.w8(32'h3bfd3236),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccac941),
	.w1(32'hbc5a1a53),
	.w2(32'h3c9d725c),
	.w3(32'hbbc0e893),
	.w4(32'hbb923f72),
	.w5(32'h3cdcd784),
	.w6(32'hbc542a57),
	.w7(32'hbc1d86c5),
	.w8(32'h3c899942),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0d73a),
	.w1(32'hbc2962cc),
	.w2(32'hbc64afa2),
	.w3(32'h3ca2571a),
	.w4(32'hbc2f058b),
	.w5(32'hbc635ada),
	.w6(32'h3cc37373),
	.w7(32'hbc24360c),
	.w8(32'hbb7a0f59),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a6149),
	.w1(32'h36df3b88),
	.w2(32'h3a848d33),
	.w3(32'h3b9d3089),
	.w4(32'hba53dacf),
	.w5(32'h3c043942),
	.w6(32'h3b209b71),
	.w7(32'hbaf53d06),
	.w8(32'hbbde430e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae62e90),
	.w1(32'h399f1108),
	.w2(32'hbb5e1ee2),
	.w3(32'h3b856b12),
	.w4(32'hbb9e03e8),
	.w5(32'hbc7fa025),
	.w6(32'hbb677c54),
	.w7(32'hbab6d5d7),
	.w8(32'hbb43ace3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03f14),
	.w1(32'hbb0b695e),
	.w2(32'hbb819447),
	.w3(32'h3b2fb112),
	.w4(32'hbc0aa22d),
	.w5(32'hbc0b400f),
	.w6(32'h3c1186df),
	.w7(32'hbc0a39b5),
	.w8(32'hbba5a76c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556b38),
	.w1(32'h3bcbdd41),
	.w2(32'h3c39968f),
	.w3(32'h3b56b257),
	.w4(32'h3bbb1318),
	.w5(32'h3af16555),
	.w6(32'h3c1ca7d8),
	.w7(32'h3b82f649),
	.w8(32'h3b0f5b33),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82686d),
	.w1(32'h3c059bc7),
	.w2(32'hbbaa0497),
	.w3(32'h3c0c9621),
	.w4(32'h3bc34197),
	.w5(32'hbc672cb8),
	.w6(32'h3c0acf01),
	.w7(32'hba375e68),
	.w8(32'hbc467ea9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc728c07),
	.w1(32'hbc760321),
	.w2(32'hbbc7d10e),
	.w3(32'hbc93f0e5),
	.w4(32'hbc54efaa),
	.w5(32'hbbc29af8),
	.w6(32'hbc1a7304),
	.w7(32'h3ab273bb),
	.w8(32'h3bb2b95d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcdbd7),
	.w1(32'h3a9d3b87),
	.w2(32'h3c0a38a1),
	.w3(32'hbb9f5174),
	.w4(32'hbbf5c440),
	.w5(32'h3b4cfe0a),
	.w6(32'hbbd5e529),
	.w7(32'hba840ef8),
	.w8(32'h3be4ed42),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c28b),
	.w1(32'h3b58f77a),
	.w2(32'h3b83c7d7),
	.w3(32'hb7e6c86a),
	.w4(32'hbb1ff739),
	.w5(32'hbc0cb838),
	.w6(32'h3b2b81aa),
	.w7(32'h3ba1f70a),
	.w8(32'h3c44d681),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a6caa),
	.w1(32'hb97a100d),
	.w2(32'hbb827456),
	.w3(32'hb9e79abb),
	.w4(32'hbbeb906a),
	.w5(32'hbc3efd1f),
	.w6(32'h3b5d259c),
	.w7(32'hbb02317c),
	.w8(32'h3bf0318d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fd6fe),
	.w1(32'hbb3aef03),
	.w2(32'hbca9199a),
	.w3(32'hba5a8edf),
	.w4(32'hbc091ba5),
	.w5(32'hbc32bc14),
	.w6(32'h3c7cdbeb),
	.w7(32'h3c8bc33e),
	.w8(32'h3cbaaf15),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d2911),
	.w1(32'h3b7e83f9),
	.w2(32'h3a0c74d4),
	.w3(32'hbc12865b),
	.w4(32'h3c0a99b6),
	.w5(32'h3b62bb28),
	.w6(32'h3be04d50),
	.w7(32'h3ae558d0),
	.w8(32'hbbd9e779),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f0ab),
	.w1(32'h3c87c34d),
	.w2(32'h3c92c4b2),
	.w3(32'hbcdec3f1),
	.w4(32'h3c39f07e),
	.w5(32'h3b98e4ce),
	.w6(32'hbca4dfe2),
	.w7(32'h3b8541de),
	.w8(32'h3c1f612c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04672e),
	.w1(32'h3b157bdc),
	.w2(32'h3aa74b2a),
	.w3(32'hbbb2b3fa),
	.w4(32'hbbb74346),
	.w5(32'hbb4a0a51),
	.w6(32'hbbad74b7),
	.w7(32'hbbbbfb99),
	.w8(32'hbb8ead06),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3816),
	.w1(32'hbc334883),
	.w2(32'hbb9ddeca),
	.w3(32'h3c0f78af),
	.w4(32'hbcb79c55),
	.w5(32'hbc9d27b1),
	.w6(32'h3c14ab99),
	.w7(32'hbca2be96),
	.w8(32'hbc723d54),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f4aa5),
	.w1(32'h3b7240d3),
	.w2(32'h39ecb304),
	.w3(32'h3ca6f171),
	.w4(32'h3b5eab44),
	.w5(32'h3c086f05),
	.w6(32'h3c517848),
	.w7(32'hbb5344d7),
	.w8(32'hb9ce3a6c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b150a49),
	.w1(32'hba88b3cb),
	.w2(32'hba3e1c04),
	.w3(32'hbcb02957),
	.w4(32'hbce7e146),
	.w5(32'hbcd3245c),
	.w6(32'hbc5eaf58),
	.w7(32'hbc12e93b),
	.w8(32'hbb8e90c7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d6b88),
	.w1(32'hbb000c46),
	.w2(32'hba826847),
	.w3(32'hbc426437),
	.w4(32'hbba7678b),
	.w5(32'hba8213c2),
	.w6(32'hbcb8427c),
	.w7(32'hbbe51334),
	.w8(32'hbb8b52e1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8217cd),
	.w1(32'h3bb84718),
	.w2(32'h3bb626f4),
	.w3(32'h3cad7c57),
	.w4(32'h3ace9165),
	.w5(32'h3b6dc26b),
	.w6(32'h3c469058),
	.w7(32'h3a88dfc0),
	.w8(32'hbb420516),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d5f4),
	.w1(32'hbbc4e398),
	.w2(32'hbb8bd868),
	.w3(32'hbbfa629f),
	.w4(32'hbb84e329),
	.w5(32'hbaea4dab),
	.w6(32'hbb4e16eb),
	.w7(32'hbb7eaf00),
	.w8(32'h3aeb7604),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f085f),
	.w1(32'h3be66f53),
	.w2(32'h3c8bce02),
	.w3(32'hbcbb2195),
	.w4(32'h3c15c692),
	.w5(32'h3bb1288a),
	.w6(32'hbc53c8de),
	.w7(32'h3c1aa259),
	.w8(32'h3c04f604),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5eca6),
	.w1(32'h3c650e4c),
	.w2(32'h3bff0ac9),
	.w3(32'hbc67b7a3),
	.w4(32'h3bed9229),
	.w5(32'hbbc30364),
	.w6(32'hbc6f916c),
	.w7(32'h3b4b74db),
	.w8(32'hb894bd48),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa641),
	.w1(32'hbb59910e),
	.w2(32'h3c0f6482),
	.w3(32'hbcaa2399),
	.w4(32'hbc6ea652),
	.w5(32'hbc6cf99c),
	.w6(32'hbc38d018),
	.w7(32'h3975199e),
	.w8(32'hb961e93e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ce4c),
	.w1(32'hbb949b95),
	.w2(32'hbb885c6f),
	.w3(32'hbc3b0a0f),
	.w4(32'hbc71c5f9),
	.w5(32'hbc918648),
	.w6(32'hbc330eb3),
	.w7(32'hbb2b8b9a),
	.w8(32'h3b93ae58),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78672a),
	.w1(32'h3c52bcea),
	.w2(32'h3c1c01ed),
	.w3(32'h3cbf9028),
	.w4(32'h3c8b0e0f),
	.w5(32'h3bc3890a),
	.w6(32'h3cb4e6ed),
	.w7(32'h3b9ab8c7),
	.w8(32'hba2b49ad),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7256d7),
	.w1(32'hbc14f0c2),
	.w2(32'h3b9325b8),
	.w3(32'hbcb94219),
	.w4(32'hbcf46e61),
	.w5(32'hbbbe5980),
	.w6(32'hbca64d1d),
	.w7(32'hbc7324b3),
	.w8(32'hb8d32976),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3302a5),
	.w1(32'hbc1c266c),
	.w2(32'hbbb14015),
	.w3(32'h3cba55db),
	.w4(32'hbc1e4f75),
	.w5(32'hbbb3c23a),
	.w6(32'h3c683abf),
	.w7(32'hbbe3c05f),
	.w8(32'hbb273b95),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcfb73),
	.w1(32'h38063b41),
	.w2(32'h3be8849c),
	.w3(32'h3bfb2b91),
	.w4(32'h3b501986),
	.w5(32'h3b9c55c4),
	.w6(32'h3b9f96e5),
	.w7(32'hbb9a3bbc),
	.w8(32'h3a0ef65f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea37a),
	.w1(32'hba026ee3),
	.w2(32'hb9025b19),
	.w3(32'hbb69e3ba),
	.w4(32'hbb7c0457),
	.w5(32'hbb0faca4),
	.w6(32'hbc0225a4),
	.w7(32'h3bc03cf7),
	.w8(32'h3cb29d49),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88db69),
	.w1(32'hba2ee06e),
	.w2(32'hbbcbb764),
	.w3(32'h3b9c2b6a),
	.w4(32'h3c0719e0),
	.w5(32'h3c39ec94),
	.w6(32'h3c82e85d),
	.w7(32'h3c8e86fe),
	.w8(32'h3cee0529),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30aec2),
	.w1(32'hbbb9ba62),
	.w2(32'hbc37ab3f),
	.w3(32'hbc50dafa),
	.w4(32'hbb8eef2b),
	.w5(32'hbc56bc12),
	.w6(32'h3a74a00e),
	.w7(32'hbbbfc378),
	.w8(32'hbb6c5014),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e1277),
	.w1(32'h3c351ca2),
	.w2(32'h3c160ff4),
	.w3(32'hbc2981f9),
	.w4(32'h3bf6fb30),
	.w5(32'h3cc69992),
	.w6(32'h3b23a300),
	.w7(32'h3ae08ec9),
	.w8(32'h3ca02c45),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7813),
	.w1(32'hba809830),
	.w2(32'hbb7a1c94),
	.w3(32'hbc2cba4c),
	.w4(32'hbb3e36c7),
	.w5(32'hbc4baf96),
	.w6(32'hbca65ddd),
	.w7(32'h3bec05e9),
	.w8(32'h3c06208b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca27e4b),
	.w1(32'hbc65383d),
	.w2(32'hbc43e975),
	.w3(32'hbca1b795),
	.w4(32'hbb42b74c),
	.w5(32'h3ae3f646),
	.w6(32'hbca1527b),
	.w7(32'h3b1c73bf),
	.w8(32'hbbeecfc7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2bd5),
	.w1(32'hbc5b82fd),
	.w2(32'hbb4f3d4c),
	.w3(32'hbbd6e615),
	.w4(32'hbc85f0b2),
	.w5(32'h3b97cd7a),
	.w6(32'hbc47ceb8),
	.w7(32'hbc96dc0d),
	.w8(32'hba72b9d0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7ffe1),
	.w1(32'hbbe0114d),
	.w2(32'h3c5d7a4d),
	.w3(32'hbd153e85),
	.w4(32'hbc8149a8),
	.w5(32'hbc4eb6cd),
	.w6(32'hbcd75dae),
	.w7(32'h3c3f1ba5),
	.w8(32'h3cd8479c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c696c47),
	.w1(32'hbbbe212f),
	.w2(32'h3c04e781),
	.w3(32'h3ba94d40),
	.w4(32'hbb92513a),
	.w5(32'h3be1fecb),
	.w6(32'hbbb26bf8),
	.w7(32'hbcd9ea6c),
	.w8(32'hbbef4793),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67e368),
	.w1(32'hbbeaa815),
	.w2(32'hbbac8e82),
	.w3(32'hbc168164),
	.w4(32'hbb024c22),
	.w5(32'hba0f6754),
	.w6(32'hbc5a32e6),
	.w7(32'hbb09f3df),
	.w8(32'hbaa37110),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd5ea),
	.w1(32'h3c1ed693),
	.w2(32'h3c0a6e9d),
	.w3(32'h3bb0f0f5),
	.w4(32'h3cabe59c),
	.w5(32'h3c869034),
	.w6(32'h3ad6fefd),
	.w7(32'h3c29df39),
	.w8(32'h3a75beee),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b935),
	.w1(32'hbb895733),
	.w2(32'h3b1a831c),
	.w3(32'hbcf6dded),
	.w4(32'hbc27d920),
	.w5(32'h3aff564b),
	.w6(32'hbccc66d0),
	.w7(32'h3a042104),
	.w8(32'h3bdff4c4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8d4d),
	.w1(32'h3b389eb4),
	.w2(32'h3c08e5d7),
	.w3(32'h3c1b5757),
	.w4(32'h3bc6bd08),
	.w5(32'h3c8ae46b),
	.w6(32'h3b1e8548),
	.w7(32'hbada4de4),
	.w8(32'h38cb251c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87fdce),
	.w1(32'hbc272e50),
	.w2(32'h393cc0e0),
	.w3(32'hbc60caa8),
	.w4(32'hbca0284b),
	.w5(32'hbba2de36),
	.w6(32'hbc54d7c7),
	.w7(32'hbc2c2c2c),
	.w8(32'hb8ee0fec),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5efe5),
	.w1(32'hbc658b61),
	.w2(32'hbcdebd1f),
	.w3(32'h3c89856e),
	.w4(32'hbc926df1),
	.w5(32'hbd3478e8),
	.w6(32'h3c51902d),
	.w7(32'h3bfb1b09),
	.w8(32'hbb81b789),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb1f80),
	.w1(32'h3c3ebaa8),
	.w2(32'hba0d1068),
	.w3(32'hbc7ab503),
	.w4(32'h3caa7bca),
	.w5(32'hbca5b3c8),
	.w6(32'h3bf8b382),
	.w7(32'h3c4ad132),
	.w8(32'hbc5c0958),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392c40),
	.w1(32'hbb7e5b27),
	.w2(32'hba3f33f9),
	.w3(32'hbca30f4c),
	.w4(32'hbb633a0b),
	.w5(32'hbc326c02),
	.w6(32'hbb4adfe0),
	.w7(32'hbbc4f67b),
	.w8(32'hbbbf3526),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a433e),
	.w1(32'h3a082646),
	.w2(32'h3c0bd272),
	.w3(32'hbc5a5e65),
	.w4(32'hbb6ff24a),
	.w5(32'h3a4b1597),
	.w6(32'hbc75e511),
	.w7(32'h3be45748),
	.w8(32'h3c0caba7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f61f1),
	.w1(32'hb8dd5b5a),
	.w2(32'hbb1a6f54),
	.w3(32'hb9d11ab8),
	.w4(32'h3a586092),
	.w5(32'hbada212a),
	.w6(32'h39645ce7),
	.w7(32'h3ba94dd2),
	.w8(32'h3b2bb220),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384246d7),
	.w1(32'hb8040ca8),
	.w2(32'h37a7575a),
	.w3(32'h389e3818),
	.w4(32'h37ac7959),
	.w5(32'h38514860),
	.w6(32'h388e7988),
	.w7(32'h3699a36d),
	.w8(32'h38107b08),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59bbf5),
	.w1(32'hbaf8783d),
	.w2(32'hbbd7cc99),
	.w3(32'hbb7759dc),
	.w4(32'h3b1cbbf2),
	.w5(32'h38bdea78),
	.w6(32'h39e1a073),
	.w7(32'h3be1a5be),
	.w8(32'h3b811069),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918c165),
	.w1(32'hb88a7d8f),
	.w2(32'hb74c06c6),
	.w3(32'h398116fd),
	.w4(32'h38801f57),
	.w5(32'h38e7a017),
	.w6(32'h398a9183),
	.w7(32'h385d3932),
	.w8(32'h377bf681),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7243b),
	.w1(32'h3b1a8018),
	.w2(32'h3b8d9950),
	.w3(32'hbb90430e),
	.w4(32'hbaa838c6),
	.w5(32'hbaf934d9),
	.w6(32'hba8504b7),
	.w7(32'h3b7f3787),
	.w8(32'h3b987a09),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95281),
	.w1(32'h3ba2ea9b),
	.w2(32'h39f8b800),
	.w3(32'h39905f36),
	.w4(32'h3bcaca7c),
	.w5(32'h3bb9f4b1),
	.w6(32'h3a77884d),
	.w7(32'h39b84794),
	.w8(32'hbada6214),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9694d3),
	.w1(32'h3bce4839),
	.w2(32'h3ba8b27b),
	.w3(32'h3a2e5fed),
	.w4(32'h3b5a774a),
	.w5(32'h3b63a5af),
	.w6(32'h3aadbb6b),
	.w7(32'h3b7eed46),
	.w8(32'h3a9da37e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813abdd),
	.w1(32'h38e30662),
	.w2(32'hba3213bd),
	.w3(32'h38914103),
	.w4(32'h370d663b),
	.w5(32'hba293988),
	.w6(32'hb9ccd364),
	.w7(32'hb9fec299),
	.w8(32'hba5c94ac),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155ef1),
	.w1(32'h3bbf3834),
	.w2(32'h3b557f93),
	.w3(32'h3b1e22ed),
	.w4(32'h3b91de0e),
	.w5(32'h3b408f09),
	.w6(32'h3c0ac4ee),
	.w7(32'h3abe4732),
	.w8(32'hbb2b87f4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd8de),
	.w1(32'hba1cb3b1),
	.w2(32'h3b66e587),
	.w3(32'hbbc25237),
	.w4(32'hbb046062),
	.w5(32'h3a65b989),
	.w6(32'hbb8bd9a8),
	.w7(32'h3a57a7f5),
	.w8(32'h3c130958),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ac1f),
	.w1(32'h3bdcba4d),
	.w2(32'h3c173319),
	.w3(32'hbbc0365c),
	.w4(32'h3b5535a3),
	.w5(32'h3b89bb0c),
	.w6(32'hbb07e9aa),
	.w7(32'h3be206a9),
	.w8(32'h3bcd5a0b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389cf915),
	.w1(32'h387a9e56),
	.w2(32'h3997dc60),
	.w3(32'h38c9114e),
	.w4(32'h37237385),
	.w5(32'h3978136e),
	.w6(32'h37f6ee51),
	.w7(32'hb8819df5),
	.w8(32'hb626c292),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d05d9),
	.w1(32'h39a93592),
	.w2(32'h39b555e1),
	.w3(32'h3a28db03),
	.w4(32'hba15507f),
	.w5(32'hbaa93bdf),
	.w6(32'h3a9caefd),
	.w7(32'h39551d03),
	.w8(32'hb9908a87),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ab16b),
	.w1(32'h3ab8bd32),
	.w2(32'h3baa24d3),
	.w3(32'hbc24a15e),
	.w4(32'hbc09bbb0),
	.w5(32'h3bb02aad),
	.w6(32'h3a77c584),
	.w7(32'h3c8282c5),
	.w8(32'h3c81fd01),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2076c9),
	.w1(32'h3b96a251),
	.w2(32'h3c022494),
	.w3(32'hbc212eec),
	.w4(32'hbc369d22),
	.w5(32'hbbd56899),
	.w6(32'hbb70b1a4),
	.w7(32'h3c8150a0),
	.w8(32'h3c6d482e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c1f1),
	.w1(32'h3c1ec6ac),
	.w2(32'h3beae66f),
	.w3(32'hbb434abc),
	.w4(32'h3b5bdd0b),
	.w5(32'h3c037119),
	.w6(32'h3ad9b640),
	.w7(32'h3c428c4f),
	.w8(32'h3c2acfa7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fec9a),
	.w1(32'hbbc8bb9d),
	.w2(32'h3c388538),
	.w3(32'hbbb21e53),
	.w4(32'hbc0d5e55),
	.w5(32'h3b15fc14),
	.w6(32'hbc19665a),
	.w7(32'hbbf2c7f7),
	.w8(32'h3bf38753),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00db7d),
	.w1(32'hbabe5bec),
	.w2(32'hbaa9e503),
	.w3(32'hbb4cd180),
	.w4(32'hba8a6993),
	.w5(32'hbb0ba78f),
	.w6(32'hbabc2f66),
	.w7(32'hba5d93d7),
	.w8(32'hbaa84037),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901adf8),
	.w1(32'h3aa2dc28),
	.w2(32'h3a96b04a),
	.w3(32'h3a00270d),
	.w4(32'hb9db2ac5),
	.w5(32'hba8de158),
	.w6(32'h3b691ff1),
	.w7(32'h3b6f4259),
	.w8(32'h3b81695d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc116732),
	.w1(32'hbc867ebf),
	.w2(32'h3b434719),
	.w3(32'hbcc08e2a),
	.w4(32'hbcb5bb9b),
	.w5(32'hbc1628d2),
	.w6(32'hbc64a078),
	.w7(32'hbb2dc8f8),
	.w8(32'h3abffa4e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc848020),
	.w1(32'hbc04b658),
	.w2(32'h3c13ac2b),
	.w3(32'hbcab3f0f),
	.w4(32'hbc86cdb4),
	.w5(32'hbc11e923),
	.w6(32'hbc0757fb),
	.w7(32'h3c14689e),
	.w8(32'h3c8f5754),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3f462),
	.w1(32'hbc4b69bb),
	.w2(32'hbb1b63dd),
	.w3(32'hbc5c1146),
	.w4(32'hbc16e2e2),
	.w5(32'hbb87bb42),
	.w6(32'hbc4af102),
	.w7(32'h3aabae73),
	.w8(32'h3c02c519),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca59f8a),
	.w1(32'h3c153506),
	.w2(32'h3b4fa339),
	.w3(32'h3bec5751),
	.w4(32'hbac827d4),
	.w5(32'hbb24c649),
	.w6(32'h3bed9a0c),
	.w7(32'hbb5e39de),
	.w8(32'hbc1b5c92),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c639568),
	.w1(32'h3bac26cf),
	.w2(32'h3a4e87bb),
	.w3(32'h3bab3ce5),
	.w4(32'h3baf74ca),
	.w5(32'h3b0c2b46),
	.w6(32'h3bd03caf),
	.w7(32'hbb693877),
	.w8(32'hbc155163),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c5b61),
	.w1(32'h37e3cbd3),
	.w2(32'h37fb876d),
	.w3(32'h384cf421),
	.w4(32'h37d4bbc4),
	.w5(32'h382384b0),
	.w6(32'h385df8ad),
	.w7(32'h37c83759),
	.w8(32'h378178ae),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38503e3e),
	.w1(32'hb73f679b),
	.w2(32'hb5d0c20b),
	.w3(32'h389c837d),
	.w4(32'h36902033),
	.w5(32'h37004118),
	.w6(32'h38837b91),
	.w7(32'hb6168b58),
	.w8(32'hb6a6e9c2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3e571),
	.w1(32'h3b747d76),
	.w2(32'h3c05d651),
	.w3(32'hbaf60bff),
	.w4(32'hbb4e2a1a),
	.w5(32'hb9449ca6),
	.w6(32'h39ed1e25),
	.w7(32'h3b13d6d0),
	.w8(32'h3bbc9362),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38011bca),
	.w1(32'hb805357b),
	.w2(32'hb7ace91c),
	.w3(32'h388162e8),
	.w4(32'hb76a492d),
	.w5(32'h360659b0),
	.w6(32'h384bb5e1),
	.w7(32'hb50ab5c9),
	.w8(32'h378ca0b0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0a5a7),
	.w1(32'hbabbab60),
	.w2(32'hbb1458b4),
	.w3(32'hbb1e412e),
	.w4(32'hbb270e85),
	.w5(32'hbb9f64a5),
	.w6(32'hbae3759d),
	.w7(32'hb84bf566),
	.w8(32'hbb18eeda),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89471c),
	.w1(32'h3a0a998e),
	.w2(32'h3bcc965a),
	.w3(32'hbbb787ea),
	.w4(32'hbba7c51e),
	.w5(32'hbab57c2b),
	.w6(32'hbb029237),
	.w7(32'h3c411973),
	.w8(32'h3c5f9154),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6898d1),
	.w1(32'h3b996fc3),
	.w2(32'h3b9ea292),
	.w3(32'hbb89e6e1),
	.w4(32'h39f9ab01),
	.w5(32'h3b170956),
	.w6(32'hbaa34e78),
	.w7(32'h3b8ba563),
	.w8(32'h3b9cc32b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385251bf),
	.w1(32'hb6c7c888),
	.w2(32'hb793c240),
	.w3(32'h38350a96),
	.w4(32'h381dee2f),
	.w5(32'h3899a1c8),
	.w6(32'h3856f42c),
	.w7(32'hb820b727),
	.w8(32'hb7436f7c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee94de),
	.w1(32'hbc26f8e5),
	.w2(32'hbbcd1818),
	.w3(32'hbcaf7713),
	.w4(32'hbc55538b),
	.w5(32'hbc2262b4),
	.w6(32'hbc66a946),
	.w7(32'h3c052cf8),
	.w8(32'h3cfea518),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5cbae),
	.w1(32'hba84a046),
	.w2(32'h3b9ed5eb),
	.w3(32'hbbdc7f5b),
	.w4(32'hbb650b82),
	.w5(32'hbaab3af1),
	.w6(32'hbb5a9206),
	.w7(32'h3b59f075),
	.w8(32'h3bca0110),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895b742),
	.w1(32'hb9099c4d),
	.w2(32'hb915ce95),
	.w3(32'hb8f7e742),
	.w4(32'hb8885d92),
	.w5(32'hb3c9b5b1),
	.w6(32'hb8246dc8),
	.w7(32'h385e1976),
	.w8(32'h389f5486),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3012e3),
	.w1(32'hbbbe8a7a),
	.w2(32'h3b58260f),
	.w3(32'hbc118fc5),
	.w4(32'hbbdde274),
	.w5(32'hbb15ccd6),
	.w6(32'hbbf2da76),
	.w7(32'hbafb9278),
	.w8(32'h3bd6916b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39110941),
	.w1(32'h38c6d8e2),
	.w2(32'h388869e7),
	.w3(32'h39236262),
	.w4(32'h39031a4c),
	.w5(32'h3905673a),
	.w6(32'h391be8c0),
	.w7(32'h38b88dfc),
	.w8(32'h389b5e30),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2171b9),
	.w1(32'hba3a25fe),
	.w2(32'hb9ae997d),
	.w3(32'hba14ae20),
	.w4(32'hba59a7ed),
	.w5(32'hb92fa0bd),
	.w6(32'hba4bce24),
	.w7(32'hb8b9031a),
	.w8(32'h3a777f78),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc0508),
	.w1(32'hb82bad6c),
	.w2(32'h38680962),
	.w3(32'h3802e57a),
	.w4(32'h37edbcc7),
	.w5(32'h3927f8a7),
	.w6(32'h37c75d1b),
	.w7(32'h386d3937),
	.w8(32'h3900d26b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b12e4),
	.w1(32'hb8583185),
	.w2(32'hb80d466a),
	.w3(32'hb7b78c21),
	.w4(32'h382a78b8),
	.w5(32'h38552356),
	.w6(32'h354267de),
	.w7(32'h37cf6b1b),
	.w8(32'h397e9b24),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9bd2b),
	.w1(32'h3b961432),
	.w2(32'h3b66e91c),
	.w3(32'h39f0730b),
	.w4(32'h39733718),
	.w5(32'hba87d50a),
	.w6(32'hb93778fa),
	.w7(32'hba8d7e75),
	.w8(32'hbb3c2de6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a20af),
	.w1(32'hbb898bbb),
	.w2(32'h3c2f6501),
	.w3(32'hbbbff3aa),
	.w4(32'h3b5d35d9),
	.w5(32'h3c22f4e1),
	.w6(32'hbc757743),
	.w7(32'hbbd3f57e),
	.w8(32'h3b0cc2b3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3573ce),
	.w1(32'hbbce2dd3),
	.w2(32'h3b4a970e),
	.w3(32'hbc36d605),
	.w4(32'hbbf71702),
	.w5(32'hbb39994d),
	.w6(32'hbbae5e3a),
	.w7(32'h3b2c392d),
	.w8(32'h3c1b1bc1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f79cb),
	.w1(32'hbb1b1863),
	.w2(32'h3c1129e9),
	.w3(32'hbc2a0d9a),
	.w4(32'hbb8d0939),
	.w5(32'h3b93804d),
	.w6(32'hbc347903),
	.w7(32'hbb30875e),
	.w8(32'h3c0800e2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b2565),
	.w1(32'h39514b64),
	.w2(32'h384bda43),
	.w3(32'h38202711),
	.w4(32'h390a76bc),
	.w5(32'h38a8881f),
	.w6(32'hb8b6ca6d),
	.w7(32'hb8cb8ae2),
	.w8(32'hb8fff3a1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fb82a),
	.w1(32'h3a73ca33),
	.w2(32'h3a682577),
	.w3(32'h3945ce74),
	.w4(32'h395a8ea9),
	.w5(32'h3994fd39),
	.w6(32'h38021041),
	.w7(32'h3a2bb325),
	.w8(32'h3aeac323),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a7349b),
	.w1(32'hb788869f),
	.w2(32'h35317032),
	.w3(32'h37cfe1a2),
	.w4(32'hb6a81373),
	.w5(32'h37a1877f),
	.w6(32'h37fab959),
	.w7(32'hb41500e7),
	.w8(32'h37827193),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b5ca0),
	.w1(32'h3582774d),
	.w2(32'hb55c2343),
	.w3(32'h386a8cc8),
	.w4(32'h3560a48c),
	.w5(32'h37719115),
	.w6(32'h386a7452),
	.w7(32'hb71bd5aa),
	.w8(32'hb68e3cdf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18c480),
	.w1(32'hbb036de8),
	.w2(32'h3c3b07d9),
	.w3(32'hbc0f2b25),
	.w4(32'hbaf9127f),
	.w5(32'h3b60efff),
	.w6(32'h3aa44e89),
	.w7(32'h3c394192),
	.w8(32'h3c88f108),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ca32a),
	.w1(32'hb9477d88),
	.w2(32'hb8bcb62e),
	.w3(32'hb95acd88),
	.w4(32'hb95ee14f),
	.w5(32'hb90302c1),
	.w6(32'hb93a8741),
	.w7(32'hb93b4f06),
	.w8(32'hb8a80dc8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905646a),
	.w1(32'h399c0418),
	.w2(32'hba704d1d),
	.w3(32'h3989e03a),
	.w4(32'h39c53976),
	.w5(32'hba376deb),
	.w6(32'hb98ac564),
	.w7(32'hb8e1e4e9),
	.w8(32'hba7f30e1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664533),
	.w1(32'hb90a292f),
	.w2(32'hbb03b785),
	.w3(32'hbba86f9a),
	.w4(32'hbafc2e5c),
	.w5(32'hba5c361c),
	.w6(32'h3a279f70),
	.w7(32'h3bb358cf),
	.w8(32'h3b13da8d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374f354c),
	.w1(32'hb791d889),
	.w2(32'h3706f914),
	.w3(32'h38459d0f),
	.w4(32'hb689d477),
	.w5(32'h37a451b3),
	.w6(32'h3855ad68),
	.w7(32'hb7ac3572),
	.w8(32'hb78a305c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fe983),
	.w1(32'hb8f857bd),
	.w2(32'h3b345678),
	.w3(32'hbb77a591),
	.w4(32'hba6e6fef),
	.w5(32'h398de9f4),
	.w6(32'hbafb6399),
	.w7(32'h3af476f6),
	.w8(32'h3b41e37f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9f1fd),
	.w1(32'hba69cb6d),
	.w2(32'hbadb4e18),
	.w3(32'h3a2889f7),
	.w4(32'h3a0b243c),
	.w5(32'hb9be61b7),
	.w6(32'h396ff999),
	.w7(32'h3a34e161),
	.w8(32'hb91c4889),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc988918),
	.w1(32'hbc3e2421),
	.w2(32'h3c376f68),
	.w3(32'hbc91ee9e),
	.w4(32'hbbbbcec0),
	.w5(32'h3c3b8405),
	.w6(32'hbc79e634),
	.w7(32'hbbc4b927),
	.w8(32'h3c1402c1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2a25e),
	.w1(32'h38471b8b),
	.w2(32'hb98bf759),
	.w3(32'hb8c5e577),
	.w4(32'hb8e582e4),
	.w5(32'hba017892),
	.w6(32'h39a0a9a6),
	.w7(32'h376600a3),
	.w8(32'hba611b8e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea17a0),
	.w1(32'h3bfc264e),
	.w2(32'h3bfa5bb8),
	.w3(32'hbc3b208d),
	.w4(32'hbc1a4992),
	.w5(32'hba6916c0),
	.w6(32'hbafa4e01),
	.w7(32'h3c2c779d),
	.w8(32'h3bd16ef6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule