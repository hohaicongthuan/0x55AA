module layer_10_featuremap_319(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4c52eae),
	.w1(32'hb6ad77df),
	.w2(32'h368c4314),
	.w3(32'hb690dcc6),
	.w4(32'h36059e13),
	.w5(32'h35e2f99c),
	.w6(32'hb72395b1),
	.w7(32'hb6adc59b),
	.w8(32'hb6e92512),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9738a),
	.w1(32'hb9830221),
	.w2(32'hb8a8bef8),
	.w3(32'hba151c41),
	.w4(32'hb91972d0),
	.w5(32'h38a71b31),
	.w6(32'hba0bf963),
	.w7(32'h38d2be4a),
	.w8(32'h394d1637),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3639cb38),
	.w1(32'hb65da645),
	.w2(32'hb730ce16),
	.w3(32'hb5e401bc),
	.w4(32'hb680cc99),
	.w5(32'hb657c5c8),
	.w6(32'hb6863bd7),
	.w7(32'hb7091ac8),
	.w8(32'hb6a7a4ba),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82bdafc),
	.w1(32'hb69f1ee6),
	.w2(32'hb8f71e3a),
	.w3(32'hb83ab454),
	.w4(32'h388181a3),
	.w5(32'hb988e050),
	.w6(32'hb7908745),
	.w7(32'h386d3af7),
	.w8(32'hb918c8ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807dffa),
	.w1(32'hb8485664),
	.w2(32'hb86c6fbb),
	.w3(32'hb803d7e6),
	.w4(32'hb83c334e),
	.w5(32'hb84be0d7),
	.w6(32'hb7ecca89),
	.w7(32'hb8027073),
	.w8(32'hb82ce221),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6991d53),
	.w1(32'hb6896954),
	.w2(32'hb47cc1e2),
	.w3(32'hb6f56ff8),
	.w4(32'h34941e80),
	.w5(32'hb68eebdb),
	.w6(32'hb737b7b5),
	.w7(32'hb67c596c),
	.w8(32'hb6fc355d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7d313),
	.w1(32'hb9fa42f6),
	.w2(32'hb9b4f167),
	.w3(32'hba1fad41),
	.w4(32'hb9f1aeb2),
	.w5(32'hb8e5c779),
	.w6(32'hb90b3cff),
	.w7(32'h39d048be),
	.w8(32'h39e0fe83),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4400f),
	.w1(32'h39ec87ee),
	.w2(32'h3a223ada),
	.w3(32'h3a55085f),
	.w4(32'h3a81c756),
	.w5(32'h392148a1),
	.w6(32'h3b02cceb),
	.w7(32'h3a4ad3a2),
	.w8(32'hb84c1b3e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39746369),
	.w1(32'h39865f19),
	.w2(32'h3999bafb),
	.w3(32'h38f766eb),
	.w4(32'h3905e124),
	.w5(32'h39ae1b95),
	.w6(32'hb93487a5),
	.w7(32'hb8d37f31),
	.w8(32'h398d401e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcfb8a),
	.w1(32'hb910416e),
	.w2(32'h3a05c979),
	.w3(32'h3959579d),
	.w4(32'hba0133e6),
	.w5(32'h3a2fed29),
	.w6(32'h3995878e),
	.w7(32'hba286f2a),
	.w8(32'h39bd0b07),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bc953),
	.w1(32'h370a9c99),
	.w2(32'hb8047625),
	.w3(32'h38d0ce8e),
	.w4(32'hb782fa1d),
	.w5(32'hb74c4226),
	.w6(32'h3828ed3d),
	.w7(32'h36e25992),
	.w8(32'h351e1eee),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb870efa1),
	.w1(32'hb92ac68d),
	.w2(32'hb982162e),
	.w3(32'hba10d084),
	.w4(32'hb9b37024),
	.w5(32'hb9ac65fb),
	.w6(32'h39c4cf5f),
	.w7(32'h399a226a),
	.w8(32'h39b8ccd5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13c3b1),
	.w1(32'h389cdfb8),
	.w2(32'h39659893),
	.w3(32'h39cccbcc),
	.w4(32'hb9d83618),
	.w5(32'h38f5559b),
	.w6(32'h3a07b5c6),
	.w7(32'hb9eb8bad),
	.w8(32'h3894bd29),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3805ffcb),
	.w1(32'hb9419f39),
	.w2(32'hb81bfb11),
	.w3(32'hb9b22e0e),
	.w4(32'hb9baea33),
	.w5(32'hb940e9ce),
	.w6(32'h392bd025),
	.w7(32'hb7bfd7e8),
	.w8(32'hb8750d9c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de06d7),
	.w1(32'hb8ae517a),
	.w2(32'h3938bd5b),
	.w3(32'hb8beddf5),
	.w4(32'hba153e28),
	.w5(32'hb8285ea0),
	.w6(32'hb9929299),
	.w7(32'hb9d5b41b),
	.w8(32'hb9312bd2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399429c0),
	.w1(32'hb8b4bcc2),
	.w2(32'h39e3666c),
	.w3(32'h397c9d86),
	.w4(32'hb944f30d),
	.w5(32'h39e3ecbf),
	.w6(32'h39a663f7),
	.w7(32'h38a91f73),
	.w8(32'h39f902a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3682f2a3),
	.w1(32'hb72770f4),
	.w2(32'hb81c9f10),
	.w3(32'hb6d5a8b8),
	.w4(32'hb7194445),
	.w5(32'h3608d2ba),
	.w6(32'h37d12e9a),
	.w7(32'h366ebe35),
	.w8(32'hb6ebdd60),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a050009),
	.w1(32'h3a0a60ad),
	.w2(32'h396c9088),
	.w3(32'h3a49133b),
	.w4(32'hb9c37e17),
	.w5(32'h3804249c),
	.w6(32'h3a669d46),
	.w7(32'hba12e95c),
	.w8(32'hba078aef),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bb616),
	.w1(32'h3a27bc8d),
	.w2(32'h3a05b2f5),
	.w3(32'h39a990f1),
	.w4(32'h383f6135),
	.w5(32'h398bded9),
	.w6(32'h3a0138ba),
	.w7(32'hb8648b4c),
	.w8(32'hb78f06af),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66948ab),
	.w1(32'hb71c0e5a),
	.w2(32'hb5c70d43),
	.w3(32'hb7a3442e),
	.w4(32'hb79a0a4b),
	.w5(32'hb74b082e),
	.w6(32'hb76a1889),
	.w7(32'h35ea5425),
	.w8(32'hb6b6eff0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f551b5),
	.w1(32'hb6d0086d),
	.w2(32'h33fed608),
	.w3(32'hb7a62e6a),
	.w4(32'h36931c48),
	.w5(32'hb6831f6c),
	.w6(32'hb7b25917),
	.w7(32'hb6bc469e),
	.w8(32'hb73860c1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b657f7),
	.w1(32'hb8c3f886),
	.w2(32'h36c677cb),
	.w3(32'hb9ba002c),
	.w4(32'hb8932137),
	.w5(32'h385c46ad),
	.w6(32'hb8fc328a),
	.w7(32'h38f870f0),
	.w8(32'h38f91560),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b077f84),
	.w1(32'h3af68183),
	.w2(32'h393c13b7),
	.w3(32'h3b0f5a98),
	.w4(32'h381cbab6),
	.w5(32'h393c39e9),
	.w6(32'h3a90fc05),
	.w7(32'hb898bf5f),
	.w8(32'h38721a62),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f356f),
	.w1(32'hb9564d47),
	.w2(32'h39afa9c0),
	.w3(32'hb97d1ec2),
	.w4(32'hba77849c),
	.w5(32'hb819174d),
	.w6(32'hb95a01f0),
	.w7(32'hba3c3365),
	.w8(32'h39235ff2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e90e62),
	.w1(32'hb953c0ba),
	.w2(32'h39799e23),
	.w3(32'hb9b5e2c1),
	.w4(32'hba4027e1),
	.w5(32'h36d3c974),
	.w6(32'hb9e9f9d6),
	.w7(32'hb794f8a8),
	.w8(32'h3a23b81d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887c09b),
	.w1(32'hb8c24fc9),
	.w2(32'hb909c82d),
	.w3(32'h38ddc2b4),
	.w4(32'hb8a05b8f),
	.w5(32'hb8c40dc9),
	.w6(32'h381b5d07),
	.w7(32'hb94637e7),
	.w8(32'hb97e9863),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be7386),
	.w1(32'hb71fb8af),
	.w2(32'hb8204fc2),
	.w3(32'hb7ab217f),
	.w4(32'hb712c905),
	.w5(32'hb7e03171),
	.w6(32'hb818066b),
	.w7(32'hb78160c6),
	.w8(32'hb81c5c4c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba227da7),
	.w1(32'hb979e785),
	.w2(32'h39c820fb),
	.w3(32'hba905afc),
	.w4(32'hb9de07e3),
	.w5(32'h3a397616),
	.w6(32'hba873bcb),
	.w7(32'hb9b19774),
	.w8(32'h3a59b3e7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940b6ab),
	.w1(32'hb93c7c03),
	.w2(32'hb91c50fe),
	.w3(32'hb92c9abf),
	.w4(32'hb93bb5d1),
	.w5(32'hb93394c1),
	.w6(32'hb7d2910f),
	.w7(32'hb8d64269),
	.w8(32'hb8c3e479),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db583c),
	.w1(32'hba0f047e),
	.w2(32'h39bc596a),
	.w3(32'hba3d32b0),
	.w4(32'hba837163),
	.w5(32'h39b1bb5b),
	.w6(32'hbabc079f),
	.w7(32'hba90ce0a),
	.w8(32'h39acbc93),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb763c599),
	.w1(32'hb6f76bd0),
	.w2(32'hb776c35b),
	.w3(32'hb6a36a4e),
	.w4(32'h36259464),
	.w5(32'hb6241963),
	.w6(32'hb66b9360),
	.w7(32'hb4d45765),
	.w8(32'hb71789fc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3747dfaa),
	.w1(32'hb7691772),
	.w2(32'hb7e321fa),
	.w3(32'h3736c04c),
	.w4(32'hb684b096),
	.w5(32'hb7d9a90c),
	.w6(32'h3799cd3e),
	.w7(32'hb608d963),
	.w8(32'hb77d0da7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c98d25),
	.w1(32'hb8c00d4f),
	.w2(32'h394947cf),
	.w3(32'h389518ed),
	.w4(32'hb9820dd5),
	.w5(32'h38f2c252),
	.w6(32'h39caf9c8),
	.w7(32'hb8cbb10e),
	.w8(32'h38224d5f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908b7b8),
	.w1(32'hb80598d4),
	.w2(32'h39116a59),
	.w3(32'hb81a3c61),
	.w4(32'hb8fbd540),
	.w5(32'h389ca64c),
	.w6(32'hb89f8cb0),
	.w7(32'hb85ce398),
	.w8(32'h38a86835),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c0c779),
	.w1(32'hb83906ed),
	.w2(32'hb81d87c1),
	.w3(32'hb81aa786),
	.w4(32'hb89293dc),
	.w5(32'hb8a1cd92),
	.w6(32'h388849d5),
	.w7(32'h3845b5de),
	.w8(32'hb7b60c71),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f0230),
	.w1(32'h37be81d4),
	.w2(32'hb863e562),
	.w3(32'h392560ed),
	.w4(32'h3932a10f),
	.w5(32'hb60485bb),
	.w6(32'h39bcd04e),
	.w7(32'h39af7e66),
	.w8(32'h39923eca),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b74a73),
	.w1(32'h39350da9),
	.w2(32'hbaa136e2),
	.w3(32'h37d477c6),
	.w4(32'h3972cfe0),
	.w5(32'hbabd4ceb),
	.w6(32'h3a1df292),
	.w7(32'h3a36dde8),
	.w8(32'hb83bf0b5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ce8f9),
	.w1(32'hba61bc31),
	.w2(32'hba5be1c9),
	.w3(32'hba2a265b),
	.w4(32'hba218808),
	.w5(32'hb80bda18),
	.w6(32'hb96ab783),
	.w7(32'h3a188141),
	.w8(32'h39ecfcdd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a093a),
	.w1(32'hba447d79),
	.w2(32'hb8d0cd64),
	.w3(32'hbb022cc0),
	.w4(32'hba092f59),
	.w5(32'h395a3c81),
	.w6(32'hbab3c621),
	.w7(32'h39c13703),
	.w8(32'h3a3c9378),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e32008),
	.w1(32'hb84ac52d),
	.w2(32'h38b066c4),
	.w3(32'hb8afc014),
	.w4(32'h389f4eb0),
	.w5(32'h396dc061),
	.w6(32'hb8f70ece),
	.w7(32'h394bde5e),
	.w8(32'h39ad9b71),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b26374),
	.w1(32'h381c5d07),
	.w2(32'h38150423),
	.w3(32'h385dba81),
	.w4(32'h38812d4f),
	.w5(32'h38505a23),
	.w6(32'h371cf6cc),
	.w7(32'h37991835),
	.w8(32'h370d6c37),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb738392b),
	.w1(32'h3640fe73),
	.w2(32'hb85e0ecd),
	.w3(32'hb7ae18b4),
	.w4(32'h36db8f7d),
	.w5(32'hb842d8d8),
	.w6(32'hb8728785),
	.w7(32'hb74ddf04),
	.w8(32'hb83a170a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807df03),
	.w1(32'hb91221bc),
	.w2(32'hb9a35a66),
	.w3(32'hb6de801b),
	.w4(32'hb9b8bd56),
	.w5(32'hb9e5368f),
	.w6(32'h3806dbfa),
	.w7(32'hb98c81ea),
	.w8(32'hb9bf716d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fdafb),
	.w1(32'h392d1067),
	.w2(32'h3a529338),
	.w3(32'h39dc3462),
	.w4(32'hb9ce45e8),
	.w5(32'h3a65a882),
	.w6(32'h3a0226e9),
	.w7(32'hba17f90a),
	.w8(32'h39871e16),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a3fc2),
	.w1(32'hb8c27198),
	.w2(32'h39e4fdf3),
	.w3(32'hb835609f),
	.w4(32'hba274415),
	.w5(32'h395edd49),
	.w6(32'hb9c8d5d5),
	.w7(32'hba373443),
	.w8(32'h38c246a0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf1cb8),
	.w1(32'hb946a39a),
	.w2(32'h399cf80c),
	.w3(32'h3913d5d3),
	.w4(32'hba460703),
	.w5(32'h386bdc8b),
	.w6(32'hb806072f),
	.w7(32'hba20441c),
	.w8(32'h38ad8ca3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a628a),
	.w1(32'h39d81d40),
	.w2(32'h3a27face),
	.w3(32'h3a06818c),
	.w4(32'h391b3a4a),
	.w5(32'h39dc63d6),
	.w6(32'h3a61cf26),
	.w7(32'h39c030e1),
	.w8(32'h3a16cd5b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3893eaa5),
	.w1(32'h39febb42),
	.w2(32'h39929720),
	.w3(32'h3a47000c),
	.w4(32'hb7c42291),
	.w5(32'hba109c77),
	.w6(32'h3aa25e24),
	.w7(32'hba1ec5a3),
	.w8(32'hba76f8fe),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f7e09),
	.w1(32'hb866e15a),
	.w2(32'h36a81985),
	.w3(32'hb89d59be),
	.w4(32'hb848efd4),
	.w5(32'hb70359b2),
	.w6(32'hb8b852d7),
	.w7(32'hb8bde856),
	.w8(32'hb8dc6276),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38804aee),
	.w1(32'h3701478f),
	.w2(32'h381b84e1),
	.w3(32'h372d2742),
	.w4(32'hb7c0061b),
	.w5(32'h380f8b60),
	.w6(32'hb91e9f20),
	.w7(32'hb923dffb),
	.w8(32'h3787b20d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f5bd2),
	.w1(32'hb8d3f3f0),
	.w2(32'hb7ca784b),
	.w3(32'hb9527e72),
	.w4(32'hb94f62fe),
	.w5(32'hb8f4809e),
	.w6(32'hb972a685),
	.w7(32'hb96b616b),
	.w8(32'hb91897c4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcc5df),
	.w1(32'h399dd4ed),
	.w2(32'h39205b60),
	.w3(32'h3981b612),
	.w4(32'hb6d36ca8),
	.w5(32'h396652f0),
	.w6(32'h39196be1),
	.w7(32'h37f23bb2),
	.w8(32'h39314003),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936891b),
	.w1(32'h392d570d),
	.w2(32'h38fe0e47),
	.w3(32'h397ce90a),
	.w4(32'h3926d4f8),
	.w5(32'h3869f974),
	.w6(32'h3924f724),
	.w7(32'h383f4850),
	.w8(32'h36bf6b2b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac0a35),
	.w1(32'h3a7a0ba3),
	.w2(32'h39bbf346),
	.w3(32'h3a9ab6b5),
	.w4(32'h38a731fb),
	.w5(32'hb9c81548),
	.w6(32'h3a770eb6),
	.w7(32'hb9b00162),
	.w8(32'hba28a204),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39777665),
	.w1(32'h39182a83),
	.w2(32'h39553bb3),
	.w3(32'h37bb74c0),
	.w4(32'hb8b8ec80),
	.w5(32'h3867239e),
	.w6(32'h3848d067),
	.w7(32'hb7fbae16),
	.w8(32'h38085e88),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ea81c6),
	.w1(32'hb7fd2dc3),
	.w2(32'h36ffb7f4),
	.w3(32'hb80de426),
	.w4(32'hb81f8aa6),
	.w5(32'hb6b18256),
	.w6(32'hb82d6a09),
	.w7(32'hb85ca401),
	.w8(32'hb782a152),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f55e21),
	.w1(32'h3604c034),
	.w2(32'h3603150f),
	.w3(32'hb661fdbf),
	.w4(32'h3674e9b5),
	.w5(32'h3609742f),
	.w6(32'hb7390929),
	.w7(32'h36191fb5),
	.w8(32'h368734b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f71179),
	.w1(32'h36a8d009),
	.w2(32'h37803bf6),
	.w3(32'hb82fc31d),
	.w4(32'hb848e5ba),
	.w5(32'h3735ba66),
	.w6(32'hb8c56f68),
	.w7(32'hb831cdef),
	.w8(32'h3833c563),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a63672),
	.w1(32'hb8fce06e),
	.w2(32'hb8d8c403),
	.w3(32'hb839eb13),
	.w4(32'hb8b78c4e),
	.w5(32'hb8c66d79),
	.w6(32'h391e31b9),
	.w7(32'h3866a1c2),
	.w8(32'hb620ac3d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7185512),
	.w1(32'h3726eea4),
	.w2(32'hb6df77c6),
	.w3(32'hb7830688),
	.w4(32'hb7b90982),
	.w5(32'hb7daf0e4),
	.w6(32'h34da3f3d),
	.w7(32'hb6df93d3),
	.w8(32'h37c62230),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a53e94),
	.w1(32'h3a1b9bca),
	.w2(32'h39a5adfc),
	.w3(32'h39cc5af0),
	.w4(32'h397355e3),
	.w5(32'h39c086c8),
	.w6(32'h39f17027),
	.w7(32'h39781d11),
	.w8(32'h398a59ba),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a370e05),
	.w1(32'h390b36a1),
	.w2(32'hb90366f0),
	.w3(32'h3a405a52),
	.w4(32'h38c854a5),
	.w5(32'h38c82a90),
	.w6(32'h39f359a7),
	.w7(32'h389628ba),
	.w8(32'h3891f698),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65716cf),
	.w1(32'hb6c3a7d3),
	.w2(32'hb7055f85),
	.w3(32'h370ae703),
	.w4(32'h36331853),
	.w5(32'hb7d0d9b5),
	.w6(32'hb6be27b9),
	.w7(32'hb6de8f64),
	.w8(32'hb8052ea6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb605b037),
	.w1(32'h36227b1c),
	.w2(32'h34846d59),
	.w3(32'hb48996a1),
	.w4(32'h34b51d6a),
	.w5(32'h3704eca2),
	.w6(32'hb7601794),
	.w7(32'hb72c42a5),
	.w8(32'hb683101a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85cf3c8),
	.w1(32'hb77a47b2),
	.w2(32'h35d84828),
	.w3(32'hb83bcb7f),
	.w4(32'hb583bdfe),
	.w5(32'h360bf18f),
	.w6(32'hb886ab00),
	.w7(32'hb7c7552f),
	.w8(32'hb7803dfc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72eaac0),
	.w1(32'h36273286),
	.w2(32'hb75324e8),
	.w3(32'h35da917a),
	.w4(32'h36bb937f),
	.w5(32'hb71dcb8c),
	.w6(32'hb74f678d),
	.w7(32'hb64889d8),
	.w8(32'hb78d272a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9104a44),
	.w1(32'h38bc07bf),
	.w2(32'h392d050f),
	.w3(32'hb9bf0e0b),
	.w4(32'hba28d205),
	.w5(32'hb9598404),
	.w6(32'h3a95c098),
	.w7(32'hb96f422d),
	.w8(32'h375f3a0e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87e3124),
	.w1(32'hb9bf0984),
	.w2(32'h384adb36),
	.w3(32'h3a251172),
	.w4(32'hb7c21a80),
	.w5(32'h3a01d0fe),
	.w6(32'h3a6185b8),
	.w7(32'h3a2d1139),
	.w8(32'h3a28e154),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a040b0e),
	.w1(32'h3a1399ec),
	.w2(32'h39c5efbc),
	.w3(32'h39ea0e38),
	.w4(32'h37c5f40f),
	.w5(32'h39c99fa1),
	.w6(32'h3a43ba62),
	.w7(32'h3a2b34d5),
	.w8(32'h3a45ae61),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b529c0),
	.w1(32'hba08b708),
	.w2(32'h39831f12),
	.w3(32'hba81ca02),
	.w4(32'hba87f9ed),
	.w5(32'hb9b29b81),
	.w6(32'hba4d8029),
	.w7(32'hb9b10174),
	.w8(32'h3a132bfe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fd363f),
	.w1(32'hb5c8112a),
	.w2(32'hb6dbdc0f),
	.w3(32'hb5ef800c),
	.w4(32'h35da5f68),
	.w5(32'hb72f6f00),
	.w6(32'hb73c59c7),
	.w7(32'hb70ea3e0),
	.w8(32'hb7b4ae9a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb781681a),
	.w1(32'hb6d7f693),
	.w2(32'hb7aa660a),
	.w3(32'hb7517105),
	.w4(32'hb612c5ce),
	.w5(32'hb78452b9),
	.w6(32'hb8078bc9),
	.w7(32'hb7a8b341),
	.w8(32'hb8001789),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3561ad3f),
	.w1(32'h37260da1),
	.w2(32'hb725d37f),
	.w3(32'hb60751df),
	.w4(32'h3743e8d8),
	.w5(32'h36d7ebe8),
	.w6(32'hb7d7db9a),
	.w7(32'hb72e4453),
	.w8(32'hb6cc075e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c0c5f),
	.w1(32'h39e3533c),
	.w2(32'h3918f168),
	.w3(32'h3872c7de),
	.w4(32'h390d054d),
	.w5(32'h390c8f2d),
	.w6(32'h39876ea3),
	.w7(32'h39c0a218),
	.w8(32'h39ada3f9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a081d),
	.w1(32'h361e886b),
	.w2(32'hb6f050c8),
	.w3(32'hb6efb5f9),
	.w4(32'h371c37df),
	.w5(32'hb67751d6),
	.w6(32'hb7e32067),
	.w7(32'hb734567a),
	.w8(32'hb78d2add),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914e48c),
	.w1(32'h39a233f0),
	.w2(32'hb8950293),
	.w3(32'hb71a1d01),
	.w4(32'hb84abd88),
	.w5(32'hba1f93aa),
	.w6(32'h399e582a),
	.w7(32'h37bde160),
	.w8(32'hb9cddf90),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9aa5b),
	.w1(32'h3a34dce5),
	.w2(32'h3a82396e),
	.w3(32'h39812a73),
	.w4(32'h3a32f049),
	.w5(32'h3a0120b3),
	.w6(32'h3aa81b1d),
	.w7(32'h3a61eec5),
	.w8(32'h39d06105),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9740524),
	.w1(32'hba06d5de),
	.w2(32'hb938ac0e),
	.w3(32'hba128271),
	.w4(32'hba3920c1),
	.w5(32'hb87ce4b9),
	.w6(32'hba05f26b),
	.w7(32'hba456bd6),
	.w8(32'hb963620d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d20c69),
	.w1(32'h39a81512),
	.w2(32'h38cf5450),
	.w3(32'h39009d7f),
	.w4(32'hb89f5c0c),
	.w5(32'hb794bb29),
	.w6(32'h38ba43be),
	.w7(32'hb925ccff),
	.w8(32'h38c3b7b9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bea2d6),
	.w1(32'hb898fe70),
	.w2(32'hb92074d3),
	.w3(32'hb989da91),
	.w4(32'hb9c4cc63),
	.w5(32'hb980a792),
	.w6(32'h3898726a),
	.w7(32'hb80a9f8a),
	.w8(32'h37aa36e7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988f3cd),
	.w1(32'hb8cb8026),
	.w2(32'h393c39fc),
	.w3(32'h37cc5de9),
	.w4(32'hb9b996f3),
	.w5(32'h3919d7cf),
	.w6(32'h38e73a6e),
	.w7(32'hb9856fd5),
	.w8(32'h38fcef0e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4c130),
	.w1(32'h399f07ea),
	.w2(32'h39604c69),
	.w3(32'h396c8d16),
	.w4(32'h382702cc),
	.w5(32'h37913a4c),
	.w6(32'h3a01282c),
	.w7(32'hb8a3c2c0),
	.w8(32'hb8457a4e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb547bfc7),
	.w1(32'hb68d36f5),
	.w2(32'hb6b0734b),
	.w3(32'hb519eaaf),
	.w4(32'h36adcbb3),
	.w5(32'h36a7603f),
	.w6(32'hb653a67f),
	.w7(32'hb59099a5),
	.w8(32'hb6927b64),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c673d5),
	.w1(32'h360253d5),
	.w2(32'hb6ad202f),
	.w3(32'hb5cf3088),
	.w4(32'hb66d5c89),
	.w5(32'hb53d09d8),
	.w6(32'hb6d6d308),
	.w7(32'hb70796a5),
	.w8(32'hb653afa5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71bba16),
	.w1(32'hb66323af),
	.w2(32'hb730d448),
	.w3(32'hb7cb1a1c),
	.w4(32'hb613245d),
	.w5(32'hb7863b33),
	.w6(32'hb7b0802e),
	.w7(32'hb6702ea7),
	.w8(32'hb74e735a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd3724),
	.w1(32'hb752b434),
	.w2(32'h37d3ae27),
	.w3(32'hb857134f),
	.w4(32'hb74b56a4),
	.w5(32'h371e452d),
	.w6(32'hb8a29007),
	.w7(32'hb7cf4716),
	.w8(32'h376bbf10),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886c0b8),
	.w1(32'hb9beeadc),
	.w2(32'hb9976c7a),
	.w3(32'hb9674ee2),
	.w4(32'hb9740ab6),
	.w5(32'h37c7f00e),
	.w6(32'hb90a5cbc),
	.w7(32'h39ae944c),
	.w8(32'h39fe92e7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85bee3c),
	.w1(32'hb84fac88),
	.w2(32'hb8f47a09),
	.w3(32'hb9210288),
	.w4(32'hb8aa7317),
	.w5(32'hb932bd21),
	.w6(32'hb7ffd142),
	.w7(32'h361928bc),
	.w8(32'hb90fc13d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1a5e2),
	.w1(32'h38fc366d),
	.w2(32'h39526e14),
	.w3(32'h39f7d312),
	.w4(32'h37df6985),
	.w5(32'hb6a8e2db),
	.w6(32'hb95285a3),
	.w7(32'hb94aed1b),
	.w8(32'h38e6fd9a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a092fd1),
	.w1(32'h3981d290),
	.w2(32'h3778515b),
	.w3(32'h3a87857c),
	.w4(32'h398f08f9),
	.w5(32'hb8e4c12f),
	.w6(32'h3aceac99),
	.w7(32'h3a331215),
	.w8(32'h37832ba9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb09da),
	.w1(32'hb9884be2),
	.w2(32'hb8fe2a93),
	.w3(32'hb9bad995),
	.w4(32'hb996fb5f),
	.w5(32'hb99c7935),
	.w6(32'hb87700bc),
	.w7(32'h38d64d38),
	.w8(32'hb86813de),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ed092),
	.w1(32'h3a28ad62),
	.w2(32'hba33a473),
	.w3(32'h3a456dca),
	.w4(32'h39160a3e),
	.w5(32'hba3e444f),
	.w6(32'h3ad0ffae),
	.w7(32'h39edda8c),
	.w8(32'h39429f0b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb9865),
	.w1(32'hb956e613),
	.w2(32'hb9780e91),
	.w3(32'hb9961dff),
	.w4(32'hb98a0a74),
	.w5(32'h38f49efd),
	.w6(32'hb9d847ff),
	.w7(32'hb8f6e4b2),
	.w8(32'h39b96eb4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdc813),
	.w1(32'h3ac18326),
	.w2(32'h3a526a2d),
	.w3(32'h3a738c75),
	.w4(32'h3a1b027e),
	.w5(32'h39cf603a),
	.w6(32'h3990b0dd),
	.w7(32'h3a0f4ea2),
	.w8(32'h3a69b9d5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b6ff9),
	.w1(32'hb9920003),
	.w2(32'h39065b17),
	.w3(32'hba16b0d8),
	.w4(32'hba1573a2),
	.w5(32'h37445588),
	.w6(32'hba15e78f),
	.w7(32'hb9fee286),
	.w8(32'h398b80af),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef7308),
	.w1(32'hb886f680),
	.w2(32'h391cdf3a),
	.w3(32'hb93ebd6b),
	.w4(32'hb9a49a26),
	.w5(32'h38a03ab1),
	.w6(32'hba0ab0c5),
	.w7(32'hb98bc097),
	.w8(32'hb716d264),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e8d31),
	.w1(32'hb8830e2b),
	.w2(32'h3822f0e8),
	.w3(32'hb8c177e5),
	.w4(32'hb8284f5d),
	.w5(32'hb7bbafd7),
	.w6(32'hb9555095),
	.w7(32'hb96f3296),
	.w8(32'hb953689b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c56c34),
	.w1(32'h39286552),
	.w2(32'h3a32ded7),
	.w3(32'h39127de1),
	.w4(32'hba3f9d46),
	.w5(32'h39ef8a09),
	.w6(32'h39824893),
	.w7(32'hba5ecc3a),
	.w8(32'hba8a036d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8893905),
	.w1(32'h3a8b362b),
	.w2(32'hba37b139),
	.w3(32'h3aa0c848),
	.w4(32'h3903ddf9),
	.w5(32'hb9d63830),
	.w6(32'h3abed4b8),
	.w7(32'hb86dda09),
	.w8(32'h3aade001),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab658e1),
	.w1(32'h3a002bd7),
	.w2(32'hb98aea90),
	.w3(32'h3a966beb),
	.w4(32'h39cd3d88),
	.w5(32'h3b2c0766),
	.w6(32'h3a3e1826),
	.w7(32'h3b443d15),
	.w8(32'h3bd2e97e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d56d),
	.w1(32'h3b35216b),
	.w2(32'hba14399e),
	.w3(32'h3b97bd9b),
	.w4(32'h3ab99970),
	.w5(32'hb9f49fb8),
	.w6(32'h3bff169d),
	.w7(32'h3b7a2509),
	.w8(32'hbac9fbaf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea81e),
	.w1(32'h390586e9),
	.w2(32'hb9f2c700),
	.w3(32'hba4ae3cd),
	.w4(32'hb9ab5de9),
	.w5(32'h3b0c0b4e),
	.w6(32'hbb7277b3),
	.w7(32'hbae67f3d),
	.w8(32'h3b8166b1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d475f),
	.w1(32'hba27e6ae),
	.w2(32'hbb84a6ff),
	.w3(32'h3b848104),
	.w4(32'hbb1907d7),
	.w5(32'hbade4408),
	.w6(32'h3a9247c6),
	.w7(32'hbb971569),
	.w8(32'hbabf56aa),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c92e),
	.w1(32'h39f28e31),
	.w2(32'h3a879f04),
	.w3(32'h3a9a3e22),
	.w4(32'h3af465e5),
	.w5(32'h3bb269df),
	.w6(32'h3b213652),
	.w7(32'h3b262309),
	.w8(32'h3b07d8da),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80ba61),
	.w1(32'h3b36c92e),
	.w2(32'h3a0103c7),
	.w3(32'h3bdaeb6a),
	.w4(32'h3bbab7ce),
	.w5(32'hb93b5a19),
	.w6(32'h3b3256ec),
	.w7(32'h3b6ad3fa),
	.w8(32'h3a03d512),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810368),
	.w1(32'h3a4eb9ba),
	.w2(32'h390a65d9),
	.w3(32'hba25e442),
	.w4(32'hbab7810c),
	.w5(32'hba85d80b),
	.w6(32'hb94a869d),
	.w7(32'hb588f9c4),
	.w8(32'h3a880c00),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8462bf),
	.w1(32'hbac967b6),
	.w2(32'h3b86d5f2),
	.w3(32'hb9fba192),
	.w4(32'h3b46b5a2),
	.w5(32'h3b94673d),
	.w6(32'hba879715),
	.w7(32'h3ba0a4ba),
	.w8(32'h3b897905),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ad73),
	.w1(32'h3a7b2942),
	.w2(32'h392e5f9c),
	.w3(32'h3b2db59e),
	.w4(32'h373ba4ab),
	.w5(32'h3b0a1e98),
	.w6(32'h3a3d7adb),
	.w7(32'hba083bff),
	.w8(32'h39e8f933),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a454aee),
	.w1(32'h3ac10bb3),
	.w2(32'h3a842a0d),
	.w3(32'h3b39290e),
	.w4(32'h3b4d924e),
	.w5(32'h3ae6e7ed),
	.w6(32'h3b1020b2),
	.w7(32'h3aa7097a),
	.w8(32'h3a147139),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954473),
	.w1(32'h3b4ab49a),
	.w2(32'h3b9e1f9a),
	.w3(32'hb939aaff),
	.w4(32'h3ab78fc6),
	.w5(32'h39bb0c4d),
	.w6(32'hbaea2c03),
	.w7(32'h3a111233),
	.w8(32'hbb189fe8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba909a78),
	.w1(32'hbaf1c221),
	.w2(32'h39f1ad58),
	.w3(32'h3a164da0),
	.w4(32'h3a4570b1),
	.w5(32'hbb3e4f4f),
	.w6(32'hbb6008f4),
	.w7(32'hba9c433c),
	.w8(32'hbb8d94ea),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88e2cf),
	.w1(32'h3b6d69ae),
	.w2(32'h3c05415a),
	.w3(32'hbb4fc108),
	.w4(32'h3be68b33),
	.w5(32'h392c7417),
	.w6(32'hbb062ba2),
	.w7(32'h3c09074c),
	.w8(32'h3a107d4d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2475ff),
	.w1(32'h3a43d47e),
	.w2(32'h3ac54095),
	.w3(32'h3a9ec6e9),
	.w4(32'h3aed5468),
	.w5(32'h3bbd4649),
	.w6(32'h3a97b535),
	.w7(32'h3a8ea511),
	.w8(32'h3c515f3e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a481),
	.w1(32'h3af6544b),
	.w2(32'h3aa82cca),
	.w3(32'h3c0ef09d),
	.w4(32'h3b9cc0e7),
	.w5(32'h3a5be063),
	.w6(32'h3c7708a8),
	.w7(32'h3c28cfc9),
	.w8(32'h39e5858c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fb532),
	.w1(32'h3af8cb0e),
	.w2(32'h3b343244),
	.w3(32'h3b64029b),
	.w4(32'hbb0427e0),
	.w5(32'h39c4ccfc),
	.w6(32'h3ad4e8e0),
	.w7(32'h3aff6354),
	.w8(32'hbb1d9954),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7409e1),
	.w1(32'h3b840eeb),
	.w2(32'h3bc18961),
	.w3(32'hbaae6c22),
	.w4(32'h3be2d7b7),
	.w5(32'h3bb3dbfd),
	.w6(32'hbb40ab59),
	.w7(32'h3bcec74c),
	.w8(32'h3c0fb003),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ad73),
	.w1(32'h3bb59959),
	.w2(32'h3aa78f72),
	.w3(32'h3ba6fb85),
	.w4(32'hb837add1),
	.w5(32'hbb1f8a3a),
	.w6(32'h3be8e051),
	.w7(32'h3b0c0cbe),
	.w8(32'hbbbe23de),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42e83),
	.w1(32'hba3c7747),
	.w2(32'h39acf389),
	.w3(32'hb9f85f6f),
	.w4(32'h39ce613d),
	.w5(32'hba4c7780),
	.w6(32'hbb1ed520),
	.w7(32'hba34f70a),
	.w8(32'hbb556198),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bbe3a),
	.w1(32'hbacb2c41),
	.w2(32'hbab8d40e),
	.w3(32'h3aff95e3),
	.w4(32'hb81e934c),
	.w5(32'hbb4abb02),
	.w6(32'hba8fa48b),
	.w7(32'hbb10e7f3),
	.w8(32'hbba1c5b7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9db67),
	.w1(32'hbbbde6d4),
	.w2(32'hbbca11e3),
	.w3(32'hbb3420c4),
	.w4(32'hbb1a3914),
	.w5(32'h398b0656),
	.w6(32'hbb9807f6),
	.w7(32'hbb80f15a),
	.w8(32'hba10ac35),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa10d4),
	.w1(32'h3b0e4db2),
	.w2(32'h3bea0c41),
	.w3(32'hbb0fae2d),
	.w4(32'h3b4c9dc1),
	.w5(32'hbb10293f),
	.w6(32'hbb485b60),
	.w7(32'h3b08834b),
	.w8(32'hbb3bf8c8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a8aaf),
	.w1(32'hba62a7a0),
	.w2(32'h3b82d603),
	.w3(32'h393e8ba2),
	.w4(32'h3bb03f3b),
	.w5(32'hbb91d85e),
	.w6(32'hb997dab5),
	.w7(32'h3b940094),
	.w8(32'hbb4b442f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13aadd),
	.w1(32'h3b483a56),
	.w2(32'h3b2b579b),
	.w3(32'hbbaaf911),
	.w4(32'hbb3dcfa7),
	.w5(32'hbaa5f218),
	.w6(32'hbb88935e),
	.w7(32'hbaf82d57),
	.w8(32'hbb577427),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c739d),
	.w1(32'hbb2101d5),
	.w2(32'h3a2ff271),
	.w3(32'h3ab5682f),
	.w4(32'h3b367387),
	.w5(32'hbb51a922),
	.w6(32'hbacb432f),
	.w7(32'h3b0bd01c),
	.w8(32'hbad26a14),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d5ac),
	.w1(32'h3b140425),
	.w2(32'h3b6d0cf6),
	.w3(32'hbb5c7693),
	.w4(32'hbac4db03),
	.w5(32'h3bb4eef4),
	.w6(32'hba8a53f8),
	.w7(32'hba9d60a8),
	.w8(32'h3afd4071),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81821),
	.w1(32'hbb3b0edd),
	.w2(32'h3af285f6),
	.w3(32'h3adcf1ee),
	.w4(32'hbab28a65),
	.w5(32'h3b65e00f),
	.w6(32'h3aa37048),
	.w7(32'h3b52475a),
	.w8(32'h3ac3612c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77f5d0),
	.w1(32'h3acf7d93),
	.w2(32'hba969c71),
	.w3(32'h3ac87367),
	.w4(32'hbac62590),
	.w5(32'h3ae2dc4a),
	.w6(32'hba43e051),
	.w7(32'hbb031205),
	.w8(32'h3b53b3d0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92f3bd),
	.w1(32'h3b7df4cd),
	.w2(32'h3b0f2390),
	.w3(32'h3a5c1b9f),
	.w4(32'hbafaf853),
	.w5(32'h3af1e931),
	.w6(32'h3be41fa7),
	.w7(32'h3b30fc5c),
	.w8(32'hb8e16a36),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812fdec),
	.w1(32'h3b2381fa),
	.w2(32'h3b7c11f4),
	.w3(32'h3b7a0f2e),
	.w4(32'h3b139f33),
	.w5(32'hbaac57d1),
	.w6(32'h3b0e80b9),
	.w7(32'h3a5c5596),
	.w8(32'hbae047b4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc8f86),
	.w1(32'hba91b420),
	.w2(32'hbb1d625e),
	.w3(32'hbb3305e7),
	.w4(32'hbafa7c9b),
	.w5(32'hbb128324),
	.w6(32'hbb2b1c26),
	.w7(32'hbad2ea14),
	.w8(32'hbac32446),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f705b),
	.w1(32'h38ef27da),
	.w2(32'h3bb14c3b),
	.w3(32'hbb70340c),
	.w4(32'h3a9f5a69),
	.w5(32'h3a00d0c3),
	.w6(32'hbae6b7c3),
	.w7(32'h3aee9648),
	.w8(32'hbade8dc4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae09508),
	.w1(32'hbb72f2d6),
	.w2(32'hbbb1b150),
	.w3(32'hbad6cb64),
	.w4(32'hbb6a9e07),
	.w5(32'h3b87e808),
	.w6(32'hbb66dcda),
	.w7(32'hbb896645),
	.w8(32'hbb44ce4f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7da1a6),
	.w1(32'h3a56bfed),
	.w2(32'h3b69fcce),
	.w3(32'h3b6af03d),
	.w4(32'h3baa202f),
	.w5(32'h3b58f9e3),
	.w6(32'hbbd60e6a),
	.w7(32'hb9f0f009),
	.w8(32'h3ab58fad),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d04a3),
	.w1(32'h38da60ce),
	.w2(32'hbacf1f4a),
	.w3(32'hba438833),
	.w4(32'hbb32b43e),
	.w5(32'h3c0109c4),
	.w6(32'hbb19e572),
	.w7(32'hbb77c958),
	.w8(32'h3c0afbcd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054b27),
	.w1(32'h3bead90f),
	.w2(32'h3adfa8cd),
	.w3(32'h3beefc9f),
	.w4(32'h3b032853),
	.w5(32'h3aa50c94),
	.w6(32'h3c1e7bc1),
	.w7(32'h3b6cf85e),
	.w8(32'h3986c013),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a540e7d),
	.w1(32'h3ac35c77),
	.w2(32'h3b624bb3),
	.w3(32'hba86b39b),
	.w4(32'hb93b61ed),
	.w5(32'h3a935e55),
	.w6(32'hbabbff51),
	.w7(32'h3b16a871),
	.w8(32'h3a3fc485),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5d41),
	.w1(32'h3ad4aa75),
	.w2(32'h3a91ed57),
	.w3(32'h3a8871af),
	.w4(32'hb945ad26),
	.w5(32'h3b2a8149),
	.w6(32'hb8fc4440),
	.w7(32'hba4ded87),
	.w8(32'h3a5abada),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b824),
	.w1(32'hba32fab2),
	.w2(32'hbb26a5c2),
	.w3(32'hb97528e6),
	.w4(32'hbb4ecc0b),
	.w5(32'h3aec889f),
	.w6(32'hbb09deda),
	.w7(32'hbb7f2fd7),
	.w8(32'h398e3575),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af37bd1),
	.w1(32'hbb16790c),
	.w2(32'hbb625a4b),
	.w3(32'hba5cf753),
	.w4(32'hbb151a98),
	.w5(32'hba6facc6),
	.w6(32'hbb36973d),
	.w7(32'hbb7f22ed),
	.w8(32'h3b8ae2d3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f47e),
	.w1(32'h3a543054),
	.w2(32'h3ae90326),
	.w3(32'h3ad3d1a6),
	.w4(32'h3ae69fb6),
	.w5(32'hb9010627),
	.w6(32'h3be3d4c9),
	.w7(32'h3b7c6793),
	.w8(32'hbaa47fdd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925a4e3),
	.w1(32'hbaf95740),
	.w2(32'h3ab8050a),
	.w3(32'hba862cab),
	.w4(32'h3a8fe70c),
	.w5(32'hbb622177),
	.w6(32'hbb728d4d),
	.w7(32'hba6ff456),
	.w8(32'hbb8312c5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2484b5),
	.w1(32'hbb446004),
	.w2(32'h3aa74487),
	.w3(32'hbb8f98b3),
	.w4(32'hbb2374c7),
	.w5(32'h3b6514e0),
	.w6(32'hbb9e0b0f),
	.w7(32'h38cc9153),
	.w8(32'h3ae236da),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cafee6),
	.w1(32'hbac03622),
	.w2(32'hbb2ee844),
	.w3(32'h3a5a9d13),
	.w4(32'hb8caf35e),
	.w5(32'h3b2c0cc7),
	.w6(32'hba18a58d),
	.w7(32'hbac17be7),
	.w8(32'h3af40a09),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194d57),
	.w1(32'h3ada73ba),
	.w2(32'h398fb4d6),
	.w3(32'h3a8ade3e),
	.w4(32'hbaa30685),
	.w5(32'h3b95e8a7),
	.w6(32'h39a53e7e),
	.w7(32'hbb5e9b63),
	.w8(32'h3b8a288a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be033),
	.w1(32'h3b4b28fe),
	.w2(32'h3a66111b),
	.w3(32'h3ad9f122),
	.w4(32'h3a991de7),
	.w5(32'h3945a064),
	.w6(32'h3ae0320d),
	.w7(32'h3a9e276a),
	.w8(32'hba85fc15),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba692004),
	.w1(32'hb7211de2),
	.w2(32'h3a380ed5),
	.w3(32'hb9a0d529),
	.w4(32'h39ae0dc7),
	.w5(32'hb8ceebbc),
	.w6(32'hba46259e),
	.w7(32'h3a2fa4ac),
	.w8(32'hb9e26422),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e73a3),
	.w1(32'h3aec2b90),
	.w2(32'hb9353191),
	.w3(32'h3a6113e2),
	.w4(32'h3a21179b),
	.w5(32'h3bc3b4e2),
	.w6(32'hb97da7d4),
	.w7(32'h38a77328),
	.w8(32'h3ade8b30),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee5bf8),
	.w1(32'hba6c6d05),
	.w2(32'h3bc8ddc7),
	.w3(32'h3b86f9c2),
	.w4(32'h3b9925fd),
	.w5(32'h3b910b10),
	.w6(32'h3b077879),
	.w7(32'h3c06cdca),
	.w8(32'h3b9d5896),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b955393),
	.w1(32'h3b039efb),
	.w2(32'hb9e4eb45),
	.w3(32'h3acd564f),
	.w4(32'hbad5815f),
	.w5(32'h3b986b40),
	.w6(32'h3b04c6a8),
	.w7(32'hbaa0cb71),
	.w8(32'h3bfa9387),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5a124),
	.w1(32'h3b8509c1),
	.w2(32'h3a2bf7ff),
	.w3(32'h3b6dd8d2),
	.w4(32'h39c10732),
	.w5(32'h3b18135d),
	.w6(32'h3bbddcee),
	.w7(32'h3a516de2),
	.w8(32'h3beb1dd4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b111883),
	.w1(32'h3b59a6cf),
	.w2(32'h3994018a),
	.w3(32'h3bebbb36),
	.w4(32'h3b3280b1),
	.w5(32'h3c06952f),
	.w6(32'h3c25d1a4),
	.w7(32'h3b4f7b7f),
	.w8(32'h3bb7c60e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cfbac),
	.w1(32'hb9d91e75),
	.w2(32'h3ae140d0),
	.w3(32'h3b01214e),
	.w4(32'hbb00c920),
	.w5(32'h388e2c3a),
	.w6(32'hbad14a2d),
	.w7(32'hbb2815f8),
	.w8(32'hbab53eca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abae0e6),
	.w1(32'hbad3d826),
	.w2(32'h3ae61bbc),
	.w3(32'hbb3094ab),
	.w4(32'h3a4ab905),
	.w5(32'h3bc77054),
	.w6(32'hbb93888b),
	.w7(32'hba1e7a76),
	.w8(32'h3b67e9ff),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856785),
	.w1(32'h3a053884),
	.w2(32'hbb354efa),
	.w3(32'h3b11c324),
	.w4(32'hb9d41694),
	.w5(32'h3bb7a5eb),
	.w6(32'h39a0d80a),
	.w7(32'hbac7e24a),
	.w8(32'h3b8b60e1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85c0d4),
	.w1(32'h3b2ea30c),
	.w2(32'h3af60b4f),
	.w3(32'h3b8c7eca),
	.w4(32'h3b7d92bb),
	.w5(32'hbb115931),
	.w6(32'h3b22e253),
	.w7(32'h3b18ae23),
	.w8(32'hbb867c24),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdb8fb),
	.w1(32'h3aef0b29),
	.w2(32'h3b8c6723),
	.w3(32'hba8d3e8c),
	.w4(32'h3ab2f45c),
	.w5(32'hbad58d4d),
	.w6(32'hbb5416b2),
	.w7(32'h3a149279),
	.w8(32'hbb890a76),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89e37),
	.w1(32'hbba8b4a7),
	.w2(32'hb6b9644d),
	.w3(32'hbb0a2c61),
	.w4(32'hbb078a87),
	.w5(32'hbb3efaba),
	.w6(32'hbb32ee79),
	.w7(32'h3af7cca2),
	.w8(32'hbb23eb78),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987e9d),
	.w1(32'hbb00dd5c),
	.w2(32'h3af5a3ce),
	.w3(32'hba5a88a6),
	.w4(32'h3b10cac6),
	.w5(32'hb93802b2),
	.w6(32'hbb00f65c),
	.w7(32'h3b3383fc),
	.w8(32'hba7c60db),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391eecc3),
	.w1(32'h3a8d8fae),
	.w2(32'h3a9a252c),
	.w3(32'h3b354237),
	.w4(32'h3b93a608),
	.w5(32'hb782c133),
	.w6(32'h3b2a0f55),
	.w7(32'h3bab6455),
	.w8(32'h3bb60508),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c8ca5),
	.w1(32'h3b300b1f),
	.w2(32'h3b877f08),
	.w3(32'h3a4e8d37),
	.w4(32'hba2aa46e),
	.w5(32'h3b83f4d1),
	.w6(32'h3be3a6bb),
	.w7(32'h3ba25799),
	.w8(32'h3b8396cd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a566),
	.w1(32'h3c162e33),
	.w2(32'h3a9a0169),
	.w3(32'h3b71616b),
	.w4(32'h3c13c131),
	.w5(32'hb998d195),
	.w6(32'h3beef44d),
	.w7(32'h3c0f20e1),
	.w8(32'hba9f08c6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad092d5),
	.w1(32'hba93e076),
	.w2(32'h39ba33c5),
	.w3(32'hba95be04),
	.w4(32'h3a28d092),
	.w5(32'h3b7f032f),
	.w6(32'hbb0452d9),
	.w7(32'h398144be),
	.w8(32'h3bc405cb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baefcc3),
	.w1(32'h3bbf360c),
	.w2(32'h3ac6e7b0),
	.w3(32'hbab92c35),
	.w4(32'hbbe70223),
	.w5(32'h3aed07d1),
	.w6(32'h3ab6f8ca),
	.w7(32'hbb855b31),
	.w8(32'h3a889699),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0c39b),
	.w1(32'h3a1343e7),
	.w2(32'h3a4b9ce5),
	.w3(32'hb95fa290),
	.w4(32'hba0ffd07),
	.w5(32'h3adb48f7),
	.w6(32'hba81e194),
	.w7(32'h37c4ff8a),
	.w8(32'h3b7a2ee1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e453a8),
	.w1(32'h3b3e7d29),
	.w2(32'h3b346365),
	.w3(32'h3b1bf5cb),
	.w4(32'h3be2390d),
	.w5(32'h3bdfd68a),
	.w6(32'h3bbcd4c7),
	.w7(32'h3bd8ccf5),
	.w8(32'h3b55b81f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4be58),
	.w1(32'h3b2106b0),
	.w2(32'hba5dcfab),
	.w3(32'h3b5c3d4b),
	.w4(32'h3a3fab5e),
	.w5(32'h3ab8baf3),
	.w6(32'h397a7e7c),
	.w7(32'hbb1795d6),
	.w8(32'hbb466da9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89edf6),
	.w1(32'hbb66f838),
	.w2(32'hbaaf57a9),
	.w3(32'h3b2a9685),
	.w4(32'h3b6b46ed),
	.w5(32'h3b413edf),
	.w6(32'hbb48fcd8),
	.w7(32'hba4cc2a8),
	.w8(32'h3b69e5fb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866212),
	.w1(32'h3b4cdec9),
	.w2(32'h39f30a1e),
	.w3(32'h3b4e1ec8),
	.w4(32'h3a78c2ea),
	.w5(32'hbad3e374),
	.w6(32'h3b7c1aa1),
	.w7(32'hb9950ed7),
	.w8(32'hba8a1505),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62d2f7),
	.w1(32'hbaa74de3),
	.w2(32'hbb00b309),
	.w3(32'h3af70130),
	.w4(32'hbb208c58),
	.w5(32'h3bb46220),
	.w6(32'h39b99848),
	.w7(32'hbb2f0923),
	.w8(32'h3b581b22),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f60bc),
	.w1(32'h39dcc743),
	.w2(32'hbb006bd5),
	.w3(32'h3a4ee624),
	.w4(32'hba43b594),
	.w5(32'h38f62441),
	.w6(32'h38e84442),
	.w7(32'hba9794df),
	.w8(32'hbb4d6a0a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9236a7),
	.w1(32'h3a3e73eb),
	.w2(32'h3ab5febf),
	.w3(32'h3aa592bd),
	.w4(32'hba6635b6),
	.w5(32'hb9c6e416),
	.w6(32'hbb325c4b),
	.w7(32'hba867ade),
	.w8(32'hbb219811),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b23a1),
	.w1(32'hb9c19f6f),
	.w2(32'h3a31a175),
	.w3(32'hba10918a),
	.w4(32'h3a56b96c),
	.w5(32'h3a71f3a5),
	.w6(32'hbb518ea0),
	.w7(32'h3947086e),
	.w8(32'hb8ebe8cd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7442f),
	.w1(32'hbad2a59e),
	.w2(32'hbb17a94f),
	.w3(32'h39e1e3b3),
	.w4(32'hb9ddaa5f),
	.w5(32'hb9ca919b),
	.w6(32'h3a8c89ed),
	.w7(32'hba210c93),
	.w8(32'hbab4478d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba165b06),
	.w1(32'h394a3dfa),
	.w2(32'h3b1d0c0b),
	.w3(32'h3a3e3492),
	.w4(32'h3afd3bc7),
	.w5(32'hba1b2cbe),
	.w6(32'h3908140e),
	.w7(32'h3b14ed96),
	.w8(32'hbb0862de),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3f0eb),
	.w1(32'hbb195ef3),
	.w2(32'hba42ed5e),
	.w3(32'hb8725e61),
	.w4(32'hb99e09f7),
	.w5(32'h3a8148e3),
	.w6(32'hba9750b8),
	.w7(32'hb9a39198),
	.w8(32'h3b0e3611),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d6416),
	.w1(32'h3a95650b),
	.w2(32'hba2ac6ec),
	.w3(32'hb9f14dcd),
	.w4(32'hbabc0b39),
	.w5(32'h3ad255c2),
	.w6(32'h39a05b62),
	.w7(32'hbaeae7b0),
	.w8(32'hba3dd1ba),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899dada),
	.w1(32'h3921f2c1),
	.w2(32'h3b29d59c),
	.w3(32'h3aa50b5b),
	.w4(32'h3ace70da),
	.w5(32'h3b92a4e8),
	.w6(32'hbaccb888),
	.w7(32'hb9ac9466),
	.w8(32'h3bda6a65),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7b812),
	.w1(32'h3b9e63e2),
	.w2(32'h3a3337b2),
	.w3(32'h3b510b03),
	.w4(32'h3a9b6a72),
	.w5(32'h3b329310),
	.w6(32'h3bb12e4b),
	.w7(32'h3b002703),
	.w8(32'h3982ec56),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaa0ee),
	.w1(32'h3c10af83),
	.w2(32'h3c63e71c),
	.w3(32'h3b6aecc1),
	.w4(32'h3c2ca821),
	.w5(32'h3b3048fe),
	.w6(32'h3b73df4b),
	.w7(32'h3c414a76),
	.w8(32'h3a1ff060),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bda8df),
	.w1(32'h3a0a1f35),
	.w2(32'hb9af0bcd),
	.w3(32'h3b022fb8),
	.w4(32'hba7c9d74),
	.w5(32'hbbd2e26a),
	.w6(32'h388cf32f),
	.w7(32'h3a5cc442),
	.w8(32'hbbf3cf0c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36071d),
	.w1(32'hbb945d8c),
	.w2(32'h3aba9ef8),
	.w3(32'hbbf4ff53),
	.w4(32'hbb8237d7),
	.w5(32'h39e4936c),
	.w6(32'hbc03f59a),
	.w7(32'hbb426d7e),
	.w8(32'hb9f163c5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410a0d),
	.w1(32'h3b096a22),
	.w2(32'h3abc8796),
	.w3(32'h3b6bfd99),
	.w4(32'h3ad9c601),
	.w5(32'h3b443ac9),
	.w6(32'h3b8b3ff3),
	.w7(32'h3a906b05),
	.w8(32'h3a9f502f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ee65a),
	.w1(32'hbaf7e72f),
	.w2(32'hba497df5),
	.w3(32'hbaa455ea),
	.w4(32'hbb714ad9),
	.w5(32'h3ab57995),
	.w6(32'hbad4bd1d),
	.w7(32'hba9ca4ed),
	.w8(32'hbb05bcb6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93dc03),
	.w1(32'hbb17b233),
	.w2(32'hbb2eb5d6),
	.w3(32'hbb07ba45),
	.w4(32'hbb954ea8),
	.w5(32'h3ba8920f),
	.w6(32'hbbc246ae),
	.w7(32'hbbedf9ef),
	.w8(32'h3bad66d5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc049ac),
	.w1(32'h3b68eb0c),
	.w2(32'h39943229),
	.w3(32'h3b550d20),
	.w4(32'hbad6626f),
	.w5(32'hba976563),
	.w6(32'h3b0e49ee),
	.w7(32'hbb5ff0f1),
	.w8(32'hbb350731),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03eaea),
	.w1(32'hbb9a8d57),
	.w2(32'h38a37e53),
	.w3(32'hbb7e7f46),
	.w4(32'h391340b3),
	.w5(32'h3bb71c11),
	.w6(32'hbbc06b77),
	.w7(32'hb9a5b88f),
	.w8(32'h3c0021ba),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6e4b4),
	.w1(32'h3bb41710),
	.w2(32'h39643e28),
	.w3(32'h3b990bfe),
	.w4(32'h3a4ab18c),
	.w5(32'h3be73c51),
	.w6(32'h3bcb642e),
	.w7(32'h3acf9e14),
	.w8(32'h3bc38e3c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2987),
	.w1(32'h3b7a4ddd),
	.w2(32'h3b97ab09),
	.w3(32'h3b91d05a),
	.w4(32'h3b47a812),
	.w5(32'h3b4bb734),
	.w6(32'h3b5a37b5),
	.w7(32'h3b2b54c4),
	.w8(32'hbabc7382),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3756ed),
	.w1(32'hbb2285f1),
	.w2(32'h3a05c0f0),
	.w3(32'h3b5867e4),
	.w4(32'h3b96542b),
	.w5(32'h3b869cfd),
	.w6(32'hbad7d9ff),
	.w7(32'h38af72a1),
	.w8(32'h3b227d2c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5de11f),
	.w1(32'h3a3e963f),
	.w2(32'h3a92e6fe),
	.w3(32'h3b3efbae),
	.w4(32'h3b12efaa),
	.w5(32'h39980ed3),
	.w6(32'h39c38a3d),
	.w7(32'h3b364ab8),
	.w8(32'hbb444541),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a79b8),
	.w1(32'h3ba3833b),
	.w2(32'h3bdc61ca),
	.w3(32'hb9a2a793),
	.w4(32'h3a9327d6),
	.w5(32'h3866f330),
	.w6(32'hbb98ae48),
	.w7(32'hbac6d0ca),
	.w8(32'hbb298afd),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17ef67),
	.w1(32'hba55815e),
	.w2(32'hbad6ec23),
	.w3(32'h3aa567c2),
	.w4(32'hbaea7df7),
	.w5(32'hbab7bc0d),
	.w6(32'hbaf19f8c),
	.w7(32'hbb1b4d91),
	.w8(32'hbb1ef76f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f6bb),
	.w1(32'hbb608e4e),
	.w2(32'hbbcae5ad),
	.w3(32'hbb96bef4),
	.w4(32'hbc1776f3),
	.w5(32'hbac69f5b),
	.w6(32'hbbddde5c),
	.w7(32'hbc08a255),
	.w8(32'hbb626c33),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb484267),
	.w1(32'hbb7686ed),
	.w2(32'hbb02fdcc),
	.w3(32'hbb2a3263),
	.w4(32'hbb4c0808),
	.w5(32'h3a8e715d),
	.w6(32'hbb9c9702),
	.w7(32'hbacaeaae),
	.w8(32'hba98aeca),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd7546),
	.w1(32'h3a871a3f),
	.w2(32'h3b8848d4),
	.w3(32'hb9d43cdf),
	.w4(32'h3ae0ae2d),
	.w5(32'hb98c003e),
	.w6(32'hbac0264b),
	.w7(32'h3a9acbdf),
	.w8(32'hba706f96),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2371ec),
	.w1(32'hbb0df098),
	.w2(32'hbb15caf3),
	.w3(32'hbb425bdb),
	.w4(32'hba52034f),
	.w5(32'h3b22c7b4),
	.w6(32'hbb8130e9),
	.w7(32'hbb15701c),
	.w8(32'h3b06f7ef),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb632),
	.w1(32'h3b364ced),
	.w2(32'h3ab7426b),
	.w3(32'h3a9c7c70),
	.w4(32'hba2c158c),
	.w5(32'h39d510c7),
	.w6(32'h3af13d6e),
	.w7(32'h3a1d2af6),
	.w8(32'h3a42217f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1c19f),
	.w1(32'h3b09f29d),
	.w2(32'hba87cf4a),
	.w3(32'h3ab7fab7),
	.w4(32'hb94665be),
	.w5(32'hbb174e61),
	.w6(32'h3ac8872e),
	.w7(32'hba04698c),
	.w8(32'hbacbb784),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7b8e4),
	.w1(32'hbaec6aa0),
	.w2(32'hbb219e0b),
	.w3(32'hbb09220d),
	.w4(32'hbb2ac92d),
	.w5(32'h39ba0721),
	.w6(32'hba8b7e68),
	.w7(32'hbb0906dc),
	.w8(32'hbb023480),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d623b),
	.w1(32'hbb487f04),
	.w2(32'hba7278a8),
	.w3(32'h3aa3125e),
	.w4(32'hb8a373d5),
	.w5(32'h3b8cc064),
	.w6(32'hb9e7e700),
	.w7(32'hbaf2f8ae),
	.w8(32'h39b34ed6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2651),
	.w1(32'hbaf5b2ed),
	.w2(32'hb9f989e9),
	.w3(32'h3b6cd463),
	.w4(32'h3b4f55db),
	.w5(32'h3ace9b16),
	.w6(32'hb9dd2a58),
	.w7(32'h3a2b8cb7),
	.w8(32'h3a8dd10b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a8372),
	.w1(32'h3b37859d),
	.w2(32'h3b389eb3),
	.w3(32'h3aec4e31),
	.w4(32'h3b2bb00f),
	.w5(32'h3b3e1d53),
	.w6(32'h3add16de),
	.w7(32'h3b4bf002),
	.w8(32'h3a7c56c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af510e1),
	.w1(32'hb9eb1cb3),
	.w2(32'hba3290ef),
	.w3(32'h3ae84231),
	.w4(32'hb9c969a3),
	.w5(32'hba998949),
	.w6(32'hb962160b),
	.w7(32'hbb3bb00b),
	.w8(32'hbb2f5086),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e45c3),
	.w1(32'hba57c577),
	.w2(32'h3b31f2b1),
	.w3(32'hb93bf164),
	.w4(32'h3ab82bcb),
	.w5(32'h3a03cc8d),
	.w6(32'hbb211817),
	.w7(32'h3ab01f64),
	.w8(32'h3b746545),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe524c),
	.w1(32'hbb603007),
	.w2(32'hbba11341),
	.w3(32'h3b76c2e0),
	.w4(32'hbaa1185d),
	.w5(32'hba71d6be),
	.w6(32'h3a8d57cf),
	.w7(32'hbb5c8159),
	.w8(32'hbb07261c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119cee),
	.w1(32'hbb191a26),
	.w2(32'hbb084212),
	.w3(32'hb99a895e),
	.w4(32'hbab32cf5),
	.w5(32'hbb0bd153),
	.w6(32'hbacd4aa5),
	.w7(32'hba5efd0e),
	.w8(32'hbb3da9ff),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d35b8),
	.w1(32'hbab80ba5),
	.w2(32'h39ee649a),
	.w3(32'hbac515cd),
	.w4(32'hb9871617),
	.w5(32'h3b993a32),
	.w6(32'hbad692ff),
	.w7(32'h3954045f),
	.w8(32'h3b69cc79),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ad5d),
	.w1(32'h3ba98b55),
	.w2(32'h3ba0b360),
	.w3(32'h3b7cb3ff),
	.w4(32'h3b8d24d3),
	.w5(32'hba97fef2),
	.w6(32'h3b55d3ed),
	.w7(32'h3b0f2c12),
	.w8(32'hba81fc9f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb000368),
	.w1(32'hba9e488c),
	.w2(32'h3a91e9f5),
	.w3(32'h3a06798c),
	.w4(32'h380a418b),
	.w5(32'h3abf187f),
	.w6(32'h3ac025cd),
	.w7(32'h3aaab1c2),
	.w8(32'h3a0cc02e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d15f0),
	.w1(32'h3ac17c6d),
	.w2(32'h3afb9f56),
	.w3(32'h3a24387f),
	.w4(32'h3ab58637),
	.w5(32'hbba8570c),
	.w6(32'h38fe456b),
	.w7(32'h3a6435f9),
	.w8(32'hbab9e60a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56a534),
	.w1(32'hbb93c190),
	.w2(32'hbbd9c76a),
	.w3(32'hba844c18),
	.w4(32'hbbb86654),
	.w5(32'h3ab71dc5),
	.w6(32'hbb41343f),
	.w7(32'hbbb16ae5),
	.w8(32'hb883069d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cb7e5),
	.w1(32'hba207ec6),
	.w2(32'hba5e5d36),
	.w3(32'h3aa429ca),
	.w4(32'h3b0c92a0),
	.w5(32'hbbc97c3b),
	.w6(32'h39bd4e77),
	.w7(32'h3a3b137e),
	.w8(32'hb9966d20),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2917b9),
	.w1(32'hbad41d7d),
	.w2(32'hbb362b49),
	.w3(32'hbb183b8e),
	.w4(32'hbb842f91),
	.w5(32'h3bb2e185),
	.w6(32'h3a8bad86),
	.w7(32'hbab9e8fe),
	.w8(32'h3b419cd1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac3b08),
	.w1(32'h3b131825),
	.w2(32'h3ba6d6ba),
	.w3(32'h3bb6fec1),
	.w4(32'h3b4acc65),
	.w5(32'h3baee331),
	.w6(32'h39e6bb7a),
	.w7(32'h3b08fb84),
	.w8(32'h3b2eadf2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96ab2d),
	.w1(32'hba824f5c),
	.w2(32'hb90374e7),
	.w3(32'h39ec1a4a),
	.w4(32'h3a6af686),
	.w5(32'h3be7203e),
	.w6(32'h3ad028af),
	.w7(32'h3af34355),
	.w8(32'hb97a79bb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1213),
	.w1(32'hbb9a6fcf),
	.w2(32'hbaece186),
	.w3(32'h3ba5871f),
	.w4(32'h3b96b7cc),
	.w5(32'h3bea05ac),
	.w6(32'hbb255d15),
	.w7(32'h3af48011),
	.w8(32'h3be4b81f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe07dc),
	.w1(32'h3be73b67),
	.w2(32'h3b8acef1),
	.w3(32'h3bc4883c),
	.w4(32'h3b8fb62b),
	.w5(32'hba1cda10),
	.w6(32'h3bd66fdd),
	.w7(32'h3b933a50),
	.w8(32'h3af53928),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b80b),
	.w1(32'h3b8d2fa1),
	.w2(32'h3b96ac9b),
	.w3(32'h3b0e1131),
	.w4(32'h3b8c6901),
	.w5(32'hbae1bb97),
	.w6(32'h3bac428b),
	.w7(32'h3bdc9ebb),
	.w8(32'h3a08f4d5),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a271188),
	.w1(32'h3a4573fd),
	.w2(32'h3ab97d54),
	.w3(32'hbaef7e8c),
	.w4(32'h3a2b9a66),
	.w5(32'h3a66e397),
	.w6(32'hb9af2c83),
	.w7(32'hbababce0),
	.w8(32'h39417cbe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af33d8c),
	.w1(32'h3b750352),
	.w2(32'h3b532730),
	.w3(32'h3b3b1b43),
	.w4(32'h3b6963a9),
	.w5(32'h3bc49441),
	.w6(32'h3b8da248),
	.w7(32'h3bc9a28c),
	.w8(32'h3bea6c99),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be45170),
	.w1(32'h3ba7e00a),
	.w2(32'h3bd2dc21),
	.w3(32'h3bc19532),
	.w4(32'h3b4cba09),
	.w5(32'hbad79f95),
	.w6(32'h3c0c6f08),
	.w7(32'h3bccc62b),
	.w8(32'hbb729222),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a446148),
	.w1(32'hbb58091f),
	.w2(32'hba2f8640),
	.w3(32'hbb7fac1c),
	.w4(32'hbb55c6d4),
	.w5(32'h3b3f0862),
	.w6(32'hbbc75027),
	.w7(32'hbb8bb0d4),
	.w8(32'h3b2cfa0d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bc2eb),
	.w1(32'h3b6e4775),
	.w2(32'h3b1403f0),
	.w3(32'h3b45cdbd),
	.w4(32'h3b5c8975),
	.w5(32'h3bab0dc9),
	.w6(32'h3b815450),
	.w7(32'h3b2a48b1),
	.w8(32'h3b7dcefb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b93a5),
	.w1(32'h3af9c717),
	.w2(32'h3b2f2685),
	.w3(32'h3bb5d5dc),
	.w4(32'h3b538420),
	.w5(32'hbb2e6a56),
	.w6(32'h3b3a1898),
	.w7(32'h3a8f00e4),
	.w8(32'hbb06bed3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1223a8),
	.w1(32'h391677c8),
	.w2(32'h39afc9ac),
	.w3(32'hba9192f1),
	.w4(32'h3a1f384b),
	.w5(32'h3c14196b),
	.w6(32'h3aa8eafc),
	.w7(32'h3a9544b2),
	.w8(32'h3c2219ba),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a964c),
	.w1(32'h3bc150c5),
	.w2(32'h3a756cdc),
	.w3(32'h3bede987),
	.w4(32'h3a270a7a),
	.w5(32'hb9a75785),
	.w6(32'h3b99653a),
	.w7(32'hba8ef6ce),
	.w8(32'hb91b3870),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b21288),
	.w1(32'hba13751e),
	.w2(32'hb9a5f4e8),
	.w3(32'hba158960),
	.w4(32'hba093602),
	.w5(32'hba0bf397),
	.w6(32'h38cd9061),
	.w7(32'h38031f6f),
	.w8(32'hba15f289),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1ba2c),
	.w1(32'hb867d40c),
	.w2(32'h39012e15),
	.w3(32'h3a2480c2),
	.w4(32'hb9c3381c),
	.w5(32'hb95aa8db),
	.w6(32'h3a8f1a83),
	.w7(32'hb98fbcad),
	.w8(32'hb9b48004),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979efa2),
	.w1(32'hba51b856),
	.w2(32'hb9b70f6d),
	.w3(32'hb725b05b),
	.w4(32'hba07ab4d),
	.w5(32'h39a1f524),
	.w6(32'hb9d51dcc),
	.w7(32'hba317c91),
	.w8(32'h399c4299),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cec68),
	.w1(32'hb9580d4b),
	.w2(32'hb9976cc7),
	.w3(32'h39e9bd94),
	.w4(32'h3a434219),
	.w5(32'hb9c6882f),
	.w6(32'h3a11904f),
	.w7(32'h38df00d9),
	.w8(32'hb8b3855f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f32f6),
	.w1(32'h39ea83e3),
	.w2(32'h3a544e52),
	.w3(32'h3a0b9711),
	.w4(32'h39ad6440),
	.w5(32'hbb06f791),
	.w6(32'h3ad7bdcf),
	.w7(32'h3a9f94a5),
	.w8(32'hba899695),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf51d5),
	.w1(32'hbacc1a58),
	.w2(32'hbb032600),
	.w3(32'hbac4c079),
	.w4(32'hbb20fcd7),
	.w5(32'h39814a7c),
	.w6(32'hb9881dc8),
	.w7(32'hbac40251),
	.w8(32'hba1df8a3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fe263),
	.w1(32'hba32cf4d),
	.w2(32'hb92a7d9d),
	.w3(32'hb75000f8),
	.w4(32'h38d2974b),
	.w5(32'hb8a6d775),
	.w6(32'hba2dd2ad),
	.w7(32'hba45a72e),
	.w8(32'hba50774f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959accc),
	.w1(32'hb9d5e6a8),
	.w2(32'hb9d83562),
	.w3(32'hb987dad4),
	.w4(32'hba5ac084),
	.w5(32'hb873c63f),
	.w6(32'hb94da610),
	.w7(32'hb9ce53a2),
	.w8(32'hb9ffe969),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5ee50),
	.w1(32'h39826eeb),
	.w2(32'h3a457bab),
	.w3(32'hb87e1992),
	.w4(32'h39c94875),
	.w5(32'hb8f65d0c),
	.w6(32'hb952b491),
	.w7(32'h3a6d0e4d),
	.w8(32'hb8e9e037),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e8ed7),
	.w1(32'hb9f967da),
	.w2(32'hb943c58a),
	.w3(32'hb98f52e7),
	.w4(32'hb8febf7c),
	.w5(32'hb95f48c4),
	.w6(32'hb938b5d3),
	.w7(32'hb9c7e4df),
	.w8(32'hb76d4d6e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930e526),
	.w1(32'hb94934a6),
	.w2(32'hb821bedb),
	.w3(32'hb9dbb341),
	.w4(32'hb995f2ea),
	.w5(32'hba1cddc3),
	.w6(32'hb7f871fa),
	.w7(32'h38db708a),
	.w8(32'hba2cb5fa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38399722),
	.w1(32'h37995922),
	.w2(32'h393e4c95),
	.w3(32'hb9ca964f),
	.w4(32'hb91bc23c),
	.w5(32'h39d41cc0),
	.w6(32'hba14e006),
	.w7(32'hb986816d),
	.w8(32'h39578c59),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8151bf),
	.w1(32'h3a8c5b86),
	.w2(32'h39cb5e90),
	.w3(32'h3a26bfce),
	.w4(32'h39e7270b),
	.w5(32'hb99f45e2),
	.w6(32'h3a557a21),
	.w7(32'h3a33107f),
	.w8(32'h3890b2e8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a580553),
	.w1(32'h3a85a37f),
	.w2(32'h3a302195),
	.w3(32'h3a21d5bb),
	.w4(32'hb9195133),
	.w5(32'h3a0f245f),
	.w6(32'h3a6cc35d),
	.w7(32'hb947b4d4),
	.w8(32'h3967f5a8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad2051),
	.w1(32'h3a7e3928),
	.w2(32'h39f5476b),
	.w3(32'h3a3366e9),
	.w4(32'hb94cff7f),
	.w5(32'h39d75cf9),
	.w6(32'h36dc7629),
	.w7(32'hba309070),
	.w8(32'hb8d82103),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ec9cc),
	.w1(32'h39e43fb3),
	.w2(32'h3a03da5f),
	.w3(32'h3929f632),
	.w4(32'hb9891777),
	.w5(32'h39c5751e),
	.w6(32'h3a4b7033),
	.w7(32'h39903467),
	.w8(32'h3a3cd8a9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57a2a4),
	.w1(32'h3a5437eb),
	.w2(32'h39934e07),
	.w3(32'h399f01e5),
	.w4(32'h39f6fd04),
	.w5(32'h38d23b9b),
	.w6(32'hb9a7f343),
	.w7(32'hb985fdfb),
	.w8(32'h39c9b4b7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22fdde),
	.w1(32'h3a1d3ef5),
	.w2(32'h39393dd4),
	.w3(32'h39f31524),
	.w4(32'h3a10fef1),
	.w5(32'h3a76e77b),
	.w6(32'h3a23424d),
	.w7(32'h39e181c4),
	.w8(32'h3a570c5d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1460f0),
	.w1(32'h3979820c),
	.w2(32'h398b186e),
	.w3(32'h3a2c6b80),
	.w4(32'h3a07c1ef),
	.w5(32'h39bb6dce),
	.w6(32'h39ee1a9a),
	.w7(32'h39c05e40),
	.w8(32'hb8112e4c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f8697),
	.w1(32'hb91b6132),
	.w2(32'h3a061e89),
	.w3(32'h39a34bdd),
	.w4(32'hb8491985),
	.w5(32'hba08328e),
	.w6(32'h3a0e21e2),
	.w7(32'hb93e364e),
	.w8(32'hba7f476a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d417ae),
	.w1(32'h3915e062),
	.w2(32'h3a6c38e9),
	.w3(32'h39ba0eda),
	.w4(32'h39f2ea07),
	.w5(32'hbb16b77b),
	.w6(32'h3921134e),
	.w7(32'hb8b0c14b),
	.w8(32'hbb1de88e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd9bc),
	.w1(32'hbb749752),
	.w2(32'hbb3cb2d9),
	.w3(32'hbb300300),
	.w4(32'hbb1b7775),
	.w5(32'h3a130560),
	.w6(32'hbb56e180),
	.w7(32'hbb0c9f62),
	.w8(32'h3a1fb82e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cddd2),
	.w1(32'h3a974ec5),
	.w2(32'h3a481411),
	.w3(32'h39d607b1),
	.w4(32'h3a4ec2d3),
	.w5(32'h37aaf4c0),
	.w6(32'h3a0bb4a7),
	.w7(32'h3a64d84c),
	.w8(32'h38e79ecf),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39829320),
	.w1(32'h3a233e81),
	.w2(32'h3a29dc37),
	.w3(32'h39b4275b),
	.w4(32'h3a32ff30),
	.w5(32'hba3595a8),
	.w6(32'hb87c2ad2),
	.w7(32'h3a2ccc9b),
	.w8(32'hb93f2924),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb7876),
	.w1(32'h39b944a1),
	.w2(32'h3a0566fa),
	.w3(32'hba34c367),
	.w4(32'hba2c7f1a),
	.w5(32'h34e9b690),
	.w6(32'h38962ffe),
	.w7(32'hb8815bf0),
	.w8(32'hb89ab385),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39521ecb),
	.w1(32'h3932be62),
	.w2(32'h3a34bc8e),
	.w3(32'h398b73e4),
	.w4(32'h3a2747eb),
	.w5(32'hb9145ec4),
	.w6(32'h39797327),
	.w7(32'h3a257ddb),
	.w8(32'h393df422),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b4ce6),
	.w1(32'h3a591a33),
	.w2(32'h398d3448),
	.w3(32'hb9235e18),
	.w4(32'hb838dba2),
	.w5(32'h3a3e681c),
	.w6(32'h39260361),
	.w7(32'h38af26b3),
	.w8(32'h3a283653),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6abaa),
	.w1(32'h3a3ed6ea),
	.w2(32'h3a2e2f52),
	.w3(32'h3a87fa6f),
	.w4(32'h396639cb),
	.w5(32'h38e8fa71),
	.w6(32'h3ab4ac51),
	.w7(32'h3a8198f9),
	.w8(32'h390ac5ee),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa05d6),
	.w1(32'hb9f98c8c),
	.w2(32'hb947edb9),
	.w3(32'hb87d20f0),
	.w4(32'hb9348c06),
	.w5(32'h3a07a857),
	.w6(32'h3796f709),
	.w7(32'hb9327e8d),
	.w8(32'h3a5a8c2e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca0d6c),
	.w1(32'h3a9834c5),
	.w2(32'h3a3d92a4),
	.w3(32'h3ad59295),
	.w4(32'h3a0f3ea6),
	.w5(32'hba28214c),
	.w6(32'h3a22ceeb),
	.w7(32'h38ac1ee8),
	.w8(32'hba4080da),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule