module layer_10_featuremap_388(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc330cba),
	.w1(32'hbb87087a),
	.w2(32'hbb45d171),
	.w3(32'hbc6e1819),
	.w4(32'hbb86fd54),
	.w5(32'hbb0aab22),
	.w6(32'hbb978159),
	.w7(32'hbae7556e),
	.w8(32'hbb2fa6f6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891499),
	.w1(32'h3c2fd423),
	.w2(32'h3c14dfd7),
	.w3(32'hbb19646a),
	.w4(32'h3c416a39),
	.w5(32'h3c88ba96),
	.w6(32'hbac00513),
	.w7(32'h3c556a3d),
	.w8(32'h3c4f4ef0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004ec5),
	.w1(32'hbc93df33),
	.w2(32'hbc6f6225),
	.w3(32'h3c1879b9),
	.w4(32'hbc258b21),
	.w5(32'h3a036d80),
	.w6(32'h3bc747d7),
	.w7(32'hbcc68a5d),
	.w8(32'hbbe5fc23),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd7f1a),
	.w1(32'hbbe73745),
	.w2(32'hbae0b2b5),
	.w3(32'h3c472ba2),
	.w4(32'hbc151997),
	.w5(32'hb955df58),
	.w6(32'h3c0987c8),
	.w7(32'hbc5d1b22),
	.w8(32'hbbf1d28c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338f36),
	.w1(32'hba9dfc34),
	.w2(32'hbb31fb06),
	.w3(32'h3b36a1cc),
	.w4(32'hbbb0cb9c),
	.w5(32'hbb85e1dc),
	.w6(32'hbb7e64b9),
	.w7(32'hba52c82b),
	.w8(32'hbb036523),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926fea),
	.w1(32'h39ed30c4),
	.w2(32'hbbb06975),
	.w3(32'h3b2b9be7),
	.w4(32'hbb00739d),
	.w5(32'hbb4ebacf),
	.w6(32'h3ae5c662),
	.w7(32'h39f5027b),
	.w8(32'hbac38e29),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883fe8),
	.w1(32'h3b260077),
	.w2(32'h39e9e540),
	.w3(32'hbbf9f583),
	.w4(32'h3aeddd7e),
	.w5(32'hbb8359e3),
	.w6(32'hbbe4b778),
	.w7(32'hbb6512ae),
	.w8(32'hbb5b7f96),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd339bd),
	.w1(32'h3c0246dd),
	.w2(32'h3c027b77),
	.w3(32'hbbc2740f),
	.w4(32'h3c53abab),
	.w5(32'h3c1b7d0f),
	.w6(32'hbbc4ca6a),
	.w7(32'h3c05d7bb),
	.w8(32'h3bba5076),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd57c),
	.w1(32'hbd0855a0),
	.w2(32'h3b9b62de),
	.w3(32'h3bee1b8c),
	.w4(32'hbd057c44),
	.w5(32'h3bf9cb35),
	.w6(32'h3a333250),
	.w7(32'hbd02b95d),
	.w8(32'h3c1af93a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359703),
	.w1(32'h3bcce301),
	.w2(32'h3aa55ef7),
	.w3(32'hbc39c909),
	.w4(32'h3ba270f4),
	.w5(32'h3a8e9a16),
	.w6(32'hbc8b9212),
	.w7(32'h3ba0aa8e),
	.w8(32'hbb8d6932),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048317),
	.w1(32'h3b1ee846),
	.w2(32'h3c07edb0),
	.w3(32'hbb86bb4c),
	.w4(32'h3b9ee470),
	.w5(32'h3b530061),
	.w6(32'hbbb66bf2),
	.w7(32'h3b27bfce),
	.w8(32'h391e2c1b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f18eac),
	.w1(32'hba832ffb),
	.w2(32'hba948f1b),
	.w3(32'hbb3ac7e5),
	.w4(32'hbbb5d1fc),
	.w5(32'hbbc01521),
	.w6(32'hbb92e2a9),
	.w7(32'hbb0e9ccc),
	.w8(32'hba72ce2e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9faa7ac),
	.w1(32'h3b078088),
	.w2(32'h39ff9ce3),
	.w3(32'hbb68aba1),
	.w4(32'h3b2ed23f),
	.w5(32'h3c1e6cda),
	.w6(32'hba367ec5),
	.w7(32'hbb3a83ea),
	.w8(32'h3b9f137e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6624b0),
	.w1(32'hbc4151df),
	.w2(32'hbc36c360),
	.w3(32'h3b783835),
	.w4(32'hbc5bafd0),
	.w5(32'hbc5da4e2),
	.w6(32'h3a5597f4),
	.w7(32'hbc260bd9),
	.w8(32'hbc393086),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ea9de),
	.w1(32'hba77eaca),
	.w2(32'hbbc67a21),
	.w3(32'hbc04ee05),
	.w4(32'hbb149298),
	.w5(32'hbbe07b22),
	.w6(32'hbc121fb1),
	.w7(32'hbb09b5d1),
	.w8(32'hbb678704),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93b31b),
	.w1(32'h3b856d69),
	.w2(32'hba75a6be),
	.w3(32'h3ac00e22),
	.w4(32'h3b8a3a38),
	.w5(32'h3ac26b61),
	.w6(32'h3b86a7f5),
	.w7(32'h3ab54a9a),
	.w8(32'hba90fc23),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48a2ad),
	.w1(32'h3a27b879),
	.w2(32'h3bbf8b2c),
	.w3(32'h3b00703b),
	.w4(32'h38cc12d7),
	.w5(32'hba876fd1),
	.w6(32'h3b138ced),
	.w7(32'h3acf0f99),
	.w8(32'h398e67d4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5460d),
	.w1(32'hbb452a2a),
	.w2(32'h3abecf17),
	.w3(32'h3824998e),
	.w4(32'hbacadb6f),
	.w5(32'h3c2e73fb),
	.w6(32'hbb377a61),
	.w7(32'hbb13ec33),
	.w8(32'h3ba81eb0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aa41d),
	.w1(32'hb9f0445b),
	.w2(32'h3bebac1c),
	.w3(32'h389fc61a),
	.w4(32'hbb906f7f),
	.w5(32'h3b0d092b),
	.w6(32'h39a50474),
	.w7(32'hbbc9955c),
	.w8(32'h3bd9b540),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf309f),
	.w1(32'h3bd92bc8),
	.w2(32'h3a0d3a5e),
	.w3(32'hbbcab80d),
	.w4(32'h3b5c2801),
	.w5(32'hbb41eba5),
	.w6(32'hbb69a9bc),
	.w7(32'hb9572f3a),
	.w8(32'hbabc8d1f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d3fc),
	.w1(32'h3a2515e2),
	.w2(32'h3b12ef2b),
	.w3(32'h3b87cf6b),
	.w4(32'hbb2d753b),
	.w5(32'hbb1cad41),
	.w6(32'h3a7597ed),
	.w7(32'h39c51efd),
	.w8(32'h3b736593),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915d264),
	.w1(32'hb5aa9ec6),
	.w2(32'h3bccceb0),
	.w3(32'hbb664098),
	.w4(32'hba6472f4),
	.w5(32'h3be02018),
	.w6(32'h3aacfaa5),
	.w7(32'h3aad8f10),
	.w8(32'h3c4b7b55),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedc72a),
	.w1(32'h3a949008),
	.w2(32'h3a2d7be9),
	.w3(32'h3a18082c),
	.w4(32'h3a902979),
	.w5(32'hba95f362),
	.w6(32'hb99ba61f),
	.w7(32'hb8870441),
	.w8(32'h3ab73ace),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fb7f3),
	.w1(32'h3c1268cc),
	.w2(32'hbbdeb19f),
	.w3(32'hba55d092),
	.w4(32'h3c055bb5),
	.w5(32'hbb2f5309),
	.w6(32'h3b093670),
	.w7(32'h3bc2ef2f),
	.w8(32'hbbea126b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225363),
	.w1(32'hb93e25de),
	.w2(32'hbbb0d8b0),
	.w3(32'h39eb137b),
	.w4(32'h3a541376),
	.w5(32'hbaec5427),
	.w6(32'hbb9f9482),
	.w7(32'hbbf8ef22),
	.w8(32'hbc142705),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8bbea),
	.w1(32'h3a3d5eed),
	.w2(32'h3b2b57da),
	.w3(32'hbb44e187),
	.w4(32'hbb0bf41d),
	.w5(32'hbb4dad3a),
	.w6(32'hbbb53f88),
	.w7(32'hbb3c20da),
	.w8(32'h39bdce12),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1790e),
	.w1(32'h3981dc2e),
	.w2(32'h3acea64a),
	.w3(32'hb884f9e2),
	.w4(32'h3a240798),
	.w5(32'h3b0835fa),
	.w6(32'h3ab80d07),
	.w7(32'hbbc2c9da),
	.w8(32'hbbcfdbce),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223f5e),
	.w1(32'hb9156bf9),
	.w2(32'hbbc75f94),
	.w3(32'hbaa2a14e),
	.w4(32'hb9fe571d),
	.w5(32'hbb53d061),
	.w6(32'hbbb82452),
	.w7(32'hbb97331e),
	.w8(32'hbbfcdc9f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a822),
	.w1(32'h3b5cdfb5),
	.w2(32'hbbeeed62),
	.w3(32'hbc1e2a91),
	.w4(32'hbb43fa36),
	.w5(32'hbb6938e0),
	.w6(32'hbc428108),
	.w7(32'hbb582099),
	.w8(32'hbb147675),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed52c2),
	.w1(32'hbc0af423),
	.w2(32'hbba94e36),
	.w3(32'hbadf7ba8),
	.w4(32'hbc274b3f),
	.w5(32'hbc169ddf),
	.w6(32'h3bc3b5e6),
	.w7(32'hbc148a0c),
	.w8(32'hbb9de2b4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9882c5),
	.w1(32'hbaf658d7),
	.w2(32'h3b8cda4e),
	.w3(32'hbb4721f5),
	.w4(32'hbb0574af),
	.w5(32'hb8ddcaf2),
	.w6(32'hbada6644),
	.w7(32'hbba193be),
	.w8(32'hb9019120),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3723d),
	.w1(32'h3b5e7ef4),
	.w2(32'h3b9c6fea),
	.w3(32'hbb9622bf),
	.w4(32'h3ca9c6ff),
	.w5(32'h3d0bcae1),
	.w6(32'hbb3e2c5b),
	.w7(32'h3c2e04b8),
	.w8(32'h3c8d6b82),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b058),
	.w1(32'hbb894d49),
	.w2(32'hbb243270),
	.w3(32'h3c8af0cd),
	.w4(32'hbc0380e2),
	.w5(32'hbbc72797),
	.w6(32'h3c42ceb8),
	.w7(32'hbbc0c4c2),
	.w8(32'hbc52e5c5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0e128),
	.w1(32'h3a43c739),
	.w2(32'h3a6c8196),
	.w3(32'hbb9acf0f),
	.w4(32'h3b2f0f3f),
	.w5(32'hba51c436),
	.w6(32'hbb8cec38),
	.w7(32'h3a222f34),
	.w8(32'hbab30913),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accdcfc),
	.w1(32'h3c16473e),
	.w2(32'h3a1f2032),
	.w3(32'hba9c82f9),
	.w4(32'h3c19ea88),
	.w5(32'h3ad53a3b),
	.w6(32'hb90a2f20),
	.w7(32'h3c18182d),
	.w8(32'hba5c01bd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ae868),
	.w1(32'hbaf7c238),
	.w2(32'h3b97a93a),
	.w3(32'h3b2d97ad),
	.w4(32'hbb002cee),
	.w5(32'h3bd87d23),
	.w6(32'hba0a5e30),
	.w7(32'hbbbc75b4),
	.w8(32'h3a837e73),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac006a4),
	.w1(32'hbc3aad84),
	.w2(32'hbbc9bff7),
	.w3(32'hbaeb92a2),
	.w4(32'hbc3c962c),
	.w5(32'hbbdb17be),
	.w6(32'hbc16b1d1),
	.w7(32'hbc572642),
	.w8(32'hbc02df7d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81556),
	.w1(32'h3aa2216c),
	.w2(32'hbc00b1b4),
	.w3(32'hbb9340c6),
	.w4(32'h3c4cab41),
	.w5(32'h3bb75795),
	.w6(32'hbb9cfd33),
	.w7(32'h3bdbbcfc),
	.w8(32'hb8eb96e8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85d594),
	.w1(32'hbb30dfd9),
	.w2(32'hbb1135b5),
	.w3(32'hbc597c20),
	.w4(32'hbab74dc1),
	.w5(32'hbbb43b95),
	.w6(32'hbc63f2f3),
	.w7(32'hbaaf1855),
	.w8(32'hbbac8f2d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4796),
	.w1(32'h3ad750f7),
	.w2(32'hbb24a48e),
	.w3(32'hbc18e5a9),
	.w4(32'h3b1f7ddb),
	.w5(32'h3b1142ba),
	.w6(32'hbc1ea823),
	.w7(32'h3a9b1d5c),
	.w8(32'hba4a7cad),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71ad1),
	.w1(32'hbcc21aee),
	.w2(32'hbc675d49),
	.w3(32'hb9bec228),
	.w4(32'hbcd762c4),
	.w5(32'h3b2d57a2),
	.w6(32'hbb4a7ba7),
	.w7(32'hbc96e1d7),
	.w8(32'hba89d637),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd632),
	.w1(32'hba1f636c),
	.w2(32'hbbdd1257),
	.w3(32'h3d108c31),
	.w4(32'hbac37314),
	.w5(32'hbb95181e),
	.w6(32'h3cce8167),
	.w7(32'hbb02b63a),
	.w8(32'hbb99d800),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d330),
	.w1(32'hbc4703a5),
	.w2(32'hbc361e9e),
	.w3(32'h3b2e7c62),
	.w4(32'hbc234883),
	.w5(32'h3aaccd94),
	.w6(32'h3c2d6aca),
	.w7(32'hbc8fcb9c),
	.w8(32'hbc25785a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892dbf),
	.w1(32'hbb8f57c5),
	.w2(32'hbab6817a),
	.w3(32'h3bdc877e),
	.w4(32'hba993979),
	.w5(32'hbb38cedf),
	.w6(32'hbadca465),
	.w7(32'h370951ca),
	.w8(32'hbb9adfb4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e0dd),
	.w1(32'hbb954a7a),
	.w2(32'hbb3d76e5),
	.w3(32'h3b527ab1),
	.w4(32'hbc0ffb15),
	.w5(32'hbac9b534),
	.w6(32'h3aa1a7a7),
	.w7(32'hbc04a7e9),
	.w8(32'h38ee5713),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dc95b),
	.w1(32'hbadc187f),
	.w2(32'hba9447e2),
	.w3(32'h37cd16c7),
	.w4(32'hbb7b0b68),
	.w5(32'h3abc9b3f),
	.w6(32'h3a00a7d5),
	.w7(32'hbb3f6623),
	.w8(32'hbb263a75),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e58bed),
	.w1(32'h3aa77f10),
	.w2(32'h3b448e83),
	.w3(32'hb99fdbf5),
	.w4(32'h3a4514bf),
	.w5(32'h392a55ae),
	.w6(32'h394cab6d),
	.w7(32'h3b1362d2),
	.w8(32'h3b96801e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0211),
	.w1(32'hbc834417),
	.w2(32'hbc658809),
	.w3(32'hba467295),
	.w4(32'hbc615b45),
	.w5(32'hbc18eaed),
	.w6(32'h39ecdf86),
	.w7(32'hbc491b46),
	.w8(32'hbc1dc789),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67ab14),
	.w1(32'hbc0e0f7e),
	.w2(32'hbbc66154),
	.w3(32'hbc424ee5),
	.w4(32'hbc9c5c95),
	.w5(32'hbc92442e),
	.w6(32'hbc476bcf),
	.w7(32'hbc76f87f),
	.w8(32'hbbd52854),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc722339),
	.w1(32'h3c856a37),
	.w2(32'h3c2c982d),
	.w3(32'hbcc376cb),
	.w4(32'h3ccf883f),
	.w5(32'h3cec2bb1),
	.w6(32'hbcacbabf),
	.w7(32'h3cd94ad9),
	.w8(32'h3cb4b540),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c960fc4),
	.w1(32'h3b6de0b6),
	.w2(32'h3b165a31),
	.w3(32'h3d044d33),
	.w4(32'h3b66f536),
	.w5(32'h3b8794b4),
	.w6(32'h3cbc2a1b),
	.w7(32'h3b85520a),
	.w8(32'h3a947f09),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9f4ac),
	.w1(32'h3bf5af4b),
	.w2(32'h3a997e5b),
	.w3(32'hba442587),
	.w4(32'h3c0a37c7),
	.w5(32'hbb3f90db),
	.w6(32'hbb42bb73),
	.w7(32'h3c0ee956),
	.w8(32'hbaafdb4c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdc677),
	.w1(32'h38b4cf24),
	.w2(32'h3ba247e7),
	.w3(32'h3ad918f5),
	.w4(32'h3a081840),
	.w5(32'h3b97a24f),
	.w6(32'h3b24d025),
	.w7(32'hb8f2b443),
	.w8(32'h3b423187),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cdf09),
	.w1(32'hbbb91649),
	.w2(32'hbb4acfb5),
	.w3(32'h3bd517dd),
	.w4(32'hba764d99),
	.w5(32'hbb75b7df),
	.w6(32'h3b6e47e9),
	.w7(32'hba99791b),
	.w8(32'hbbc9c901),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47dbf2),
	.w1(32'hbba35c9d),
	.w2(32'hbc22e1af),
	.w3(32'hbae09aee),
	.w4(32'h3a532e9e),
	.w5(32'hba3e9f26),
	.w6(32'hbb70a548),
	.w7(32'h3a1f169a),
	.w8(32'hbbd17779),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4329a),
	.w1(32'h3ae79155),
	.w2(32'h3b3f7825),
	.w3(32'hba8d000c),
	.w4(32'hb8cd0737),
	.w5(32'h3c192858),
	.w6(32'hbb950b4c),
	.w7(32'hb9cae11e),
	.w8(32'h3bde0609),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26b56b),
	.w1(32'h3a57e6d7),
	.w2(32'h3a0e861f),
	.w3(32'hbacafcbc),
	.w4(32'hbb4267d0),
	.w5(32'hbb5e0cbb),
	.w6(32'hbb3d1cb6),
	.w7(32'hbb0bf721),
	.w8(32'hb9394cad),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cdf83),
	.w1(32'h3b0ae652),
	.w2(32'hbae8df87),
	.w3(32'hbb09bfd2),
	.w4(32'h3b8bff21),
	.w5(32'hbaeae522),
	.w6(32'h3a8ea442),
	.w7(32'hb9f6295a),
	.w8(32'hbb5a821d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4b72),
	.w1(32'hbb74dc71),
	.w2(32'hbc3b9afe),
	.w3(32'hbb3da03b),
	.w4(32'hbb77e6f8),
	.w5(32'hbc4d6818),
	.w6(32'hbbb0a399),
	.w7(32'hbb09db87),
	.w8(32'hbc5f5698),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8f1c7),
	.w1(32'hbaa2ec53),
	.w2(32'h3ab821dc),
	.w3(32'hbb9f54de),
	.w4(32'hba4668a4),
	.w5(32'hbb4cf85c),
	.w6(32'hbbc7485b),
	.w7(32'hba7ab195),
	.w8(32'hba868ece),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2276a),
	.w1(32'h3b61eaee),
	.w2(32'h3a912dea),
	.w3(32'hbb2c211f),
	.w4(32'h3b56897c),
	.w5(32'hb9fa2075),
	.w6(32'hbb9a6bfe),
	.w7(32'h3b290c93),
	.w8(32'h3a856a70),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3ef0f),
	.w1(32'hbb725ddc),
	.w2(32'hbb984af7),
	.w3(32'hbbf6e484),
	.w4(32'hbae38688),
	.w5(32'hbaea40c5),
	.w6(32'hbabe75e9),
	.w7(32'hbb0d63d9),
	.w8(32'h398ef13d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30fd56),
	.w1(32'h3b7667c6),
	.w2(32'hbb143b5c),
	.w3(32'h3b009ed6),
	.w4(32'h3bb05b6d),
	.w5(32'h3c34498e),
	.w6(32'h3bc4f7b4),
	.w7(32'h3a1bf175),
	.w8(32'hbbda60c8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6efb17),
	.w1(32'hba632872),
	.w2(32'hbab1af39),
	.w3(32'h3cdebbbe),
	.w4(32'hbb88f3c4),
	.w5(32'hbbaf67da),
	.w6(32'h3c898ae9),
	.w7(32'hbb2d7872),
	.w8(32'hbafd81a5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07366b),
	.w1(32'h3ba2a83e),
	.w2(32'h3b391852),
	.w3(32'hbafce0f5),
	.w4(32'h3a8b6c80),
	.w5(32'hb898c974),
	.w6(32'h3b4772f6),
	.w7(32'h3ad05f88),
	.w8(32'h3996af90),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67f4a3),
	.w1(32'hbb92c1ef),
	.w2(32'h3afa65c9),
	.w3(32'h3a5a018e),
	.w4(32'hbbeec70f),
	.w5(32'hbaee2436),
	.w6(32'h3ac255cf),
	.w7(32'hbbc89fc3),
	.w8(32'hbaba614a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb77ecd),
	.w1(32'hbb5b3e4f),
	.w2(32'h3b808afc),
	.w3(32'hbc02417a),
	.w4(32'hbb54db6c),
	.w5(32'h3b78e0eb),
	.w6(32'hbbb7854a),
	.w7(32'hb9c89de5),
	.w8(32'h3bb70cec),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49c714),
	.w1(32'h3baffce3),
	.w2(32'hba5bc317),
	.w3(32'hbbff7e0d),
	.w4(32'hb99fa3ea),
	.w5(32'h3b1d2708),
	.w6(32'hbbe3923a),
	.w7(32'h3b820785),
	.w8(32'h3b9488ac),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ea578),
	.w1(32'hbb1bb503),
	.w2(32'hbbccb419),
	.w3(32'h3bd1cb9e),
	.w4(32'hbba17a1b),
	.w5(32'hbb20e15a),
	.w6(32'h3bd0caae),
	.w7(32'hbae11a77),
	.w8(32'hbbb6b3c1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41234f),
	.w1(32'hb9b31c20),
	.w2(32'h390068d5),
	.w3(32'h3ac9c80a),
	.w4(32'hb6aa129b),
	.w5(32'h39a72cca),
	.w6(32'h3b0ff9a7),
	.w7(32'hba36ce3b),
	.w8(32'h39095194),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373ec0ee),
	.w1(32'hb7a11459),
	.w2(32'h3695b65b),
	.w3(32'hb8208db9),
	.w4(32'hb6d489d2),
	.w5(32'h3782fe55),
	.w6(32'hb8255d2a),
	.w7(32'hb60b492f),
	.w8(32'h3730eb74),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37417d86),
	.w1(32'h366e67a1),
	.w2(32'hb792820c),
	.w3(32'h36117a53),
	.w4(32'h37306200),
	.w5(32'h367415f1),
	.w6(32'h371fc8de),
	.w7(32'h37c1c6a0),
	.w8(32'h3798dbbe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372e4fc4),
	.w1(32'hb7b0d416),
	.w2(32'h3780f8d3),
	.w3(32'hb7636082),
	.w4(32'hb7369595),
	.w5(32'h372ec8df),
	.w6(32'hb58fa19d),
	.w7(32'h3609b2b3),
	.w8(32'h370c031d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815eb67),
	.w1(32'hb813c906),
	.w2(32'hb7895395),
	.w3(32'hb83a786b),
	.w4(32'hb7f0f9f7),
	.w5(32'hb71d533b),
	.w6(32'hb85b578f),
	.w7(32'hb7aea33a),
	.w8(32'hb758264e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3719ad1c),
	.w1(32'h37ceac46),
	.w2(32'h37349c56),
	.w3(32'h371c6d81),
	.w4(32'h3773fc3a),
	.w5(32'h3506ccbf),
	.w6(32'hb71f065c),
	.w7(32'h3815017c),
	.w8(32'h37221a42),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937010f),
	.w1(32'hb8f129d6),
	.w2(32'hb7ff8156),
	.w3(32'hb8a16624),
	.w4(32'h331bf6f4),
	.w5(32'h370811c0),
	.w6(32'hb983c7da),
	.w7(32'hb8c0bacf),
	.w8(32'hb81c5878),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abf375),
	.w1(32'hb8c81d4d),
	.w2(32'hb79dfe2d),
	.w3(32'hb744a4ce),
	.w4(32'h36875e56),
	.w5(32'h37e01ed2),
	.w6(32'hb9f20f19),
	.w7(32'hb9ab20d8),
	.w8(32'hb8aaa83c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9447226),
	.w1(32'hb8f0ca17),
	.w2(32'h38e2d1d4),
	.w3(32'hb930ed60),
	.w4(32'hb7bb3968),
	.w5(32'h39422547),
	.w6(32'hb9bda826),
	.w7(32'hb9a8dc15),
	.w8(32'h38c2d58e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957bf98),
	.w1(32'hb8c8beff),
	.w2(32'hb78e6d5d),
	.w3(32'hb8f93c54),
	.w4(32'hb87e57f8),
	.w5(32'h37d8431a),
	.w6(32'hb9961d8c),
	.w7(32'hb92d7ab4),
	.w8(32'hb7803590),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f9627),
	.w1(32'hb82f2481),
	.w2(32'hb69d4ce1),
	.w3(32'hb87f4b60),
	.w4(32'hb79b84aa),
	.w5(32'h380e8f72),
	.w6(32'hb918db0e),
	.w7(32'hb9070fa0),
	.w8(32'hb7ccbca8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888daee),
	.w1(32'hb80f605a),
	.w2(32'h379f3958),
	.w3(32'hb860c778),
	.w4(32'h379cf8fe),
	.w5(32'h38ad597e),
	.w6(32'hb919c9ff),
	.w7(32'hb8f93aa1),
	.w8(32'h384b7898),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91adc1b),
	.w1(32'hb894bf60),
	.w2(32'hb8057d0f),
	.w3(32'hb88004d1),
	.w4(32'hb87f339a),
	.w5(32'hb7bd57c7),
	.w6(32'hb95af318),
	.w7(32'hb905416a),
	.w8(32'hb858d2cc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3533cb55),
	.w1(32'hb5a5ef90),
	.w2(32'hb74657af),
	.w3(32'hb6eadd57),
	.w4(32'hb6a1429b),
	.w5(32'hb720c26f),
	.w6(32'h36d9a029),
	.w7(32'hb682cf7f),
	.w8(32'h364a1da3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75e4444),
	.w1(32'hb83c7db5),
	.w2(32'hb76f63f8),
	.w3(32'hb7a718e6),
	.w4(32'hb652db01),
	.w5(32'h37f575b7),
	.w6(32'hb72597bb),
	.w7(32'h3703d64b),
	.w8(32'h36da8cad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62919c3),
	.w1(32'hb8087bf4),
	.w2(32'h373c17b6),
	.w3(32'h36ae5f95),
	.w4(32'hb58a5d1b),
	.w5(32'h37924465),
	.w6(32'hb7036bbc),
	.w7(32'hb7f3301a),
	.w8(32'h370abeb6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53c71db),
	.w1(32'h37408e8a),
	.w2(32'h36bbb35b),
	.w3(32'hb6335114),
	.w4(32'h381a14f2),
	.w5(32'hb766af0c),
	.w6(32'hb7008e2b),
	.w7(32'hb6c67464),
	.w8(32'h37657655),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b292),
	.w1(32'hb905ac2d),
	.w2(32'h38af36e1),
	.w3(32'hb91bc722),
	.w4(32'hb836bacd),
	.w5(32'h39155448),
	.w6(32'hb99d435f),
	.w7(32'hb974d8bd),
	.w8(32'h38bff429),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787a926),
	.w1(32'h37a3cb0c),
	.w2(32'h370f2185),
	.w3(32'h38177a4e),
	.w4(32'h37f09b41),
	.w5(32'h3754ccf8),
	.w6(32'hb797bbfc),
	.w7(32'hb7b3fe81),
	.w8(32'h3761ccdd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946fa9d),
	.w1(32'hb92e524f),
	.w2(32'hb84048de),
	.w3(32'hb8f58d39),
	.w4(32'hb8b8b000),
	.w5(32'h380516d0),
	.w6(32'hb98b0424),
	.w7(32'hb951ade3),
	.w8(32'hb8455f52),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a001db),
	.w1(32'hb7fb3696),
	.w2(32'hb8e42b5a),
	.w3(32'hb954b99d),
	.w4(32'hb81170b8),
	.w5(32'hb8f55a31),
	.w6(32'hba414307),
	.w7(32'hb97cf0de),
	.w8(32'hb960a664),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb834d4d7),
	.w1(32'h378c8717),
	.w2(32'h3809f0d9),
	.w3(32'h3907cc8e),
	.w4(32'h391d83e1),
	.w5(32'h390c4a2b),
	.w6(32'hb7456a9f),
	.w7(32'hb87b00c7),
	.w8(32'h3863db82),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f933e),
	.w1(32'hb92e3c4c),
	.w2(32'h3813c7e6),
	.w3(32'hb8be854f),
	.w4(32'h37e75631),
	.w5(32'h38e05034),
	.w6(32'hb9b47ba1),
	.w7(32'hb9b982a8),
	.w8(32'hb881262d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b284f),
	.w1(32'hb8fd264e),
	.w2(32'hb8570c3e),
	.w3(32'hb8ff7227),
	.w4(32'hb8228897),
	.w5(32'h385669a4),
	.w6(32'hb93b64bd),
	.w7(32'hb8f41146),
	.w8(32'h37e1a026),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980b429),
	.w1(32'hb9337b78),
	.w2(32'h38464f1a),
	.w3(32'hb91df9df),
	.w4(32'hb798e01e),
	.w5(32'h390431b2),
	.w6(32'hb9b416bb),
	.w7(32'hb9955cfd),
	.w8(32'h37f1deed),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932d500),
	.w1(32'hb956e8e5),
	.w2(32'hb88403cf),
	.w3(32'hb92bbe5b),
	.w4(32'hb8db6d94),
	.w5(32'h37a05fc1),
	.w6(32'hb98c13e4),
	.w7(32'hb9603196),
	.w8(32'hb8c56132),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9387a40),
	.w1(32'hb9025b35),
	.w2(32'hb68ddf94),
	.w3(32'hb87baa61),
	.w4(32'h3711b4bf),
	.w5(32'h38f26492),
	.w6(32'hb95f0acc),
	.w7(32'hb98c6fdf),
	.w8(32'h375dd899),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b39738),
	.w1(32'hb6d409ea),
	.w2(32'hb6520d42),
	.w3(32'h373ecc00),
	.w4(32'h370c30f5),
	.w5(32'hb75ed291),
	.w6(32'h3705140a),
	.w7(32'hb49b3e77),
	.w8(32'hb74e9a6f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d1af8),
	.w1(32'hb8fbe69e),
	.w2(32'hb53bfcd0),
	.w3(32'hb901f59c),
	.w4(32'hb829be59),
	.w5(32'h38b7addb),
	.w6(32'hb9d0c4e4),
	.w7(32'hb9b64126),
	.w8(32'h34371eec),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b04ca7),
	.w1(32'hb93a9a23),
	.w2(32'hb890e6c6),
	.w3(32'hb883eeb8),
	.w4(32'hb80faca7),
	.w5(32'h38770a56),
	.w6(32'hb9481332),
	.w7(32'hb9834480),
	.w8(32'hb7895524),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba012e83),
	.w1(32'hb8fea777),
	.w2(32'hb863d5ef),
	.w3(32'hb989d831),
	.w4(32'hb8ec9152),
	.w5(32'hb901526e),
	.w6(32'hba0d7698),
	.w7(32'hb9ad73d2),
	.w8(32'hb93b0257),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a18de6),
	.w1(32'hb9c06601),
	.w2(32'hb8369488),
	.w3(32'h380ef2c5),
	.w4(32'h390e379a),
	.w5(32'h3966e471),
	.w6(32'hb936dd1c),
	.w7(32'hb9de73ba),
	.w8(32'h3803988e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999fe2e),
	.w1(32'hb9438740),
	.w2(32'h38098bb6),
	.w3(32'hb959bdcd),
	.w4(32'hb82a43e5),
	.w5(32'h39346e61),
	.w6(32'hb9f45f52),
	.w7(32'hb9d1317a),
	.w8(32'h38143354),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968812a),
	.w1(32'hb9042d04),
	.w2(32'hb8bffda4),
	.w3(32'hb9345ef0),
	.w4(32'hb8066070),
	.w5(32'hb7c52fda),
	.w6(32'hb97edb2d),
	.w7(32'hb94ae4f4),
	.w8(32'hb8c8e263),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cfaab5),
	.w1(32'hb7718e06),
	.w2(32'h3727fe76),
	.w3(32'h3832f20f),
	.w4(32'hb7bdff41),
	.w5(32'hb728e835),
	.w6(32'h3820c137),
	.w7(32'hb6f2b463),
	.w8(32'hb797fe88),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949a758),
	.w1(32'hb84a4a4d),
	.w2(32'hb8a6881e),
	.w3(32'hb8f0a933),
	.w4(32'h386d3d6a),
	.w5(32'hb89f552c),
	.w6(32'hb9f40fc7),
	.w7(32'hb969cfaf),
	.w8(32'hb8a689b7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81aa88e),
	.w1(32'hb8a3d97d),
	.w2(32'hb84d80c4),
	.w3(32'hb89ed38e),
	.w4(32'hb827c1a3),
	.w5(32'h380c9b63),
	.w6(32'hb873a7cd),
	.w7(32'hb97374b3),
	.w8(32'h371128c1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742855a),
	.w1(32'hb601e731),
	.w2(32'h373b185f),
	.w3(32'h365ba368),
	.w4(32'h35dccd03),
	.w5(32'h36870965),
	.w6(32'h3725bbc8),
	.w7(32'h36795f12),
	.w8(32'h36ea2804),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b024f7),
	.w1(32'hb83948f0),
	.w2(32'hb7165a32),
	.w3(32'hb8d16291),
	.w4(32'hb8858b77),
	.w5(32'h38121b87),
	.w6(32'hb8ee350e),
	.w7(32'hb8977d51),
	.w8(32'hb72825fc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923f9c7),
	.w1(32'hb84e9f3b),
	.w2(32'h3836b6e9),
	.w3(32'hb8b1718d),
	.w4(32'h37632eab),
	.w5(32'h3912789d),
	.w6(32'hb98a49cd),
	.w7(32'hb9731a75),
	.w8(32'h38837a32),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912b298),
	.w1(32'hb8bda115),
	.w2(32'h37e4c524),
	.w3(32'hb901b778),
	.w4(32'h379c0dd7),
	.w5(32'h3910c79d),
	.w6(32'hb990fe67),
	.w7(32'hb9800b6d),
	.w8(32'h384d35a6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38107454),
	.w1(32'hb619e19a),
	.w2(32'h389dee5e),
	.w3(32'hb6474bfd),
	.w4(32'h3921b8d2),
	.w5(32'h391089fb),
	.w6(32'hb92b9666),
	.w7(32'hb8b4ce2d),
	.w8(32'h380e8b7d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ff45e),
	.w1(32'hb8b77d89),
	.w2(32'h381bc1a0),
	.w3(32'hb9048f95),
	.w4(32'hb7fe7ad7),
	.w5(32'h389a3ffb),
	.w6(32'hb9748439),
	.w7(32'hb94c1657),
	.w8(32'hb7c81ae0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9d76e),
	.w1(32'hb8305f01),
	.w2(32'hb7b87d0c),
	.w3(32'h37dbe7d0),
	.w4(32'h38067fa1),
	.w5(32'hb6369c2a),
	.w6(32'hb88b313b),
	.w7(32'hb85c2c7e),
	.w8(32'hb688c63a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e41b45),
	.w1(32'hb84fca1a),
	.w2(32'h358be82c),
	.w3(32'hb86d34d7),
	.w4(32'hb7e1b508),
	.w5(32'h388e9ff2),
	.w6(32'hb9404db5),
	.w7(32'hb928e552),
	.w8(32'hb78dc04f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6c7d4),
	.w1(32'hb867e315),
	.w2(32'h38136a53),
	.w3(32'hb8994ca8),
	.w4(32'h37713826),
	.w5(32'h38ee404f),
	.w6(32'hb96d468b),
	.w7(32'hb93cd84c),
	.w8(32'h38002998),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c04121),
	.w1(32'hb75fee0a),
	.w2(32'hb6edfe3e),
	.w3(32'h36840e9f),
	.w4(32'h3694fc55),
	.w5(32'hb6829c4b),
	.w6(32'hb5e8ccae),
	.w7(32'h36f26c0f),
	.w8(32'hb56e0078),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7188053),
	.w1(32'h37ef3cf7),
	.w2(32'hb71e760a),
	.w3(32'hb72ef3fa),
	.w4(32'h3793424c),
	.w5(32'hb77b9a66),
	.w6(32'hb764167a),
	.w7(32'h37a165d5),
	.w8(32'hb6f6424f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d425a6),
	.w1(32'hb73a7b51),
	.w2(32'h370366a2),
	.w3(32'hb78b73ca),
	.w4(32'h370a9dc9),
	.w5(32'hb6efa722),
	.w6(32'hb60b1bad),
	.w7(32'hb55e44bc),
	.w8(32'hb735f7e7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806741e),
	.w1(32'h37c00dbb),
	.w2(32'h34993a1d),
	.w3(32'hb8241383),
	.w4(32'hb6d1aa26),
	.w5(32'hb75e2927),
	.w6(32'hb63b6fe0),
	.w7(32'hb7643352),
	.w8(32'hb654b507),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bdde8),
	.w1(32'hb8bf7158),
	.w2(32'h37b1f42f),
	.w3(32'hb8e504a5),
	.w4(32'hb797ae90),
	.w5(32'h38d61a14),
	.w6(32'hb98e3c66),
	.w7(32'hb976e99f),
	.w8(32'h3887bd87),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361c589e),
	.w1(32'hb747b79c),
	.w2(32'hb788e550),
	.w3(32'h372106ae),
	.w4(32'hb704a0fd),
	.w5(32'h368e20ee),
	.w6(32'h38092ea7),
	.w7(32'hb662a338),
	.w8(32'hb62ac06d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c71bd),
	.w1(32'hb853d23e),
	.w2(32'hb7aa7d00),
	.w3(32'hb6961796),
	.w4(32'hb8565101),
	.w5(32'hb8555e63),
	.w6(32'hb8cb3074),
	.w7(32'hb8b45e76),
	.w8(32'hb8137e84),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9601a14),
	.w1(32'hb8b0cc71),
	.w2(32'hb817f01a),
	.w3(32'hb96d355f),
	.w4(32'hb83073f8),
	.w5(32'h375e922d),
	.w6(32'hb97686e7),
	.w7(32'hb9af556a),
	.w8(32'hb8aeb1cc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57aca92),
	.w1(32'h36d1ce5d),
	.w2(32'hb7b37105),
	.w3(32'h376e4e3b),
	.w4(32'hb70ca219),
	.w5(32'hb7ea252c),
	.w6(32'h37d137ad),
	.w7(32'h3618b6a8),
	.w8(32'hb7d4d742),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3733821d),
	.w1(32'hb5f4b291),
	.w2(32'hb7635373),
	.w3(32'h37535ed7),
	.w4(32'h37ce0547),
	.w5(32'hb612f5a4),
	.w6(32'h381210a0),
	.w7(32'hb6850a34),
	.w8(32'h372387a3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ab25f),
	.w1(32'hb7299c2c),
	.w2(32'h370ab576),
	.w3(32'hb795e193),
	.w4(32'h372a292d),
	.w5(32'h37853172),
	.w6(32'h3630907e),
	.w7(32'h37c6cf61),
	.w8(32'h371c8b1e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7723b22),
	.w1(32'hb7c89c22),
	.w2(32'h37d3af23),
	.w3(32'hb8258596),
	.w4(32'h376f2f80),
	.w5(32'h37b14e48),
	.w6(32'hb8258db6),
	.w7(32'hb7a24eeb),
	.w8(32'hb7605a3d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9288b65),
	.w1(32'hb87210c7),
	.w2(32'h373e6c48),
	.w3(32'hb8c5d7f6),
	.w4(32'h37a53a1f),
	.w5(32'h380d1a71),
	.w6(32'hb98447b8),
	.w7(32'hb926c9c0),
	.w8(32'h37a4552a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ece02),
	.w1(32'hb8dca16d),
	.w2(32'hb7d55278),
	.w3(32'hb93bb453),
	.w4(32'hb87ea521),
	.w5(32'h37d415a3),
	.w6(32'hb9a6c84b),
	.w7(32'hb972c60d),
	.w8(32'hb802c5fa),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ae6950),
	.w1(32'hb72d6674),
	.w2(32'hb77c7061),
	.w3(32'h3528476c),
	.w4(32'h35f454a8),
	.w5(32'hb5836be9),
	.w6(32'h3657d87d),
	.w7(32'h372a4f35),
	.w8(32'hb59450c0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb822c3f0),
	.w1(32'hb7a50b2b),
	.w2(32'h38821ae7),
	.w3(32'h3866e595),
	.w4(32'h382daa77),
	.w5(32'h3806acb7),
	.w6(32'hb8c698d3),
	.w7(32'hb7d96c96),
	.w8(32'hb739da84),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87094a5),
	.w1(32'hb88eb2dc),
	.w2(32'h36da87d8),
	.w3(32'hb80762cf),
	.w4(32'hb56f2e1b),
	.w5(32'h38410106),
	.w6(32'hb8cd5e3e),
	.w7(32'hb8ac73bd),
	.w8(32'h37672533),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885ddde),
	.w1(32'hb608cb8e),
	.w2(32'h363daad8),
	.w3(32'hb88546f2),
	.w4(32'h37869546),
	.w5(32'h380e7f32),
	.w6(32'hb93ee77b),
	.w7(32'hb8a4badf),
	.w8(32'hb70d8807),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e4a6e),
	.w1(32'hb8f0e4fa),
	.w2(32'hb7e8757d),
	.w3(32'hb9b6fe5c),
	.w4(32'hb8f98a85),
	.w5(32'hb6d1134a),
	.w6(32'hb9b027a8),
	.w7(32'hb92d6e43),
	.w8(32'hb885d00a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b9b33),
	.w1(32'hb8ebaa7a),
	.w2(32'hb70807d4),
	.w3(32'hb8d37af5),
	.w4(32'hb85cf648),
	.w5(32'h382d72b9),
	.w6(32'hb9c18310),
	.w7(32'hb98c055d),
	.w8(32'hb8844522),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9156b),
	.w1(32'hb91406f3),
	.w2(32'h363e0a52),
	.w3(32'hb859ab58),
	.w4(32'h371a11c0),
	.w5(32'h38a4fbe8),
	.w6(32'hb9600654),
	.w7(32'hb9823c6a),
	.w8(32'h36e54a59),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91380ca),
	.w1(32'hb9409954),
	.w2(32'hb8858d44),
	.w3(32'hb90aa53d),
	.w4(32'hb8d1f47f),
	.w5(32'h34932d32),
	.w6(32'hb98f25a7),
	.w7(32'hb9826e7b),
	.w8(32'hb8bc7499),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978c6f3),
	.w1(32'hb90a7a83),
	.w2(32'hb8f4dc3c),
	.w3(32'hb9157d89),
	.w4(32'hb8dc26ca),
	.w5(32'hb8bc5ad9),
	.w6(32'hb9b886b5),
	.w7(32'hb957d67a),
	.w8(32'hb904c8aa),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fb55a),
	.w1(32'hb901e0af),
	.w2(32'hb7d4cfff),
	.w3(32'hb908b9e3),
	.w4(32'hb7bd6818),
	.w5(32'h38414417),
	.w6(32'hb96fc660),
	.w7(32'hb939d0f7),
	.w8(32'h36ab24ec),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9161258),
	.w1(32'hb8c0dca0),
	.w2(32'hb76b7ec6),
	.w3(32'hb8b95b0e),
	.w4(32'hb70703f6),
	.w5(32'h382a3a27),
	.w6(32'hb93866b1),
	.w7(32'hb923fd9b),
	.w8(32'hb750c420),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e27fdb),
	.w1(32'hb88e737b),
	.w2(32'hb72dc3ad),
	.w3(32'hb781e875),
	.w4(32'hb74690ab),
	.w5(32'h378214ab),
	.w6(32'hb899a89a),
	.w7(32'hb8064876),
	.w8(32'h373ca873),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c51332),
	.w1(32'hb942bbb9),
	.w2(32'h37ad38fc),
	.w3(32'hb970ca52),
	.w4(32'hb5dfa424),
	.w5(32'h3947880b),
	.w6(32'hb9c85d06),
	.w7(32'hb9c71a8c),
	.w8(32'h36a1e3c3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c07fff),
	.w1(32'hb883bf37),
	.w2(32'hb7e8a4b5),
	.w3(32'hb85d6988),
	.w4(32'hb780c802),
	.w5(32'hb790ed7a),
	.w6(32'hb8cb0f62),
	.w7(32'hb8b30d92),
	.w8(32'hb84d8a93),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3682561d),
	.w1(32'hb6cc3b18),
	.w2(32'h361ce136),
	.w3(32'h35d306eb),
	.w4(32'h3764506d),
	.w5(32'h35e97849),
	.w6(32'h373cb322),
	.w7(32'hb7064222),
	.w8(32'h351bfb2e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a506fd),
	.w1(32'h37af1c85),
	.w2(32'h36ddef23),
	.w3(32'hb7887b06),
	.w4(32'hb68a06eb),
	.w5(32'h3665811e),
	.w6(32'hb7dd21b1),
	.w7(32'hb5dbe220),
	.w8(32'hb6a5d98d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83e5895),
	.w1(32'hb8201211),
	.w2(32'h37f2cb4c),
	.w3(32'hb77db9e6),
	.w4(32'hb7b50b57),
	.w5(32'h38264f2f),
	.w6(32'hb89c74fb),
	.w7(32'hb8dc6212),
	.w8(32'h3813cc09),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9207e75),
	.w1(32'hb8d34ef9),
	.w2(32'h35b0534e),
	.w3(32'hb6af1375),
	.w4(32'h385b445b),
	.w5(32'h39009eb6),
	.w6(32'hb936e876),
	.w7(32'hb94ad378),
	.w8(32'h37ce9df6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9ca00),
	.w1(32'hb8c421e7),
	.w2(32'h38cf6813),
	.w3(32'hb8d2c5c0),
	.w4(32'hb80bc08e),
	.w5(32'h392395da),
	.w6(32'hb9b6cf0a),
	.w7(32'hb9b08b2e),
	.w8(32'h38376dba),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3706b8ed),
	.w1(32'hb5ab2c74),
	.w2(32'hb741c636),
	.w3(32'h37ebbf7f),
	.w4(32'h37578833),
	.w5(32'hb63dcf3d),
	.w6(32'h373485f0),
	.w7(32'h3781f4eb),
	.w8(32'hb5445aa2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935e416),
	.w1(32'hb8f3cfd0),
	.w2(32'h37f0ee3f),
	.w3(32'hb908ab95),
	.w4(32'hb7a8ca28),
	.w5(32'h38b821e5),
	.w6(32'hb9a1a514),
	.w7(32'hb985d84f),
	.w8(32'hb675b676),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9d2b8),
	.w1(32'hb90b5684),
	.w2(32'h37fcab49),
	.w3(32'hb8b9432c),
	.w4(32'hb8377475),
	.w5(32'h38a764a0),
	.w6(32'hb95f8951),
	.w7(32'hb971836d),
	.w8(32'h3824d8a1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90334e8),
	.w1(32'hb8c69fdc),
	.w2(32'hb883a03e),
	.w3(32'hb8b8343d),
	.w4(32'hb80e7839),
	.w5(32'hb7a3f30d),
	.w6(32'hb95a41f2),
	.w7(32'hb8edb2fd),
	.w8(32'hb86021be),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f44f6),
	.w1(32'hb94f180e),
	.w2(32'h3836bf38),
	.w3(32'hb910eb66),
	.w4(32'hb8e9608a),
	.w5(32'h3959d129),
	.w6(32'hb9aeeee6),
	.w7(32'hb9bd7869),
	.w8(32'h388336d3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a11c9d),
	.w1(32'hb82089e7),
	.w2(32'h38212f62),
	.w3(32'hb8830501),
	.w4(32'hb7be213d),
	.w5(32'h36a9cc23),
	.w6(32'hb80c9f3c),
	.w7(32'hb83c1b3c),
	.w8(32'h375691c6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f884d8),
	.w1(32'h374ba920),
	.w2(32'hb655c59c),
	.w3(32'h36839a50),
	.w4(32'h36a28b8b),
	.w5(32'hb7605e7f),
	.w6(32'h38351c43),
	.w7(32'hb65b45d8),
	.w8(32'hb7255e80),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742e6d8),
	.w1(32'hb7a11ab4),
	.w2(32'h37d1d16d),
	.w3(32'h388a303d),
	.w4(32'h38a02480),
	.w5(32'h3882f474),
	.w6(32'hb833bb1c),
	.w7(32'hb8b38194),
	.w8(32'h382162ad),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8faa5ba),
	.w1(32'hb8c619d1),
	.w2(32'hb81e3cf9),
	.w3(32'hb5e6946b),
	.w4(32'h37f6728a),
	.w5(32'h37e74e08),
	.w6(32'hb87e34d2),
	.w7(32'hb8667fe1),
	.w8(32'hb7abe972),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37825de0),
	.w1(32'h374072ff),
	.w2(32'h36d57b6b),
	.w3(32'h38841a03),
	.w4(32'h388e7971),
	.w5(32'h3785f901),
	.w6(32'h37ed1279),
	.w7(32'h37588a4e),
	.w8(32'h37cedbb7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896a6bb),
	.w1(32'hb757ac7b),
	.w2(32'hb7a18f31),
	.w3(32'h36952ba3),
	.w4(32'h38144309),
	.w5(32'h3828a674),
	.w6(32'hb8c3d2be),
	.w7(32'hb83b75cc),
	.w8(32'hb7c89bd5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dce652),
	.w1(32'hb65db7d7),
	.w2(32'h3745825c),
	.w3(32'hb5cc09c5),
	.w4(32'hb7179cbb),
	.w5(32'hb7a82c1a),
	.w6(32'hb7bb5aa0),
	.w7(32'hb66a7451),
	.w8(32'hb67e3b26),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9386992),
	.w1(32'hb89a85bc),
	.w2(32'hb6fc5c99),
	.w3(32'hb908ef50),
	.w4(32'hb802c2f9),
	.w5(32'h38587a5c),
	.w6(32'hb98fed09),
	.w7(32'hb93a8bd9),
	.w8(32'hb8012167),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8291e52),
	.w1(32'hb6f67ee2),
	.w2(32'hb769d08b),
	.w3(32'hb780f64e),
	.w4(32'h35f686d6),
	.w5(32'hb6acbf9b),
	.w6(32'hb807e866),
	.w7(32'hb6ae29ff),
	.w8(32'hb5d3b8a9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd5662),
	.w1(32'hb8a1be22),
	.w2(32'hb7c1f9a4),
	.w3(32'hb8a69c6e),
	.w4(32'hb7c7797d),
	.w5(32'h38700e6d),
	.w6(32'hb91d7b3f),
	.w7(32'hb9111f81),
	.w8(32'h38918360),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369b09e0),
	.w1(32'h3727ccad),
	.w2(32'h36f29e09),
	.w3(32'h36c7e4ae),
	.w4(32'hb665c19a),
	.w5(32'h3711f0ed),
	.w6(32'h36c9319d),
	.w7(32'hb721c9df),
	.w8(32'hb556aa84),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80844e0),
	.w1(32'hb6e5ab14),
	.w2(32'h38146646),
	.w3(32'hb78a8b65),
	.w4(32'hb630641d),
	.w5(32'h381053fa),
	.w6(32'h35814914),
	.w7(32'h3835ec68),
	.w8(32'h384182bd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b1aa7),
	.w1(32'h36227a7d),
	.w2(32'h3607613e),
	.w3(32'h37ac0da7),
	.w4(32'h37477f8b),
	.w5(32'hb73ba9d8),
	.w6(32'h378a8d26),
	.w7(32'h380a45d0),
	.w8(32'hb56d8d82),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a58b3e),
	.w1(32'h372c2dd1),
	.w2(32'hb72c9e69),
	.w3(32'hb5796791),
	.w4(32'hb6fb9348),
	.w5(32'hb7ce6e90),
	.w6(32'hb7beb1d6),
	.w7(32'h3690a18e),
	.w8(32'hb66d06c4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b5b84),
	.w1(32'hb8520fe1),
	.w2(32'h37eed349),
	.w3(32'h3876a10c),
	.w4(32'h38a3a658),
	.w5(32'h3878b727),
	.w6(32'h361e4517),
	.w7(32'hb8b98f92),
	.w8(32'h371041bb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977bff1),
	.w1(32'hb90dface),
	.w2(32'hb7212850),
	.w3(32'hb829dc00),
	.w4(32'h38a2a701),
	.w5(32'h38cebb9d),
	.w6(32'hba19d656),
	.w7(32'hb9c74984),
	.w8(32'hb842dbd2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf1393),
	.w1(32'h382b213f),
	.w2(32'hb74824ce),
	.w3(32'h37fb9c93),
	.w4(32'h3835430b),
	.w5(32'hb75a5baf),
	.w6(32'h383779f9),
	.w7(32'h3788bb47),
	.w8(32'h370747e5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f587a),
	.w1(32'hb90a490b),
	.w2(32'h388384e5),
	.w3(32'hb8bd6268),
	.w4(32'h36b330c1),
	.w5(32'h392e9416),
	.w6(32'hb9776b8b),
	.w7(32'hb982385a),
	.w8(32'h388f5528),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805489b),
	.w1(32'hb7a585c5),
	.w2(32'hb7062374),
	.w3(32'hb7c972ed),
	.w4(32'hb743aab2),
	.w5(32'hb5f6aa1f),
	.w6(32'hb88483fe),
	.w7(32'hb859a09f),
	.w8(32'hb7430b91),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b7f1c),
	.w1(32'hb964c3ec),
	.w2(32'hb8e274ae),
	.w3(32'hb93094a1),
	.w4(32'hb8d0e528),
	.w5(32'h3843e618),
	.w6(32'hb9e57fb2),
	.w7(32'hb9a47e84),
	.w8(32'hb79d3092),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957206b),
	.w1(32'hb8eec314),
	.w2(32'h37e47a2a),
	.w3(32'hb90ae75d),
	.w4(32'hb73d9af3),
	.w5(32'h38ca84da),
	.w6(32'hb9ac9eca),
	.w7(32'hb98dc1a6),
	.w8(32'hb6ad77cc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cf13b),
	.w1(32'hb918ace2),
	.w2(32'hb8a214d1),
	.w3(32'hb96042e8),
	.w4(32'hb8b162fe),
	.w5(32'hb71fe992),
	.w6(32'hb9f77df7),
	.w7(32'hb980fa75),
	.w8(32'hb8940c63),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3778419f),
	.w1(32'h37fa3901),
	.w2(32'h37b284e1),
	.w3(32'hb7b3e5c9),
	.w4(32'h37915c49),
	.w5(32'h35dd1fc6),
	.w6(32'hb778f232),
	.w7(32'h3784e7e8),
	.w8(32'h35a0c960),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904a7e0),
	.w1(32'hb8e1c7f3),
	.w2(32'hb862e2a3),
	.w3(32'hb8e9b320),
	.w4(32'hb85becb7),
	.w5(32'hb6c373e8),
	.w6(32'hb939662b),
	.w7(32'hb930d1c6),
	.w8(32'hb842bd2e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc90ad),
	.w1(32'h38483057),
	.w2(32'hb69eaaea),
	.w3(32'h379cf82a),
	.w4(32'h37836a76),
	.w5(32'hb767b0e5),
	.w6(32'h37c10364),
	.w7(32'h37297233),
	.w8(32'h379e501c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85bce7a),
	.w1(32'hb762b50d),
	.w2(32'h368eafb1),
	.w3(32'hb70eb33e),
	.w4(32'h36caf858),
	.w5(32'h380cb6b9),
	.w6(32'hb883c467),
	.w7(32'hb86aacfc),
	.w8(32'hb7689024),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb698342e),
	.w1(32'hb5e3d8c7),
	.w2(32'h36a63482),
	.w3(32'h3821f062),
	.w4(32'h3835d4c5),
	.w5(32'h37cff323),
	.w6(32'h37af97b4),
	.w7(32'hb720b18c),
	.w8(32'hb64f8fea),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90899e3),
	.w1(32'hb84b32c5),
	.w2(32'h37edb216),
	.w3(32'hb8b1354b),
	.w4(32'hb7ab3ab6),
	.w5(32'h387c2115),
	.w6(32'hb965d4c5),
	.w7(32'hb9229bd4),
	.w8(32'hb588f9f9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fa5a3f),
	.w1(32'hb7db6409),
	.w2(32'hb78b517e),
	.w3(32'h371cce46),
	.w4(32'hb754a300),
	.w5(32'hb70963d3),
	.w6(32'h349682fd),
	.w7(32'h35af7931),
	.w8(32'h37bca09b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7763300),
	.w1(32'hb7b573ee),
	.w2(32'h3807ad4d),
	.w3(32'h3799bf23),
	.w4(32'hb78ac6c0),
	.w5(32'hb6c1ba49),
	.w6(32'hb7765a81),
	.w7(32'h35a530a9),
	.w8(32'h37268eba),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83d028e),
	.w1(32'hb76cf5d6),
	.w2(32'h384c421e),
	.w3(32'hb6b7ce81),
	.w4(32'h3722bf8c),
	.w5(32'h385897f5),
	.w6(32'hb8e5de7d),
	.w7(32'hb80bf3f9),
	.w8(32'h3820df5b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9270332),
	.w1(32'hb8df2662),
	.w2(32'h385b19ab),
	.w3(32'hb87b64b5),
	.w4(32'hb6d148f8),
	.w5(32'h38ce932e),
	.w6(32'hb9ae1719),
	.w7(32'hb9793e10),
	.w8(32'h37c8fcfc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791ea24),
	.w1(32'h38716b63),
	.w2(32'h3743e815),
	.w3(32'hb786736c),
	.w4(32'h37ded915),
	.w5(32'h37bd0b4f),
	.w6(32'hb6c4f68a),
	.w7(32'h380a015b),
	.w8(32'hb71922e2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb724b29f),
	.w1(32'hb7f4d834),
	.w2(32'h38014a2c),
	.w3(32'h37c55246),
	.w4(32'h378c13a8),
	.w5(32'h38065df9),
	.w6(32'hb84d369e),
	.w7(32'hb7842464),
	.w8(32'h37a807d5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ec6e5),
	.w1(32'hb9835775),
	.w2(32'hb940a2af),
	.w3(32'hb9669fb6),
	.w4(32'hb960fd95),
	.w5(32'hb7ea0419),
	.w6(32'hba09efde),
	.w7(32'hb9c2570f),
	.w8(32'hb8263df7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945c7ba),
	.w1(32'hb9272078),
	.w2(32'h37ba2df1),
	.w3(32'hb816553d),
	.w4(32'h37bb8d94),
	.w5(32'h3915f920),
	.w6(32'hb9801ddc),
	.w7(32'hb9b92876),
	.w8(32'hb7911cee),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65a3f0e),
	.w1(32'h358c7491),
	.w2(32'hb77f06d4),
	.w3(32'hb6726026),
	.w4(32'hb5e5fd2f),
	.w5(32'hb79cf56e),
	.w6(32'h3799d7a8),
	.w7(32'h359c3464),
	.w8(32'hb77e81ad),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fa66c6),
	.w1(32'hb7cc2f66),
	.w2(32'h37b3eed3),
	.w3(32'h369aff6c),
	.w4(32'hb7b8f300),
	.w5(32'h37928c3d),
	.w6(32'h370a9ccd),
	.w7(32'hb72b1c11),
	.w8(32'h3785c647),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3507d978),
	.w1(32'hb799f802),
	.w2(32'hb7b74824),
	.w3(32'h370ea375),
	.w4(32'hb791497f),
	.w5(32'hb747b6a6),
	.w6(32'hb6adde96),
	.w7(32'h368a6f6f),
	.w8(32'hb70235fb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb688d3a1),
	.w1(32'hb6d724c0),
	.w2(32'hb7661a1f),
	.w3(32'hb6881eab),
	.w4(32'hb697cfbf),
	.w5(32'hb63ec439),
	.w6(32'h3682c8c0),
	.w7(32'hb6b87300),
	.w8(32'hb57808a9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8321e51),
	.w1(32'hb6c247e6),
	.w2(32'hb51954a4),
	.w3(32'hb76a2ae3),
	.w4(32'h374b4aed),
	.w5(32'h37966af8),
	.w6(32'hb7b96ef1),
	.w7(32'hb787d970),
	.w8(32'hb68161ed),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cfaa0f),
	.w1(32'hb8d88d7e),
	.w2(32'hb85909c6),
	.w3(32'h353a925b),
	.w4(32'h386ed30f),
	.w5(32'h37c7c5b4),
	.w6(32'hb92ebe46),
	.w7(32'hb90e73e0),
	.w8(32'hb88f0eda),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9116df4),
	.w1(32'hb8c86b65),
	.w2(32'h37859731),
	.w3(32'hb9017052),
	.w4(32'hb72e7463),
	.w5(32'h38c1323a),
	.w6(32'hb99eccc5),
	.w7(32'hb979d53b),
	.w8(32'h38239316),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6ed13),
	.w1(32'h378e3d0e),
	.w2(32'h380f3789),
	.w3(32'h3815054d),
	.w4(32'h3815bbd3),
	.w5(32'h382a148b),
	.w6(32'h3708d54f),
	.w7(32'hb6ac8d53),
	.w8(32'h370a5b5f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9410f36),
	.w1(32'hbbb29607),
	.w2(32'hbb3a4c58),
	.w3(32'hb8f63f5c),
	.w4(32'hbb335d12),
	.w5(32'h3b3d5f80),
	.w6(32'hb9c10cc2),
	.w7(32'hbb095443),
	.w8(32'hba78b784),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc3234),
	.w1(32'hbb0aadd7),
	.w2(32'h3b0efde4),
	.w3(32'hbbcb64c5),
	.w4(32'hbb325a1c),
	.w5(32'h3bb3428a),
	.w6(32'hbbc2499f),
	.w7(32'h3a5fa38b),
	.w8(32'h3bf168aa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6fbae),
	.w1(32'h3add75b3),
	.w2(32'hbb9c9707),
	.w3(32'hbb2aba76),
	.w4(32'hbb91b2d0),
	.w5(32'hbb394812),
	.w6(32'h3ad57bc8),
	.w7(32'hbbb9f0a4),
	.w8(32'h3b0383bc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e6a1),
	.w1(32'h3acfa071),
	.w2(32'hba2fe57c),
	.w3(32'h37939d40),
	.w4(32'hba3c4499),
	.w5(32'hb9ed26b2),
	.w6(32'hbbb03f0e),
	.w7(32'hbb4422a3),
	.w8(32'hbb388e0e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6bbb1),
	.w1(32'h3ad1e863),
	.w2(32'hb913666e),
	.w3(32'hbb96edc6),
	.w4(32'h3c084f08),
	.w5(32'hbafe5089),
	.w6(32'h3994f3cd),
	.w7(32'h3bea579d),
	.w8(32'hbbcaed90),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7ae4),
	.w1(32'hbb8f1a89),
	.w2(32'hbbd33260),
	.w3(32'hbb39fb61),
	.w4(32'hbbac6386),
	.w5(32'hbbd7836c),
	.w6(32'hbb69b152),
	.w7(32'hbc151056),
	.w8(32'hbbc5e3a5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18fb33),
	.w1(32'h3b4f716d),
	.w2(32'h3bc00e9d),
	.w3(32'hbbc68e3d),
	.w4(32'h3a000454),
	.w5(32'h3a700b64),
	.w6(32'h38d34fe6),
	.w7(32'h3b4ce129),
	.w8(32'h3b5781dc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9903e7d),
	.w1(32'hbb4be848),
	.w2(32'h3932684d),
	.w3(32'h3ab20125),
	.w4(32'h3a2a5bcf),
	.w5(32'h3af0dae4),
	.w6(32'h3af03a93),
	.w7(32'h3bbd5362),
	.w8(32'hbac9d36b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945ec9),
	.w1(32'hbb1d6b40),
	.w2(32'h3afbee5b),
	.w3(32'h3895d271),
	.w4(32'hbb005cd2),
	.w5(32'h39833dd9),
	.w6(32'hbb83f65e),
	.w7(32'hb9baac7c),
	.w8(32'h3bb63e48),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a3c9),
	.w1(32'hbb777321),
	.w2(32'h3a31d52f),
	.w3(32'h3b7ed8dc),
	.w4(32'hbab6e47e),
	.w5(32'h3c2b144d),
	.w6(32'h39e74e24),
	.w7(32'h3afc387b),
	.w8(32'h3c237cdf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f6cf),
	.w1(32'hbaa317cc),
	.w2(32'h3add5dfd),
	.w3(32'h3b58c65a),
	.w4(32'hbacfbf45),
	.w5(32'hbabf3ea3),
	.w6(32'h3b82fded),
	.w7(32'h3b954ff0),
	.w8(32'hbac276d9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31eaeb),
	.w1(32'h3a8a6614),
	.w2(32'hbb017bc5),
	.w3(32'h3ac0ae6b),
	.w4(32'h38b950ef),
	.w5(32'h3a61f9c8),
	.w6(32'hb9f3ce4a),
	.w7(32'h39b5b11d),
	.w8(32'hba994217),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad55ca7),
	.w1(32'hb980d2a1),
	.w2(32'h3b0f5801),
	.w3(32'h3a86b4aa),
	.w4(32'hba2892b3),
	.w5(32'h3a3a350e),
	.w6(32'h37824ea7),
	.w7(32'hb9183f41),
	.w8(32'hb9cbc0a2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07a197),
	.w1(32'h3a82e5ea),
	.w2(32'h3adc8b92),
	.w3(32'hbab5771f),
	.w4(32'hbb93ab59),
	.w5(32'h3b580254),
	.w6(32'hba498258),
	.w7(32'hbbcc7486),
	.w8(32'h3b8d10d0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44ac9c),
	.w1(32'h3b5333d5),
	.w2(32'hbc1281e9),
	.w3(32'h3b92399c),
	.w4(32'h3b02ee2a),
	.w5(32'hbb201c89),
	.w6(32'h38d3be28),
	.w7(32'h39fbbdb5),
	.w8(32'hbb81fbac),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fa9ca),
	.w1(32'h3bc03ad2),
	.w2(32'hb812a28a),
	.w3(32'hbbaccd68),
	.w4(32'h3b086bb6),
	.w5(32'hbbc20661),
	.w6(32'h3a814462),
	.w7(32'hbb49ad93),
	.w8(32'hbb34d45a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ae5e4),
	.w1(32'hbb304fb5),
	.w2(32'h3b19a7dd),
	.w3(32'hba98a3f1),
	.w4(32'h3b55c68b),
	.w5(32'h3989bc52),
	.w6(32'hbaffd66c),
	.w7(32'h3a6ca383),
	.w8(32'hbae231cc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cee42),
	.w1(32'hbb993811),
	.w2(32'hbbcace62),
	.w3(32'h3aceaf23),
	.w4(32'hb927fd9a),
	.w5(32'hbbe12767),
	.w6(32'h3aadafb8),
	.w7(32'h3bcf932e),
	.w8(32'h3c03b587),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb283daf),
	.w1(32'hbb22f6f6),
	.w2(32'hbb9f5957),
	.w3(32'h3b249d33),
	.w4(32'h3bfaaf32),
	.w5(32'hbb93967e),
	.w6(32'h3b109139),
	.w7(32'h3c172373),
	.w8(32'hba880cae),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae77db),
	.w1(32'h3acb23c9),
	.w2(32'hba40a8a9),
	.w3(32'h3a936805),
	.w4(32'h3a5e6c9a),
	.w5(32'hbacc4f3b),
	.w6(32'h3bb8d7e9),
	.w7(32'h3b6a3968),
	.w8(32'hbb5c120c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2834),
	.w1(32'hbaf9f270),
	.w2(32'h395d6568),
	.w3(32'hbb65a076),
	.w4(32'h39ec567b),
	.w5(32'hbb3550d3),
	.w6(32'h3b34c1ec),
	.w7(32'h3aa8b534),
	.w8(32'hbb1e8912),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f21d0),
	.w1(32'hbbcf2b22),
	.w2(32'h38b0bdca),
	.w3(32'hbb161078),
	.w4(32'hbb6f4147),
	.w5(32'h3ae680e2),
	.w6(32'h3a39c5ca),
	.w7(32'hbb01838d),
	.w8(32'hbb33f42f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ac240),
	.w1(32'hbaed6992),
	.w2(32'hbb0d6700),
	.w3(32'hbbb09e12),
	.w4(32'h3af8d7b3),
	.w5(32'hba167ad8),
	.w6(32'hbb97b110),
	.w7(32'h3b0b8973),
	.w8(32'hba2910af),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951e787),
	.w1(32'hba19056b),
	.w2(32'hba3b2140),
	.w3(32'h3b861995),
	.w4(32'hbbb9a209),
	.w5(32'h3ab4143c),
	.w6(32'h3aee518d),
	.w7(32'hbba00862),
	.w8(32'hbaf5231f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdde03d),
	.w1(32'hb88b1889),
	.w2(32'hbb4ae66e),
	.w3(32'h3b6e9262),
	.w4(32'h3ac1734d),
	.w5(32'hbadeda9a),
	.w6(32'h3ac1175f),
	.w7(32'h3b4cc04f),
	.w8(32'hbb3f7408),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f24f5),
	.w1(32'h3b258cd0),
	.w2(32'h3b2492c3),
	.w3(32'hba8f9a73),
	.w4(32'h3ab7a8d3),
	.w5(32'h38b45ab4),
	.w6(32'h399f6d0b),
	.w7(32'h3c3bf014),
	.w8(32'h3bbfb007),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fc6e0),
	.w1(32'hba242e84),
	.w2(32'h3b4719ab),
	.w3(32'h3b341c71),
	.w4(32'h3b99db7c),
	.w5(32'hbb74fe1c),
	.w6(32'h3c128244),
	.w7(32'h3bc9e748),
	.w8(32'hbbf1fe67),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdb698),
	.w1(32'h3aef0b88),
	.w2(32'h3c1ad147),
	.w3(32'hba2a1941),
	.w4(32'h3c3f69ce),
	.w5(32'h3b8702b3),
	.w6(32'hbb685fba),
	.w7(32'h3bd4a76f),
	.w8(32'hbbc8f996),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64f9d),
	.w1(32'hbba1787c),
	.w2(32'hbb22c1d2),
	.w3(32'hbb2f2b30),
	.w4(32'hbb1aaa82),
	.w5(32'hbbbe4419),
	.w6(32'h3b0f7a39),
	.w7(32'hbb9d9966),
	.w8(32'hbaf1c037),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ce65),
	.w1(32'hbaafb603),
	.w2(32'h3abf703f),
	.w3(32'hbac78e49),
	.w4(32'hbb4e4599),
	.w5(32'hba45dde0),
	.w6(32'hbac21ef3),
	.w7(32'hbaa8bc07),
	.w8(32'hbaf81b23),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305e96),
	.w1(32'h3b599dd9),
	.w2(32'hbac19c5f),
	.w3(32'hbb56aade),
	.w4(32'hbb3326a0),
	.w5(32'hbb8793c8),
	.w6(32'hb9d1ec8a),
	.w7(32'h3a9085f2),
	.w8(32'h3be27874),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76ea79),
	.w1(32'hbb77affe),
	.w2(32'hbb216ccc),
	.w3(32'hba7bc782),
	.w4(32'h3bad90e5),
	.w5(32'hb9ebd071),
	.w6(32'h3b088078),
	.w7(32'h3c01359d),
	.w8(32'hbaa2afa6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf7fab),
	.w1(32'h3bc1ffe3),
	.w2(32'h3bf2548b),
	.w3(32'hb935ca3a),
	.w4(32'h3b50b78b),
	.w5(32'hbb150189),
	.w6(32'h3aa90adf),
	.w7(32'hbb391b49),
	.w8(32'hbb554ab2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a211fa4),
	.w1(32'h3b9397cb),
	.w2(32'h3b1daf4d),
	.w3(32'hb9b7d691),
	.w4(32'hba566ea4),
	.w5(32'hbb112771),
	.w6(32'h3b2a81d5),
	.w7(32'hba45200f),
	.w8(32'h3a97117b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37160a),
	.w1(32'h3b870197),
	.w2(32'h3a043195),
	.w3(32'h3bea8b0e),
	.w4(32'h3b9ec9d0),
	.w5(32'hbb3672df),
	.w6(32'h3b84202c),
	.w7(32'h3b54cde8),
	.w8(32'h3a68171f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867250),
	.w1(32'hba25a469),
	.w2(32'h3ab7c432),
	.w3(32'h3b486c78),
	.w4(32'hbb78365c),
	.w5(32'h3be7ed82),
	.w6(32'h3b98b505),
	.w7(32'hbbf2b0d1),
	.w8(32'h3b72adf5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519d3a),
	.w1(32'hbb3800fd),
	.w2(32'h393f4d5a),
	.w3(32'h3b9fdd6a),
	.w4(32'hbb47cccf),
	.w5(32'hbb58760b),
	.w6(32'h3b2232e9),
	.w7(32'hba229fe1),
	.w8(32'hbb86b8e0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac8a1),
	.w1(32'hbb7e9f68),
	.w2(32'h3b2ad9be),
	.w3(32'hbbb5024a),
	.w4(32'hbb5085f0),
	.w5(32'h3bb4222d),
	.w6(32'hbb47c89f),
	.w7(32'hbb0a15e6),
	.w8(32'h3be80c0f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6c37),
	.w1(32'hbaa095ee),
	.w2(32'hbaf012dd),
	.w3(32'h3b6027f8),
	.w4(32'h39d51c37),
	.w5(32'hb936c612),
	.w6(32'h3a6b07f3),
	.w7(32'hbb7dde9a),
	.w8(32'h3a6d3d0b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e3f76),
	.w1(32'h3abb1c77),
	.w2(32'hbb854026),
	.w3(32'h39d9bd5d),
	.w4(32'h396d546c),
	.w5(32'hbbae151d),
	.w6(32'h3bfc943a),
	.w7(32'hbbb4c12f),
	.w8(32'hbb1e6b2a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b96541),
	.w1(32'h3a686a05),
	.w2(32'h3b858329),
	.w3(32'h3b6f78cc),
	.w4(32'hbb045d1c),
	.w5(32'hbb258d91),
	.w6(32'h3b95c1f4),
	.w7(32'hbbc53100),
	.w8(32'hbbac9101),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29b635),
	.w1(32'h3b45898d),
	.w2(32'h3ad5dcc3),
	.w3(32'h3b530118),
	.w4(32'h3b4b4f27),
	.w5(32'hbb2ae84a),
	.w6(32'hba84e5b1),
	.w7(32'hbb63dad1),
	.w8(32'hbbbf9d82),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44aced),
	.w1(32'hb99b0f37),
	.w2(32'h3ba8f4bc),
	.w3(32'h3b0e26d9),
	.w4(32'hba521092),
	.w5(32'hb8db8519),
	.w6(32'h39a5452a),
	.w7(32'hbacd510e),
	.w8(32'hbb485613),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2699d1),
	.w1(32'h399b8645),
	.w2(32'hb9bab3b3),
	.w3(32'hbb0bb52b),
	.w4(32'h3b51511d),
	.w5(32'hbb3f621a),
	.w6(32'h3a901ccf),
	.w7(32'h390ce3ed),
	.w8(32'hbbeda89f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f75a),
	.w1(32'hbb13cf19),
	.w2(32'h3abcdb79),
	.w3(32'hbafc6c36),
	.w4(32'h39776477),
	.w5(32'hb9512c1d),
	.w6(32'h3a19b284),
	.w7(32'h3b34979e),
	.w8(32'hbb7ec219),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaf7a2),
	.w1(32'hbb8e2d4a),
	.w2(32'hbbc4b567),
	.w3(32'h3baf9709),
	.w4(32'hbbc3baa7),
	.w5(32'h3b0f338b),
	.w6(32'h3b0f3391),
	.w7(32'hbb7f7190),
	.w8(32'h3bc22d4a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43f82),
	.w1(32'h3941e179),
	.w2(32'hba8adf9b),
	.w3(32'hb931bfc3),
	.w4(32'h39ab1f35),
	.w5(32'h3b3c9230),
	.w6(32'hb92b73e3),
	.w7(32'h3ab29a23),
	.w8(32'h3ae0476d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb498f56),
	.w1(32'hbb0fafae),
	.w2(32'hbb357266),
	.w3(32'hbbdbcc65),
	.w4(32'hbad6d8a7),
	.w5(32'h3ac8c039),
	.w6(32'hbb19952e),
	.w7(32'hbb1b61e0),
	.w8(32'hb9e52640),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf1c6),
	.w1(32'hbb6f1ec4),
	.w2(32'hbb5c02a4),
	.w3(32'hbb5814fb),
	.w4(32'hbc1266b6),
	.w5(32'hbb0ffb3c),
	.w6(32'hbae37e19),
	.w7(32'hbbe265b8),
	.w8(32'hbb06b813),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11363b),
	.w1(32'h3b7ec16d),
	.w2(32'h3b3b7b7f),
	.w3(32'h3b181f45),
	.w4(32'h3c213b07),
	.w5(32'h39bd28f6),
	.w6(32'hbb1244f4),
	.w7(32'h3b97bd21),
	.w8(32'hbb3cadc7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b1ea0),
	.w1(32'hb90fdb9d),
	.w2(32'hbbabda7a),
	.w3(32'h3b4735d6),
	.w4(32'hbb1cc15a),
	.w5(32'hbb963043),
	.w6(32'h3ad61af6),
	.w7(32'hbb7aa616),
	.w8(32'h3a79b18c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5cc2b),
	.w1(32'h3a396537),
	.w2(32'hbb10b1a5),
	.w3(32'h3bcb0cbe),
	.w4(32'h39e0e66b),
	.w5(32'h3b3bdc0d),
	.w6(32'h3b096707),
	.w7(32'h3b1d41d5),
	.w8(32'h3a553a6d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc7126),
	.w1(32'hbac3edaa),
	.w2(32'hbb7a3e64),
	.w3(32'hbac46291),
	.w4(32'hbb0c9fae),
	.w5(32'hb999b426),
	.w6(32'hbbb30387),
	.w7(32'hbb090843),
	.w8(32'h3b0e3073),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cc50f),
	.w1(32'h3a5d9392),
	.w2(32'h3adf5a59),
	.w3(32'hbb3daeaa),
	.w4(32'h3bdf27e4),
	.w5(32'h3b27d091),
	.w6(32'h3b4c8fa9),
	.w7(32'h3b319ce8),
	.w8(32'h3a04fad7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacdd94),
	.w1(32'h3bf089b8),
	.w2(32'h3ba00ff0),
	.w3(32'hbac0b4f1),
	.w4(32'h3c232576),
	.w5(32'hbbce3ae6),
	.w6(32'h3a94bf25),
	.w7(32'h3b1e1837),
	.w8(32'hbc1a9d3a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b66de),
	.w1(32'h3c01a40f),
	.w2(32'hbb023d31),
	.w3(32'hbc035b15),
	.w4(32'hbb6e26ab),
	.w5(32'hbc08878a),
	.w6(32'hbad616c3),
	.w7(32'hbb914c7d),
	.w8(32'hba84e549),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b535162),
	.w1(32'hb8c7c8cb),
	.w2(32'hbb1893f3),
	.w3(32'h3aa52ee4),
	.w4(32'hbba73b10),
	.w5(32'h3b56be79),
	.w6(32'h3aeeee7e),
	.w7(32'hbb1e0fc8),
	.w8(32'h3b3f8f6f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cf848),
	.w1(32'hbbb54a70),
	.w2(32'hbbe2eaa9),
	.w3(32'h3b433780),
	.w4(32'hbc2b897e),
	.w5(32'hbc01217a),
	.w6(32'hb925323d),
	.w7(32'hbbed0b47),
	.w8(32'hbbc2fb93),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96724d),
	.w1(32'hbb0fc5fb),
	.w2(32'hbb7e7b8a),
	.w3(32'hbbb7abdb),
	.w4(32'hbb284efa),
	.w5(32'hba8b13be),
	.w6(32'hbb8efebc),
	.w7(32'hbb337b62),
	.w8(32'hba823729),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule