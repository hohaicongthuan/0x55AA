module layer_10_featuremap_438(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c813be),
	.w1(32'h36fb7c6d),
	.w2(32'h3733ec03),
	.w3(32'h37c625e2),
	.w4(32'h36ac993b),
	.w5(32'h36edc3c7),
	.w6(32'h37dee79b),
	.w7(32'h378088c3),
	.w8(32'h3734a471),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a7006),
	.w1(32'h3b1e03a3),
	.w2(32'h3b0b34a0),
	.w3(32'h39a7cffb),
	.w4(32'h3b0357d8),
	.w5(32'h3a3e0197),
	.w6(32'h394cce8d),
	.w7(32'h3a8ec237),
	.w8(32'h3abcb546),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3777c149),
	.w1(32'h3748081d),
	.w2(32'h37634060),
	.w3(32'h374ed312),
	.w4(32'h371f90ac),
	.w5(32'h373e5d1d),
	.w6(32'h374a1c9f),
	.w7(32'h3717d736),
	.w8(32'h377002f5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f3322),
	.w1(32'h3a7ba381),
	.w2(32'h391409ae),
	.w3(32'h3a31b2af),
	.w4(32'h3a7d9d1a),
	.w5(32'h39da4be2),
	.w6(32'h3a2a54a5),
	.w7(32'h3a8792fa),
	.w8(32'h397a104d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e53bf0),
	.w1(32'h39add1b7),
	.w2(32'hb94a7317),
	.w3(32'h39d6b3fa),
	.w4(32'h39a9ff36),
	.w5(32'hb8735970),
	.w6(32'h39dccfe2),
	.w7(32'h39e27855),
	.w8(32'h389b4209),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ab7019),
	.w1(32'h377cc4c4),
	.w2(32'h378da0b9),
	.w3(32'h37c009b4),
	.w4(32'h378b37c3),
	.w5(32'h375d0e1b),
	.w6(32'h37b8921a),
	.w7(32'h37b5afb0),
	.w8(32'h37d788dc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b212fc3),
	.w1(32'h38e2cc91),
	.w2(32'hbac22bc0),
	.w3(32'h3b4ced0f),
	.w4(32'h3a459b1a),
	.w5(32'hbac0f55f),
	.w6(32'h3b04d374),
	.w7(32'hb9ceaa41),
	.w8(32'hbb5fdb1e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97f35a),
	.w1(32'hbb31c44b),
	.w2(32'hbbe618f6),
	.w3(32'hbb8bd7c0),
	.w4(32'hbbc761d2),
	.w5(32'hbb97fd94),
	.w6(32'hbb0c4be9),
	.w7(32'hbbba495e),
	.w8(32'hbbce12ab),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e88192),
	.w1(32'h3759e802),
	.w2(32'hb947b388),
	.w3(32'h3a2707de),
	.w4(32'h3976c29c),
	.w5(32'hb992c501),
	.w6(32'h3a33be68),
	.w7(32'h375fa291),
	.w8(32'hba0fac41),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845318),
	.w1(32'hbacaf7f2),
	.w2(32'h3b3376d0),
	.w3(32'h390df438),
	.w4(32'hba6786b3),
	.w5(32'h39907b2d),
	.w6(32'h3a0b27cd),
	.w7(32'hba81ce93),
	.w8(32'hbaeba298),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921ad2a),
	.w1(32'hb9e2ce47),
	.w2(32'hba2965ba),
	.w3(32'hb9486e17),
	.w4(32'hb98d4b1a),
	.w5(32'hb9b88118),
	.w6(32'h3906905c),
	.w7(32'hb92764dd),
	.w8(32'hb9023fc2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e8890),
	.w1(32'h3acf4ac4),
	.w2(32'hbb3af74a),
	.w3(32'h3b30ba65),
	.w4(32'h3b1b55e1),
	.w5(32'hba15930b),
	.w6(32'h3ac54707),
	.w7(32'h3a342b42),
	.w8(32'hbb89cad4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca6878),
	.w1(32'hbaa39aa5),
	.w2(32'h3889a4ae),
	.w3(32'h3a96c209),
	.w4(32'hbaab91b3),
	.w5(32'hbaa07bb1),
	.w6(32'h3b485292),
	.w7(32'hb990970d),
	.w8(32'hbb222be3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31374f),
	.w1(32'h39a3c3ab),
	.w2(32'hba8aa180),
	.w3(32'hb85e4bba),
	.w4(32'hba02b2be),
	.w5(32'hba5cabe8),
	.w6(32'hb9edfb0c),
	.w7(32'hba7c167c),
	.w8(32'hba4019c9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05dcd4),
	.w1(32'hb947e37f),
	.w2(32'hb863b565),
	.w3(32'h398d7700),
	.w4(32'h3a82d39a),
	.w5(32'hb9fdf728),
	.w6(32'h3a58641e),
	.w7(32'h399e9421),
	.w8(32'hb93a7ee3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9986bb1),
	.w1(32'hb8d9daf5),
	.w2(32'h3a9f930a),
	.w3(32'hba6a02b3),
	.w4(32'hb9e88c19),
	.w5(32'hb982026e),
	.w6(32'hbadfca0a),
	.w7(32'hbb1e8dbc),
	.w8(32'hbaa5bff9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39222721),
	.w1(32'h3932f157),
	.w2(32'h392fdb5d),
	.w3(32'h3697248c),
	.w4(32'h393421ff),
	.w5(32'h391b9106),
	.w6(32'h37dd2406),
	.w7(32'h390743a0),
	.w8(32'h393f1158),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0974ad),
	.w1(32'hbc28b55a),
	.w2(32'hbc3d215e),
	.w3(32'hbbeaef2f),
	.w4(32'hbc11f660),
	.w5(32'hbc06e316),
	.w6(32'hbbc86deb),
	.w7(32'hbc3803d0),
	.w8(32'hbc4ec1f1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3841fc02),
	.w1(32'hbb86488c),
	.w2(32'hbb6e3456),
	.w3(32'hbabed054),
	.w4(32'hbb545820),
	.w5(32'hbb076295),
	.w6(32'hbad9d2f7),
	.w7(32'hbb75ed8c),
	.w8(32'hbb9245b7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e4ab7),
	.w1(32'h3833a142),
	.w2(32'h385baff8),
	.w3(32'h38299300),
	.w4(32'h38800df3),
	.w5(32'h37cddbdb),
	.w6(32'h37f66378),
	.w7(32'h380d1f66),
	.w8(32'hb7e013ac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d3511),
	.w1(32'hb87da53e),
	.w2(32'hb6dde8c3),
	.w3(32'h3861d6c1),
	.w4(32'hb88a1ee4),
	.w5(32'hb59fca6a),
	.w6(32'h38745c4a),
	.w7(32'hb783c654),
	.w8(32'h38e5d2ff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf338e),
	.w1(32'h3ae622a0),
	.w2(32'h38e8cffc),
	.w3(32'h3b04380d),
	.w4(32'h3b0e2d15),
	.w5(32'h3a2d30f5),
	.w6(32'h3ac38d37),
	.w7(32'h3af11ab8),
	.w8(32'h3a2bd41f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c4448),
	.w1(32'hbc3d705c),
	.w2(32'hbc49f091),
	.w3(32'hbbb68dd9),
	.w4(32'hbbdf0a7c),
	.w5(32'hbc123fdd),
	.w6(32'hbc23506f),
	.w7(32'hbb9b679f),
	.w8(32'hbc612bf4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0477b9),
	.w1(32'hba1de275),
	.w2(32'h3b91883c),
	.w3(32'hb9af02ad),
	.w4(32'h38d23fc8),
	.w5(32'h3abb988b),
	.w6(32'hb9e9fb45),
	.w7(32'h39cd2063),
	.w8(32'h3a72fb66),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b5d73),
	.w1(32'h3ab6a8e8),
	.w2(32'h3ba7e59b),
	.w3(32'hba5dd859),
	.w4(32'h3b959733),
	.w5(32'h3af70487),
	.w6(32'hba8a5138),
	.w7(32'h3b17613c),
	.w8(32'h3ade40fd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915a8db),
	.w1(32'h395f4a77),
	.w2(32'h38345a44),
	.w3(32'h391ee14e),
	.w4(32'h382e22d7),
	.w5(32'hb943ef44),
	.w6(32'h399d701a),
	.w7(32'hb66fe561),
	.w8(32'hb99c6fd4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383dc85d),
	.w1(32'h38998950),
	.w2(32'h38bb8412),
	.w3(32'h384fcfca),
	.w4(32'h386166ec),
	.w5(32'h383a266b),
	.w6(32'h3856f701),
	.w7(32'h389012bf),
	.w8(32'h38ec137f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990038f),
	.w1(32'h3b07dbcc),
	.w2(32'hba150b89),
	.w3(32'h3ad0a2e6),
	.w4(32'h3b8bd7a2),
	.w5(32'h3a6c0a2a),
	.w6(32'h3b08366f),
	.w7(32'h3acadf29),
	.w8(32'h39cc573b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508dcd),
	.w1(32'h3aa901f0),
	.w2(32'h3a294ad0),
	.w3(32'h3a140532),
	.w4(32'h3a978489),
	.w5(32'h3a4707af),
	.w6(32'h3969c961),
	.w7(32'h3987127e),
	.w8(32'h39bed6f6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36662e),
	.w1(32'h3b3879c7),
	.w2(32'h3b974a41),
	.w3(32'h3b3082f3),
	.w4(32'h3b7e154d),
	.w5(32'h3b30b59e),
	.w6(32'h3b6e400d),
	.w7(32'h3b647359),
	.w8(32'h3b326c15),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38001a2a),
	.w1(32'h37ea26e3),
	.w2(32'h3826419a),
	.w3(32'h37b43db1),
	.w4(32'h37b4333e),
	.w5(32'h37e6d018),
	.w6(32'h37b2646b),
	.w7(32'h37830c7f),
	.w8(32'h37c61fe7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377d1c5e),
	.w1(32'h37a7053a),
	.w2(32'h38813686),
	.w3(32'hb5c9365b),
	.w4(32'h37030a65),
	.w5(32'h38623504),
	.w6(32'h375e8da7),
	.w7(32'h37fed52a),
	.w8(32'h389c117f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31868c),
	.w1(32'hbaaf2a20),
	.w2(32'hba49029f),
	.w3(32'hba2cf7ff),
	.w4(32'hbab49670),
	.w5(32'hbaa70cff),
	.w6(32'hba2d8e56),
	.w7(32'hbac0ddb6),
	.w8(32'hbae9874f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df11a),
	.w1(32'h3aa68be5),
	.w2(32'h3aaf423f),
	.w3(32'h398cb0b6),
	.w4(32'h3a4ce486),
	.w5(32'h39ef9698),
	.w6(32'h38d9e829),
	.w7(32'h3a274a46),
	.w8(32'h39f489ea),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eda7d0),
	.w1(32'hb8930dec),
	.w2(32'hb894c11d),
	.w3(32'h392f396e),
	.w4(32'h393f2e52),
	.w5(32'h392aa058),
	.w6(32'hb692083d),
	.w7(32'hb9b3334d),
	.w8(32'hb994c4c5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a945e),
	.w1(32'hb980475a),
	.w2(32'hb9e3df5b),
	.w3(32'hb8653a5e),
	.w4(32'hba34f1a7),
	.w5(32'hba5741db),
	.w6(32'hb89ccd52),
	.w7(32'h3a015937),
	.w8(32'hbafd4387),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018a56),
	.w1(32'h3b2e5621),
	.w2(32'hbb1ea33f),
	.w3(32'h3b5375a1),
	.w4(32'hba072e8c),
	.w5(32'h3b6f89ca),
	.w6(32'h3ab7236a),
	.w7(32'h3b22cb5d),
	.w8(32'hba3d3605),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae627f1),
	.w1(32'h3c2aa084),
	.w2(32'h3bdc5d6a),
	.w3(32'h3bfa8536),
	.w4(32'h3c525c3d),
	.w5(32'h3bc0d509),
	.w6(32'h3b424f11),
	.w7(32'h3bead024),
	.w8(32'h3beae83d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb03b),
	.w1(32'h3c0cf220),
	.w2(32'h3b5d052f),
	.w3(32'h3ba7bf7a),
	.w4(32'h3c1c1325),
	.w5(32'h3b38790a),
	.w6(32'h3b9b5c22),
	.w7(32'h3bc4200a),
	.w8(32'h3b92c5eb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1be9e5),
	.w1(32'h3aeac899),
	.w2(32'h3aa05e2a),
	.w3(32'h3b13a309),
	.w4(32'h3b1659c4),
	.w5(32'h3ab4d14b),
	.w6(32'h3abd787c),
	.w7(32'h3aff7173),
	.w8(32'h3acec55c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38780d3b),
	.w1(32'h35fcf751),
	.w2(32'h384f8edc),
	.w3(32'h37fc9905),
	.w4(32'hb8081ae4),
	.w5(32'h37f92412),
	.w6(32'h38435dec),
	.w7(32'hb708fb54),
	.w8(32'h3808f35b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2c9c4),
	.w1(32'h39240704),
	.w2(32'h3954c3e6),
	.w3(32'h390341af),
	.w4(32'h3933e9f4),
	.w5(32'h395a2a9e),
	.w6(32'h38e0a642),
	.w7(32'h38db0b29),
	.w8(32'h397380a2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30aefb),
	.w1(32'h39c7f391),
	.w2(32'hbaa30afb),
	.w3(32'hba07ba25),
	.w4(32'h387fcfaa),
	.w5(32'hba3767d3),
	.w6(32'hba03b2d8),
	.w7(32'hba1dfd45),
	.w8(32'hba9a2d3d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cdfd5),
	.w1(32'hbad29df6),
	.w2(32'h3a1364fd),
	.w3(32'hbb083792),
	.w4(32'hbaf313fe),
	.w5(32'hba942075),
	.w6(32'hbaa984d9),
	.w7(32'hbb7eed91),
	.w8(32'hbb538cb1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e6ff1),
	.w1(32'hba154561),
	.w2(32'h3b060391),
	.w3(32'hba83972b),
	.w4(32'h3a538550),
	.w5(32'h39c3ac2c),
	.w6(32'hb908bc81),
	.w7(32'h3a70fc38),
	.w8(32'h39b64947),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb447cd2),
	.w1(32'hba2f03ef),
	.w2(32'h3b92b831),
	.w3(32'hba0e89a8),
	.w4(32'hb947cb35),
	.w5(32'h3a9d7b22),
	.w6(32'hba870a87),
	.w7(32'h3a167f78),
	.w8(32'h3a866132),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15315),
	.w1(32'h39858387),
	.w2(32'h38043cbe),
	.w3(32'hba18fa38),
	.w4(32'hb819e027),
	.w5(32'h39b27cd8),
	.w6(32'hbb3bf987),
	.w7(32'hbae3abc3),
	.w8(32'hbaef82a0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21d6aa),
	.w1(32'hbbd1a004),
	.w2(32'hbc46ab5e),
	.w3(32'hbb47e3df),
	.w4(32'hbbc86d54),
	.w5(32'hbbc2114d),
	.w6(32'hbb80f200),
	.w7(32'hbbc7685e),
	.w8(32'hbc2db375),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b7b2d),
	.w1(32'h36caa8cf),
	.w2(32'h3735fea5),
	.w3(32'h38b30454),
	.w4(32'hb639ef81),
	.w5(32'h3824a09d),
	.w6(32'h38ee9cc5),
	.w7(32'h3799dc4e),
	.w8(32'h381290e1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996ee32),
	.w1(32'hb910b17e),
	.w2(32'h3a0ca00e),
	.w3(32'h3990a853),
	.w4(32'h38c66afc),
	.w5(32'h3a27a370),
	.w6(32'h39a79437),
	.w7(32'hb89d24a1),
	.w8(32'hb8fc9008),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acf290),
	.w1(32'hb8c185d9),
	.w2(32'hb5bbc59d),
	.w3(32'h37e4d622),
	.w4(32'hb819c742),
	.w5(32'hb80fff0c),
	.w6(32'h38893b69),
	.w7(32'hb8170664),
	.w8(32'hb854693e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd6ab7),
	.w1(32'hbb069d7e),
	.w2(32'hba925a60),
	.w3(32'hba8909b8),
	.w4(32'hb9e35247),
	.w5(32'hba8bf3a5),
	.w6(32'hbac35d48),
	.w7(32'hba984b69),
	.w8(32'hbaeb037e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c929e6),
	.w1(32'hba46a532),
	.w2(32'hbaa89a90),
	.w3(32'hba85e5a9),
	.w4(32'hbaabd33e),
	.w5(32'hba7478a1),
	.w6(32'hba91f0e2),
	.w7(32'hba91525f),
	.w8(32'hbab8109b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27ea0b),
	.w1(32'hbbe1be31),
	.w2(32'hbbd0ceb6),
	.w3(32'hbbae926d),
	.w4(32'hbbeda238),
	.w5(32'hbb952966),
	.w6(32'hbb9746fd),
	.w7(32'hbc002ebb),
	.w8(32'hbc1fc4e6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ee088),
	.w1(32'hb93d77d2),
	.w2(32'hbaa95950),
	.w3(32'hb9cd481d),
	.w4(32'hb900f652),
	.w5(32'hba4603b5),
	.w6(32'hb907ca4c),
	.w7(32'hb9181459),
	.w8(32'hba9d2b7e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f44686),
	.w1(32'h388d1279),
	.w2(32'h36f67d56),
	.w3(32'h394888ac),
	.w4(32'h38f0eca0),
	.w5(32'h37df3248),
	.w6(32'h388f04b0),
	.w7(32'hb804fce2),
	.w8(32'hb8990508),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c3c83),
	.w1(32'hb7401e83),
	.w2(32'h3744c67b),
	.w3(32'h3738321a),
	.w4(32'hb59eebc9),
	.w5(32'h3790a49b),
	.w6(32'h37c6f15f),
	.w7(32'h375d09eb),
	.w8(32'h37cb1d7e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f875c8),
	.w1(32'hb97bf5a7),
	.w2(32'hb74d96f2),
	.w3(32'h3903a760),
	.w4(32'hb834d934),
	.w5(32'hb80ceb05),
	.w6(32'h393742f4),
	.w7(32'hb756d9fa),
	.w8(32'h391c09ba),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a066528),
	.w1(32'h3a2ec71a),
	.w2(32'hb920bd36),
	.w3(32'h3a27c82f),
	.w4(32'h3a680d4d),
	.w5(32'h3930deb2),
	.w6(32'h398a2c3a),
	.w7(32'h3a0ba7d3),
	.w8(32'hb8d08fc8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b09724),
	.w1(32'hb7f8be77),
	.w2(32'hb8c03fed),
	.w3(32'hb92e6544),
	.w4(32'hb87c8fb9),
	.w5(32'hb90e5b56),
	.w6(32'h38f14fac),
	.w7(32'hb95e9fcf),
	.w8(32'hb9333dc6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba748d9a),
	.w1(32'hbb5ecd9f),
	.w2(32'hbb765aac),
	.w3(32'hbb49d949),
	.w4(32'hbb2b0959),
	.w5(32'hbb19eb57),
	.w6(32'hbacb4288),
	.w7(32'hbb370276),
	.w8(32'hbb88a9b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a14c5),
	.w1(32'hbba436c0),
	.w2(32'hbb1b7ebf),
	.w3(32'hbbad33a2),
	.w4(32'hbb3e5a4c),
	.w5(32'hbb830b0a),
	.w6(32'hbb751825),
	.w7(32'hbb863514),
	.w8(32'hbb953e84),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ea1e34),
	.w1(32'h37df1ce7),
	.w2(32'h38acd9ab),
	.w3(32'hb8724c0a),
	.w4(32'h378c8d36),
	.w5(32'h3898b05a),
	.w6(32'hb78465da),
	.w7(32'h375d6cf9),
	.w8(32'h38941310),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59a3240),
	.w1(32'hb7214dee),
	.w2(32'h37eb443b),
	.w3(32'hb68fecbb),
	.w4(32'hb72b0ae2),
	.w5(32'h3799c2ab),
	.w6(32'h378af60d),
	.w7(32'h361b9f4c),
	.w8(32'h37e9f79e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382fe09e),
	.w1(32'h382aaf85),
	.w2(32'h37bbc52d),
	.w3(32'h38258dc5),
	.w4(32'h381783de),
	.w5(32'h3780190b),
	.w6(32'h3809bcb1),
	.w7(32'h37f1e1a0),
	.w8(32'h37d0c58a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c89af8),
	.w1(32'h378e2ef2),
	.w2(32'h38443999),
	.w3(32'h36e5a6e5),
	.w4(32'h36c76a57),
	.w5(32'h37b6aea5),
	.w6(32'h37b3c09a),
	.w7(32'h37871a4f),
	.w8(32'h3884c3fb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9f707),
	.w1(32'hbadd80f0),
	.w2(32'hbb02120f),
	.w3(32'hba8db921),
	.w4(32'hbaf34717),
	.w5(32'hbaaf890b),
	.w6(32'hbb051819),
	.w7(32'hbba4f551),
	.w8(32'hbb98ce47),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacace83),
	.w1(32'h3a657ec2),
	.w2(32'h3a894f88),
	.w3(32'hbab0765b),
	.w4(32'hbaa4c63b),
	.w5(32'hbb00c4cd),
	.w6(32'hbaf357bb),
	.w7(32'hba1e8f90),
	.w8(32'hbb27113f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b3fa),
	.w1(32'hbbda9a9a),
	.w2(32'hbbec2aea),
	.w3(32'hbbb2fb61),
	.w4(32'hbbac68ac),
	.w5(32'hbc0b8bbc),
	.w6(32'hbbf85821),
	.w7(32'hbc075685),
	.w8(32'hbc1e68af),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcafa84),
	.w1(32'h3b3c9548),
	.w2(32'h38a35aa7),
	.w3(32'h3aa1c7c4),
	.w4(32'h3afa596d),
	.w5(32'hba0b1159),
	.w6(32'h39b523fb),
	.w7(32'h3c6a3d8b),
	.w8(32'h3c2dbee8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0249d1),
	.w1(32'hbb461beb),
	.w2(32'hb9e06d01),
	.w3(32'h3c177401),
	.w4(32'hbbb92eb1),
	.w5(32'h3b0fa266),
	.w6(32'h3c1773e3),
	.w7(32'hbb33704a),
	.w8(32'hbbab2637),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba616318),
	.w1(32'h3abf8dd1),
	.w2(32'h3c93decf),
	.w3(32'hb97e59c7),
	.w4(32'h3bac121d),
	.w5(32'hbd0895d5),
	.w6(32'hbbbc7148),
	.w7(32'h3b8b1416),
	.w8(32'h3cba4a1b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5c0b),
	.w1(32'h3a3c597a),
	.w2(32'h3b1fbefe),
	.w3(32'h3b4d506c),
	.w4(32'hbc02221e),
	.w5(32'hbc0d65de),
	.w6(32'h3bf3f8a2),
	.w7(32'h3b1618a3),
	.w8(32'hbb4adf64),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e574),
	.w1(32'hbbb43c76),
	.w2(32'hbc294504),
	.w3(32'hbb679e77),
	.w4(32'h3b837a47),
	.w5(32'h3d1ec337),
	.w6(32'h3a16338c),
	.w7(32'hbb9a1609),
	.w8(32'hbc0acd58),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90a9c3),
	.w1(32'hbaf105fa),
	.w2(32'h3ba49b1a),
	.w3(32'hbb9e8a11),
	.w4(32'hbc157353),
	.w5(32'hbc7b0638),
	.w6(32'hbc1896ee),
	.w7(32'hba918c71),
	.w8(32'hbabfc91f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9682),
	.w1(32'h3b4e8096),
	.w2(32'hbc1b933b),
	.w3(32'hbc08f27c),
	.w4(32'hbaab65b6),
	.w5(32'h3c749d4c),
	.w6(32'hbbca35a8),
	.w7(32'hbc4541f4),
	.w8(32'hbc77b318),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c2b3),
	.w1(32'hbbb557f7),
	.w2(32'hbcce4bab),
	.w3(32'hbb54a265),
	.w4(32'hbbe28621),
	.w5(32'hba3365e9),
	.w6(32'hbc023064),
	.w7(32'hbb0ac561),
	.w8(32'hbb776067),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd517a),
	.w1(32'hbac6ba6c),
	.w2(32'h3bd300ba),
	.w3(32'h3c5b565c),
	.w4(32'hbbd77826),
	.w5(32'h3cad12fe),
	.w6(32'h3c69f767),
	.w7(32'hba03b8fd),
	.w8(32'hbc0c90ea),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eed1b),
	.w1(32'hbb805bce),
	.w2(32'hbb0a67c9),
	.w3(32'hbc571127),
	.w4(32'hbc358544),
	.w5(32'hba3817b2),
	.w6(32'hbc3dc46e),
	.w7(32'hbbeac058),
	.w8(32'h3b4c299f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc25e),
	.w1(32'hbba42265),
	.w2(32'hbc2c2df4),
	.w3(32'hbbbd92ce),
	.w4(32'h3b2aa278),
	.w5(32'hbc47fc2b),
	.w6(32'h3b35548c),
	.w7(32'h3c08830e),
	.w8(32'h3bea982b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a2da3),
	.w1(32'h3c4d6a81),
	.w2(32'h3c590e5b),
	.w3(32'h3b3c042e),
	.w4(32'h3cad9d6b),
	.w5(32'h3c5ba8e4),
	.w6(32'h3b012c5c),
	.w7(32'h3cd746eb),
	.w8(32'h3c88f2ba),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a0326),
	.w1(32'hbc0f343e),
	.w2(32'hbc1df755),
	.w3(32'h3c2779da),
	.w4(32'hbbe44c0b),
	.w5(32'hbadf6d96),
	.w6(32'h3c8ac19a),
	.w7(32'hbc17ba13),
	.w8(32'hbb94126a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587b56),
	.w1(32'h3a315bae),
	.w2(32'hb9b43f0f),
	.w3(32'h396a3bf7),
	.w4(32'hbc35e939),
	.w5(32'hbd22c1d5),
	.w6(32'hba4edfea),
	.w7(32'h3b84145d),
	.w8(32'h3c46e295),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f4f5f),
	.w1(32'h3bbe6f23),
	.w2(32'hbc69328c),
	.w3(32'hbc1dbe44),
	.w4(32'h3b9eb5cb),
	.w5(32'hbab0d4e7),
	.w6(32'h3c1956bf),
	.w7(32'hbacd842e),
	.w8(32'h3850f645),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079c72),
	.w1(32'hba373498),
	.w2(32'h3c573991),
	.w3(32'h3b069f32),
	.w4(32'h3b965425),
	.w5(32'hbbf331c9),
	.w6(32'h3bb2b11b),
	.w7(32'hbba1384f),
	.w8(32'hbb3f6a7d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8b257),
	.w1(32'h3b827463),
	.w2(32'h3b87cca7),
	.w3(32'hbb6b5b5d),
	.w4(32'hbbaa3ab4),
	.w5(32'h3b285a51),
	.w6(32'hba9b41de),
	.w7(32'h3b390ef4),
	.w8(32'hbb056fd7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4018e0),
	.w1(32'hbba0c6ab),
	.w2(32'h3b992281),
	.w3(32'hbbe06e64),
	.w4(32'hbc6aead3),
	.w5(32'h3c52da08),
	.w6(32'h3ab836b4),
	.w7(32'hba9f9422),
	.w8(32'hbafae727),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e17d9),
	.w1(32'hbc305171),
	.w2(32'hbba83e32),
	.w3(32'hb9f6e51d),
	.w4(32'hbc90070a),
	.w5(32'h3cef29dc),
	.w6(32'hbb790da7),
	.w7(32'hbc5a54ee),
	.w8(32'hbb9d1823),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fb0e4),
	.w1(32'hbc5d9d51),
	.w2(32'hbc28cb40),
	.w3(32'hbc56e6cd),
	.w4(32'hbb7e0b52),
	.w5(32'h3b4c3178),
	.w6(32'hbc7cad8f),
	.w7(32'hbbbabb46),
	.w8(32'hbbee1452),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb786e67),
	.w1(32'hbc43c4d1),
	.w2(32'hbab445f5),
	.w3(32'hbcafa72e),
	.w4(32'hbcb01d84),
	.w5(32'hbc80f827),
	.w6(32'hbc0c7552),
	.w7(32'hbc54bc84),
	.w8(32'hbcb6d5f1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24df82),
	.w1(32'hbb811056),
	.w2(32'hbb7ed298),
	.w3(32'h3c09c546),
	.w4(32'hb80f33ea),
	.w5(32'h3b52f6b9),
	.w6(32'hbbafeeea),
	.w7(32'hbb621265),
	.w8(32'hbbd2c4d8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb121c5),
	.w1(32'hbb1f8bcd),
	.w2(32'hbc7149a8),
	.w3(32'h3b1777f3),
	.w4(32'hbc5beedd),
	.w5(32'hbc534a99),
	.w6(32'hbb917639),
	.w7(32'h3ae2f473),
	.w8(32'hbb8bf96e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88d2ed),
	.w1(32'hbba662b6),
	.w2(32'hbb6408d3),
	.w3(32'hbbb6fd74),
	.w4(32'hbc6063ce),
	.w5(32'hbd118f57),
	.w6(32'h3be32d89),
	.w7(32'h3b746baa),
	.w8(32'h3bb106c9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dfc8c),
	.w1(32'h3b7f9b8f),
	.w2(32'h3bb2c9e8),
	.w3(32'hbca36474),
	.w4(32'hbb98678f),
	.w5(32'h3c61fb26),
	.w6(32'hbb539b8b),
	.w7(32'h3b077b09),
	.w8(32'hbbe022de),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6aeda4),
	.w1(32'hba6e60b5),
	.w2(32'hbc534db3),
	.w3(32'h3a5a4ce3),
	.w4(32'h3ad5539b),
	.w5(32'h3c38a7dc),
	.w6(32'h3be05376),
	.w7(32'h3c396da8),
	.w8(32'h3bc421a3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278dfe),
	.w1(32'h3bc29737),
	.w2(32'h3b2086b3),
	.w3(32'h3c3986f0),
	.w4(32'h3b897c68),
	.w5(32'h3bd7edde),
	.w6(32'h3c2f8dbf),
	.w7(32'hbc33dba6),
	.w8(32'hba43e9f6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37de59),
	.w1(32'hbad4fac3),
	.w2(32'hbcb83c69),
	.w3(32'hbc5ada02),
	.w4(32'hbbd56c1b),
	.w5(32'h3cad1561),
	.w6(32'hbbbe515f),
	.w7(32'hbc3d203a),
	.w8(32'hbad088ef),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22a405),
	.w1(32'h3af44314),
	.w2(32'hbac16fec),
	.w3(32'hbb8d480e),
	.w4(32'hbb93ddda),
	.w5(32'hbbfa93ed),
	.w6(32'hbc20baad),
	.w7(32'h3b56a45e),
	.w8(32'hbbff886a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc22c5),
	.w1(32'hbc04c6d4),
	.w2(32'hbcad4073),
	.w3(32'h3c1de922),
	.w4(32'hbbb8d1bc),
	.w5(32'hbc6fd00f),
	.w6(32'h3bc93f99),
	.w7(32'hbb2db409),
	.w8(32'hbc6d8abd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4253dd),
	.w1(32'hbc61105d),
	.w2(32'hbc25016e),
	.w3(32'hbc5ce6f6),
	.w4(32'hbc3ad7ae),
	.w5(32'hbcc8232b),
	.w6(32'hbc49c558),
	.w7(32'hbb9f0a48),
	.w8(32'hbbf35a6c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e2c27),
	.w1(32'h3b245cd4),
	.w2(32'hbae019de),
	.w3(32'h3c23bef1),
	.w4(32'h3c6f8fd9),
	.w5(32'h3d578269),
	.w6(32'h3c0fa0d7),
	.w7(32'hbbd0c8a9),
	.w8(32'hbb9faa38),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e0f10),
	.w1(32'hbc6ad335),
	.w2(32'hbb37efd4),
	.w3(32'h3b4b27b1),
	.w4(32'hbb40daf4),
	.w5(32'hbc20b382),
	.w6(32'hba9f96a8),
	.w7(32'hbcb898ef),
	.w8(32'hbc06f4e4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc730407),
	.w1(32'h3a9f938b),
	.w2(32'hbb347775),
	.w3(32'hbbf494ab),
	.w4(32'h393d4e95),
	.w5(32'h3c3e6706),
	.w6(32'hbbd75e66),
	.w7(32'hbafafd6a),
	.w8(32'hbbf6bdc7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5213ee),
	.w1(32'hbbf83c6a),
	.w2(32'h3995848a),
	.w3(32'hb90bd45a),
	.w4(32'hbbeed64d),
	.w5(32'hbc315abd),
	.w6(32'h3a24fe33),
	.w7(32'hba90bbdf),
	.w8(32'hbbbbf1bd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397155e8),
	.w1(32'hbc4ca0a7),
	.w2(32'hbcd7b566),
	.w3(32'hbc2c5e79),
	.w4(32'hbc585df7),
	.w5(32'hbce6f462),
	.w6(32'hbbb84d6a),
	.w7(32'h3c3d3bdf),
	.w8(32'h3c12cac4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb513e4a),
	.w1(32'h3a006706),
	.w2(32'hba7e0188),
	.w3(32'h3bfafe24),
	.w4(32'hbb93286b),
	.w5(32'hbc5027d7),
	.w6(32'h3c3e1243),
	.w7(32'h3bb49fbe),
	.w8(32'h3b0c4aeb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46fdc5),
	.w1(32'h3bb6fc09),
	.w2(32'hbaf0fa54),
	.w3(32'h3ae98e0f),
	.w4(32'h3b012b7a),
	.w5(32'h3c07f63c),
	.w6(32'hbb4bd8b4),
	.w7(32'h3aa7da3d),
	.w8(32'h3bd44c88),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f127e),
	.w1(32'h3b496aba),
	.w2(32'h3c0d935d),
	.w3(32'h3b063d8d),
	.w4(32'hba454c68),
	.w5(32'hbb5f3133),
	.w6(32'h38da3c3b),
	.w7(32'h3b3ec260),
	.w8(32'hba980a42),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fed5b),
	.w1(32'hbb363376),
	.w2(32'h3b16eef8),
	.w3(32'h3ba0c560),
	.w4(32'h3b753610),
	.w5(32'hbca61f0d),
	.w6(32'hbad489b5),
	.w7(32'h3be82086),
	.w8(32'h3c9f21a2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea643),
	.w1(32'hbba8b4e9),
	.w2(32'h3c7f1e30),
	.w3(32'h3c11c0b1),
	.w4(32'h3bf97684),
	.w5(32'hbb33cba2),
	.w6(32'hba912a43),
	.w7(32'hbc1ef638),
	.w8(32'h3b08c3f2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526119),
	.w1(32'h3add8329),
	.w2(32'hbbf149bd),
	.w3(32'h3ba4c30d),
	.w4(32'h3c388b07),
	.w5(32'h3b214a0f),
	.w6(32'hb8c497c1),
	.w7(32'hbb28b29f),
	.w8(32'h38e895d4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a127fe9),
	.w1(32'h3bd3543d),
	.w2(32'hba843987),
	.w3(32'h3bb0af14),
	.w4(32'h3c2993a8),
	.w5(32'h3b0dbf94),
	.w6(32'h3c3018af),
	.w7(32'h3bf600b4),
	.w8(32'hba02f391),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6fab3),
	.w1(32'hbb28c722),
	.w2(32'hbc214de0),
	.w3(32'h3b657c9d),
	.w4(32'h3bfbbeb7),
	.w5(32'h3d0f3093),
	.w6(32'h3b8926e3),
	.w7(32'hbb9b14a6),
	.w8(32'hbc90b58f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be32ace),
	.w1(32'h3b0ec68a),
	.w2(32'hbb19b02b),
	.w3(32'hbaa76104),
	.w4(32'hbc484a77),
	.w5(32'h3ad3c8b5),
	.w6(32'hbc862960),
	.w7(32'hbc6b2e88),
	.w8(32'hbbcfa1a3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd6913),
	.w1(32'h3be810b2),
	.w2(32'h3bbff60b),
	.w3(32'hbbeca4e8),
	.w4(32'h3b8754d9),
	.w5(32'hbb6c9583),
	.w6(32'hbbf7aa9d),
	.w7(32'h3be97ca3),
	.w8(32'h39c2514f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba166cc),
	.w1(32'h3abd0dbb),
	.w2(32'h3b2dc668),
	.w3(32'h3bc8bc4f),
	.w4(32'hb8ec542f),
	.w5(32'h3b5c4efe),
	.w6(32'h3bfe1d57),
	.w7(32'h3b5ca851),
	.w8(32'h3b597633),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca3f69),
	.w1(32'h3b35153e),
	.w2(32'h3b323b6c),
	.w3(32'hbba06ce4),
	.w4(32'hba3a7a57),
	.w5(32'hbc2d5a33),
	.w6(32'hbb808c6c),
	.w7(32'hbb1d6930),
	.w8(32'hbbb2c0dc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28d970),
	.w1(32'h3b80b007),
	.w2(32'hbb7e8273),
	.w3(32'hba38f44a),
	.w4(32'h3bef92f3),
	.w5(32'hbca10f64),
	.w6(32'hbb763a74),
	.w7(32'h3c71e821),
	.w8(32'h3ae65d18),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144603),
	.w1(32'hbb8ddc41),
	.w2(32'h3bff473b),
	.w3(32'h398f38a4),
	.w4(32'hbc6727fc),
	.w5(32'h3ca7594a),
	.w6(32'h3bad48b4),
	.w7(32'hbc44e600),
	.w8(32'h3946d214),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a817e3b),
	.w1(32'h39ef0ab2),
	.w2(32'h3ad6d46f),
	.w3(32'hbc83c542),
	.w4(32'hbbf8dd1f),
	.w5(32'hbc3ae424),
	.w6(32'hbc2e96b3),
	.w7(32'h3b78d31a),
	.w8(32'hbbc99a54),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f7e78),
	.w1(32'hbb934d19),
	.w2(32'hbc88f348),
	.w3(32'hbbb6bf0c),
	.w4(32'hbb2f2dba),
	.w5(32'h3acc3be6),
	.w6(32'h3a91f118),
	.w7(32'h3afae794),
	.w8(32'h3afec3d3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a67c),
	.w1(32'h3bcfadf3),
	.w2(32'hbc1ef7bf),
	.w3(32'hbb9589ff),
	.w4(32'h3bd7f5dc),
	.w5(32'h3ba83fc0),
	.w6(32'h3b2324b3),
	.w7(32'h3ac97ca4),
	.w8(32'hbbe21bea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f6614),
	.w1(32'hbbf706fd),
	.w2(32'hbbb21ebd),
	.w3(32'hbb70451d),
	.w4(32'h3b534cd4),
	.w5(32'h3cde6ec0),
	.w6(32'h3a689f27),
	.w7(32'h3991c950),
	.w8(32'h3a67dea3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b300790),
	.w1(32'hbbf9192b),
	.w2(32'hb96439ff),
	.w3(32'h3aa6f4d9),
	.w4(32'h3b72ffde),
	.w5(32'hbc432728),
	.w6(32'hbbe7be51),
	.w7(32'h3b9230e3),
	.w8(32'hba93f3c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c82d7),
	.w1(32'hbc05696c),
	.w2(32'h3bfeb3da),
	.w3(32'hbb8c751f),
	.w4(32'h3bd16bc4),
	.w5(32'hbcaece1d),
	.w6(32'hbb9d7d60),
	.w7(32'h3a1a6aa4),
	.w8(32'h3c4a3370),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a02d),
	.w1(32'hbb6fa169),
	.w2(32'h3a84f024),
	.w3(32'h3b3cf74b),
	.w4(32'h3aeb0daa),
	.w5(32'hbb8a865c),
	.w6(32'hba9f5c4c),
	.w7(32'hbb30521a),
	.w8(32'hbb92a1d3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b48c),
	.w1(32'hbc0314e4),
	.w2(32'h3bee7c73),
	.w3(32'h3c2f460e),
	.w4(32'hbbee3213),
	.w5(32'hbbb012c6),
	.w6(32'hbafe9e99),
	.w7(32'hbc12dcfe),
	.w8(32'hbc05a16a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6256d2),
	.w1(32'h3b955d5e),
	.w2(32'h3b177094),
	.w3(32'h3b143444),
	.w4(32'hbb0c4643),
	.w5(32'hbc350a35),
	.w6(32'hbb6c9aa8),
	.w7(32'h393f4ed9),
	.w8(32'h3b6fda9e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0bfce),
	.w1(32'hbbe61c44),
	.w2(32'h3a5c748d),
	.w3(32'hbb74243e),
	.w4(32'hbb52cc53),
	.w5(32'hb98e585d),
	.w6(32'h3b81fb94),
	.w7(32'hbb009625),
	.w8(32'h3b14cb92),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1a62a),
	.w1(32'hbb453db2),
	.w2(32'h3a14b595),
	.w3(32'hb9e3f02f),
	.w4(32'hbc46ee5e),
	.w5(32'hbcac3dfd),
	.w6(32'h3ba65ec1),
	.w7(32'hbaa9282d),
	.w8(32'hbc045c5e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de4cc),
	.w1(32'hbaf70d37),
	.w2(32'hbca4ee72),
	.w3(32'h3ba64b30),
	.w4(32'hb953c4fc),
	.w5(32'h3d04bcb9),
	.w6(32'hbc3cb4dc),
	.w7(32'hbc3dd9a8),
	.w8(32'hbca65d20),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2230b0),
	.w1(32'hbac527c8),
	.w2(32'hba4cd11e),
	.w3(32'hbba14521),
	.w4(32'hbc0c936b),
	.w5(32'hbc83145a),
	.w6(32'hbbe96436),
	.w7(32'hbab07a7c),
	.w8(32'hba88265f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea7987),
	.w1(32'hbb8624be),
	.w2(32'hbb68f91b),
	.w3(32'h3bfeb822),
	.w4(32'h3c2f912a),
	.w5(32'h3b34a640),
	.w6(32'hbb63936f),
	.w7(32'h3a9fc851),
	.w8(32'h3bf58f47),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5e50e),
	.w1(32'hbb88268f),
	.w2(32'h3b9726c0),
	.w3(32'hba75a20d),
	.w4(32'hbbd31736),
	.w5(32'hbbb9f209),
	.w6(32'h3a383c2d),
	.w7(32'hbbd6610a),
	.w8(32'hb9b20615),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdf98d),
	.w1(32'hbbccc4f5),
	.w2(32'hbcd152fb),
	.w3(32'hbb3d32b1),
	.w4(32'hbc044b09),
	.w5(32'h3cfc2dcd),
	.w6(32'hbb4929f3),
	.w7(32'hbc8c3b59),
	.w8(32'hbc8f8535),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e309c),
	.w1(32'h3bbd1fec),
	.w2(32'h3c2b9950),
	.w3(32'hbc462461),
	.w4(32'hbb0aed91),
	.w5(32'h3d345cb6),
	.w6(32'hba351778),
	.w7(32'hbc4e1aa0),
	.w8(32'hbc520756),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0af89),
	.w1(32'hba20cbf1),
	.w2(32'hbc394a05),
	.w3(32'h3ba0dc4c),
	.w4(32'h39dc7958),
	.w5(32'hbbdbe6cd),
	.w6(32'h38d189aa),
	.w7(32'h3c192d26),
	.w8(32'hbbcdaa95),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b4fd7),
	.w1(32'h3c4d511c),
	.w2(32'h3b4a6260),
	.w3(32'hbc6b506f),
	.w4(32'h3b24792f),
	.w5(32'hbb61ddb1),
	.w6(32'hbc33d7ac),
	.w7(32'h3b97242a),
	.w8(32'h3b52ec9c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd1ad7),
	.w1(32'h3bbeaa18),
	.w2(32'h3bab21a2),
	.w3(32'h3c29c9d5),
	.w4(32'h3b9f007f),
	.w5(32'h3a67e328),
	.w6(32'h3a0abee8),
	.w7(32'h39e2d632),
	.w8(32'h3c595b99),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34d006),
	.w1(32'hb854b2ee),
	.w2(32'hbb9d8e5a),
	.w3(32'h3bba7572),
	.w4(32'h3c1f2a61),
	.w5(32'h3bcf2601),
	.w6(32'h3a6a7f32),
	.w7(32'hbb46db20),
	.w8(32'h3bb56794),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99adc1),
	.w1(32'h3b3751a2),
	.w2(32'h3bb62f06),
	.w3(32'hbb45552f),
	.w4(32'hba3ae091),
	.w5(32'hbc2d05ee),
	.w6(32'hbaf00775),
	.w7(32'h3bd78e59),
	.w8(32'hbb0111aa),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d88c62),
	.w1(32'hbc2809ae),
	.w2(32'h3aa70390),
	.w3(32'h3c5846c4),
	.w4(32'h3c04cf91),
	.w5(32'hbc22b569),
	.w6(32'h3bb48c6c),
	.w7(32'h3bb1ae1a),
	.w8(32'h3b5476b8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9898),
	.w1(32'hbbf16984),
	.w2(32'h3b46d217),
	.w3(32'hbbfe9025),
	.w4(32'h3b087f3f),
	.w5(32'hbc8e81e8),
	.w6(32'hba2d9d37),
	.w7(32'hbb4c74bb),
	.w8(32'h3b4d0902),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9719e7),
	.w1(32'hbba01fe1),
	.w2(32'h3b09e151),
	.w3(32'h3a4c3863),
	.w4(32'h3c0537bb),
	.w5(32'h3b517374),
	.w6(32'h3b03cb78),
	.w7(32'h3bcf11cd),
	.w8(32'h3c000697),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574e79),
	.w1(32'h39f935b4),
	.w2(32'hbbe1e0db),
	.w3(32'hbbb1e4ea),
	.w4(32'h3baacae5),
	.w5(32'hb9ae97d5),
	.w6(32'hbaf093ea),
	.w7(32'h3bb02d2a),
	.w8(32'h3bc292f1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc495161),
	.w1(32'hb99583ef),
	.w2(32'hbb7519ca),
	.w3(32'hba7d49c8),
	.w4(32'hbbbff8e9),
	.w5(32'h3a01751e),
	.w6(32'h3c0b428f),
	.w7(32'hbbd09a94),
	.w8(32'h3a62deeb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcafee4),
	.w1(32'h3b9f0fca),
	.w2(32'hbc119667),
	.w3(32'h3a94d229),
	.w4(32'h3ba1bb34),
	.w5(32'h3a749b9a),
	.w6(32'hbadb3eff),
	.w7(32'hbb2d8929),
	.w8(32'h3aff8c91),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8efba9),
	.w1(32'hbb6cf2b5),
	.w2(32'hbbf39ac7),
	.w3(32'hbbc1202f),
	.w4(32'h3b7cff1b),
	.w5(32'hbab2c8e2),
	.w6(32'hbb9306fd),
	.w7(32'h3be223ff),
	.w8(32'h3c081c2e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c136d96),
	.w1(32'h3ab0c423),
	.w2(32'h3ab39fa7),
	.w3(32'hbb64b59e),
	.w4(32'h3bb9d1ed),
	.w5(32'h3bfb7f08),
	.w6(32'h3b3d7e41),
	.w7(32'h3c01ae78),
	.w8(32'h3b0fe7a5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89778),
	.w1(32'h3b7c1871),
	.w2(32'h3b824992),
	.w3(32'hb9a1a360),
	.w4(32'hbb233bea),
	.w5(32'hbb8b7f45),
	.w6(32'hbb59cda2),
	.w7(32'hba9f6740),
	.w8(32'hbb8828b3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a41ee),
	.w1(32'hbbb6480b),
	.w2(32'h3a432886),
	.w3(32'h3c3eedda),
	.w4(32'hbbadb55a),
	.w5(32'hbc8001f0),
	.w6(32'h3b28322f),
	.w7(32'h3a8c9c68),
	.w8(32'hbb17bdee),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f9953),
	.w1(32'hbb9b6f9b),
	.w2(32'h393dcc8d),
	.w3(32'h3bac8cab),
	.w4(32'hbaebb9fd),
	.w5(32'hb9a55028),
	.w6(32'hbb49a3f9),
	.w7(32'hbb545d67),
	.w8(32'hbb108852),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cdbeb),
	.w1(32'hba75fbfe),
	.w2(32'h3b9c7169),
	.w3(32'h3b515201),
	.w4(32'hba4c1f09),
	.w5(32'hbad17573),
	.w6(32'h3c3b4316),
	.w7(32'h3b89dc3f),
	.w8(32'hbba410f7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b7c57),
	.w1(32'h3b1ea507),
	.w2(32'hbb4837d5),
	.w3(32'hbbbac935),
	.w4(32'hbb334adc),
	.w5(32'hbc126c79),
	.w6(32'hbb297904),
	.w7(32'h3bb3d5f1),
	.w8(32'h3c0abac1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d97f),
	.w1(32'h3c569d63),
	.w2(32'hbc0a11d7),
	.w3(32'hba25e759),
	.w4(32'hbba472bd),
	.w5(32'hbbdafeab),
	.w6(32'h3bae7484),
	.w7(32'hbaccb271),
	.w8(32'h3a4201fb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcc458),
	.w1(32'h3c45c87e),
	.w2(32'h3be3353b),
	.w3(32'hbb9fa77e),
	.w4(32'hba86dad1),
	.w5(32'hba41ee0e),
	.w6(32'h3bc19aeb),
	.w7(32'hbb6a25e2),
	.w8(32'hbc4dff09),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0da797),
	.w1(32'h3b745949),
	.w2(32'hb9bf6bab),
	.w3(32'hbbc67ec1),
	.w4(32'h3b0dd21d),
	.w5(32'hbb3b6f0c),
	.w6(32'hbb7c287e),
	.w7(32'hba7bcbb8),
	.w8(32'h3c0005d9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc43156),
	.w1(32'h3b1d538a),
	.w2(32'h3ae8eb67),
	.w3(32'hbafa5d11),
	.w4(32'h3bab7530),
	.w5(32'h3bf9cb19),
	.w6(32'h3a9a6570),
	.w7(32'hbb8e413f),
	.w8(32'h3b5333a6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3e163),
	.w1(32'hbb45c3e4),
	.w2(32'hbbe50e19),
	.w3(32'h3b4f4857),
	.w4(32'hbb0eaa74),
	.w5(32'hbc6d40e5),
	.w6(32'hbc0a4455),
	.w7(32'hb9b33787),
	.w8(32'h3be1bd73),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff84cb),
	.w1(32'h3bf3cb8c),
	.w2(32'hbad723e8),
	.w3(32'hbb5ef307),
	.w4(32'hbc2aa9bd),
	.w5(32'hba2b9d6e),
	.w6(32'h3bbb80f0),
	.w7(32'hbc398002),
	.w8(32'hbc4c56c7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb743636),
	.w1(32'h3c319108),
	.w2(32'hbb960ab1),
	.w3(32'h3b9a64f9),
	.w4(32'hbadf20a4),
	.w5(32'h3d4919db),
	.w6(32'h3b2bc11a),
	.w7(32'hbc066690),
	.w8(32'hbccc68e9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa35f6),
	.w1(32'h3b25375c),
	.w2(32'hbaae17b4),
	.w3(32'h3cbc4e5d),
	.w4(32'h3b0657df),
	.w5(32'h3cdd1cde),
	.w6(32'hba7c06a2),
	.w7(32'hbb9e6d33),
	.w8(32'hbc673c5d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d223b),
	.w1(32'hbb6ebafa),
	.w2(32'h3b51645d),
	.w3(32'hbae7926c),
	.w4(32'hbb0226f9),
	.w5(32'hbcf0458f),
	.w6(32'h3acf7994),
	.w7(32'h3c763f09),
	.w8(32'h3c991225),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ac0a),
	.w1(32'h3b69594e),
	.w2(32'hba31e421),
	.w3(32'hbbdc49fe),
	.w4(32'hbaf7d9ba),
	.w5(32'hbc34c1ae),
	.w6(32'hbb2bfb37),
	.w7(32'hbb7b6b27),
	.w8(32'h3b98e6da),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06fb9d),
	.w1(32'h3c802b33),
	.w2(32'hb9e57865),
	.w3(32'hbb98e964),
	.w4(32'h3c434ce4),
	.w5(32'hbb4056b9),
	.w6(32'h3bc62da9),
	.w7(32'h3c27c383),
	.w8(32'h3c1d3651),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c19a4),
	.w1(32'h3c0618f0),
	.w2(32'h3ad2b368),
	.w3(32'h3aa140bd),
	.w4(32'hbbc34d3c),
	.w5(32'h3c4c075b),
	.w6(32'h3c19e5a8),
	.w7(32'h3aed8850),
	.w8(32'h3bf7cecd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3032bc),
	.w1(32'hba848f42),
	.w2(32'h3bbe25d5),
	.w3(32'h3c15a4c2),
	.w4(32'hbb3281ff),
	.w5(32'hbbca5fc2),
	.w6(32'h3c1f9754),
	.w7(32'hbb91deda),
	.w8(32'h3b6b750d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83c42e),
	.w1(32'hbba491ea),
	.w2(32'hbb6ffe4a),
	.w3(32'h3b0f71cb),
	.w4(32'hbbd68284),
	.w5(32'h3bcd7685),
	.w6(32'hb82c2062),
	.w7(32'h3ac8d437),
	.w8(32'h3bbfea26),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2576d3),
	.w1(32'hbc13147f),
	.w2(32'h3d00bc35),
	.w3(32'h3b8e884b),
	.w4(32'hbb66a2fc),
	.w5(32'hbc81f773),
	.w6(32'h3b233800),
	.w7(32'h3c2f8f4c),
	.w8(32'h3904d2f5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29fe0d),
	.w1(32'hbbaaf3b9),
	.w2(32'hbc5b5579),
	.w3(32'h3b485351),
	.w4(32'hbb81e8d1),
	.w5(32'hbc232194),
	.w6(32'h3c3030af),
	.w7(32'hbc57a7bd),
	.w8(32'hbb6fae49),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17d1c0),
	.w1(32'hbb8a567c),
	.w2(32'h3c094ea3),
	.w3(32'hbc1c7d90),
	.w4(32'hbb99d964),
	.w5(32'hbc67cd6d),
	.w6(32'hbbc96e20),
	.w7(32'hbb41751a),
	.w8(32'hbbf813ac),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68551),
	.w1(32'h3c0a7322),
	.w2(32'h3bfd1214),
	.w3(32'h3c210727),
	.w4(32'h3adb50f2),
	.w5(32'hba41e976),
	.w6(32'hbb530661),
	.w7(32'h3c13dfee),
	.w8(32'h3c038272),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae6f39),
	.w1(32'h3adaedf2),
	.w2(32'hbb281517),
	.w3(32'h3a819d2b),
	.w4(32'h3bdb6fd7),
	.w5(32'h3c247dab),
	.w6(32'h3b13ec41),
	.w7(32'hba70a03a),
	.w8(32'hbc3e49fe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd15df),
	.w1(32'hbb866c69),
	.w2(32'h3a408907),
	.w3(32'hbba2a707),
	.w4(32'h3b5a1eac),
	.w5(32'hbc1f3243),
	.w6(32'hbbe7a62d),
	.w7(32'h3b1024b9),
	.w8(32'h3b92b114),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7b4d),
	.w1(32'hbb84be75),
	.w2(32'h3c1d148d),
	.w3(32'hbc197c39),
	.w4(32'hbb919561),
	.w5(32'hbc8fbc38),
	.w6(32'hbbf408f8),
	.w7(32'hbc1d6b50),
	.w8(32'hbc15b1e0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5467),
	.w1(32'hbb1256a0),
	.w2(32'h3b3348ba),
	.w3(32'hba5d6286),
	.w4(32'hbc210733),
	.w5(32'hbb209b02),
	.w6(32'h3b040cdc),
	.w7(32'hbb14b19e),
	.w8(32'h39e3fd3c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc19c3),
	.w1(32'hbc4b0184),
	.w2(32'h3ba0540e),
	.w3(32'h3bca25a0),
	.w4(32'hba144e34),
	.w5(32'hbbf24301),
	.w6(32'h3bea4bf3),
	.w7(32'h3a859ab7),
	.w8(32'hbc07fc86),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c203573),
	.w1(32'h3bd76d20),
	.w2(32'h3c34665d),
	.w3(32'hbc2f094d),
	.w4(32'hbb96766d),
	.w5(32'hbbee4061),
	.w6(32'hbc05cf76),
	.w7(32'hbc533634),
	.w8(32'hbc344040),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82951a),
	.w1(32'hbb0864cf),
	.w2(32'hbc238723),
	.w3(32'hbc3ff714),
	.w4(32'h3ac5d4de),
	.w5(32'hb7539708),
	.w6(32'h38ccb08e),
	.w7(32'h3b76535e),
	.w8(32'h3aaa9811),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb042431),
	.w1(32'hba887125),
	.w2(32'h3b9dd28e),
	.w3(32'hba261f72),
	.w4(32'hbaca6c86),
	.w5(32'h3a466a6c),
	.w6(32'h3b782c15),
	.w7(32'h3a8442f8),
	.w8(32'h3b529e61),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38692),
	.w1(32'hbbbfa8cd),
	.w2(32'h3bf8636e),
	.w3(32'h3c04c3d8),
	.w4(32'h3ab9c559),
	.w5(32'h3cd41e0c),
	.w6(32'h3bec9e33),
	.w7(32'hbc199825),
	.w8(32'hba5fc95e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20849),
	.w1(32'h3b7bfbdf),
	.w2(32'h3be2502d),
	.w3(32'hbbb3327b),
	.w4(32'h3a8cde74),
	.w5(32'h3d48791a),
	.w6(32'hbc100057),
	.w7(32'hbc2e25f6),
	.w8(32'hbbdde6c4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149d5e),
	.w1(32'hbc20d9c2),
	.w2(32'hbc8f0c11),
	.w3(32'h3c4111ce),
	.w4(32'hbb71dc9f),
	.w5(32'hbb8d0bf7),
	.w6(32'hbc333e5b),
	.w7(32'h3c049a55),
	.w8(32'h3c1b1938),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4181e4),
	.w1(32'h3b928fe0),
	.w2(32'h3b128598),
	.w3(32'hbb9a72e3),
	.w4(32'hbc2979d0),
	.w5(32'hb9288b20),
	.w6(32'hbc07d0e4),
	.w7(32'hba528e10),
	.w8(32'hbb6acbfc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1018a1),
	.w1(32'h39bd225f),
	.w2(32'hbb394ac2),
	.w3(32'h3b0e8aea),
	.w4(32'h3b932bd2),
	.w5(32'h3b6a052c),
	.w6(32'hbbfd3c52),
	.w7(32'h3b415aca),
	.w8(32'h3b1bcb1a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395af8),
	.w1(32'h3b824417),
	.w2(32'hb90baaa3),
	.w3(32'h3b999e2b),
	.w4(32'h3b8cad27),
	.w5(32'hbb897b84),
	.w6(32'hb8b4de3f),
	.w7(32'h3c33f0c1),
	.w8(32'h3baf0533),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335a35),
	.w1(32'hba2a1b82),
	.w2(32'h3baddefc),
	.w3(32'hbb9c8984),
	.w4(32'h3bf3681c),
	.w5(32'h3b8da548),
	.w6(32'h3adde45e),
	.w7(32'h3b893998),
	.w8(32'h3c042f0d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22247),
	.w1(32'hbbecc792),
	.w2(32'hbc3bfb66),
	.w3(32'h3b3feb69),
	.w4(32'hbc15f8b8),
	.w5(32'hbb05f527),
	.w6(32'hbab5b1ba),
	.w7(32'hbb36efc6),
	.w8(32'hbb9e6fd0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e26cd),
	.w1(32'h3b04fbb5),
	.w2(32'hbc1bf1a8),
	.w3(32'h3a2d0c00),
	.w4(32'h3b6d593e),
	.w5(32'hba66272e),
	.w6(32'h3a2c76bd),
	.w7(32'h3bcea32a),
	.w8(32'h3a83428e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6a24c),
	.w1(32'h3bc90c09),
	.w2(32'hbb2e848a),
	.w3(32'h3b53585e),
	.w4(32'h3b911b30),
	.w5(32'hbc3a2843),
	.w6(32'h3a51a880),
	.w7(32'h3bdabb90),
	.w8(32'hbb180fbe),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c2c54),
	.w1(32'hbb6a04e2),
	.w2(32'h3ba0f41e),
	.w3(32'hb993773b),
	.w4(32'hbc221909),
	.w5(32'hbc3ff3b4),
	.w6(32'hbb1103f6),
	.w7(32'hbace3649),
	.w8(32'hbbe49af3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23e85f),
	.w1(32'h3b7df74b),
	.w2(32'hbbdf666a),
	.w3(32'hbbc148e9),
	.w4(32'h3a84e3f6),
	.w5(32'h3b7e1440),
	.w6(32'hbc50d454),
	.w7(32'h3b899dd0),
	.w8(32'h3b827244),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57f0f0),
	.w1(32'h3be610ff),
	.w2(32'h3a182104),
	.w3(32'h3a9bd2ec),
	.w4(32'h3bfd358f),
	.w5(32'h3b8255b0),
	.w6(32'hb9ae5f0e),
	.w7(32'h3c671a23),
	.w8(32'h3bf19bcc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b043a0e),
	.w1(32'hbb095144),
	.w2(32'h3b98b746),
	.w3(32'h3bd9c791),
	.w4(32'h3ac741b2),
	.w5(32'h3b639846),
	.w6(32'h3bcc4907),
	.w7(32'hbadb6def),
	.w8(32'h3bb44147),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b759f0e),
	.w1(32'hbaeb551d),
	.w2(32'hbb4aef18),
	.w3(32'hbbc99f59),
	.w4(32'hbc56bd21),
	.w5(32'hbc42808b),
	.w6(32'hbbaab6c6),
	.w7(32'hbc13c02c),
	.w8(32'hbc47d275),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2348d0),
	.w1(32'hbc0bd02b),
	.w2(32'h3bc25357),
	.w3(32'h3b144704),
	.w4(32'hb6db0e28),
	.w5(32'hbac0707e),
	.w6(32'hbac312ca),
	.w7(32'h3a0c8007),
	.w8(32'hbc6959dd),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa491d6),
	.w1(32'h3c4bd1a4),
	.w2(32'hba066cf2),
	.w3(32'hbb15a32d),
	.w4(32'h3bda7391),
	.w5(32'hbb66564e),
	.w6(32'hbc0222fe),
	.w7(32'h3b9a65c5),
	.w8(32'hbb852f48),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc2a61),
	.w1(32'hba1ef8e5),
	.w2(32'hbaa6cc67),
	.w3(32'h3a93fa03),
	.w4(32'hb67b44da),
	.w5(32'hbaf8d15f),
	.w6(32'h3c138624),
	.w7(32'hb9a93b64),
	.w8(32'hbb31f8cc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39459f68),
	.w1(32'h3af0e56c),
	.w2(32'h3904eca2),
	.w3(32'h3a03dea1),
	.w4(32'h3aaf99a5),
	.w5(32'hb9800bb7),
	.w6(32'hb9c1c1fc),
	.w7(32'h3a6c015e),
	.w8(32'hb9200c2e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef2e12),
	.w1(32'h39e2c095),
	.w2(32'h39935910),
	.w3(32'h3a0da184),
	.w4(32'h39b6b789),
	.w5(32'h398efbdc),
	.w6(32'h398a255e),
	.w7(32'h3a300f97),
	.w8(32'h3a11dd0a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f76cf),
	.w1(32'hbad2dd3d),
	.w2(32'hbb10b2ae),
	.w3(32'hba81f130),
	.w4(32'hbae2738a),
	.w5(32'hba8f735c),
	.w6(32'hb9eefb4c),
	.w7(32'hba1e802e),
	.w8(32'hba92353b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8efe5c),
	.w1(32'hb9670d66),
	.w2(32'hb9ab1ef8),
	.w3(32'hbabff0db),
	.w4(32'hb9ff6c8b),
	.w5(32'hba1e492b),
	.w6(32'hbac643e9),
	.w7(32'hb9e03e29),
	.w8(32'hba133e9a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bc9c9),
	.w1(32'hbadccb3b),
	.w2(32'hbb31fef4),
	.w3(32'hba993f14),
	.w4(32'hba0a94f8),
	.w5(32'hba97f0f9),
	.w6(32'hbac72ff7),
	.w7(32'hbaa109d9),
	.w8(32'hbb0040f3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882e1a),
	.w1(32'h3b288bcd),
	.w2(32'h3b3f57b0),
	.w3(32'h37b8fc6d),
	.w4(32'h3b562b1a),
	.w5(32'h3a892150),
	.w6(32'hbae84c2f),
	.w7(32'hb958a06e),
	.w8(32'h3a0c5525),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bd6a5),
	.w1(32'h3a9601cd),
	.w2(32'h3b04ac71),
	.w3(32'hb91c3444),
	.w4(32'h3acf666b),
	.w5(32'h3a74bd02),
	.w6(32'hb85dc898),
	.w7(32'h3aede216),
	.w8(32'h3aaa92d7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03ce52),
	.w1(32'h3a4b86d1),
	.w2(32'hb9fb39b0),
	.w3(32'h3ab25900),
	.w4(32'h3a1c796c),
	.w5(32'hba8b716c),
	.w6(32'h3a2c5ee5),
	.w7(32'hb7ec89ba),
	.w8(32'hba846f65),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e1716),
	.w1(32'h3b75cdf4),
	.w2(32'h3b692f5d),
	.w3(32'h3b200e3c),
	.w4(32'h3ba7001c),
	.w5(32'h3b2dec59),
	.w6(32'h3ac63eb7),
	.w7(32'h3b92706e),
	.w8(32'h3b62b409),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928771a),
	.w1(32'hba54af4e),
	.w2(32'h3a93ba25),
	.w3(32'hb99a0295),
	.w4(32'hbab68357),
	.w5(32'h392be59f),
	.w6(32'hb9c90c01),
	.w7(32'hbaad448c),
	.w8(32'hba7aaacb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d062f3),
	.w1(32'h3ac93f80),
	.w2(32'h3b1b698e),
	.w3(32'h3ab16613),
	.w4(32'h3a3ea30a),
	.w5(32'h38865904),
	.w6(32'h3b77175d),
	.w7(32'h3b0115a1),
	.w8(32'h38e786ef),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a459683),
	.w1(32'h35a80c97),
	.w2(32'h39ea177c),
	.w3(32'h39beba48),
	.w4(32'hb82edc7b),
	.w5(32'h39dd408b),
	.w6(32'h394a1f16),
	.w7(32'hb8911309),
	.w8(32'h393aa7cd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bec92),
	.w1(32'h3a1058cb),
	.w2(32'h3988f342),
	.w3(32'h39975ccc),
	.w4(32'h391abad0),
	.w5(32'h3973dece),
	.w6(32'h39a7ef1f),
	.w7(32'hb945f399),
	.w8(32'h38ad168e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf8655),
	.w1(32'h3b5c897a),
	.w2(32'h3afcd97c),
	.w3(32'h3b5ac2d4),
	.w4(32'h3a9709b2),
	.w5(32'hb8ac72d6),
	.w6(32'h3aa61395),
	.w7(32'h3afa0c0c),
	.w8(32'h39854f62),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a8525),
	.w1(32'hbb6f8591),
	.w2(32'hbb14fa31),
	.w3(32'hbb233d8a),
	.w4(32'hbb9d2d7c),
	.w5(32'hbb108aa3),
	.w6(32'hbbd1f8d4),
	.w7(32'hbbb14fca),
	.w8(32'hbbf65fb5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aacda),
	.w1(32'h3a9769ac),
	.w2(32'h3b620637),
	.w3(32'hba41ca03),
	.w4(32'h3abb552c),
	.w5(32'h3aac0dae),
	.w6(32'hba87092f),
	.w7(32'h3a96ab12),
	.w8(32'h3a9f4281),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ababd2a),
	.w1(32'h3a6e1012),
	.w2(32'h39bdfba1),
	.w3(32'h3a4faac5),
	.w4(32'h3b2b12c3),
	.w5(32'h3a635cce),
	.w6(32'h3985b517),
	.w7(32'hbac76f4d),
	.w8(32'hbb2b07d3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc0bcf),
	.w1(32'h39c6a697),
	.w2(32'h39df4a4e),
	.w3(32'hb92aa01d),
	.w4(32'hb9541128),
	.w5(32'hb93f930e),
	.w6(32'hb8f9e7f9),
	.w7(32'hb99c25d4),
	.w8(32'h38199c44),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1482),
	.w1(32'h3a47e91b),
	.w2(32'h3a206bb1),
	.w3(32'h3a2e7721),
	.w4(32'h39c5c0be),
	.w5(32'h3a1d46e6),
	.w6(32'h3a035564),
	.w7(32'h3969a3a4),
	.w8(32'h3999f7ea),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51e8a2),
	.w1(32'h3b894792),
	.w2(32'hbb224aab),
	.w3(32'h3b626a1e),
	.w4(32'h3afbc7e4),
	.w5(32'hbac713bd),
	.w6(32'h3afb6e19),
	.w7(32'h3b831ebd),
	.w8(32'hbaf7a63b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885b63),
	.w1(32'hbbca2422),
	.w2(32'hbbad3416),
	.w3(32'hbb883980),
	.w4(32'hbbc0e8ba),
	.w5(32'hbb84f572),
	.w6(32'hbb3befed),
	.w7(32'hbbc10db4),
	.w8(32'hbbfd0611),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c4daf),
	.w1(32'h39b868d9),
	.w2(32'hbb95ef05),
	.w3(32'h3a267c2b),
	.w4(32'hbb311449),
	.w5(32'hbb0e05db),
	.w6(32'hbb5cb17c),
	.w7(32'hba50e3be),
	.w8(32'hbb2c6ca1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabf8b9),
	.w1(32'h3b42d3b3),
	.w2(32'h3b09e651),
	.w3(32'h3a513795),
	.w4(32'h3b5a2e7e),
	.w5(32'h3ae07911),
	.w6(32'h39ba083f),
	.w7(32'h3adec9be),
	.w8(32'h3aa95ba2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bdd69),
	.w1(32'h3b2a4ef0),
	.w2(32'h3b4df80d),
	.w3(32'hba08ec98),
	.w4(32'h3b73d051),
	.w5(32'h3af02e49),
	.w6(32'hba6ff257),
	.w7(32'h3a48270d),
	.w8(32'h3a6978a2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8fa51),
	.w1(32'hb9bec1c3),
	.w2(32'hb98400ac),
	.w3(32'h398e4e84),
	.w4(32'hb92c66b5),
	.w5(32'hb911a1ae),
	.w6(32'h37f6045d),
	.w7(32'hb98cb123),
	.w8(32'hb999f945),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967a7ec),
	.w1(32'hb9bf4c3a),
	.w2(32'hb72c7917),
	.w3(32'hb8af64d3),
	.w4(32'hba7782d5),
	.w5(32'h384c5372),
	.w6(32'h3800f81a),
	.w7(32'hba42c5b9),
	.w8(32'hb9946a7c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39f53f),
	.w1(32'hb888b1ad),
	.w2(32'hb9d6e546),
	.w3(32'h398e46a8),
	.w4(32'hb863be52),
	.w5(32'hb9bc3a17),
	.w6(32'hb96b5330),
	.w7(32'hb9dd1ead),
	.w8(32'hb97fc62a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97400d3),
	.w1(32'hb94a092d),
	.w2(32'h38ef401b),
	.w3(32'hb91c5a4f),
	.w4(32'hb94535c7),
	.w5(32'h3a81765d),
	.w6(32'hb9a0ee3a),
	.w7(32'hb8d3f5c3),
	.w8(32'h39b4a0a7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6099a2),
	.w1(32'h3a449f01),
	.w2(32'hb94c7c13),
	.w3(32'h3ae067aa),
	.w4(32'h39b724fb),
	.w5(32'h3a1b73ed),
	.w6(32'h3a9f355e),
	.w7(32'h389b63b6),
	.w8(32'hb9b9c62e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0726d3),
	.w1(32'hba95ffd3),
	.w2(32'hbb0641d1),
	.w3(32'h391fdc23),
	.w4(32'hbaaba85e),
	.w5(32'hbb6e157c),
	.w6(32'hba845287),
	.w7(32'hb98fce6b),
	.w8(32'hbb96c1ee),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2cf2c),
	.w1(32'h3add0fd2),
	.w2(32'h3ac61423),
	.w3(32'h3a9fe3a6),
	.w4(32'h3b200aeb),
	.w5(32'h3a9cab0f),
	.w6(32'h3af978b6),
	.w7(32'h3acfd3d1),
	.w8(32'h38804dfc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa4c62),
	.w1(32'hb7f7d415),
	.w2(32'h35abbcd9),
	.w3(32'h3992f526),
	.w4(32'hb9227691),
	.w5(32'h391331a2),
	.w6(32'hb8bc560c),
	.w7(32'hb7807c25),
	.w8(32'h390563fa),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b379926),
	.w1(32'hbaa3470b),
	.w2(32'hbbff487f),
	.w3(32'h38487597),
	.w4(32'hbb655c39),
	.w5(32'hbb61ae3f),
	.w6(32'hbb49af73),
	.w7(32'hbb30bde4),
	.w8(32'hbbf10b80),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58fc1e),
	.w1(32'hbb175c32),
	.w2(32'hbb030e77),
	.w3(32'hbb040115),
	.w4(32'hbae7a2c8),
	.w5(32'hbaf2132c),
	.w6(32'hbaf5b93c),
	.w7(32'hbb124f32),
	.w8(32'hbb1f785e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18e969),
	.w1(32'h387dd0c8),
	.w2(32'h3a044363),
	.w3(32'hba0ed199),
	.w4(32'hb7aed56c),
	.w5(32'h38dc407d),
	.w6(32'hb9f1e5df),
	.w7(32'hb922c7c7),
	.w8(32'h3803fcfa),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2127),
	.w1(32'hbac2bf29),
	.w2(32'hbb0725be),
	.w3(32'hb9fffe28),
	.w4(32'hbaca1bed),
	.w5(32'hbaafbe50),
	.w6(32'hba418c05),
	.w7(32'hbae64f0f),
	.w8(32'hbb382f49),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04b69b),
	.w1(32'h39b26f7f),
	.w2(32'h3a190698),
	.w3(32'h39c20d5a),
	.w4(32'h39a06fe8),
	.w5(32'h3a471450),
	.w6(32'h3a150c71),
	.w7(32'h3a400af9),
	.w8(32'h3a8617f0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a450a38),
	.w1(32'hba89351d),
	.w2(32'hba70e989),
	.w3(32'h3a80c65e),
	.w4(32'hba1cf25a),
	.w5(32'hb9f5b049),
	.w6(32'h3a6724aa),
	.w7(32'hba9229c7),
	.w8(32'hba81c3cc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60ae47),
	.w1(32'hb9ae5e1b),
	.w2(32'hb90c25e0),
	.w3(32'hba279f9a),
	.w4(32'hb743112d),
	.w5(32'h3a69eb02),
	.w6(32'hba98b0d7),
	.w7(32'h38f64c74),
	.w8(32'h39e41e67),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d01412),
	.w1(32'hb98b27f0),
	.w2(32'h3876e850),
	.w3(32'hb8d3ceef),
	.w4(32'hba7e990f),
	.w5(32'hba2918ee),
	.w6(32'h39dd7fe2),
	.w7(32'hba7f163a),
	.w8(32'hba22c1a6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce8597),
	.w1(32'h3a506d06),
	.w2(32'h3a3a1a4b),
	.w3(32'hb8d8f28c),
	.w4(32'h3ab71d22),
	.w5(32'h3acef3a2),
	.w6(32'hba80a432),
	.w7(32'h3a866794),
	.w8(32'h3a814d2d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22f9b9),
	.w1(32'hbb3487e4),
	.w2(32'hbaa53de8),
	.w3(32'hbb3cc084),
	.w4(32'hbb47d2b3),
	.w5(32'hbb2a64bf),
	.w6(32'hbb7a5e72),
	.w7(32'hbb9fb95c),
	.w8(32'hbba247aa),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d322),
	.w1(32'hbb0e1907),
	.w2(32'hba4b5439),
	.w3(32'hbabe4c9b),
	.w4(32'hbb2c31ef),
	.w5(32'hba8cd4d9),
	.w6(32'hba90ef34),
	.w7(32'hbb272127),
	.w8(32'hbb5cfd06),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b16286),
	.w1(32'hbb4edcf4),
	.w2(32'hbadb0b7a),
	.w3(32'hba19d252),
	.w4(32'hbb349814),
	.w5(32'hbacb1b1c),
	.w6(32'hba0ece76),
	.w7(32'hbb86542f),
	.w8(32'hbb7b09a0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61f7e5),
	.w1(32'h3a485fea),
	.w2(32'h39d1cffb),
	.w3(32'hba9b4615),
	.w4(32'h3acd48c8),
	.w5(32'h3a23d890),
	.w6(32'hba894918),
	.w7(32'h3a6e417a),
	.w8(32'h3a19b22a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c12d6),
	.w1(32'h3a81e2f7),
	.w2(32'h3a5529ef),
	.w3(32'h3957e078),
	.w4(32'h39fd7504),
	.w5(32'h38ee9cea),
	.w6(32'h39b2dcc1),
	.w7(32'h39fa1265),
	.w8(32'h398088e3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9c26),
	.w1(32'h395be494),
	.w2(32'h3a46d9aa),
	.w3(32'h391a5b9b),
	.w4(32'h391438f3),
	.w5(32'h3a85545e),
	.w6(32'h39610136),
	.w7(32'h38ecfc59),
	.w8(32'h396a6716),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384f914d),
	.w1(32'h3aada59d),
	.w2(32'h3aae90d7),
	.w3(32'h39c74d7f),
	.w4(32'h3a64e667),
	.w5(32'h39f19bf8),
	.w6(32'h3972a788),
	.w7(32'hb873bc69),
	.w8(32'hb9d73592),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab1381),
	.w1(32'hbb1703f3),
	.w2(32'hbb744642),
	.w3(32'hbadeed47),
	.w4(32'hbb337f9e),
	.w5(32'hbb622524),
	.w6(32'hbae5d2b1),
	.w7(32'hbb5b29a0),
	.w8(32'hbb9605bf),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910485a),
	.w1(32'h3a3e3129),
	.w2(32'h3a0b2f8e),
	.w3(32'h38a46ad0),
	.w4(32'h39677d84),
	.w5(32'h3a0693fe),
	.w6(32'hb9548768),
	.w7(32'h399d379c),
	.w8(32'h39bf91bd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3be3e6),
	.w1(32'h3ab99712),
	.w2(32'hb99b5526),
	.w3(32'h3a3a88f3),
	.w4(32'h39fc82c1),
	.w5(32'hba8b4005),
	.w6(32'h394b091e),
	.w7(32'h38d769e9),
	.w8(32'hb9d485ea),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5e26f),
	.w1(32'hb8b32e69),
	.w2(32'hba71f070),
	.w3(32'hbab44f04),
	.w4(32'h39548f17),
	.w5(32'h39d0b89e),
	.w6(32'hba312247),
	.w7(32'h3a46346f),
	.w8(32'h3a22ef37),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911ba53),
	.w1(32'hb8a9bdf3),
	.w2(32'hb91be681),
	.w3(32'hb957990d),
	.w4(32'hb93ccc85),
	.w5(32'hb9b4c063),
	.w6(32'hb86944af),
	.w7(32'hb818b939),
	.w8(32'hb9b26d9f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68be32),
	.w1(32'hb950dad4),
	.w2(32'hba3ae426),
	.w3(32'h3a97ce8b),
	.w4(32'hb8e58063),
	.w5(32'hb927805e),
	.w6(32'h3a812707),
	.w7(32'h39bf9382),
	.w8(32'hb9aa21f1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a74587),
	.w1(32'h390dcb5e),
	.w2(32'h379aaf18),
	.w3(32'hb968d51a),
	.w4(32'hb88f9523),
	.w5(32'hb925cb77),
	.w6(32'h383ea0c2),
	.w7(32'hb9c34e43),
	.w8(32'hb9ee373a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad872fa),
	.w1(32'hbb82eeae),
	.w2(32'hbb9d9f22),
	.w3(32'hbb9b5328),
	.w4(32'hbbac6f52),
	.w5(32'hbbcac4b3),
	.w6(32'hbbbf1038),
	.w7(32'hbc0d0f73),
	.w8(32'hbbd1e60b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50a211),
	.w1(32'hba623175),
	.w2(32'hbaa60b97),
	.w3(32'hba0962ff),
	.w4(32'hba1004d0),
	.w5(32'hbab02f95),
	.w6(32'hb9caf5b0),
	.w7(32'hba1adaad),
	.w8(32'hba6eed78),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb692ab4),
	.w1(32'h387846a2),
	.w2(32'h3b5d71f7),
	.w3(32'hbb3e0e03),
	.w4(32'hb9b3f338),
	.w5(32'h3a566d7f),
	.w6(32'hbbe8242d),
	.w7(32'hbaf3420d),
	.w8(32'hba75068d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule