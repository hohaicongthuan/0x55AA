module layer_10_featuremap_244(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbdfb),
	.w1(32'hbbc822a1),
	.w2(32'hbb9c8efa),
	.w3(32'h3b6cdf0e),
	.w4(32'hb94479f0),
	.w5(32'hbae5df08),
	.w6(32'hb8327d43),
	.w7(32'hbb3f7575),
	.w8(32'hbb3044c0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7736c),
	.w1(32'hba3d1d14),
	.w2(32'hbaef7505),
	.w3(32'h3afa423d),
	.w4(32'h39379a9e),
	.w5(32'hbb6deff0),
	.w6(32'hbad5ace6),
	.w7(32'h3bde4ad7),
	.w8(32'hbba87c55),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aa3e9),
	.w1(32'h3af576e8),
	.w2(32'h3bd9e61d),
	.w3(32'hbb392b6c),
	.w4(32'hbae19300),
	.w5(32'h3a559eb6),
	.w6(32'hba8ccb8a),
	.w7(32'hbb6ac3ac),
	.w8(32'h3b8c4992),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dc0ad),
	.w1(32'hbab4d286),
	.w2(32'hbb8213e9),
	.w3(32'h3a898077),
	.w4(32'h3aa427c0),
	.w5(32'hbb746932),
	.w6(32'h3c0137b7),
	.w7(32'h3a967e35),
	.w8(32'hbbf4f3a5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c604d53),
	.w1(32'h3bdf782f),
	.w2(32'h3b0d56f4),
	.w3(32'hbc0312c5),
	.w4(32'hbc0eadb4),
	.w5(32'h3b36aa7e),
	.w6(32'hbc937235),
	.w7(32'hbc06cf22),
	.w8(32'h3aa9990b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a271),
	.w1(32'hbb7e26bc),
	.w2(32'hbb936c45),
	.w3(32'h3bc7e433),
	.w4(32'h3b4c5f61),
	.w5(32'h3b5b7b11),
	.w6(32'h3bf0bb91),
	.w7(32'h3b26c397),
	.w8(32'h3b84ca52),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239451),
	.w1(32'hbb3e644a),
	.w2(32'hbbaab466),
	.w3(32'h3ba39ca5),
	.w4(32'h3b86b35b),
	.w5(32'h3a994bf5),
	.w6(32'h3bb081a7),
	.w7(32'h3b88bb4f),
	.w8(32'h3bea0859),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81aa70),
	.w1(32'h3b03843f),
	.w2(32'h3af0bd36),
	.w3(32'h392210e3),
	.w4(32'hbaec349b),
	.w5(32'h3b894100),
	.w6(32'h3c04479d),
	.w7(32'hbb6e254d),
	.w8(32'h3b169adf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace6519),
	.w1(32'h3a56416b),
	.w2(32'h3be41319),
	.w3(32'h3b649f50),
	.w4(32'h3b92e5d1),
	.w5(32'h3af12e58),
	.w6(32'h3bc567e8),
	.w7(32'h3bbaa5dc),
	.w8(32'h3ac6d7a1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45902e),
	.w1(32'h38aa64ce),
	.w2(32'hba93272c),
	.w3(32'h3bacd1a8),
	.w4(32'h3b07f254),
	.w5(32'h3b51e625),
	.w6(32'h3c0157bd),
	.w7(32'h3b1b3ab9),
	.w8(32'h3bf1ce25),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb38265),
	.w1(32'hbb31f38d),
	.w2(32'hbb91ddc6),
	.w3(32'h3baacbb9),
	.w4(32'h3b2cbfbc),
	.w5(32'hba802d78),
	.w6(32'h3c35f8b5),
	.w7(32'h3ab7bdb8),
	.w8(32'hbb8dd54a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00602f),
	.w1(32'hbb825284),
	.w2(32'hbb2d5930),
	.w3(32'h3b1e8373),
	.w4(32'hbb4a14d9),
	.w5(32'hbb0366af),
	.w6(32'h39585780),
	.w7(32'hbbe77fa6),
	.w8(32'h3b83385f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007ce1),
	.w1(32'h3bf1298a),
	.w2(32'h3c238614),
	.w3(32'hbad1624d),
	.w4(32'hbb27009b),
	.w5(32'hb8a0d9c3),
	.w6(32'h3b601692),
	.w7(32'h3a51cb36),
	.w8(32'h381e1fdd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ef0ea),
	.w1(32'h3af07772),
	.w2(32'hbb91eb16),
	.w3(32'h3b23e3dd),
	.w4(32'hbb1345c4),
	.w5(32'h3aeb1496),
	.w6(32'h3bad8c8f),
	.w7(32'h3bd084ca),
	.w8(32'h3b7789cb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ea986),
	.w1(32'hbb30382f),
	.w2(32'hbac9e599),
	.w3(32'h3b6cb0b2),
	.w4(32'h3adb00d7),
	.w5(32'hbb3c291d),
	.w6(32'h3c266729),
	.w7(32'h3a55fa3e),
	.w8(32'hbb7e1668),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f9e6),
	.w1(32'h3b1f616c),
	.w2(32'h3a18755a),
	.w3(32'hbb3b5a59),
	.w4(32'hba80f278),
	.w5(32'hbb28c578),
	.w6(32'h3b0bdb8b),
	.w7(32'h3ae23fcc),
	.w8(32'hbbbe91ac),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8992),
	.w1(32'hbc489198),
	.w2(32'hbc1bb94d),
	.w3(32'hbac783bd),
	.w4(32'h39e8d73e),
	.w5(32'hbafa29d7),
	.w6(32'h3ba25b11),
	.w7(32'hbae793aa),
	.w8(32'h3a1214b5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952bb4),
	.w1(32'h3ba265d7),
	.w2(32'h3c0db0c7),
	.w3(32'hb9412be3),
	.w4(32'hbb79c0ff),
	.w5(32'h3b4d041a),
	.w6(32'hbb60766b),
	.w7(32'hbbb9c43d),
	.w8(32'h3b06222e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d3761),
	.w1(32'h3c860ac0),
	.w2(32'h3bb4b6ce),
	.w3(32'h3b453ffe),
	.w4(32'h3ae9d337),
	.w5(32'hbbfc3e9d),
	.w6(32'h3b761091),
	.w7(32'h3bc95159),
	.w8(32'h3aa32c43),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088520),
	.w1(32'h3c0a6aa3),
	.w2(32'hba600db0),
	.w3(32'hba465218),
	.w4(32'hbbe14fd3),
	.w5(32'h3aab87ad),
	.w6(32'hbb8df423),
	.w7(32'hbba4bcee),
	.w8(32'h3a0d8960),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290b45),
	.w1(32'h3b17a6ac),
	.w2(32'hbbb071e3),
	.w3(32'hbb37bd76),
	.w4(32'hb99d4f5c),
	.w5(32'h3b51c417),
	.w6(32'h3b0466e6),
	.w7(32'h3c0af9c9),
	.w8(32'h3ac256a2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8922c),
	.w1(32'hbb9a6f75),
	.w2(32'hbb54717b),
	.w3(32'hbb9a918f),
	.w4(32'h3989a2cc),
	.w5(32'hbbe9fdc4),
	.w6(32'hba737243),
	.w7(32'hb883e75c),
	.w8(32'hbb9a54e5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd6c7a),
	.w1(32'h3b182913),
	.w2(32'h3b1df68b),
	.w3(32'hbc14ceda),
	.w4(32'hba901723),
	.w5(32'hb9d49b87),
	.w6(32'hbbfb3084),
	.w7(32'hbb499272),
	.w8(32'h3a7e3ff2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245496),
	.w1(32'h3a873d32),
	.w2(32'h39e1f1d2),
	.w3(32'h3b98bc79),
	.w4(32'hbb54a93c),
	.w5(32'hbc07bea1),
	.w6(32'h3bf226af),
	.w7(32'hbb790f75),
	.w8(32'hbc0e0827),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e73d8),
	.w1(32'h3c91207f),
	.w2(32'h3c16a15a),
	.w3(32'hbbc87699),
	.w4(32'hbb11c606),
	.w5(32'h3b5c44f6),
	.w6(32'hbca611d6),
	.w7(32'hbb808f8a),
	.w8(32'h3be01f8c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68dfb3),
	.w1(32'hb91ff7b2),
	.w2(32'hbb9d7140),
	.w3(32'hbaea2e78),
	.w4(32'hba24f9a7),
	.w5(32'h3a6895e5),
	.w6(32'h3bf70508),
	.w7(32'hba857bfe),
	.w8(32'hbb0866d9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7da447),
	.w1(32'hbbb18cc9),
	.w2(32'hbb97211d),
	.w3(32'hb9f18ecb),
	.w4(32'h3a9a1797),
	.w5(32'h3a8dd33e),
	.w6(32'h3baa6ad7),
	.w7(32'h3a8b9f96),
	.w8(32'hbba61fb2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3c50),
	.w1(32'hbb3c6cd2),
	.w2(32'h3ae17e45),
	.w3(32'h3b14f290),
	.w4(32'h3aecf412),
	.w5(32'hbbf100e9),
	.w6(32'hbb172111),
	.w7(32'h3b805adb),
	.w8(32'hba30973d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16ce04),
	.w1(32'h3ab0201c),
	.w2(32'hbab4da46),
	.w3(32'hbb198e0b),
	.w4(32'h3914647e),
	.w5(32'hbba5d692),
	.w6(32'hbc081f7f),
	.w7(32'hbb38c53a),
	.w8(32'hbb31dcb7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897103),
	.w1(32'h3b1ee788),
	.w2(32'hbb0e15c7),
	.w3(32'h3a411094),
	.w4(32'h3a1c192d),
	.w5(32'h3b22f20f),
	.w6(32'h3b309efd),
	.w7(32'h3a8dc35e),
	.w8(32'hbbe84b15),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133ad6),
	.w1(32'h3cbca853),
	.w2(32'h3bd82f0d),
	.w3(32'h3b2d5567),
	.w4(32'hbb4f9316),
	.w5(32'hbbba6c50),
	.w6(32'hbcabd579),
	.w7(32'hbbfeb596),
	.w8(32'hbc5c0a7e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7491e1),
	.w1(32'h36e7fe56),
	.w2(32'h3b0dcbef),
	.w3(32'hba98ed52),
	.w4(32'hbb4dd9f1),
	.w5(32'h3a9e6051),
	.w6(32'hbad407ed),
	.w7(32'hbc1a5226),
	.w8(32'h3a3857a0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedaf88),
	.w1(32'h3c3ca40d),
	.w2(32'hbad06bea),
	.w3(32'h3b8739c9),
	.w4(32'h3af4fa38),
	.w5(32'hb81514e3),
	.w6(32'hbc8ceb52),
	.w7(32'h3ab21e04),
	.w8(32'h3b871596),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4200d),
	.w1(32'hbba0ccfc),
	.w2(32'h3b4e253d),
	.w3(32'h3a1c02de),
	.w4(32'hbaa302d6),
	.w5(32'h3bae6a72),
	.w6(32'hbbb519c2),
	.w7(32'hbab83404),
	.w8(32'h3c94fa8d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6133b5),
	.w1(32'h3c170b3c),
	.w2(32'h3a3ffc48),
	.w3(32'hbb0b94c3),
	.w4(32'hba417087),
	.w5(32'hbb876c0a),
	.w6(32'h39cb540a),
	.w7(32'hbbf7e8d3),
	.w8(32'h3b860397),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8792d8),
	.w1(32'hbae10fd6),
	.w2(32'h3c3cbba0),
	.w3(32'hbba04f01),
	.w4(32'hbbb6c66c),
	.w5(32'h3a99897a),
	.w6(32'hbb097122),
	.w7(32'h3c1b1b96),
	.w8(32'hbbd43290),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4437e7),
	.w1(32'h3c7671bd),
	.w2(32'h3c0481dc),
	.w3(32'h3bc792e1),
	.w4(32'h3ab9bd3c),
	.w5(32'h3c1130a7),
	.w6(32'hbcf6e11f),
	.w7(32'hbad31469),
	.w8(32'h3b8d51fc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6dd2),
	.w1(32'h398547cf),
	.w2(32'h3b575182),
	.w3(32'h3b9f9069),
	.w4(32'h3b8a06ea),
	.w5(32'hba4f3787),
	.w6(32'h3c641bcc),
	.w7(32'h3c4f6cdc),
	.w8(32'hbb3e4cae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d6d7),
	.w1(32'h3ab1ca45),
	.w2(32'hba04fbf8),
	.w3(32'h3bdacaf6),
	.w4(32'h3ac59d20),
	.w5(32'h3a53f404),
	.w6(32'hbbe6ab0f),
	.w7(32'hbb2349bb),
	.w8(32'h3af0431a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc358efe),
	.w1(32'hbc40d81a),
	.w2(32'hbbe4d00c),
	.w3(32'hbc1ecb60),
	.w4(32'h393528ec),
	.w5(32'hbb1b82ac),
	.w6(32'h3b21aa90),
	.w7(32'h37329af7),
	.w8(32'hbb4fdc01),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b646b77),
	.w1(32'hbab0021b),
	.w2(32'h3c16eb96),
	.w3(32'hba587792),
	.w4(32'hbb5435b1),
	.w5(32'hb985b57f),
	.w6(32'hbc0241d1),
	.w7(32'h3b8af739),
	.w8(32'h3b4d8d73),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0dcff),
	.w1(32'hbb7ec80d),
	.w2(32'hbbb5af8f),
	.w3(32'hbb9cfedb),
	.w4(32'h3969e5ca),
	.w5(32'hb915c008),
	.w6(32'h3badc1d3),
	.w7(32'hbacf8f08),
	.w8(32'h3b27cce0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cd7b3),
	.w1(32'h3c5124b5),
	.w2(32'h3c7b099d),
	.w3(32'hbb88df8d),
	.w4(32'hbaece7b2),
	.w5(32'h3aa46407),
	.w6(32'h3b80c51d),
	.w7(32'h3bbe7b9a),
	.w8(32'h3b1a2585),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a036),
	.w1(32'h3b503e85),
	.w2(32'hbbbc0580),
	.w3(32'h3a99319a),
	.w4(32'hbba9e88d),
	.w5(32'h3ba1592a),
	.w6(32'h3cc1e364),
	.w7(32'h3bf5cf2f),
	.w8(32'h3bf66042),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83d597),
	.w1(32'hba3701d7),
	.w2(32'h3b916bab),
	.w3(32'h3bc2263f),
	.w4(32'h3c12377a),
	.w5(32'h3b5e3e78),
	.w6(32'h3c1c1df1),
	.w7(32'h3c2c0597),
	.w8(32'h3aa8e6e7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29e0c3),
	.w1(32'hbc305657),
	.w2(32'hbc06b2d6),
	.w3(32'h3bdd40d7),
	.w4(32'h39032054),
	.w5(32'h3bc9bf3d),
	.w6(32'h3bb36fc2),
	.w7(32'hbae9d85c),
	.w8(32'h3b9fb0b0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d17a),
	.w1(32'hbc16a84c),
	.w2(32'hbb6f89db),
	.w3(32'h3bdbf153),
	.w4(32'h3a1e8e26),
	.w5(32'h3b1d2be8),
	.w6(32'h3c489bc4),
	.w7(32'h3bd86cf7),
	.w8(32'hbb5f4251),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe685c),
	.w1(32'h3a954f76),
	.w2(32'h3bcbb9e1),
	.w3(32'h3b40baec),
	.w4(32'h3bd93942),
	.w5(32'h3af20f23),
	.w6(32'h3a94a845),
	.w7(32'h3b40f8f5),
	.w8(32'h3bacc950),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75381),
	.w1(32'h3a860b57),
	.w2(32'h3b627751),
	.w3(32'hbac16c96),
	.w4(32'hbb96bf9d),
	.w5(32'h3bc77cf2),
	.w6(32'h3be38b9f),
	.w7(32'h3bc080c4),
	.w8(32'h3b9dc421),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ef97e),
	.w1(32'hbb2241cd),
	.w2(32'hbae7aafb),
	.w3(32'hbafe6333),
	.w4(32'h3b6409c4),
	.w5(32'hbbae7c44),
	.w6(32'hba9affa4),
	.w7(32'h3b292709),
	.w8(32'hbc3384a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31fa12),
	.w1(32'h3be6d6b7),
	.w2(32'h3c0a84bd),
	.w3(32'hbb072a29),
	.w4(32'h3b1b3120),
	.w5(32'hbbebaa85),
	.w6(32'hbc529cf1),
	.w7(32'h39dca234),
	.w8(32'hbb006810),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835d38),
	.w1(32'h3b9d994b),
	.w2(32'hbb85198b),
	.w3(32'hbbd9767c),
	.w4(32'hbaba7491),
	.w5(32'hb9f21624),
	.w6(32'h3a0c37f2),
	.w7(32'h3ac0b3bb),
	.w8(32'hbb831b8b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940cb83),
	.w1(32'h3c0bcc31),
	.w2(32'h3be95d99),
	.w3(32'hbaab598d),
	.w4(32'hbb89731a),
	.w5(32'hbb868923),
	.w6(32'hbbd192c8),
	.w7(32'h3b9547bc),
	.w8(32'hbb3be472),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91fdab),
	.w1(32'h3b5c7280),
	.w2(32'hb96dc4a6),
	.w3(32'h3bf059e0),
	.w4(32'h3bd055de),
	.w5(32'hbc27c0fb),
	.w6(32'h3be769d7),
	.w7(32'h3aaf580d),
	.w8(32'hbb564cb3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90e31f),
	.w1(32'h3c06a94e),
	.w2(32'hbbace8fb),
	.w3(32'hbbeb75ce),
	.w4(32'hbc1125e6),
	.w5(32'hbb1e3b03),
	.w6(32'hbc26689d),
	.w7(32'hbc332d63),
	.w8(32'h3ac87703),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07745c),
	.w1(32'h3b1794c3),
	.w2(32'h3aec5184),
	.w3(32'hbb888c88),
	.w4(32'hbb639231),
	.w5(32'hbb30d097),
	.w6(32'hbc0d5946),
	.w7(32'hbc1c1ba3),
	.w8(32'hbaeb7986),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841a3a),
	.w1(32'hbb3b8a94),
	.w2(32'h3b7260e2),
	.w3(32'hbaaf6b55),
	.w4(32'hb89a4ee6),
	.w5(32'hbc03d254),
	.w6(32'hbb8f0f71),
	.w7(32'h39038b22),
	.w8(32'hbaa3a1b5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b182),
	.w1(32'h3c0f97ba),
	.w2(32'h3afe872f),
	.w3(32'h3bde36db),
	.w4(32'h3be18e99),
	.w5(32'h3bb7fbf8),
	.w6(32'h3c346e11),
	.w7(32'h3bb6becd),
	.w8(32'h3b9fbbce),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb5a05),
	.w1(32'hba8e65cd),
	.w2(32'hb8191241),
	.w3(32'hbaf358eb),
	.w4(32'hb8331fb8),
	.w5(32'h3bed605c),
	.w6(32'h39a06f17),
	.w7(32'h3a28acee),
	.w8(32'hb9f69967),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90139),
	.w1(32'hbb72d0e6),
	.w2(32'hbb88e5fc),
	.w3(32'hbb3bedc5),
	.w4(32'h3b7a6151),
	.w5(32'h3ab0378e),
	.w6(32'hbb2cffc4),
	.w7(32'h3bf76119),
	.w8(32'hba7f6e85),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9e1aa),
	.w1(32'hba9a1c0c),
	.w2(32'hbaa9ee7e),
	.w3(32'h3c248f74),
	.w4(32'h3b9a3805),
	.w5(32'h3a85c639),
	.w6(32'hba68cfa7),
	.w7(32'h3a855963),
	.w8(32'h3b5b5b98),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46c21f),
	.w1(32'hbb722496),
	.w2(32'hbc22a95f),
	.w3(32'h3b99e443),
	.w4(32'h3b522a92),
	.w5(32'h3a306d2d),
	.w6(32'h3c24ff80),
	.w7(32'h3a8d9f6e),
	.w8(32'h3c49ca93),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c588627),
	.w1(32'h3ccff26c),
	.w2(32'h3b80b9ec),
	.w3(32'hbc41eb74),
	.w4(32'hbc0ebf68),
	.w5(32'hbbbaa41c),
	.w6(32'hbbd976f6),
	.w7(32'h3af9f1a7),
	.w8(32'h3b45135a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acef196),
	.w1(32'h3afd7e2e),
	.w2(32'h3b51ab5a),
	.w3(32'hbbcc3417),
	.w4(32'hba82fd74),
	.w5(32'h3bb419cf),
	.w6(32'hbbf631b6),
	.w7(32'hbbd2d3cc),
	.w8(32'h3c9bdac5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e7ccc),
	.w1(32'h3c7e643a),
	.w2(32'h3ad4084b),
	.w3(32'h3b1689a6),
	.w4(32'hbac16f92),
	.w5(32'hbbf9eb71),
	.w6(32'hba859376),
	.w7(32'hbbbd6507),
	.w8(32'hbc0635ef),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094e25),
	.w1(32'h3c70af30),
	.w2(32'h3b38a0cf),
	.w3(32'hbb808c2b),
	.w4(32'hbc0d0bfc),
	.w5(32'hb9b34913),
	.w6(32'hbc6cf5df),
	.w7(32'hbb46df1e),
	.w8(32'h3bb455c9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e1c6f),
	.w1(32'hbb23516e),
	.w2(32'hbbca3802),
	.w3(32'h3b5fc334),
	.w4(32'h3b6c056f),
	.w5(32'h3acdb1bd),
	.w6(32'h3be1ffd4),
	.w7(32'hbb8fb277),
	.w8(32'h3b87a199),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2cde9),
	.w1(32'hbc458be2),
	.w2(32'hbbcc570b),
	.w3(32'h3b92bd51),
	.w4(32'hbabbce84),
	.w5(32'hba939c7b),
	.w6(32'h3c9396f4),
	.w7(32'h394d92eb),
	.w8(32'h3b2a9961),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3470),
	.w1(32'hbbb75ae7),
	.w2(32'hbbc3d322),
	.w3(32'h394fa7c8),
	.w4(32'hbc0d5756),
	.w5(32'h3b8d892a),
	.w6(32'hb73c3b54),
	.w7(32'hbb8b5655),
	.w8(32'h3b217813),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29de20),
	.w1(32'hbbbc55ec),
	.w2(32'h3c0ddadd),
	.w3(32'h3b99d42c),
	.w4(32'h3bb6c806),
	.w5(32'hbb0fa703),
	.w6(32'h3c7757fa),
	.w7(32'h3bb5f052),
	.w8(32'h3ba1b180),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b558174),
	.w1(32'hbb91cb93),
	.w2(32'h372a5042),
	.w3(32'h3a8dab95),
	.w4(32'hba9c0549),
	.w5(32'h38bf8732),
	.w6(32'h3a96ceeb),
	.w7(32'h3b5aab65),
	.w8(32'hbb5e804f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7c98b),
	.w1(32'hbaa97e55),
	.w2(32'hbc0ed3b2),
	.w3(32'hbb8d89c4),
	.w4(32'h39bdeef2),
	.w5(32'hba3cac9b),
	.w6(32'h3a6435bb),
	.w7(32'hbb9c45cb),
	.w8(32'h3be6371b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1334a),
	.w1(32'h39a9049d),
	.w2(32'hbb556e56),
	.w3(32'h3b31dab2),
	.w4(32'h3bc747d7),
	.w5(32'hbbaf99bc),
	.w6(32'h3b850b8c),
	.w7(32'h3b11f516),
	.w8(32'h3a27a4aa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5d5e0),
	.w1(32'h3af0ba69),
	.w2(32'h39f1c75f),
	.w3(32'h3a879eed),
	.w4(32'h3a780c87),
	.w5(32'hba91dd0d),
	.w6(32'hbb3fa9f5),
	.w7(32'h3afdf5ab),
	.w8(32'h3b7958db),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19dbe2),
	.w1(32'hbbcd3155),
	.w2(32'hbbcfb98b),
	.w3(32'h3b8544eb),
	.w4(32'h3b4f6672),
	.w5(32'hbb7a3612),
	.w6(32'h3c183766),
	.w7(32'hba39dafa),
	.w8(32'h39d98691),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf35be3),
	.w1(32'h3bcdf571),
	.w2(32'h3c2fea39),
	.w3(32'hbb5e37e2),
	.w4(32'hbb72ca37),
	.w5(32'hbb08b1da),
	.w6(32'h3a45cc8e),
	.w7(32'h3a7f6292),
	.w8(32'hbb897163),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1869e3),
	.w1(32'h3c0ae8e2),
	.w2(32'h3b9cbdaa),
	.w3(32'hba93af03),
	.w4(32'hbb694807),
	.w5(32'h3a83be67),
	.w6(32'hbbc7c184),
	.w7(32'hba3f0f10),
	.w8(32'h3a9b1d2a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c245b3e),
	.w1(32'h3bd5d508),
	.w2(32'hba753d27),
	.w3(32'h3c1d08de),
	.w4(32'hbb25efe1),
	.w5(32'h3b9206bb),
	.w6(32'h3bffb2cd),
	.w7(32'h3a765690),
	.w8(32'h3b82d3d0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03e97d),
	.w1(32'hbc158df1),
	.w2(32'hbbff7c70),
	.w3(32'h3a8a4f9c),
	.w4(32'h3b211968),
	.w5(32'h3b557b8f),
	.w6(32'h3c19a0bb),
	.w7(32'h3ac4d54d),
	.w8(32'h3b1ef1ab),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8138),
	.w1(32'hbc0b2541),
	.w2(32'hbb9b382c),
	.w3(32'h3bb92cd0),
	.w4(32'h3bb021e4),
	.w5(32'h3b54e756),
	.w6(32'h3be76c9b),
	.w7(32'h3a183d1b),
	.w8(32'h3c38b491),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae524),
	.w1(32'hbbaf3966),
	.w2(32'hbba530c5),
	.w3(32'hbbabfaa2),
	.w4(32'h3b651cb9),
	.w5(32'hba5ce87a),
	.w6(32'h3c8eac14),
	.w7(32'h3bd62405),
	.w8(32'hba7d2899),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93408a),
	.w1(32'h3bafc1a6),
	.w2(32'h3c213b9a),
	.w3(32'hbae2dee4),
	.w4(32'hb9cef12a),
	.w5(32'h3b90ec9c),
	.w6(32'hbba20cae),
	.w7(32'h3b25a2ea),
	.w8(32'h3bcf9219),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7017c9),
	.w1(32'h3b34e491),
	.w2(32'h3b40008f),
	.w3(32'h3ba555b1),
	.w4(32'hbbca0658),
	.w5(32'h3be55f2e),
	.w6(32'h39c5e307),
	.w7(32'hbb983a47),
	.w8(32'h3b8d9e52),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f25bb),
	.w1(32'hbb564f01),
	.w2(32'hbb6ec556),
	.w3(32'h3b92c87c),
	.w4(32'h3b6f8f06),
	.w5(32'hbb573774),
	.w6(32'h3c926754),
	.w7(32'h3ad24875),
	.w8(32'hbb73e369),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936c684),
	.w1(32'h3a8a3a03),
	.w2(32'h3bb86201),
	.w3(32'hba401594),
	.w4(32'hbb911319),
	.w5(32'h3bc25474),
	.w6(32'hbc047f21),
	.w7(32'hbba2f39f),
	.w8(32'h3b9262bd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38b93e),
	.w1(32'hbc43c2a7),
	.w2(32'hbc5c5c80),
	.w3(32'h3bde86ff),
	.w4(32'hbb29e215),
	.w5(32'hbb20ad93),
	.w6(32'h3be83295),
	.w7(32'h3ba3a9fa),
	.w8(32'h3b4de701),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf847ca),
	.w1(32'hbb89112d),
	.w2(32'hbba7e5c1),
	.w3(32'h3ba06847),
	.w4(32'h3b83e631),
	.w5(32'hbc51c729),
	.w6(32'h3c779fae),
	.w7(32'hba7f7eba),
	.w8(32'hbaaef8e9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e9d71),
	.w1(32'h3c66688e),
	.w2(32'h3b42c1a9),
	.w3(32'hbc470d8b),
	.w4(32'hbc1c8c89),
	.w5(32'h3b3e1015),
	.w6(32'hbb289ace),
	.w7(32'hbb4ba57c),
	.w8(32'hb99e3d7d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ad31),
	.w1(32'hbb060347),
	.w2(32'h3adffdcd),
	.w3(32'h3bcd41db),
	.w4(32'h3bc5f2d2),
	.w5(32'h39422387),
	.w6(32'h3bbfc313),
	.w7(32'h3b8ec4a2),
	.w8(32'h3a52a69a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c780d),
	.w1(32'hba28bd12),
	.w2(32'h3b1d8826),
	.w3(32'hbba5def0),
	.w4(32'hbba46f2e),
	.w5(32'hbabb3509),
	.w6(32'h3abc8053),
	.w7(32'h3baa83fb),
	.w8(32'h3b574016),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89f5b6),
	.w1(32'hbbad704a),
	.w2(32'h3a80741e),
	.w3(32'hba157bab),
	.w4(32'hba7c2c68),
	.w5(32'h3bc3af5e),
	.w6(32'h3ac711c2),
	.w7(32'h3acb3677),
	.w8(32'h3be1bffd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08613),
	.w1(32'h388dd1b3),
	.w2(32'hbc156569),
	.w3(32'h3b801ead),
	.w4(32'hba70b1fa),
	.w5(32'hb9f661d5),
	.w6(32'h3bba91ea),
	.w7(32'hbb8021cb),
	.w8(32'hbbe2306e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41e457),
	.w1(32'hbaf7c15a),
	.w2(32'hbaf25f9b),
	.w3(32'h3b650298),
	.w4(32'hbbde7536),
	.w5(32'hb8de34fa),
	.w6(32'hbbc89339),
	.w7(32'hbbd7b0e9),
	.w8(32'h3b27ce1a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306488),
	.w1(32'hbc3a060d),
	.w2(32'hbc6614f3),
	.w3(32'hbb1ec509),
	.w4(32'hbb273f28),
	.w5(32'h3bc2f9d0),
	.w6(32'h3b28da12),
	.w7(32'hbac42475),
	.w8(32'h3c1b2d42),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f5c1),
	.w1(32'h3b3f0247),
	.w2(32'h3ac69818),
	.w3(32'h3af6749e),
	.w4(32'hbaf73007),
	.w5(32'h3a939605),
	.w6(32'h3c2a0715),
	.w7(32'h3bda9ed9),
	.w8(32'hbc713a23),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a193341),
	.w1(32'hba9760ac),
	.w2(32'h3b5a4ae0),
	.w3(32'h3a18f583),
	.w4(32'hb8856687),
	.w5(32'h3b6b8e79),
	.w6(32'hbb68c2b4),
	.w7(32'hbc3898f1),
	.w8(32'h3a80c27d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba76e84),
	.w1(32'hbc3af721),
	.w2(32'hbc2df6ed),
	.w3(32'h3ad68721),
	.w4(32'h3c035386),
	.w5(32'hb949b7b3),
	.w6(32'h3b62a7c4),
	.w7(32'h3b59df24),
	.w8(32'hbb3fbb4e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc50d30),
	.w1(32'h3c531888),
	.w2(32'hb9cb74f8),
	.w3(32'h3c188007),
	.w4(32'hbae85aed),
	.w5(32'h3b0e4814),
	.w6(32'hbbf7e7c2),
	.w7(32'hbba79151),
	.w8(32'h3ada2c82),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b664304),
	.w1(32'h3afeddf8),
	.w2(32'h3a6f911c),
	.w3(32'h3aef85dc),
	.w4(32'h3adcaf15),
	.w5(32'hb96dbf81),
	.w6(32'h3a895be2),
	.w7(32'h399ed1ba),
	.w8(32'hba5b4c82),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb132705),
	.w1(32'h3aa08580),
	.w2(32'h3abef885),
	.w3(32'hba9229fe),
	.w4(32'hbb015fa0),
	.w5(32'h3a95354c),
	.w6(32'hbb5a6ee0),
	.w7(32'h3a1f4102),
	.w8(32'h3b219b6b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f0f9c),
	.w1(32'hba930c78),
	.w2(32'hbb085b66),
	.w3(32'h3ac35490),
	.w4(32'hb9ec7f4c),
	.w5(32'h3aa71cd9),
	.w6(32'h3b4af413),
	.w7(32'h3aa4b9aa),
	.w8(32'h38936456),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ccbc1),
	.w1(32'h3b107728),
	.w2(32'h3b4081fe),
	.w3(32'hb8d678bb),
	.w4(32'hba53798b),
	.w5(32'hbaa6c5e1),
	.w6(32'h3a0753dd),
	.w7(32'hba2258db),
	.w8(32'hb9243496),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7359d),
	.w1(32'h3b4f49a7),
	.w2(32'h3a37dc52),
	.w3(32'hb999aab2),
	.w4(32'h3b4bc14d),
	.w5(32'hbae330d0),
	.w6(32'h3b7fc8c5),
	.w7(32'h3b46797c),
	.w8(32'hbafaa6cd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab78303),
	.w1(32'hbafc434d),
	.w2(32'hb9ce928f),
	.w3(32'hba8b5daa),
	.w4(32'hba45e963),
	.w5(32'h3aca87be),
	.w6(32'hbb45bc82),
	.w7(32'hba73c590),
	.w8(32'h39ac06ba),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a825ac5),
	.w1(32'h3ad56fc9),
	.w2(32'h3b0e8acd),
	.w3(32'h3ae024ce),
	.w4(32'h3a88567f),
	.w5(32'h3b025e30),
	.w6(32'h3a30140c),
	.w7(32'h3af4091e),
	.w8(32'hb91cfb37),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec2349),
	.w1(32'h3aa964d7),
	.w2(32'h3aa31dfc),
	.w3(32'h3a3b387c),
	.w4(32'h3934c1ad),
	.w5(32'hb8fbe2ef),
	.w6(32'hb9357e54),
	.w7(32'h3a0e37f7),
	.w8(32'h3a8686d0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995aba8),
	.w1(32'hbaa3ba68),
	.w2(32'hbb119ab2),
	.w3(32'h3ac93ff2),
	.w4(32'h38be16da),
	.w5(32'h39639f72),
	.w6(32'h3ae49428),
	.w7(32'hbaf1bc34),
	.w8(32'h39b130a1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58cd20),
	.w1(32'hba38d641),
	.w2(32'h3998356f),
	.w3(32'hb9bbe635),
	.w4(32'h3ae56a28),
	.w5(32'h3b9fe5fb),
	.w6(32'h3a3e5dfa),
	.w7(32'h3a57c70f),
	.w8(32'h3b9c64a7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73a21),
	.w1(32'h3b4325a4),
	.w2(32'h3b422cd8),
	.w3(32'h3b684f2a),
	.w4(32'h3b4ed680),
	.w5(32'h3a6322dc),
	.w6(32'h3b383b73),
	.w7(32'h3b0448ce),
	.w8(32'h3a25da67),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c370b),
	.w1(32'hbaaf357b),
	.w2(32'hb7ebd390),
	.w3(32'h3a8bb819),
	.w4(32'h3aba963c),
	.w5(32'hba916c69),
	.w6(32'hbad743e9),
	.w7(32'hbac8d164),
	.w8(32'hbab9f60e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ac498),
	.w1(32'hba63c7f8),
	.w2(32'hba3f1996),
	.w3(32'hba5688bf),
	.w4(32'hba902d51),
	.w5(32'hba5c4f30),
	.w6(32'hbb647730),
	.w7(32'hba0c63e7),
	.w8(32'hba857bae),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24bfe),
	.w1(32'hba997192),
	.w2(32'hb7f932ef),
	.w3(32'hba62b771),
	.w4(32'hba68654d),
	.w5(32'h3a8fe019),
	.w6(32'h3a08cd3d),
	.w7(32'hba31c96f),
	.w8(32'h39fa57a0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63d524),
	.w1(32'h39decac6),
	.w2(32'hba905a25),
	.w3(32'hb81a409d),
	.w4(32'h3a49ce52),
	.w5(32'hba6f60ed),
	.w6(32'h3a69925a),
	.w7(32'hb8441650),
	.w8(32'hba614c49),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b6a4),
	.w1(32'h3b24a5d7),
	.w2(32'h3b090233),
	.w3(32'h3a07d3d9),
	.w4(32'h3b0eeb88),
	.w5(32'h3b20a281),
	.w6(32'h3b05af22),
	.w7(32'h3aa0a60f),
	.w8(32'h3a84b2c6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c7e44),
	.w1(32'h398c214a),
	.w2(32'h382ad87a),
	.w3(32'h3ae457f4),
	.w4(32'hb734cd06),
	.w5(32'hbabb69cb),
	.w6(32'h3a4ff99e),
	.w7(32'hb90e3740),
	.w8(32'hbb261dd5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a374a),
	.w1(32'hbb137465),
	.w2(32'h39333d4d),
	.w3(32'hbb18bed7),
	.w4(32'hbb38f806),
	.w5(32'h3521431c),
	.w6(32'hba86265b),
	.w7(32'hbafd5767),
	.w8(32'h3a55fdc0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb89f),
	.w1(32'h3ac2e2cc),
	.w2(32'h3a70f27a),
	.w3(32'h3a42a681),
	.w4(32'h3a8ce720),
	.w5(32'hba13f378),
	.w6(32'h3aa79300),
	.w7(32'h3a7b8743),
	.w8(32'hbad6d69d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46705b),
	.w1(32'hbb2b681d),
	.w2(32'hba9e646d),
	.w3(32'hba9132ce),
	.w4(32'hba215306),
	.w5(32'hbb2eada2),
	.w6(32'hbada8579),
	.w7(32'hbaeba0f4),
	.w8(32'hbb228b98),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0664b8),
	.w1(32'hba61252a),
	.w2(32'hbafc1440),
	.w3(32'hbb061f0e),
	.w4(32'hbaaf6155),
	.w5(32'h3b170437),
	.w6(32'hba8896fb),
	.w7(32'hbae17e51),
	.w8(32'h3b0bb9fb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7edc2c),
	.w1(32'h3b250ffa),
	.w2(32'h3abba973),
	.w3(32'h3b396dbb),
	.w4(32'h3af347b8),
	.w5(32'hba42cf1f),
	.w6(32'h3b762a4c),
	.w7(32'hb880cc22),
	.w8(32'h3a636487),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388181e0),
	.w1(32'h38506587),
	.w2(32'h37ae9d43),
	.w3(32'hbae07573),
	.w4(32'hb9e2c5e6),
	.w5(32'h3ab4bf15),
	.w6(32'h3ae4d706),
	.w7(32'h3aa3f229),
	.w8(32'h3ac96cb6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cb21),
	.w1(32'h3ad24d6f),
	.w2(32'hb8ea1676),
	.w3(32'h394e8c2d),
	.w4(32'h3b08895d),
	.w5(32'h3b02df2d),
	.w6(32'h3b03ab24),
	.w7(32'h383e4023),
	.w8(32'h3a734b53),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96461e),
	.w1(32'h38b1f959),
	.w2(32'hba85950e),
	.w3(32'h3b8a7d23),
	.w4(32'h3b56e49b),
	.w5(32'hb7dd8837),
	.w6(32'h3b73ecba),
	.w7(32'h3a0c2b1b),
	.w8(32'hbaee2128),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08f3c8),
	.w1(32'hba8bc6ba),
	.w2(32'hbabbb5ea),
	.w3(32'hbb115889),
	.w4(32'hb95ac983),
	.w5(32'h39ed4093),
	.w6(32'hbb5e7a2c),
	.w7(32'hba8b0a75),
	.w8(32'h3a179ad6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992056a),
	.w1(32'hb97bddb5),
	.w2(32'h39ae8b0e),
	.w3(32'h3b3c6be5),
	.w4(32'h3b40a64e),
	.w5(32'hba899b38),
	.w6(32'h3b056afe),
	.w7(32'hb93fd843),
	.w8(32'hbb05a270),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba366d47),
	.w1(32'hbb21f28f),
	.w2(32'hbae6b475),
	.w3(32'hbb42c52f),
	.w4(32'hbb0c763e),
	.w5(32'h3a90e25d),
	.w6(32'hbbafceac),
	.w7(32'hbb19c8dc),
	.w8(32'h3a3c8733),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27afa3),
	.w1(32'h3a2e4b37),
	.w2(32'h3a873301),
	.w3(32'h3aa96f8c),
	.w4(32'h3afef206),
	.w5(32'h39bc672a),
	.w6(32'h3a347259),
	.w7(32'h39fe5a5e),
	.w8(32'hb9bac953),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0295b8),
	.w1(32'hb98e6dcf),
	.w2(32'hb98efa33),
	.w3(32'h3910b960),
	.w4(32'h398dfc41),
	.w5(32'h3aa02274),
	.w6(32'hb8561e6e),
	.w7(32'hba53ac1e),
	.w8(32'h3aec5074),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2f384),
	.w1(32'h3b5534aa),
	.w2(32'h3b5f1a3d),
	.w3(32'h3afe697d),
	.w4(32'h3ba910dc),
	.w5(32'h3a33b8f3),
	.w6(32'h3b6ca6be),
	.w7(32'h3b5df7c7),
	.w8(32'h39480700),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf724a),
	.w1(32'hb92cf7bb),
	.w2(32'hba0fc023),
	.w3(32'h393d2f1c),
	.w4(32'hb975c424),
	.w5(32'hba912db1),
	.w6(32'h3ad87cb1),
	.w7(32'hb9505347),
	.w8(32'h3a28df21),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad94700),
	.w1(32'hbb0d345b),
	.w2(32'h3a959d4d),
	.w3(32'hba8fac81),
	.w4(32'h3915a2a5),
	.w5(32'h3a14a05a),
	.w6(32'h3a449e0d),
	.w7(32'hba72fbdb),
	.w8(32'h390b9f5c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacabc5),
	.w1(32'h3a493997),
	.w2(32'h3985590c),
	.w3(32'h3a656251),
	.w4(32'h3aa8979f),
	.w5(32'h3af08cc8),
	.w6(32'h3a91ef30),
	.w7(32'hb9144a5e),
	.w8(32'hba59a97e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a248144),
	.w1(32'hbacf6dd7),
	.w2(32'hb799f17d),
	.w3(32'h394e784c),
	.w4(32'h3a9940fb),
	.w5(32'h39df4017),
	.w6(32'hbadcdca7),
	.w7(32'hba9eaca2),
	.w8(32'h39949ca4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f975fb),
	.w1(32'h395ce957),
	.w2(32'h3a800dc6),
	.w3(32'h39633c45),
	.w4(32'h3b0ba77a),
	.w5(32'h3b1cd22b),
	.w6(32'hba082c47),
	.w7(32'hb73e4994),
	.w8(32'h3a93cdf5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8953),
	.w1(32'h3b47746c),
	.w2(32'h3b90980a),
	.w3(32'h3b212ce1),
	.w4(32'h3b176e43),
	.w5(32'h3b35efb4),
	.w6(32'h3b378daf),
	.w7(32'h3b01c949),
	.w8(32'h3b813616),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde90fc),
	.w1(32'h3b910a8f),
	.w2(32'h3a842918),
	.w3(32'h3b82536d),
	.w4(32'h3bb903b8),
	.w5(32'h3acc8637),
	.w6(32'h3bd3d4d6),
	.w7(32'h3b73cedf),
	.w8(32'h3a834316),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bfde0),
	.w1(32'h3b19aeea),
	.w2(32'h3addc0bf),
	.w3(32'h3ad59bb1),
	.w4(32'h3b332291),
	.w5(32'h3929e173),
	.w6(32'h3ab63358),
	.w7(32'h3b2c92c6),
	.w8(32'h3a63a32f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e968),
	.w1(32'h3ab03902),
	.w2(32'h3a919460),
	.w3(32'h3a2e3a63),
	.w4(32'h3b3104f2),
	.w5(32'h3af975b7),
	.w6(32'h392e829a),
	.w7(32'h39c939fb),
	.w8(32'h3ac279b3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18d7c4),
	.w1(32'h39737dc4),
	.w2(32'hba48f2da),
	.w3(32'h391037f7),
	.w4(32'h3b54bbc8),
	.w5(32'hba59fa00),
	.w6(32'h3b056046),
	.w7(32'h3a9eec0f),
	.w8(32'h3ab780eb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b688404),
	.w1(32'h3ae9105d),
	.w2(32'h3b0eab00),
	.w3(32'h3ae6478d),
	.w4(32'h3b4981cd),
	.w5(32'hba26db97),
	.w6(32'h3beb968f),
	.w7(32'h3b5d481e),
	.w8(32'hb9cb32ae),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6140b1),
	.w1(32'h399a1e27),
	.w2(32'hb9c1755e),
	.w3(32'hb9b6584b),
	.w4(32'h3a3bf964),
	.w5(32'h36b0196b),
	.w6(32'hba3fcab7),
	.w7(32'h3a2f26a5),
	.w8(32'h3af9a4c8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e9dc8),
	.w1(32'h3a5df93f),
	.w2(32'hbaf773ac),
	.w3(32'hb99187fe),
	.w4(32'hba6634a4),
	.w5(32'hba2f081b),
	.w6(32'h3b18a34e),
	.w7(32'hb9f93de1),
	.w8(32'hba547da3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a783098),
	.w1(32'h38e2537e),
	.w2(32'hb8a78ab0),
	.w3(32'h35b78aed),
	.w4(32'h382f6f49),
	.w5(32'hbaaff3ae),
	.w6(32'hbaaacd31),
	.w7(32'hb9961b5f),
	.w8(32'hba8b794a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf7107),
	.w1(32'h3934db9f),
	.w2(32'h3aa8d8b6),
	.w3(32'hbaf4f9de),
	.w4(32'h3ab7d04c),
	.w5(32'h3b0decaa),
	.w6(32'h39da967f),
	.w7(32'h3b1af8db),
	.w8(32'h39e6cf72),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79882d),
	.w1(32'hba7a91a1),
	.w2(32'h39a5d924),
	.w3(32'h3a8041e9),
	.w4(32'h396570ec),
	.w5(32'hb950f764),
	.w6(32'hb94e2352),
	.w7(32'h3a2cccae),
	.w8(32'hb995e76e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dd269),
	.w1(32'h38afbb89),
	.w2(32'h3996dc81),
	.w3(32'hb90e9bf7),
	.w4(32'hba5a108b),
	.w5(32'h39e50692),
	.w6(32'hb9048a90),
	.w7(32'hba299b8d),
	.w8(32'hba0de639),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dac329),
	.w1(32'h3a6b6e03),
	.w2(32'h3ae0f340),
	.w3(32'hb8f5cf48),
	.w4(32'hb9bd120c),
	.w5(32'hb8cbcb9a),
	.w6(32'hb99493cf),
	.w7(32'h3b476905),
	.w8(32'hbaf59c07),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a931949),
	.w1(32'h3916dd30),
	.w2(32'h3b09f3a1),
	.w3(32'h3ad4a613),
	.w4(32'h3a569767),
	.w5(32'h3a247a20),
	.w6(32'hbac3b3df),
	.w7(32'h39bb95f7),
	.w8(32'h394f9d43),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a8c8f),
	.w1(32'hbaa119ac),
	.w2(32'h38fedc27),
	.w3(32'hbacfaf91),
	.w4(32'hba0b1a4e),
	.w5(32'h39909da1),
	.w6(32'hbaa56b44),
	.w7(32'h3a87be09),
	.w8(32'h3aae076a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eae77),
	.w1(32'h3b4d7a26),
	.w2(32'h3b0ada48),
	.w3(32'h3b23da51),
	.w4(32'h3b01eb23),
	.w5(32'hb9d386d5),
	.w6(32'h3ab6eed8),
	.w7(32'h3a3b75ea),
	.w8(32'hb799d2cc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6736ca),
	.w1(32'h3b814ac0),
	.w2(32'h3ab71026),
	.w3(32'hb84e5e40),
	.w4(32'h3b26b393),
	.w5(32'hbae05a77),
	.w6(32'h3b8f6cb9),
	.w7(32'h3b1b03bc),
	.w8(32'hba81c9ee),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881b41),
	.w1(32'h3b1af1eb),
	.w2(32'h3b817836),
	.w3(32'hbad93720),
	.w4(32'h3b8ad3fc),
	.w5(32'h329b3ae8),
	.w6(32'h3b546d61),
	.w7(32'h3b814de1),
	.w8(32'hb99ce0ad),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2286c),
	.w1(32'hba60892c),
	.w2(32'h39f296ee),
	.w3(32'hbb148e11),
	.w4(32'hbb92d738),
	.w5(32'h3994c1da),
	.w6(32'hb90400ae),
	.w7(32'hbb67d26b),
	.w8(32'hbae5d8e6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67830b),
	.w1(32'hbacfc4fb),
	.w2(32'hb9297555),
	.w3(32'hb98dbb4d),
	.w4(32'h394268ab),
	.w5(32'h3b420f21),
	.w6(32'hba1d16d9),
	.w7(32'h3aa7f6e6),
	.w8(32'h3b6eaa5f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72b26d),
	.w1(32'h3a28c58b),
	.w2(32'h3aad4df8),
	.w3(32'h3ae3c087),
	.w4(32'h3a94311d),
	.w5(32'h3a9a858a),
	.w6(32'h3aefd2be),
	.w7(32'h3ab4e312),
	.w8(32'h3a38e212),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2406),
	.w1(32'hbb34b808),
	.w2(32'hbab81b6c),
	.w3(32'hba4a5ebb),
	.w4(32'h3951d11c),
	.w5(32'h397dafbf),
	.w6(32'hbb19ee0c),
	.w7(32'hbaafda68),
	.w8(32'h3a1c96e4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a756727),
	.w1(32'h3a7671f3),
	.w2(32'hba237eb8),
	.w3(32'hba8893d7),
	.w4(32'hbb20c485),
	.w5(32'h3a5f4858),
	.w6(32'hb9fded32),
	.w7(32'hba3afd22),
	.w8(32'h3b02f1b3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba7265),
	.w1(32'hbb24d44e),
	.w2(32'hbb46767f),
	.w3(32'hba8ac5d1),
	.w4(32'hbaa59818),
	.w5(32'h3a918fe0),
	.w6(32'hb95f05ec),
	.w7(32'hbb10c6de),
	.w8(32'h3b391f8a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b68a),
	.w1(32'h3a90b3cc),
	.w2(32'h3af23545),
	.w3(32'h3b94bfc1),
	.w4(32'h3b94e206),
	.w5(32'h39d7165a),
	.w6(32'h3b97ca2b),
	.w7(32'h3addbd95),
	.w8(32'h3abda17e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac92f99),
	.w1(32'hbb07f362),
	.w2(32'h3a47360e),
	.w3(32'h39eed4ca),
	.w4(32'hb9d2b99f),
	.w5(32'h3a2323b6),
	.w6(32'h39602d32),
	.w7(32'hba3f1eb5),
	.w8(32'hbb17ddb2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c24af),
	.w1(32'h3a9dab94),
	.w2(32'h3aabc4b4),
	.w3(32'hbb2f54d5),
	.w4(32'hba6fdd3e),
	.w5(32'h396faac3),
	.w6(32'h3adddb6d),
	.w7(32'h3aa88125),
	.w8(32'h38a91541),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1568f0),
	.w1(32'h398fc5ab),
	.w2(32'hba208039),
	.w3(32'h39bdc8dd),
	.w4(32'hb936a959),
	.w5(32'hb9f5cfa9),
	.w6(32'h3a400740),
	.w7(32'hb9f0b1d7),
	.w8(32'hbaa5dc1e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384ea916),
	.w1(32'hba4167eb),
	.w2(32'hba96c2d0),
	.w3(32'hbb08745d),
	.w4(32'hbb37f643),
	.w5(32'hb9b3d5d2),
	.w6(32'hbb64d028),
	.w7(32'hbb322891),
	.w8(32'hba8fb371),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ca0a7),
	.w1(32'h3ac5518b),
	.w2(32'h3ae338c7),
	.w3(32'h387bba61),
	.w4(32'h3a245fbe),
	.w5(32'hba073d8a),
	.w6(32'h3b0926cf),
	.w7(32'h3b2392d7),
	.w8(32'hba9d8781),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c5393),
	.w1(32'hbae43951),
	.w2(32'hbb08a239),
	.w3(32'hbb24816f),
	.w4(32'hbb471457),
	.w5(32'hb9874620),
	.w6(32'hba1ff65b),
	.w7(32'hbafa35cc),
	.w8(32'hba34b058),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f3f14),
	.w1(32'hba5bc0dc),
	.w2(32'h392d7fe9),
	.w3(32'hb8c21c3b),
	.w4(32'h3a0be811),
	.w5(32'h39aee6c3),
	.w6(32'hb9047a38),
	.w7(32'h391a0ba4),
	.w8(32'hbae61c02),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18b0b8),
	.w1(32'h3b1a0baf),
	.w2(32'h3b1771ac),
	.w3(32'hba179f20),
	.w4(32'h39842ba7),
	.w5(32'hbaf77a27),
	.w6(32'hba800601),
	.w7(32'hb8c37784),
	.w8(32'hba9b8b7e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11c3a0),
	.w1(32'hbb6a6d96),
	.w2(32'hbbab6d81),
	.w3(32'hba9b1d2b),
	.w4(32'hbb3a2db7),
	.w5(32'hba49457c),
	.w6(32'hbb5a01a8),
	.w7(32'hbb535383),
	.w8(32'h3b523e43),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5cf57),
	.w1(32'h3bcf51b9),
	.w2(32'h3b739b6c),
	.w3(32'h3b7af395),
	.w4(32'h3baf2ee0),
	.w5(32'h3a2dc80a),
	.w6(32'h3c0c28c7),
	.w7(32'h3bab517f),
	.w8(32'h3a90958a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2238ec),
	.w1(32'hbad96846),
	.w2(32'h37592cd5),
	.w3(32'hb8850a09),
	.w4(32'h38fb98e1),
	.w5(32'h3b0d58f6),
	.w6(32'h396cdd63),
	.w7(32'h38a380fa),
	.w8(32'h3b1bb715),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32fe45),
	.w1(32'h3b24bfe6),
	.w2(32'h3b3c7762),
	.w3(32'h3b1283bb),
	.w4(32'h3a9a8633),
	.w5(32'hbaa5bf73),
	.w6(32'h3ac7682e),
	.w7(32'h3ac17062),
	.w8(32'hba774596),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7832c4),
	.w1(32'hbb623140),
	.w2(32'hbb7d71a5),
	.w3(32'hbadf7e4f),
	.w4(32'hbb531686),
	.w5(32'hbad42d21),
	.w6(32'hbaae7c7f),
	.w7(32'hbafef50f),
	.w8(32'hba8bc0fb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047766),
	.w1(32'h3a069777),
	.w2(32'hba1b48b0),
	.w3(32'h3b1ab3d6),
	.w4(32'hba1215a3),
	.w5(32'h3b09a342),
	.w6(32'h3a86ca10),
	.w7(32'hbb2383e6),
	.w8(32'h3a86cd49),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9af2e6),
	.w1(32'h3a965fb5),
	.w2(32'h3b50ed08),
	.w3(32'h3b54d665),
	.w4(32'h3b1407be),
	.w5(32'h3aa5b31e),
	.w6(32'h3a50d619),
	.w7(32'h3ac93537),
	.w8(32'h3b1515a0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c4ecd),
	.w1(32'h3b3b1e57),
	.w2(32'h3b6fa81f),
	.w3(32'h3b355b03),
	.w4(32'h3b09e3c3),
	.w5(32'h3b32e5c1),
	.w6(32'h3aec2139),
	.w7(32'h3a960d85),
	.w8(32'h3af799a5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7242e),
	.w1(32'h3afc683c),
	.w2(32'h3ab9da06),
	.w3(32'h3990206b),
	.w4(32'h3af5e255),
	.w5(32'hba80946d),
	.w6(32'h3a3ab290),
	.w7(32'h3adafc52),
	.w8(32'hba96168b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e674),
	.w1(32'h3a23fab7),
	.w2(32'hb9a1b9bb),
	.w3(32'hb7cf61d5),
	.w4(32'h3ab8803a),
	.w5(32'h3a6b13a1),
	.w6(32'hba0d2545),
	.w7(32'hb9b5882f),
	.w8(32'h3b04e619),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc236c),
	.w1(32'h3a3f79f5),
	.w2(32'h3a2407ab),
	.w3(32'h3a6b4c5f),
	.w4(32'h3a83fba7),
	.w5(32'hba1a26fa),
	.w6(32'h3a9c46f1),
	.w7(32'h392809f1),
	.w8(32'hb9e42c85),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2cb7f),
	.w1(32'hba9778ea),
	.w2(32'h3a91d0b3),
	.w3(32'hb932de76),
	.w4(32'hbb0bd180),
	.w5(32'h39b99a75),
	.w6(32'hbb4e96a0),
	.w7(32'hba2b587d),
	.w8(32'hba3e7c9b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c4533),
	.w1(32'hba75a629),
	.w2(32'hb99134e3),
	.w3(32'h39d603b1),
	.w4(32'h399c299a),
	.w5(32'hbb4427b7),
	.w6(32'hba1733f6),
	.w7(32'hb9d52826),
	.w8(32'h3ab78478),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42dd9f),
	.w1(32'h3a8a57a6),
	.w2(32'hba4075dd),
	.w3(32'hb9dddc5a),
	.w4(32'h3b4c693f),
	.w5(32'h391ef16a),
	.w6(32'h3bcea77a),
	.w7(32'h3b28edaf),
	.w8(32'h3a86f328),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638891),
	.w1(32'h39d4b46e),
	.w2(32'h3a77e913),
	.w3(32'h3aea1efc),
	.w4(32'h39f32a4b),
	.w5(32'h3abdf12d),
	.w6(32'h3b62042a),
	.w7(32'h3a3662c1),
	.w8(32'hb9aeee2d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafff94b),
	.w1(32'hba4b68ea),
	.w2(32'h3abfccb4),
	.w3(32'h3b05aaa6),
	.w4(32'h3a267c4e),
	.w5(32'hb9f75829),
	.w6(32'hba13a575),
	.w7(32'h3adfcff1),
	.w8(32'hba7f0e3f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd1d8d),
	.w1(32'hb9015da5),
	.w2(32'hba82f5e0),
	.w3(32'hba93e7b5),
	.w4(32'hb9f45280),
	.w5(32'h3a29657c),
	.w6(32'hbb07b83e),
	.w7(32'hbaf6dc86),
	.w8(32'h3a230698),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26261a),
	.w1(32'h3afbee33),
	.w2(32'h3aabd0f1),
	.w3(32'h3aa3c843),
	.w4(32'h3b019b85),
	.w5(32'h3a33b4b8),
	.w6(32'h39dea09a),
	.w7(32'h3aa73dfa),
	.w8(32'h3b0123c8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c844),
	.w1(32'h3abafea9),
	.w2(32'hba8a576f),
	.w3(32'h3a7ef294),
	.w4(32'h3a57b4ba),
	.w5(32'h3a0e0c56),
	.w6(32'h3b229b4e),
	.w7(32'h36dc1994),
	.w8(32'h3a462258),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ac905),
	.w1(32'h395ede7a),
	.w2(32'h3a6220a4),
	.w3(32'h39a9b395),
	.w4(32'h3a37ee88),
	.w5(32'h3b24c7c6),
	.w6(32'h3a660b10),
	.w7(32'h39e95176),
	.w8(32'h3af68e1e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139e94),
	.w1(32'h3c0039c3),
	.w2(32'h3bce265b),
	.w3(32'h3c2241e9),
	.w4(32'h3bbd39ee),
	.w5(32'h3adf2ffa),
	.w6(32'h3b7c41e8),
	.w7(32'h3b1d8761),
	.w8(32'hba924453),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15cd5a),
	.w1(32'h3a5faf6b),
	.w2(32'h3883ab5d),
	.w3(32'h36aeaaeb),
	.w4(32'hba6ca061),
	.w5(32'h3a92556f),
	.w6(32'hba6061ca),
	.w7(32'hb9e0c2b5),
	.w8(32'h394503b2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5f9c8),
	.w1(32'h3a98d5d6),
	.w2(32'h3b09832e),
	.w3(32'h3b00c26d),
	.w4(32'h3b5c18cd),
	.w5(32'hba3edb9d),
	.w6(32'h3aba3cff),
	.w7(32'h3ae7351f),
	.w8(32'hbb205548),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14965b),
	.w1(32'hbb2fd1d3),
	.w2(32'hbaf38484),
	.w3(32'hba4a79cc),
	.w4(32'hbae88bd6),
	.w5(32'hb9e6c871),
	.w6(32'hbb18ed99),
	.w7(32'hbaed07ad),
	.w8(32'hb9d72aee),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779fdb),
	.w1(32'hb8930eed),
	.w2(32'hbac479ce),
	.w3(32'hbac8b388),
	.w4(32'hba72c10e),
	.w5(32'hbab4b3a6),
	.w6(32'hbad45be0),
	.w7(32'hbaf59945),
	.w8(32'hbb431f0d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b443),
	.w1(32'hbb1b1e48),
	.w2(32'hbb05b034),
	.w3(32'hba89dba6),
	.w4(32'hbad56156),
	.w5(32'hba38cd2b),
	.w6(32'hbb3fa10b),
	.w7(32'hbac28488),
	.w8(32'hb99ac214),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25fe44),
	.w1(32'h3a31a0ec),
	.w2(32'h39f9c2df),
	.w3(32'h3b3c936f),
	.w4(32'h3b4588f6),
	.w5(32'h3ac34499),
	.w6(32'h3b8e9002),
	.w7(32'h3b264c90),
	.w8(32'h3a4aabae),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a358),
	.w1(32'h3b7c2a02),
	.w2(32'h3a5fefef),
	.w3(32'h3b5f9af8),
	.w4(32'h3b804b21),
	.w5(32'h3971ed70),
	.w6(32'h3b635f9f),
	.w7(32'h3a99860d),
	.w8(32'hba4c644d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388747ce),
	.w1(32'hb8b95462),
	.w2(32'hb80cec8a),
	.w3(32'hb8315b31),
	.w4(32'hb6e8de41),
	.w5(32'h3945fcaf),
	.w6(32'hba3b5fe0),
	.w7(32'hba4e6656),
	.w8(32'hbb0019eb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16721e),
	.w1(32'hbad25712),
	.w2(32'hba052ff3),
	.w3(32'hbb0ab09c),
	.w4(32'hbae65581),
	.w5(32'hba22522e),
	.w6(32'hbaa9442a),
	.w7(32'h3970bdae),
	.w8(32'hb93eee00),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08bbcb),
	.w1(32'h3a6f7c9d),
	.w2(32'h3a38eefe),
	.w3(32'h3a759be1),
	.w4(32'h39e5e781),
	.w5(32'h3acacf0e),
	.w6(32'hbacf27ac),
	.w7(32'hb98f311c),
	.w8(32'h3a6e22af),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b196686),
	.w1(32'h3b10644e),
	.w2(32'h3b12aa1f),
	.w3(32'h39c27017),
	.w4(32'h3a6f7d37),
	.w5(32'h3a1a15d2),
	.w6(32'h3b0124ed),
	.w7(32'h3ad01dd9),
	.w8(32'hba90caac),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b9050),
	.w1(32'hb998199b),
	.w2(32'h3ac306ab),
	.w3(32'h39541746),
	.w4(32'h382ab02f),
	.w5(32'h394665f1),
	.w6(32'hb9e08f02),
	.w7(32'h3a42ad42),
	.w8(32'hba6bbb63),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe39e),
	.w1(32'hba4a8c26),
	.w2(32'h39c9a714),
	.w3(32'hbaa011cd),
	.w4(32'hb83d879f),
	.w5(32'hba69907b),
	.w6(32'hba9183d7),
	.w7(32'hba8e857d),
	.w8(32'hbad521bb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0b73),
	.w1(32'hba84f3c5),
	.w2(32'hbac21b0e),
	.w3(32'hb9a1892c),
	.w4(32'h39a0af1d),
	.w5(32'h3abf392b),
	.w6(32'hbae58a6a),
	.w7(32'hb9cf3d53),
	.w8(32'h3a8782c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ff9c3),
	.w1(32'h3aa2e738),
	.w2(32'hba08f435),
	.w3(32'h3ad186b9),
	.w4(32'h3af1dcad),
	.w5(32'hbaf141d0),
	.w6(32'h3b800eed),
	.w7(32'h3a71bc24),
	.w8(32'hbb15ed30),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6bf7f),
	.w1(32'hba032aae),
	.w2(32'hb998c48e),
	.w3(32'h3a1aa891),
	.w4(32'hb88a9a29),
	.w5(32'hbb363879),
	.w6(32'hb9eebae6),
	.w7(32'h3a2426e7),
	.w8(32'h3a81e3b8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96959e),
	.w1(32'h3b769bd1),
	.w2(32'h3aaa1584),
	.w3(32'h3a08b605),
	.w4(32'h3b8af45c),
	.w5(32'h39aa78ba),
	.w6(32'h3bf92e77),
	.w7(32'h3b53ff44),
	.w8(32'hb816e11a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacefd13),
	.w1(32'hbae2d11f),
	.w2(32'hba9e4704),
	.w3(32'h3a255299),
	.w4(32'h39cc8a84),
	.w5(32'hba07ae9c),
	.w6(32'hb96b9aa7),
	.w7(32'hb93b6632),
	.w8(32'h39a7dc64),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917e4e),
	.w1(32'h3b1f0018),
	.w2(32'h3aca62bc),
	.w3(32'h3b10224a),
	.w4(32'h3b455087),
	.w5(32'h3b27ff76),
	.w6(32'h3b371f99),
	.w7(32'h3adeed85),
	.w8(32'h3a8068be),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273544),
	.w1(32'h3b388a5f),
	.w2(32'h3b47913b),
	.w3(32'h3b6f1a8a),
	.w4(32'h3b793548),
	.w5(32'hb8b62a3b),
	.w6(32'h3ad04ca9),
	.w7(32'h3a869ced),
	.w8(32'h3aad3094),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbbee5),
	.w1(32'h3bad112a),
	.w2(32'h3b47e4ce),
	.w3(32'h3b9585b4),
	.w4(32'h3b78a8c3),
	.w5(32'h3a02ee36),
	.w6(32'h3b181be4),
	.w7(32'h3affb651),
	.w8(32'hba006cc7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39048609),
	.w1(32'h3a220c72),
	.w2(32'hb90f7751),
	.w3(32'h39253bb3),
	.w4(32'h37fdb5dc),
	.w5(32'hbaa8ef59),
	.w6(32'hba71f07a),
	.w7(32'hb99da15a),
	.w8(32'hbb10ffb3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcbfda),
	.w1(32'h3aebc7e0),
	.w2(32'hb95db0f3),
	.w3(32'hbb0df752),
	.w4(32'h39decda0),
	.w5(32'h3b2c00c3),
	.w6(32'h3ad277c6),
	.w7(32'h3ac2bc7d),
	.w8(32'h3b2f16ed),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd00e8),
	.w1(32'hb923e19f),
	.w2(32'hba5044d8),
	.w3(32'h3aacad5f),
	.w4(32'h3a55c084),
	.w5(32'hbab21775),
	.w6(32'h3a226cf7),
	.w7(32'h3a1b0454),
	.w8(32'hbb092713),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e17b2),
	.w1(32'h3aebda36),
	.w2(32'h38dff647),
	.w3(32'hba290c1e),
	.w4(32'hba32351c),
	.w5(32'h3aba44d6),
	.w6(32'h3aac0264),
	.w7(32'hb9d480be),
	.w8(32'h3ac88c0d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b870744),
	.w1(32'h3b50568b),
	.w2(32'h3b8d7185),
	.w3(32'h3b931ceb),
	.w4(32'h3bbf0faa),
	.w5(32'hba4607cc),
	.w6(32'h3b8e302e),
	.w7(32'h3b57378f),
	.w8(32'h3a0f4858),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f4691),
	.w1(32'hbae19c63),
	.w2(32'h397b9f61),
	.w3(32'h3a0b96eb),
	.w4(32'hba9f2f00),
	.w5(32'hba61920a),
	.w6(32'h3a2edd7d),
	.w7(32'hbaf298ff),
	.w8(32'hba0428eb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9620f3),
	.w1(32'h3a1e2b48),
	.w2(32'h3a34a2f5),
	.w3(32'hba359159),
	.w4(32'h391a5641),
	.w5(32'h3afa5dee),
	.w6(32'hba30b8fe),
	.w7(32'h3928f29b),
	.w8(32'h3a81bdf3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccc70f),
	.w1(32'h3a319998),
	.w2(32'h3ae40e8b),
	.w3(32'h3a89d095),
	.w4(32'h3a874417),
	.w5(32'h3b4f83ab),
	.w6(32'h3a2b33a8),
	.w7(32'h3a8f1ce6),
	.w8(32'h3bb29dc6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb55b4c),
	.w1(32'h3aa89931),
	.w2(32'hb980cc38),
	.w3(32'h3b867b79),
	.w4(32'h3b486d4f),
	.w5(32'hb9bfbfe6),
	.w6(32'h3b8cb21e),
	.w7(32'h3a1dc84a),
	.w8(32'hba746ff3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ef0f),
	.w1(32'h3b046751),
	.w2(32'h3b205fc7),
	.w3(32'h3b4e652c),
	.w4(32'h3b3c5dd9),
	.w5(32'h3b004f8f),
	.w6(32'h3a97c70f),
	.w7(32'h3a0222c8),
	.w8(32'h3aa76553),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e3842),
	.w1(32'h3ab1a365),
	.w2(32'hb9d0947e),
	.w3(32'hb98ba126),
	.w4(32'hba103264),
	.w5(32'h3a629a6b),
	.w6(32'h3a8a7058),
	.w7(32'hb92720fd),
	.w8(32'hba34a29b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bec22),
	.w1(32'hbb732832),
	.w2(32'hbb116bfe),
	.w3(32'hba8e79a7),
	.w4(32'hbb04676b),
	.w5(32'hb89ac1d4),
	.w6(32'h39fb174e),
	.w7(32'hbb0c158f),
	.w8(32'h3a0df6ce),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39860f79),
	.w1(32'h38b8a2cd),
	.w2(32'hba4a1682),
	.w3(32'hb9bfb1a3),
	.w4(32'hba01f0cb),
	.w5(32'h3a9854b4),
	.w6(32'hb9e053d9),
	.w7(32'hba8dbe4a),
	.w8(32'h3ad28e45),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81358f),
	.w1(32'hba963a3a),
	.w2(32'hba783e2e),
	.w3(32'hb8b5dd84),
	.w4(32'hb99bc8a1),
	.w5(32'h3aefec59),
	.w6(32'hb990c528),
	.w7(32'hba2deda7),
	.w8(32'h3ad0433b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3118e),
	.w1(32'h3a16cfe8),
	.w2(32'h3b296058),
	.w3(32'h3a28e086),
	.w4(32'h39531743),
	.w5(32'hbb4b9726),
	.w6(32'h3a1d10e7),
	.w7(32'h3aaeb7a9),
	.w8(32'hbad34fce),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43c3df),
	.w1(32'hb9362115),
	.w2(32'h38c0d6d2),
	.w3(32'hba799d2f),
	.w4(32'h39b649fc),
	.w5(32'h39d669e8),
	.w6(32'hbb41e0b8),
	.w7(32'hb90e73fa),
	.w8(32'h3b814f3a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804cfb),
	.w1(32'h3b53dbac),
	.w2(32'h3b5ed225),
	.w3(32'h3ad61ec8),
	.w4(32'h3bb855b1),
	.w5(32'h3893aa2d),
	.w6(32'h3bea0f76),
	.w7(32'h3bd663f6),
	.w8(32'hbb2425b3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08d02e),
	.w1(32'h3b94793b),
	.w2(32'h39d2b926),
	.w3(32'h3b284d26),
	.w4(32'h390f2099),
	.w5(32'hbb4974f2),
	.w6(32'hb9acf8da),
	.w7(32'h3acc8fb9),
	.w8(32'hbaec47b2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b0ac),
	.w1(32'h3bb45753),
	.w2(32'h39ced2be),
	.w3(32'h3c058ed0),
	.w4(32'h3ad5ef24),
	.w5(32'h3b55676c),
	.w6(32'h3c4da967),
	.w7(32'h3bfe66d3),
	.w8(32'h3b799b8d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0e61),
	.w1(32'h3b7a64f8),
	.w2(32'hbafbea5a),
	.w3(32'h3b7283d6),
	.w4(32'hba873eba),
	.w5(32'h3a09b952),
	.w6(32'h3b374833),
	.w7(32'hbb156e97),
	.w8(32'hbb33eab4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16a063),
	.w1(32'hbbae9e9b),
	.w2(32'h3c31972c),
	.w3(32'hbc4b40fb),
	.w4(32'hba4b6218),
	.w5(32'hbc1573ea),
	.w6(32'hbbe001a7),
	.w7(32'h3bb315d9),
	.w8(32'hbc7a87dc),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917aff),
	.w1(32'hbc181e5d),
	.w2(32'hba5b3d7f),
	.w3(32'hbc1995a2),
	.w4(32'hbaf33c0b),
	.w5(32'h3b022c21),
	.w6(32'hbc23dfb8),
	.w7(32'hbbcdb424),
	.w8(32'h3bc90f63),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f019c),
	.w1(32'h3b0abe24),
	.w2(32'hbbe9a7c7),
	.w3(32'h3b0bfc07),
	.w4(32'hbbc5297d),
	.w5(32'hbb86a433),
	.w6(32'h3b092346),
	.w7(32'hbbb31fa5),
	.w8(32'hbbf781f7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae11610),
	.w1(32'hbb84bcfa),
	.w2(32'hbaa3385a),
	.w3(32'hbb00ad9e),
	.w4(32'hb8120cd0),
	.w5(32'hbb0a1099),
	.w6(32'hba4b0f3c),
	.w7(32'hbb0621ed),
	.w8(32'hba34d871),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ec384),
	.w1(32'h3b0cd57c),
	.w2(32'hbb04c480),
	.w3(32'hbb1cd9d9),
	.w4(32'h3b6d15a6),
	.w5(32'hbb9ce35a),
	.w6(32'hbac8b808),
	.w7(32'hbb3ebe7e),
	.w8(32'hbb68c0da),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba475942),
	.w1(32'h38815ddd),
	.w2(32'hbbe67abc),
	.w3(32'hba97f46f),
	.w4(32'hbbeaa655),
	.w5(32'h3c1189a4),
	.w6(32'h3bc1c196),
	.w7(32'hbbfe6626),
	.w8(32'h3bf40974),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5b33),
	.w1(32'h3ba307d3),
	.w2(32'h3ba01af5),
	.w3(32'h3b494b66),
	.w4(32'h3bbd8faa),
	.w5(32'hbb582b0c),
	.w6(32'h3c08fc23),
	.w7(32'h3b9f5dd1),
	.w8(32'hbba9d3be),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857d03),
	.w1(32'h3c27dd39),
	.w2(32'h3a4f0e41),
	.w3(32'h3bd253fa),
	.w4(32'h3a5f2332),
	.w5(32'h3b83e9c4),
	.w6(32'h3ad72d9d),
	.w7(32'h3b1af3c8),
	.w8(32'h392b1c6b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1099c),
	.w1(32'hbbd34a3f),
	.w2(32'hbb084f27),
	.w3(32'hb993985d),
	.w4(32'h3b902c77),
	.w5(32'hbafc365c),
	.w6(32'hbbc2cf55),
	.w7(32'hbb562ede),
	.w8(32'hba6de144),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c85224),
	.w1(32'h3a42f0b6),
	.w2(32'h3b1a6082),
	.w3(32'h3b2a296d),
	.w4(32'hbb3ed884),
	.w5(32'hbc3f4e52),
	.w6(32'hba763878),
	.w7(32'hba8437ec),
	.w8(32'hbb594440),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b0f2),
	.w1(32'h3ad33f8a),
	.w2(32'hbc49136d),
	.w3(32'h3c41d848),
	.w4(32'hbb89fe24),
	.w5(32'hba36d682),
	.w6(32'h3cc13a3c),
	.w7(32'hbb796894),
	.w8(32'hbb1537b8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54dcc1),
	.w1(32'h3acc3e40),
	.w2(32'h3b09fac2),
	.w3(32'h3b4c2607),
	.w4(32'h3b2bc928),
	.w5(32'hbac487b9),
	.w6(32'h3aa6103a),
	.w7(32'hb8cffd82),
	.w8(32'h3b8043a5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f19ac),
	.w1(32'h3bbf1b69),
	.w2(32'hbc245540),
	.w3(32'hbb5af7bb),
	.w4(32'hbc047a81),
	.w5(32'h3ab65565),
	.w6(32'hbbe9e344),
	.w7(32'hbc4dfd36),
	.w8(32'hbaf7684a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db59e),
	.w1(32'h3c045c43),
	.w2(32'hbad7653d),
	.w3(32'h3b1b2f32),
	.w4(32'h3a81e291),
	.w5(32'hbc08b624),
	.w6(32'h3ba02b1c),
	.w7(32'h3a16f529),
	.w8(32'hbbbc9be6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fd2bc),
	.w1(32'hbc345f36),
	.w2(32'hbcc46034),
	.w3(32'hbbff8e6e),
	.w4(32'hbc84c77a),
	.w5(32'h3a4ce2d4),
	.w6(32'h3af89715),
	.w7(32'hbc803ad4),
	.w8(32'hba647de5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18327e),
	.w1(32'hbaa87aa7),
	.w2(32'h3a7d2ce3),
	.w3(32'h3adc4e38),
	.w4(32'h3b8646fe),
	.w5(32'h3b17e952),
	.w6(32'hbb06d35c),
	.w7(32'h3a53b5c9),
	.w8(32'h3a2304b2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f66a66),
	.w1(32'hbbbb6c12),
	.w2(32'hbb24afeb),
	.w3(32'hbb2177cd),
	.w4(32'hbbc1afa0),
	.w5(32'h3a9208bc),
	.w6(32'h3ba29de3),
	.w7(32'hba720f9a),
	.w8(32'hbaef4322),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b097f0b),
	.w1(32'h3a96a1e4),
	.w2(32'h3a30be00),
	.w3(32'h3bbf62ed),
	.w4(32'h3bd1af7e),
	.w5(32'hbb7a98f2),
	.w6(32'h3aacdb12),
	.w7(32'h3abb76d6),
	.w8(32'hbc310561),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8268),
	.w1(32'h3b822562),
	.w2(32'h3afcfe93),
	.w3(32'h3b2ef1d0),
	.w4(32'hbb8e7e43),
	.w5(32'hbc2ce476),
	.w6(32'h39de7e6e),
	.w7(32'h3b0bf58b),
	.w8(32'hbba92341),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce0b0b),
	.w1(32'hba804560),
	.w2(32'h3c15cae0),
	.w3(32'hbb00a0d0),
	.w4(32'h3c5f4584),
	.w5(32'hba9837fb),
	.w6(32'h3c36f8d0),
	.w7(32'h3c9380ff),
	.w8(32'hbae475a1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7bca),
	.w1(32'h3b5a1f2e),
	.w2(32'h3bdbae9a),
	.w3(32'h3acbd367),
	.w4(32'h3b1e7aa4),
	.w5(32'hb9364f9f),
	.w6(32'h3bc3b066),
	.w7(32'h3be6e3fc),
	.w8(32'h3965b00c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04fc9e),
	.w1(32'h3a270c33),
	.w2(32'hbbaf5781),
	.w3(32'hbbaad0dc),
	.w4(32'hbb68855d),
	.w5(32'h3b1d2107),
	.w6(32'hbad60c66),
	.w7(32'hbbeb0730),
	.w8(32'hbb0842cc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60823c),
	.w1(32'h33866f19),
	.w2(32'hbaf71232),
	.w3(32'hba2fdbd8),
	.w4(32'hbb53051a),
	.w5(32'hb93bdcb1),
	.w6(32'h3be06693),
	.w7(32'hbb98b8db),
	.w8(32'hba871d95),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c448d),
	.w1(32'hbac1495f),
	.w2(32'hbba2a0c5),
	.w3(32'hbb9e8a6f),
	.w4(32'hbbe7e657),
	.w5(32'h3aa4cd50),
	.w6(32'hbb3f3939),
	.w7(32'hbb6a7836),
	.w8(32'h39eac9a2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c048c),
	.w1(32'h3c240161),
	.w2(32'h3c789431),
	.w3(32'hbb0d4013),
	.w4(32'h3b39c0c0),
	.w5(32'h3a70faaf),
	.w6(32'h3bb28893),
	.w7(32'h3c44622c),
	.w8(32'h389ab87e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa77ab2),
	.w1(32'hbac23ba4),
	.w2(32'hbb8d2c06),
	.w3(32'hbaace269),
	.w4(32'hbb0273a2),
	.w5(32'h3b20ba9a),
	.w6(32'h3a96909c),
	.w7(32'hbbb8ce68),
	.w8(32'h3c247823),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac060a),
	.w1(32'h3c4e3997),
	.w2(32'hbb830820),
	.w3(32'h3c265d8c),
	.w4(32'hbb020970),
	.w5(32'hbb9325ce),
	.w6(32'h3b6096e1),
	.w7(32'hbbf6efa9),
	.w8(32'hbb6d84ce),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule