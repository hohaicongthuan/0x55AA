module layer_8_featuremap_134(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27d40),
	.w1(32'h3ac4b4af),
	.w2(32'hbb37a308),
	.w3(32'h3bb14f3d),
	.w4(32'h3c6203e0),
	.w5(32'h3ba0797e),
	.w6(32'h3c939369),
	.w7(32'h3c4d1593),
	.w8(32'hb9fe8ee8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d5e0d),
	.w1(32'hb9cdf0a5),
	.w2(32'h3bb052f0),
	.w3(32'hbbedf4fb),
	.w4(32'hb9ad9406),
	.w5(32'hbbcc3891),
	.w6(32'hbc5e8dea),
	.w7(32'h3a88c0a7),
	.w8(32'hbbd9eb2e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe880af),
	.w1(32'hbbe87baa),
	.w2(32'h3b3b3db3),
	.w3(32'h3a5cb4d1),
	.w4(32'hbb62248d),
	.w5(32'h3cf1da8b),
	.w6(32'hbbbea30e),
	.w7(32'h3bde00e8),
	.w8(32'h3d213c2e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc059),
	.w1(32'h3c3870e1),
	.w2(32'hbaf4ca08),
	.w3(32'hbca7c198),
	.w4(32'hbb5a0cef),
	.w5(32'hbc788291),
	.w6(32'h3d0dae15),
	.w7(32'h3c37f920),
	.w8(32'hbc45fe18),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c505eea),
	.w1(32'hbcbe1429),
	.w2(32'hbc136aec),
	.w3(32'h3cd43028),
	.w4(32'h3bf9f1bc),
	.w5(32'hbb9fe362),
	.w6(32'h3b278a0a),
	.w7(32'hba034c05),
	.w8(32'hba867e64),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c4db7),
	.w1(32'h3cad5f39),
	.w2(32'h3c5e144d),
	.w3(32'h3c729e17),
	.w4(32'h3c083edf),
	.w5(32'hbcc9a1c6),
	.w6(32'h3c2bea4c),
	.w7(32'h3c0127f2),
	.w8(32'hbd420386),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e8de8),
	.w1(32'h3af50bf9),
	.w2(32'h3bb77fa1),
	.w3(32'h3b8972c1),
	.w4(32'h3b9953ae),
	.w5(32'hbc7a38cd),
	.w6(32'hbc13a220),
	.w7(32'h3c3bff5a),
	.w8(32'h3b217659),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4635c0),
	.w1(32'hbb9d9e7f),
	.w2(32'hbaa39976),
	.w3(32'h368482e5),
	.w4(32'hbbd68e30),
	.w5(32'hbc46dc4e),
	.w6(32'hbc3e4b52),
	.w7(32'h3b6ae46f),
	.w8(32'hbc953ab8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c291),
	.w1(32'h3cd935c3),
	.w2(32'h3b29d8b4),
	.w3(32'hbb9475a1),
	.w4(32'h3c89b035),
	.w5(32'h3c001f7a),
	.w6(32'hbba5aae8),
	.w7(32'h3c3936fa),
	.w8(32'h3bd63f05),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7f9f0),
	.w1(32'hbc8d7765),
	.w2(32'hbc820417),
	.w3(32'hbc325dcc),
	.w4(32'h39ce1796),
	.w5(32'h3d08b150),
	.w6(32'hbc2a11ec),
	.w7(32'h3c02d938),
	.w8(32'hbbd78823),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca67277),
	.w1(32'h3c0dee69),
	.w2(32'hbb42fd4c),
	.w3(32'hbc583db9),
	.w4(32'hbc56f357),
	.w5(32'h3b94a67c),
	.w6(32'h3cacceba),
	.w7(32'hbc20f429),
	.w8(32'h3ccdffdd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9852a9),
	.w1(32'hbc614f2d),
	.w2(32'hbc0873c3),
	.w3(32'h3bbd7d9d),
	.w4(32'h3c4d0270),
	.w5(32'h3abda86d),
	.w6(32'hb8c8428a),
	.w7(32'h3c26082f),
	.w8(32'hbc832d24),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bc990),
	.w1(32'h3bff37f3),
	.w2(32'hba056764),
	.w3(32'hbb90b4b0),
	.w4(32'h3ac9101f),
	.w5(32'h3b33ea6a),
	.w6(32'hbca6fc48),
	.w7(32'hbba81545),
	.w8(32'h3b77d9de),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfef3c),
	.w1(32'hba1b783c),
	.w2(32'hbaab894e),
	.w3(32'h39d047e3),
	.w4(32'hbbb2541b),
	.w5(32'h398f9927),
	.w6(32'h3b97fb9f),
	.w7(32'hbbbea547),
	.w8(32'hb9f011a3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac376c),
	.w1(32'h3b8eaa5c),
	.w2(32'h3aef4ebc),
	.w3(32'h3b873209),
	.w4(32'hbabe3022),
	.w5(32'h3acc8f57),
	.w6(32'h3b8afcdb),
	.w7(32'hbb83e05b),
	.w8(32'h35aec157),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07573e),
	.w1(32'hba7480bb),
	.w2(32'hbb9b0c2c),
	.w3(32'hba06caff),
	.w4(32'h3c663bb4),
	.w5(32'h3c3ee7ff),
	.w6(32'hba980c27),
	.w7(32'hbb8b3830),
	.w8(32'hbc3b6295),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc55f8),
	.w1(32'hbbdbd208),
	.w2(32'h3bae8b17),
	.w3(32'h3bbcfad5),
	.w4(32'hbad47124),
	.w5(32'hbbdb7ff9),
	.w6(32'hbbdaf6c3),
	.w7(32'hbc92508d),
	.w8(32'hbcc3f73a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7c99d),
	.w1(32'hbbd86527),
	.w2(32'hba2af936),
	.w3(32'hba89fe6d),
	.w4(32'h3c0ca8bd),
	.w5(32'h3bb2df45),
	.w6(32'hbc36f70f),
	.w7(32'hbbd65ed2),
	.w8(32'hbca22c6a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b363b),
	.w1(32'hbd0690d1),
	.w2(32'h3af59758),
	.w3(32'hbbad3dd7),
	.w4(32'hbd143a4c),
	.w5(32'h3ba7ca6f),
	.w6(32'h3c47c38b),
	.w7(32'h3d13b202),
	.w8(32'h3c29c4a5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9470793),
	.w1(32'hbb98646c),
	.w2(32'hbc45cbf8),
	.w3(32'h3c580326),
	.w4(32'hbb8824d0),
	.w5(32'hbca6b192),
	.w6(32'hbc07e53b),
	.w7(32'h3c1a0b73),
	.w8(32'h3b99e5a9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c867113),
	.w1(32'hba8155a4),
	.w2(32'hbcbf5b2e),
	.w3(32'h3c1b5512),
	.w4(32'h3c4cc085),
	.w5(32'hbc40c469),
	.w6(32'h3cc185fd),
	.w7(32'h3c8031c0),
	.w8(32'h3c8bc152),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46e835),
	.w1(32'h3b4c36a4),
	.w2(32'hbcb19482),
	.w3(32'h3ad1ca3a),
	.w4(32'hbb1e1ece),
	.w5(32'h3bfbfcbd),
	.w6(32'hbcc0f8cd),
	.w7(32'h3c81cf02),
	.w8(32'h3c8efb5b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4625ad),
	.w1(32'hbcbd9aa4),
	.w2(32'h3ada8123),
	.w3(32'h3c4af97d),
	.w4(32'hbcc76bab),
	.w5(32'hbc04d13b),
	.w6(32'h3c404147),
	.w7(32'h3b86c337),
	.w8(32'h3cbb2056),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3edb87),
	.w1(32'hbb5a04c4),
	.w2(32'h3b33d0a2),
	.w3(32'hbbd959b6),
	.w4(32'h3bb4787f),
	.w5(32'h3c3d04b3),
	.w6(32'h3bb20464),
	.w7(32'hbb0eeed8),
	.w8(32'hbb43c58e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113db1),
	.w1(32'h3c0b5af5),
	.w2(32'h3bff6bd5),
	.w3(32'h3b839133),
	.w4(32'h3bb36109),
	.w5(32'hbb07719e),
	.w6(32'h3b085cfe),
	.w7(32'hbb40f5b9),
	.w8(32'hbc0278f0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8bc3c),
	.w1(32'hbbdf4e67),
	.w2(32'hbb145a81),
	.w3(32'hbb7fc5ef),
	.w4(32'hbafa1dfc),
	.w5(32'hbc1ed946),
	.w6(32'h3a36515c),
	.w7(32'h3c40da3c),
	.w8(32'h3c66be9e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccb0b1),
	.w1(32'h3c90df21),
	.w2(32'hbc87533f),
	.w3(32'hbbac7d5c),
	.w4(32'hba9cf6ee),
	.w5(32'h3bbc27b0),
	.w6(32'hbbed5dd6),
	.w7(32'h3c3f1da5),
	.w8(32'h3c950fec),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcd765a),
	.w1(32'hbd3c1aa8),
	.w2(32'hbd48eeaa),
	.w3(32'h3d50537c),
	.w4(32'hbdedffb3),
	.w5(32'hbe247cc4),
	.w6(32'hbc89a198),
	.w7(32'h3c8cb6b4),
	.w8(32'h3c9807de),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30040d),
	.w1(32'hbc0d12f0),
	.w2(32'h3ca5da18),
	.w3(32'hbd03218f),
	.w4(32'hb9980637),
	.w5(32'hbc33bdeb),
	.w6(32'h3c8dd074),
	.w7(32'hbb9e218c),
	.w8(32'h3cb01543),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab419),
	.w1(32'hbb238135),
	.w2(32'h3ceb62fb),
	.w3(32'h3c89f4e7),
	.w4(32'h3b79939e),
	.w5(32'h3d0a80ee),
	.w6(32'hbc2222de),
	.w7(32'hbcececd8),
	.w8(32'hbdc41fd9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d048c9d),
	.w1(32'h3b483d1b),
	.w2(32'h3991618f),
	.w3(32'h3c9c4bfb),
	.w4(32'hb9837cf8),
	.w5(32'h3b6183b3),
	.w6(32'hbd020287),
	.w7(32'hbbb36c31),
	.w8(32'hbad7df5d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2327a7),
	.w1(32'h3c0d82b6),
	.w2(32'hbc46fc1f),
	.w3(32'h3c10bedf),
	.w4(32'h3ba0ab7c),
	.w5(32'hbb847144),
	.w6(32'h38790b5f),
	.w7(32'hbb8a1b6f),
	.w8(32'h3ca4e3b4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07028),
	.w1(32'hbc5a4049),
	.w2(32'hbcd9a34b),
	.w3(32'hbc6d0108),
	.w4(32'h3c5087f6),
	.w5(32'h3d0877c9),
	.w6(32'hbb2c7eff),
	.w7(32'hbc37bc98),
	.w8(32'hbc1691bf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1dbee2),
	.w1(32'hbc524c56),
	.w2(32'hbb714111),
	.w3(32'h3c2c3dcd),
	.w4(32'hba010174),
	.w5(32'h3b98d229),
	.w6(32'h3b9de6d8),
	.w7(32'hbbadda56),
	.w8(32'hbc4cf69c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63ce9b),
	.w1(32'h3c266874),
	.w2(32'h3b05959f),
	.w3(32'h3c3cf315),
	.w4(32'h3caf1cbc),
	.w5(32'h3ba6907b),
	.w6(32'hbc0147cd),
	.w7(32'h3c4c8811),
	.w8(32'h3be7945f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61716d),
	.w1(32'hbc3c999d),
	.w2(32'hbc273f14),
	.w3(32'hbc12ab4e),
	.w4(32'hbb803e0f),
	.w5(32'hbc0506d0),
	.w6(32'hbb90aa40),
	.w7(32'hbcb9261e),
	.w8(32'h3d0ca3b3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc781865),
	.w1(32'hb833225a),
	.w2(32'hbc448de7),
	.w3(32'hbc5a65b6),
	.w4(32'hbc6eaa79),
	.w5(32'hbc4105b8),
	.w6(32'h3d5205c1),
	.w7(32'h3c92381b),
	.w8(32'h3d5173eb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29bd21),
	.w1(32'hbb9fcb62),
	.w2(32'h3a840363),
	.w3(32'hbc121866),
	.w4(32'h3bc2dfee),
	.w5(32'h3b73bc50),
	.w6(32'h3af246ad),
	.w7(32'h3c0d5855),
	.w8(32'hbc91ea73),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32a9a8),
	.w1(32'hbc7ed8e7),
	.w2(32'h3c948a45),
	.w3(32'h3adbad25),
	.w4(32'h3c048689),
	.w5(32'hbc3d3853),
	.w6(32'hbc5726fe),
	.w7(32'h38f71393),
	.w8(32'h3b991164),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e4faa),
	.w1(32'hb8a7d66a),
	.w2(32'hbb9bda93),
	.w3(32'hbbfdb1f1),
	.w4(32'h39e72c8b),
	.w5(32'hbb9e22a9),
	.w6(32'hbb945f52),
	.w7(32'hbc0a354c),
	.w8(32'hba16020b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7008c),
	.w1(32'hbb5ee09e),
	.w2(32'hbb6e835a),
	.w3(32'hbbb70ad1),
	.w4(32'h3bf3daff),
	.w5(32'hbca335ab),
	.w6(32'h3bc2e204),
	.w7(32'h3c9c67ff),
	.w8(32'hbd0130e9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af30805),
	.w1(32'h3c111a12),
	.w2(32'h3b55fa6c),
	.w3(32'h3b125dbb),
	.w4(32'hbb5b540b),
	.w5(32'hbb600a02),
	.w6(32'hbcbbb2c4),
	.w7(32'h3c18844f),
	.w8(32'h3cc9a769),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d0d4c),
	.w1(32'hbb57be8e),
	.w2(32'hbc30f087),
	.w3(32'hbc9d7651),
	.w4(32'h3c7cbb07),
	.w5(32'h3c96c501),
	.w6(32'h3c0df610),
	.w7(32'h3c10aab5),
	.w8(32'h3c5342da),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc745cb3),
	.w1(32'hbc88a699),
	.w2(32'hbb9d29e2),
	.w3(32'h3b508e09),
	.w4(32'hbc3962e5),
	.w5(32'hbbc7c7fd),
	.w6(32'h3c93e65f),
	.w7(32'hbbff5fc6),
	.w8(32'h3ba021b9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66a906),
	.w1(32'hbc3299cb),
	.w2(32'h3ccaf9c1),
	.w3(32'h3a44cf80),
	.w4(32'hbc31a3fe),
	.w5(32'hbc61a30e),
	.w6(32'h3c3b1569),
	.w7(32'h3b3f5d89),
	.w8(32'hbb3ad9f9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5b199),
	.w1(32'hbbc25919),
	.w2(32'hba963adf),
	.w3(32'hbc2bf75f),
	.w4(32'hbcb1a887),
	.w5(32'hba229e6a),
	.w6(32'hbc3d4da3),
	.w7(32'hbd0059fe),
	.w8(32'h3c310d3c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1d7ad),
	.w1(32'hbb9e2b9c),
	.w2(32'hbc9606f3),
	.w3(32'h3b75ca80),
	.w4(32'h3917e8ba),
	.w5(32'hbb6d60aa),
	.w6(32'h3bf6e5de),
	.w7(32'hbc0d471d),
	.w8(32'h3b29b5c3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc9fa),
	.w1(32'hbbdc7abe),
	.w2(32'h3bfea66e),
	.w3(32'hbc66ec54),
	.w4(32'hbc7ad894),
	.w5(32'h3ba6249b),
	.w6(32'hbc1fd472),
	.w7(32'h3c31b9f7),
	.w8(32'hba487f89),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4728de),
	.w1(32'h3c86fe8d),
	.w2(32'h3ba88b05),
	.w3(32'h3cabacc6),
	.w4(32'h3c54f4d3),
	.w5(32'h3c7f4fd3),
	.w6(32'hbc935ae8),
	.w7(32'hbb9dad50),
	.w8(32'hbc269434),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca65a0a),
	.w1(32'hbcadb5a8),
	.w2(32'h3aac4fd8),
	.w3(32'h3b1edbd7),
	.w4(32'hbc73f2de),
	.w5(32'h398be093),
	.w6(32'h3c1e0c77),
	.w7(32'hbc5d9eae),
	.w8(32'hbcd3b7c8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c926d46),
	.w1(32'h3c5c4e55),
	.w2(32'h3d08822d),
	.w3(32'h3be66a79),
	.w4(32'h3ca0aa94),
	.w5(32'h3afd3d04),
	.w6(32'hbc8ceb88),
	.w7(32'h3d022d7f),
	.w8(32'hbd29cf2a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d0b35),
	.w1(32'h3b998f1b),
	.w2(32'hbc212cc3),
	.w3(32'hbbbc337e),
	.w4(32'hbd263696),
	.w5(32'hbcbd4819),
	.w6(32'hbcc0bc1c),
	.w7(32'h3d14551a),
	.w8(32'h3cc114b1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0128ca),
	.w1(32'hbbb002f5),
	.w2(32'hbb08feef),
	.w3(32'h3c006e24),
	.w4(32'hbc0aec79),
	.w5(32'h3ba16e71),
	.w6(32'h3b09607d),
	.w7(32'h3c2ff216),
	.w8(32'hbc314b0b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b98e0),
	.w1(32'hbb801a0e),
	.w2(32'hbc50ca7e),
	.w3(32'h3b1ccc24),
	.w4(32'hbab07d6f),
	.w5(32'h3c244f0d),
	.w6(32'hbb582a3f),
	.w7(32'hbba57d49),
	.w8(32'h3c1bea64),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0054bc),
	.w1(32'h3b2d357f),
	.w2(32'h3b81e377),
	.w3(32'h39dec1c7),
	.w4(32'hbc1868f5),
	.w5(32'hbc9cf0cf),
	.w6(32'h3b3a97e1),
	.w7(32'h3bb06a78),
	.w8(32'h3d459528),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06d510),
	.w1(32'hbd5b3d8d),
	.w2(32'hbca3f327),
	.w3(32'h3af2dfa0),
	.w4(32'hbc6b3153),
	.w5(32'hbcb10e97),
	.w6(32'h3abf663d),
	.w7(32'h3c59baab),
	.w8(32'h3c81a589),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5da1cf),
	.w1(32'h3beacc9e),
	.w2(32'hba957697),
	.w3(32'h3b139e7a),
	.w4(32'h3bb97971),
	.w5(32'h3c2ff43b),
	.w6(32'h3bd7b196),
	.w7(32'h398facfc),
	.w8(32'h3c4d296a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736f67),
	.w1(32'h3b9e768e),
	.w2(32'h3d153009),
	.w3(32'hbba34387),
	.w4(32'hbd04edb8),
	.w5(32'hbc9f16af),
	.w6(32'hbb3a79b2),
	.w7(32'hbbb413e0),
	.w8(32'hbd07490c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cecea6a),
	.w1(32'h3b8eac08),
	.w2(32'hbbaa68db),
	.w3(32'h3b39c32a),
	.w4(32'hbc896281),
	.w5(32'hbc10605f),
	.w6(32'hbcbe3bdd),
	.w7(32'hbc770cb6),
	.w8(32'h3a0f1cda),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a97f),
	.w1(32'h3ae0cf43),
	.w2(32'hbc291d38),
	.w3(32'h3a97fd13),
	.w4(32'h3a36ef18),
	.w5(32'hbb9d7b7d),
	.w6(32'hbab57de2),
	.w7(32'h3c0ffce2),
	.w8(32'hbb02afff),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc703f10),
	.w1(32'hba53037f),
	.w2(32'h3b878763),
	.w3(32'h3c26e935),
	.w4(32'h3c15bd26),
	.w5(32'hbc1ae086),
	.w6(32'h3c21363b),
	.w7(32'h3a8ae8b2),
	.w8(32'hbb0c3977),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36f397),
	.w1(32'h3c953e2d),
	.w2(32'h3bd97c65),
	.w3(32'hbbee4524),
	.w4(32'hbb63162c),
	.w5(32'hbb2c4877),
	.w6(32'h3bb98b00),
	.w7(32'hbb6bc9da),
	.w8(32'h3be02528),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c2574),
	.w1(32'hbb0b2bd7),
	.w2(32'hb90d9c6b),
	.w3(32'hb986b43e),
	.w4(32'hb95da270),
	.w5(32'h3c0fff79),
	.w6(32'h3c37f433),
	.w7(32'h3b8b54de),
	.w8(32'hbc6b9ebf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b0f4),
	.w1(32'hbbef610c),
	.w2(32'h3c5e51ba),
	.w3(32'h3c3fa2d3),
	.w4(32'h3c08c8bf),
	.w5(32'h3b7341d9),
	.w6(32'hbc40767a),
	.w7(32'hba5baa0b),
	.w8(32'h3c718866),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c056eeb),
	.w1(32'hbadb5e37),
	.w2(32'hbb94d5c7),
	.w3(32'hbb2d709f),
	.w4(32'hba78b1da),
	.w5(32'h3c0a355e),
	.w6(32'h3c345876),
	.w7(32'hbcbbbc64),
	.w8(32'h3c43d553),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75008b),
	.w1(32'hbc0dcf3e),
	.w2(32'h3c987c7c),
	.w3(32'hbb8dc33d),
	.w4(32'h3b0d7b77),
	.w5(32'h3cace476),
	.w6(32'hbc7798d4),
	.w7(32'hbc2cbd89),
	.w8(32'hbc9582de),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf28688),
	.w1(32'h3cbf42dd),
	.w2(32'h3c1ce5b4),
	.w3(32'h3c430fe5),
	.w4(32'hbb417bcd),
	.w5(32'hbb9b8b66),
	.w6(32'hba321c08),
	.w7(32'hbb3d6100),
	.w8(32'hbcba70b0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd22be2),
	.w1(32'hbbaee64c),
	.w2(32'hbd3496b0),
	.w3(32'h3a0be755),
	.w4(32'h3c09abc1),
	.w5(32'h3c82ed00),
	.w6(32'h3b8ca77b),
	.w7(32'h3c1555fe),
	.w8(32'h3d2fb560),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd21398),
	.w1(32'hbb9461f2),
	.w2(32'hbc930513),
	.w3(32'h3b30dd88),
	.w4(32'hbaf8f831),
	.w5(32'hbb1261f9),
	.w6(32'h3ca6207c),
	.w7(32'h3adf0cce),
	.w8(32'h3c789650),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc674084),
	.w1(32'hbc6e4f1e),
	.w2(32'h3cb5a3cf),
	.w3(32'hbac7f7c5),
	.w4(32'hbd0cad89),
	.w5(32'h3bcdebbf),
	.w6(32'hbbd76fbc),
	.w7(32'hbcd90e04),
	.w8(32'hbcfdd515),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cc1e3),
	.w1(32'hb9f40d2e),
	.w2(32'h3c79d322),
	.w3(32'h3c9cce7a),
	.w4(32'h3bd63ef9),
	.w5(32'h3c8cf3d8),
	.w6(32'h393038ff),
	.w7(32'h3a3a039f),
	.w8(32'hbc451f83),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfadc26),
	.w1(32'h3c8147a4),
	.w2(32'h3bb2ab3a),
	.w3(32'h3ca63010),
	.w4(32'h3a5ebf58),
	.w5(32'h3c9de245),
	.w6(32'hbb3c6b1b),
	.w7(32'hbcb0ae9f),
	.w8(32'hbca438ba),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14ea64),
	.w1(32'hbb9d130d),
	.w2(32'hbc382623),
	.w3(32'hbbba579f),
	.w4(32'hbb976803),
	.w5(32'h3b6fad75),
	.w6(32'h3a748028),
	.w7(32'hbc898d25),
	.w8(32'h3c61b27b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4e05),
	.w1(32'hbc970573),
	.w2(32'hbade4732),
	.w3(32'hbc49901e),
	.w4(32'h3bb2547f),
	.w5(32'hbc16a10e),
	.w6(32'hbc3543a6),
	.w7(32'h3cb7137b),
	.w8(32'h3c4309e7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35a9c9),
	.w1(32'h3c00a740),
	.w2(32'hbbd6e11b),
	.w3(32'hbb11d0fd),
	.w4(32'h3a0f9ae4),
	.w5(32'h3cf5557e),
	.w6(32'h3c0a213c),
	.w7(32'h39812789),
	.w8(32'hbcca29a7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc232ea),
	.w1(32'hbb0e7f34),
	.w2(32'h3c30b743),
	.w3(32'h3c2c057b),
	.w4(32'h3baab538),
	.w5(32'h3c284a20),
	.w6(32'hbc8205fa),
	.w7(32'hbbfe6bf0),
	.w8(32'hbae9f656),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c445a0f),
	.w1(32'h3ba57457),
	.w2(32'h3a7cb83e),
	.w3(32'h3ad06bb3),
	.w4(32'hba3f27a2),
	.w5(32'hbb2abf96),
	.w6(32'h3c8770c8),
	.w7(32'h3b94ada6),
	.w8(32'h3c448b18),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf7896),
	.w1(32'hbb698eb6),
	.w2(32'h3b62f863),
	.w3(32'h3b3747c0),
	.w4(32'hbbb251a1),
	.w5(32'hbbe2d5cf),
	.w6(32'h3bbc1bfa),
	.w7(32'h3c39ebf1),
	.w8(32'h3b7f2813),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50c1a3),
	.w1(32'hbc6abfb9),
	.w2(32'h3b98b838),
	.w3(32'hbb5ce003),
	.w4(32'h3b895e0d),
	.w5(32'h3ab63563),
	.w6(32'hbbb2caf8),
	.w7(32'h3bf8fb9c),
	.w8(32'h3c0f8331),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891909),
	.w1(32'h3bb8ea53),
	.w2(32'h394c7c5a),
	.w3(32'h3be85b5a),
	.w4(32'hba51da26),
	.w5(32'h3bf23453),
	.w6(32'h3b380185),
	.w7(32'hb9a126c7),
	.w8(32'hbc8fc7b5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b3d94),
	.w1(32'hbc2f1c88),
	.w2(32'h3c196867),
	.w3(32'h3a0962d6),
	.w4(32'h3b01c8cc),
	.w5(32'hbc0bb9fb),
	.w6(32'h3bafd774),
	.w7(32'h3ac6d1cc),
	.w8(32'h3c3c2f3d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43475d),
	.w1(32'h3bfac58b),
	.w2(32'h3c0516a4),
	.w3(32'h3c54f676),
	.w4(32'hb9f35256),
	.w5(32'h3c6eb8fd),
	.w6(32'h3be71dd0),
	.w7(32'hbcb0f732),
	.w8(32'hbbefad3e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e984),
	.w1(32'hbbd84085),
	.w2(32'h3a8a6050),
	.w3(32'h3c319665),
	.w4(32'hbb51b730),
	.w5(32'hbbf7edee),
	.w6(32'h3c2a32cc),
	.w7(32'hbbd6b7dc),
	.w8(32'h3c8bf1f6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d42b8),
	.w1(32'hbc5087a0),
	.w2(32'hbc8d4224),
	.w3(32'hbc1957d7),
	.w4(32'hbb1c6f14),
	.w5(32'hbc22366a),
	.w6(32'h3cbe5cf9),
	.w7(32'h3bd30bc1),
	.w8(32'hbc00dff2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c88de),
	.w1(32'hbcf90101),
	.w2(32'hbb47084a),
	.w3(32'h3c19d88e),
	.w4(32'hbc750f21),
	.w5(32'hbcdde116),
	.w6(32'h3cb76157),
	.w7(32'h3b953ca4),
	.w8(32'h3d00d3a9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1b7ef),
	.w1(32'h3b800b32),
	.w2(32'hbd248bfe),
	.w3(32'hbb2437a1),
	.w4(32'hbc738d1f),
	.w5(32'hbc1f84c5),
	.w6(32'h3bab2fa2),
	.w7(32'hbc85cc44),
	.w8(32'h39d94666),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8969e2),
	.w1(32'h3b9d4418),
	.w2(32'h3c54c7bf),
	.w3(32'h3c85f0a6),
	.w4(32'h3c115c3f),
	.w5(32'h3bdbb881),
	.w6(32'hbd0b9239),
	.w7(32'hbb941fb3),
	.w8(32'hbc5ab749),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5f36),
	.w1(32'hbbb1a1e3),
	.w2(32'h3a9d786b),
	.w3(32'h3c684ac1),
	.w4(32'hbb491aed),
	.w5(32'h3bbbc3ac),
	.w6(32'hbc833200),
	.w7(32'hbb856f88),
	.w8(32'hbc5ee806),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3f17e),
	.w1(32'h3acfc624),
	.w2(32'h3a9f6dcd),
	.w3(32'hb9e374d7),
	.w4(32'hbb079cc6),
	.w5(32'hbc30d177),
	.w6(32'hbbc6a5b5),
	.w7(32'hbb03d47e),
	.w8(32'hbb278b95),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122672),
	.w1(32'hbb81a0cd),
	.w2(32'hbbf7b03a),
	.w3(32'hb7dc4804),
	.w4(32'hbc9a58a5),
	.w5(32'hbb273b3f),
	.w6(32'hbc1b63f9),
	.w7(32'h3c8715af),
	.w8(32'hbc13e071),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14c965),
	.w1(32'hbc4c4c98),
	.w2(32'hbc42654d),
	.w3(32'h3c243b30),
	.w4(32'h3b1cf62c),
	.w5(32'hbc0195c8),
	.w6(32'h3c150530),
	.w7(32'hbc45440b),
	.w8(32'hbcd19884),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba71c9),
	.w1(32'h3b89044e),
	.w2(32'hbbfe3d22),
	.w3(32'h3a9464ff),
	.w4(32'hbc84f735),
	.w5(32'hbaa46582),
	.w6(32'hbbf34e89),
	.w7(32'h3c5deed9),
	.w8(32'hbb8bf408),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c529841),
	.w1(32'hbb8b4537),
	.w2(32'h3bf0be1f),
	.w3(32'hba21c033),
	.w4(32'hbba49014),
	.w5(32'h39c90ee4),
	.w6(32'hbc0d987d),
	.w7(32'hbcc00203),
	.w8(32'h3d725c9f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2bc2b),
	.w1(32'hbc7931e1),
	.w2(32'h3c1d3415),
	.w3(32'hbb401aea),
	.w4(32'h3b89ee65),
	.w5(32'h3bfc1a65),
	.w6(32'hb98e262d),
	.w7(32'hbca74b85),
	.w8(32'hba94ae9c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed70cd),
	.w1(32'hbcd1a411),
	.w2(32'hb8583f40),
	.w3(32'hbc0f8624),
	.w4(32'h3c1e9180),
	.w5(32'hb9b84215),
	.w6(32'h3cd59b9a),
	.w7(32'h3b72cce1),
	.w8(32'hbb4aea9f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33ddae),
	.w1(32'hbbc6d5a1),
	.w2(32'hbc582a73),
	.w3(32'h3c0693fa),
	.w4(32'hbca4f584),
	.w5(32'hbc852748),
	.w6(32'h3b92b52c),
	.w7(32'hbaf016d2),
	.w8(32'h3cf3cb4e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc818e93),
	.w1(32'hbc312ec7),
	.w2(32'hbaa1f10c),
	.w3(32'hbbf16dcd),
	.w4(32'hb82d4ee6),
	.w5(32'hbb59fcff),
	.w6(32'hbc96610d),
	.w7(32'hbb034e8a),
	.w8(32'h3c81af3f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67deb5),
	.w1(32'h3be59053),
	.w2(32'h3c237647),
	.w3(32'hbb8c2291),
	.w4(32'h3ba4c019),
	.w5(32'hbb4f9dba),
	.w6(32'h3c2b8f09),
	.w7(32'hbc2db4df),
	.w8(32'h3c84508b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccbaa8),
	.w1(32'h3ca98476),
	.w2(32'hbbc9a54f),
	.w3(32'h3c1883c4),
	.w4(32'hbb35a75e),
	.w5(32'hbb08ec6e),
	.w6(32'hbc9d2f58),
	.w7(32'hbba98bce),
	.w8(32'h3b938c85),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7249b3),
	.w1(32'h3bbeca83),
	.w2(32'h38e20ae1),
	.w3(32'hb94ad1f1),
	.w4(32'hbc24095a),
	.w5(32'hbb9c498b),
	.w6(32'h3af0c48a),
	.w7(32'hbc103324),
	.w8(32'h3aedb755),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4413c),
	.w1(32'h3c92a636),
	.w2(32'h3b9fd64f),
	.w3(32'h3bf99a32),
	.w4(32'hbacaf111),
	.w5(32'h3af5ce7e),
	.w6(32'hbc7caaae),
	.w7(32'h3c5dbfea),
	.w8(32'h3c343709),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c174796),
	.w1(32'h3c2bbd32),
	.w2(32'hbb36fc21),
	.w3(32'hbb0d41eb),
	.w4(32'h3befee02),
	.w5(32'h3bb5277c),
	.w6(32'hbccf8710),
	.w7(32'h3c4f1e40),
	.w8(32'hbb54df9c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bee6e),
	.w1(32'h3bfdabbf),
	.w2(32'hbbd771c1),
	.w3(32'hbc076459),
	.w4(32'hbc0f9954),
	.w5(32'hbcafe117),
	.w6(32'hbb7726a5),
	.w7(32'hbc6362bc),
	.w8(32'h3d2837b3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4ab2b),
	.w1(32'h3c52ce3d),
	.w2(32'h3c3ac2af),
	.w3(32'h3b8bdc09),
	.w4(32'h3bb69998),
	.w5(32'hbb3e4454),
	.w6(32'hbcb9cdf7),
	.w7(32'hbb49d949),
	.w8(32'h3c13184f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7394b),
	.w1(32'hbb42a23e),
	.w2(32'h3c53e309),
	.w3(32'h39d7416d),
	.w4(32'h3ba058d2),
	.w5(32'h3bfe242b),
	.w6(32'hbbdc2105),
	.w7(32'hbbce0638),
	.w8(32'hbc8f3537),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ad01e),
	.w1(32'hbc58d67a),
	.w2(32'hbc54a882),
	.w3(32'hbbed455e),
	.w4(32'hbcb92c10),
	.w5(32'h3c2bc1c1),
	.w6(32'h3b8dbd3a),
	.w7(32'h3c4e5840),
	.w8(32'hbd5cf2e7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80a77e),
	.w1(32'hbc9066f8),
	.w2(32'h3adb7093),
	.w3(32'hbc0eb221),
	.w4(32'h3c565b38),
	.w5(32'hbc939b6a),
	.w6(32'h3cd89074),
	.w7(32'hbcaed9a5),
	.w8(32'h3d71df8e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a05e1),
	.w1(32'h3ce1232b),
	.w2(32'h3ac506da),
	.w3(32'h3bc181fa),
	.w4(32'h3b7b182c),
	.w5(32'hb93315b0),
	.w6(32'hbca8552a),
	.w7(32'h3b4852b7),
	.w8(32'h3be7d384),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c84ad),
	.w1(32'h3b2095a2),
	.w2(32'h3b6820da),
	.w3(32'h3aaea937),
	.w4(32'h3a5f1157),
	.w5(32'hbbcc4740),
	.w6(32'hbb19a6c0),
	.w7(32'hbc312e46),
	.w8(32'h3c9465dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce61717),
	.w1(32'hbbe46e26),
	.w2(32'h3b1fff85),
	.w3(32'hbc0e1e12),
	.w4(32'hbc9c9fea),
	.w5(32'h3d136d1d),
	.w6(32'h3c2e359c),
	.w7(32'h3caae9ac),
	.w8(32'hbd386ba5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc21984),
	.w1(32'hbc876e25),
	.w2(32'hbced4d7d),
	.w3(32'hb8869b75),
	.w4(32'hbacfa9d8),
	.w5(32'hbcec94c1),
	.w6(32'h3cacff66),
	.w7(32'h3c1ab8b7),
	.w8(32'h3ce18f75),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae74b7),
	.w1(32'hbc097500),
	.w2(32'h3b9bbcc8),
	.w3(32'h3be7dcb0),
	.w4(32'hbbe38263),
	.w5(32'h3b3195c7),
	.w6(32'h3b3882c5),
	.w7(32'hbb806fcc),
	.w8(32'h3bcad6d2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914bc52),
	.w1(32'h3b4741c0),
	.w2(32'hbb7a1449),
	.w3(32'h3bcc84a0),
	.w4(32'h3b8abb1b),
	.w5(32'h3b95e209),
	.w6(32'h3b20f1fa),
	.w7(32'hbc93e3c2),
	.w8(32'hbc679a80),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cda13),
	.w1(32'hbbad5937),
	.w2(32'hbc83cc6e),
	.w3(32'hbcc53968),
	.w4(32'hbbad8d17),
	.w5(32'hbbb6f840),
	.w6(32'hbc06bcdf),
	.w7(32'hbc6f0156),
	.w8(32'hbc299144),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829adb),
	.w1(32'hbc2e8b9b),
	.w2(32'hbc95796b),
	.w3(32'hbc361c0a),
	.w4(32'hbcdf5ea4),
	.w5(32'h3d28fb69),
	.w6(32'hbc34e076),
	.w7(32'h3d2cd5d9),
	.w8(32'hbde9d546),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8f53f4),
	.w1(32'hbcb25fe2),
	.w2(32'hbc3981d8),
	.w3(32'h39e61cf9),
	.w4(32'hbbab204f),
	.w5(32'h3b4a5f10),
	.w6(32'h3d30f691),
	.w7(32'h3cade5a5),
	.w8(32'h399abed1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe0553),
	.w1(32'hbc4c5bd7),
	.w2(32'h3b0eec9b),
	.w3(32'hbc02a2e4),
	.w4(32'h3b395fa9),
	.w5(32'h3b6c03a4),
	.w6(32'h3c5358a3),
	.w7(32'h3c2a6ce0),
	.w8(32'hbc372205),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75bc4f),
	.w1(32'h3bb77749),
	.w2(32'hbb1a0bb2),
	.w3(32'hbbadd242),
	.w4(32'hbbac714d),
	.w5(32'hbc2b67bd),
	.w6(32'hbb81664c),
	.w7(32'h3bd0f828),
	.w8(32'h3b5d06c8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13b2b6),
	.w1(32'h3a421fac),
	.w2(32'h3c46d002),
	.w3(32'h3a5ff4ac),
	.w4(32'hbc20ede6),
	.w5(32'hbb785c6d),
	.w6(32'hba758fe4),
	.w7(32'hbbf55c8d),
	.w8(32'h3c3ceebb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89e267),
	.w1(32'h3c85cabe),
	.w2(32'h3b9b824d),
	.w3(32'hbced8001),
	.w4(32'hbb5d522d),
	.w5(32'h3b888e5d),
	.w6(32'h3b0cc86a),
	.w7(32'hbca22103),
	.w8(32'hbbd636c1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbba586),
	.w1(32'h3ae6f886),
	.w2(32'h3b9e9d1a),
	.w3(32'hbc7b7155),
	.w4(32'h3b7de734),
	.w5(32'h3c2a7424),
	.w6(32'h3abd5f63),
	.w7(32'hbc0a93f3),
	.w8(32'h3b197485),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98d184),
	.w1(32'hb95f2cf3),
	.w2(32'h3c86a539),
	.w3(32'hbb109c89),
	.w4(32'hbc4e251a),
	.w5(32'hba1954a2),
	.w6(32'hbb237d2c),
	.w7(32'hbad77587),
	.w8(32'h3a894ddd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c789),
	.w1(32'hbc0d2ee6),
	.w2(32'h3a57afba),
	.w3(32'h3c296fb8),
	.w4(32'h3b388f57),
	.w5(32'hbb22e08d),
	.w6(32'h3c3c5ef6),
	.w7(32'h3b29f6e2),
	.w8(32'h3b72fb54),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b1552),
	.w1(32'h3aa5ea93),
	.w2(32'hbb137ade),
	.w3(32'h3acc6e1b),
	.w4(32'hbc3ad933),
	.w5(32'hbb82f8d8),
	.w6(32'hbb07e551),
	.w7(32'h3c98492e),
	.w8(32'h3b990f85),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9dd25),
	.w1(32'h3c8bbc6c),
	.w2(32'h3c3b3929),
	.w3(32'hbb308473),
	.w4(32'h3b433a46),
	.w5(32'h3cc12ae5),
	.w6(32'hbc905c70),
	.w7(32'h3c12692e),
	.w8(32'hbcfe0a0f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c884c48),
	.w1(32'hbcd372c8),
	.w2(32'hbbf91ebc),
	.w3(32'hbc1a6d71),
	.w4(32'h39884a91),
	.w5(32'hb858a850),
	.w6(32'h3cd79079),
	.w7(32'h3bcf2254),
	.w8(32'h3bc76d9c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07efca),
	.w1(32'hbb1cf94b),
	.w2(32'h3b820423),
	.w3(32'h3b1b2593),
	.w4(32'h3beb0580),
	.w5(32'hbba44f0e),
	.w6(32'h3bdd22af),
	.w7(32'h3b198ca8),
	.w8(32'hbb5995ae),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4407a),
	.w1(32'h3b8e8c67),
	.w2(32'hbc0b1ee2),
	.w3(32'h39ef843d),
	.w4(32'hbc019f71),
	.w5(32'hbc5dd19c),
	.w6(32'hbbb40d05),
	.w7(32'hbbd22f40),
	.w8(32'h3bd72a3e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule