module layer_8_featuremap_253(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a293b),
	.w1(32'hbb6a6b16),
	.w2(32'h3bff2f37),
	.w3(32'hbc40b9a5),
	.w4(32'hbbf49d52),
	.w5(32'h3c1afaf0),
	.w6(32'hbcdb02af),
	.w7(32'hbc19d5b8),
	.w8(32'h3b4a6e9a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dac6a),
	.w1(32'hba8770bd),
	.w2(32'hbb8c590b),
	.w3(32'h3b34cdc3),
	.w4(32'h3baeb6a7),
	.w5(32'h3b035be7),
	.w6(32'h3b8e9faf),
	.w7(32'h3bb186da),
	.w8(32'h3b9c19a6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac972ab),
	.w1(32'h3c3530c8),
	.w2(32'h3ca9a84c),
	.w3(32'h3b926672),
	.w4(32'h3ba3aeb5),
	.w5(32'h3c41aa94),
	.w6(32'h3b87d376),
	.w7(32'h3b76e683),
	.w8(32'hbb346cdf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2da18),
	.w1(32'h3c5e4a6b),
	.w2(32'h3c65d93f),
	.w3(32'h3b81cde1),
	.w4(32'h3ac390d1),
	.w5(32'h3c85af75),
	.w6(32'hbccd250e),
	.w7(32'hbcdee4d2),
	.w8(32'hbcb11eec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8295fb),
	.w1(32'h3bc4e8f3),
	.w2(32'h3bbad65e),
	.w3(32'h3c72068f),
	.w4(32'hbae4610d),
	.w5(32'hbbad4a19),
	.w6(32'h3b8bb2fd),
	.w7(32'h3b03214b),
	.w8(32'h3aa4fb7b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb53ab4),
	.w1(32'h3bba668d),
	.w2(32'hba893d3d),
	.w3(32'h3c588c2c),
	.w4(32'hba8ec42f),
	.w5(32'hbc46da18),
	.w6(32'h3c1a730e),
	.w7(32'h3ae33d1b),
	.w8(32'hbc85659b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcde023),
	.w1(32'h3b209433),
	.w2(32'h3b9f8bf1),
	.w3(32'hbbeaedf4),
	.w4(32'hbbe2bb29),
	.w5(32'hbb7d182c),
	.w6(32'hba7715bd),
	.w7(32'hbb0e4d6a),
	.w8(32'hbb09c229),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2271),
	.w1(32'hbb2b92fd),
	.w2(32'hbb5c69ac),
	.w3(32'h398e7666),
	.w4(32'h3c92eb51),
	.w5(32'h3ca955f2),
	.w6(32'h3ba4a151),
	.w7(32'h3c2fa169),
	.w8(32'h3c71e727),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe333e),
	.w1(32'h3b2e8a4e),
	.w2(32'h39a4edef),
	.w3(32'h3c531c17),
	.w4(32'hbb5a7edf),
	.w5(32'hbc28fde9),
	.w6(32'hbbb7cd43),
	.w7(32'hbc319b70),
	.w8(32'hbc1a1bdb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebe9d6),
	.w1(32'h3b8bbb67),
	.w2(32'h3d077e52),
	.w3(32'hbc3010b2),
	.w4(32'hbc82a507),
	.w5(32'hbc481810),
	.w6(32'hbc437040),
	.w7(32'hbb6d26f6),
	.w8(32'h3b8aa22e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95024e),
	.w1(32'h3c758d17),
	.w2(32'h3c488d6b),
	.w3(32'hbcedc1a8),
	.w4(32'h3b73f554),
	.w5(32'h3cda1a4b),
	.w6(32'hbc060ffc),
	.w7(32'hbc212ee7),
	.w8(32'hb8e63c6f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6e5a),
	.w1(32'h3a967869),
	.w2(32'h3c52510b),
	.w3(32'h3b48ecf2),
	.w4(32'hbc1ce50a),
	.w5(32'hbb4608c0),
	.w6(32'hbc8fb1c6),
	.w7(32'hbca06ec1),
	.w8(32'hbc90faf2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b014),
	.w1(32'h3980a9ac),
	.w2(32'h3bf30403),
	.w3(32'h3b27ab29),
	.w4(32'h3bb39e52),
	.w5(32'h3c679f9a),
	.w6(32'hbca9b8fd),
	.w7(32'hbca2c343),
	.w8(32'hbc996d89),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4051fc),
	.w1(32'hbba1e677),
	.w2(32'h3a3d92f5),
	.w3(32'h3c2fff7b),
	.w4(32'hbc83f92c),
	.w5(32'hbc6cfd51),
	.w6(32'h3c0be54d),
	.w7(32'h3bcc5fc2),
	.w8(32'h3bdf4ff6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba330bc),
	.w1(32'hba60e872),
	.w2(32'h3b4a2e27),
	.w3(32'hbc82c187),
	.w4(32'hbc0dd16a),
	.w5(32'hbc10bfc5),
	.w6(32'hbbc12b9b),
	.w7(32'hbc230cf1),
	.w8(32'hbbefcd63),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64cee9),
	.w1(32'h3b6fec5b),
	.w2(32'h3bb0e8be),
	.w3(32'hbc0cfd48),
	.w4(32'h3bb64c73),
	.w5(32'hba45fe7d),
	.w6(32'h3b124e87),
	.w7(32'h3b8febdd),
	.w8(32'h3b1db52f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f1db1),
	.w1(32'hba8d89eb),
	.w2(32'hbb163153),
	.w3(32'hbbc6abc8),
	.w4(32'hbb9bd905),
	.w5(32'h3b1a56e5),
	.w6(32'h3ac54cfe),
	.w7(32'h3c008a98),
	.w8(32'h3bb028f6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8685de),
	.w1(32'h3bbb9ac6),
	.w2(32'h3c858035),
	.w3(32'hba862614),
	.w4(32'hbb02b7f3),
	.w5(32'hbbaf1887),
	.w6(32'hbc8a68e9),
	.w7(32'hbba095cb),
	.w8(32'hbc2c47e3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14ade3),
	.w1(32'h3d38ca23),
	.w2(32'h3daa6743),
	.w3(32'hbc9f93c9),
	.w4(32'h3bf21089),
	.w5(32'h3d4aca5b),
	.w6(32'hbd3aeaaa),
	.w7(32'hbbd8f8bb),
	.w8(32'h3d00332d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c970485),
	.w1(32'h3be1282a),
	.w2(32'h3c6ca0a8),
	.w3(32'hbc96d39d),
	.w4(32'hbcaee78b),
	.w5(32'hbc9df427),
	.w6(32'hbc056e24),
	.w7(32'hbc16486b),
	.w8(32'hbaaa502c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b40e9),
	.w1(32'h3cafc0a0),
	.w2(32'h3d637ef3),
	.w3(32'hbc58364c),
	.w4(32'hbd0519e1),
	.w5(32'hbd081062),
	.w6(32'h3c8033e7),
	.w7(32'h3bcb155e),
	.w8(32'hbb34d73d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc66396),
	.w1(32'h3a9be800),
	.w2(32'h3a7585e9),
	.w3(32'hbc0dc77b),
	.w4(32'hba5e52e6),
	.w5(32'hbbf3e7c1),
	.w6(32'h3b81c56c),
	.w7(32'hb91c9461),
	.w8(32'h3bf7e269),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4f4b83),
	.w1(32'hbc476e5d),
	.w2(32'h3d20c206),
	.w3(32'hbd1893d5),
	.w4(32'hbd03dcfb),
	.w5(32'h3ca056a1),
	.w6(32'hbd11563b),
	.w7(32'hbb650d68),
	.w8(32'h3ccf698c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a6630),
	.w1(32'h3cbdeb24),
	.w2(32'h3c2b5161),
	.w3(32'h3c3783e2),
	.w4(32'hb9912d27),
	.w5(32'hbbc70b10),
	.w6(32'h3c383e8b),
	.w7(32'h3bfa7c45),
	.w8(32'h3a1e2ea7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948a882),
	.w1(32'hbc694b8f),
	.w2(32'hbc9398ad),
	.w3(32'h3a29c8d7),
	.w4(32'hbbe64b72),
	.w5(32'hbbd46bb3),
	.w6(32'h3aace54a),
	.w7(32'hbb247642),
	.w8(32'hb8e8fdc9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1d929),
	.w1(32'hbb5012bb),
	.w2(32'h3ae5377c),
	.w3(32'hbc826fd2),
	.w4(32'hbb16cd29),
	.w5(32'h3c654715),
	.w6(32'hbb24a869),
	.w7(32'h3c4d8942),
	.w8(32'h38aa959c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f98a),
	.w1(32'hbc58e0ba),
	.w2(32'hbc67489e),
	.w3(32'h3bc9e3c8),
	.w4(32'hbb09d172),
	.w5(32'h3aef124b),
	.w6(32'h3a396f30),
	.w7(32'h3c3759a1),
	.w8(32'h3bb54abd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdca33fa),
	.w1(32'h3c31ec98),
	.w2(32'h3df8ce84),
	.w3(32'hbb4df578),
	.w4(32'h3c092cf3),
	.w5(32'h3d1ecdd7),
	.w6(32'hbcce7f0d),
	.w7(32'hbbd7d75a),
	.w8(32'h3d37f792),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18b25f),
	.w1(32'h3c2e0d32),
	.w2(32'h3c9611fb),
	.w3(32'hbcce7bbd),
	.w4(32'h3ba36e52),
	.w5(32'h3c85d798),
	.w6(32'hbc6a532a),
	.w7(32'hbc8dfe94),
	.w8(32'hbc445dca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba132e60),
	.w1(32'hbbc1484a),
	.w2(32'hbb673004),
	.w3(32'hba6ffe5d),
	.w4(32'hbba1b9b0),
	.w5(32'hbbf2185b),
	.w6(32'hbb33797f),
	.w7(32'hbb78cea1),
	.w8(32'h3bbeae64),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add8749),
	.w1(32'h3b36b074),
	.w2(32'h3c177077),
	.w3(32'h3b2bc464),
	.w4(32'h3c8e1c32),
	.w5(32'h3cd38aab),
	.w6(32'hbc8b6e3f),
	.w7(32'hbce77823),
	.w8(32'hbc86836a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac49f2d),
	.w1(32'hbc70ab52),
	.w2(32'hbccaf886),
	.w3(32'h3c959059),
	.w4(32'h3b0ab6e6),
	.w5(32'hbbcf9535),
	.w6(32'h3c22fce7),
	.w7(32'h3c35f427),
	.w8(32'h3b05e9fb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ca4a5),
	.w1(32'h3c010bab),
	.w2(32'h3aacc93f),
	.w3(32'hba93e34c),
	.w4(32'hbc35d0c8),
	.w5(32'hbc8c2815),
	.w6(32'hbc3d303c),
	.w7(32'hbb171792),
	.w8(32'hb7ae4eea),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2387f9),
	.w1(32'h3c491da8),
	.w2(32'h3bc4e3d1),
	.w3(32'hbc8b4567),
	.w4(32'h3be11b60),
	.w5(32'h3986317d),
	.w6(32'hb9258c02),
	.w7(32'h3bf3285d),
	.w8(32'h3b9f87ce),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc717),
	.w1(32'hbc6e11c7),
	.w2(32'hbc693612),
	.w3(32'h3b0c9627),
	.w4(32'hbc417a1d),
	.w5(32'hbc968566),
	.w6(32'h3c1680b7),
	.w7(32'hbafb5fd6),
	.w8(32'hbbba4399),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7821bd),
	.w1(32'h3af2728b),
	.w2(32'h3cce4faf),
	.w3(32'hbb4fdbbd),
	.w4(32'h3c2710fb),
	.w5(32'h3cdf8f2b),
	.w6(32'h3a980b48),
	.w7(32'h3ba47ff5),
	.w8(32'h3c5988fe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05180),
	.w1(32'hbb30691d),
	.w2(32'hbb18688e),
	.w3(32'h3b4abb3a),
	.w4(32'hbb0aa66e),
	.w5(32'hba560e26),
	.w6(32'h3a3a4ef5),
	.w7(32'h3aeee9d4),
	.w8(32'h3ac12b05),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e874),
	.w1(32'h3b8666a8),
	.w2(32'h3a8f347b),
	.w3(32'h3b7dfd3d),
	.w4(32'h3b21ee19),
	.w5(32'hbaacc65b),
	.w6(32'hbafddb06),
	.w7(32'hbbff5c40),
	.w8(32'hbbfa20bb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6d617),
	.w1(32'h3b3ebec6),
	.w2(32'h3c006215),
	.w3(32'hba1eec43),
	.w4(32'h3b2d3560),
	.w5(32'h3b00a8ae),
	.w6(32'hbb653863),
	.w7(32'hb99c095e),
	.w8(32'hbaa9426a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66e85),
	.w1(32'h3c004a8c),
	.w2(32'h3b933335),
	.w3(32'h3c277d92),
	.w4(32'h39da5487),
	.w5(32'hb95212f2),
	.w6(32'h3a3eb950),
	.w7(32'h3b5a8b94),
	.w8(32'h3a6a8693),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c632b97),
	.w1(32'h3b6e095e),
	.w2(32'h3c30615b),
	.w3(32'hbc41de1f),
	.w4(32'hbcb4bab9),
	.w5(32'hbc9e0fcb),
	.w6(32'hbd134ed3),
	.w7(32'hbd319d62),
	.w8(32'hbcddc50c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14c122),
	.w1(32'h3c65aa32),
	.w2(32'h3c7c5c44),
	.w3(32'h3aa96965),
	.w4(32'h397d8c8a),
	.w5(32'h3bc4315f),
	.w6(32'h3bf1e69c),
	.w7(32'h3b92bcb6),
	.w8(32'h3bb71ca8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cad1),
	.w1(32'hba48bab8),
	.w2(32'h3b1a0166),
	.w3(32'h3b871651),
	.w4(32'hbbce6c0f),
	.w5(32'hbb9345ad),
	.w6(32'h3ad483e4),
	.w7(32'h3c0ada01),
	.w8(32'h39248b29),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fa56e),
	.w1(32'h3c14fbae),
	.w2(32'h3c1226c2),
	.w3(32'hbc38b2f3),
	.w4(32'hbc1af161),
	.w5(32'h3a30062d),
	.w6(32'hbc6cfc2d),
	.w7(32'hbbb171be),
	.w8(32'h3c04b4da),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a54bf),
	.w1(32'h3c59cb7e),
	.w2(32'h3cd612e7),
	.w3(32'hbc006b78),
	.w4(32'h3a8e25ca),
	.w5(32'h3c811855),
	.w6(32'hbc613057),
	.w7(32'hbc16e2fa),
	.w8(32'h3c26d12b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c9750),
	.w1(32'h3c395cf4),
	.w2(32'h3ccdc6de),
	.w3(32'h3af78ea9),
	.w4(32'h3bfbda59),
	.w5(32'h3c8a9f31),
	.w6(32'h3ae7617c),
	.w7(32'h3bd98a26),
	.w8(32'h3c94bddd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd959a1),
	.w1(32'h3bd24451),
	.w2(32'h3ce1a242),
	.w3(32'hbaa937b0),
	.w4(32'hbc5a9ab3),
	.w5(32'hbc0d0247),
	.w6(32'hbaf30afa),
	.w7(32'h3b593907),
	.w8(32'h3ace7083),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf88649),
	.w1(32'h3b7ec042),
	.w2(32'h3ce936f7),
	.w3(32'hbc266eac),
	.w4(32'h3ac1c6ee),
	.w5(32'h3c92a67d),
	.w6(32'hbb528529),
	.w7(32'h3b97b82a),
	.w8(32'h3c0fb46a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c76ac),
	.w1(32'h3b19c841),
	.w2(32'h3c94ef85),
	.w3(32'hbb1e8c96),
	.w4(32'hbad4a835),
	.w5(32'hbc18cea3),
	.w6(32'h3b4ff150),
	.w7(32'hbbb9f330),
	.w8(32'hbba4bef9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5bf14),
	.w1(32'h3992abd1),
	.w2(32'h3cccab98),
	.w3(32'hbc2437f6),
	.w4(32'hbca7315c),
	.w5(32'hbc86e30a),
	.w6(32'h3aa79686),
	.w7(32'h3b2ba644),
	.w8(32'h3b0f98cb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a305e),
	.w1(32'h3be359bb),
	.w2(32'h3a5e9610),
	.w3(32'h3a37188b),
	.w4(32'h3bf60aa0),
	.w5(32'hbc3d7e90),
	.w6(32'h3c8de02d),
	.w7(32'hba8d3555),
	.w8(32'hbc8c9cb0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac709c),
	.w1(32'h3cf90715),
	.w2(32'h3d37f32f),
	.w3(32'hbc2b5b54),
	.w4(32'h3c07c072),
	.w5(32'h3cf7c4cc),
	.w6(32'hbd08ab3c),
	.w7(32'hbc5b4d91),
	.w8(32'h3ce58769),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c192347),
	.w1(32'h3adb1cdc),
	.w2(32'hbb1a557c),
	.w3(32'hbc0277ea),
	.w4(32'h3b01d844),
	.w5(32'h3ae602b9),
	.w6(32'hbc09f11c),
	.w7(32'hbc20e839),
	.w8(32'hbaa2bccb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22dc29),
	.w1(32'h3ba24181),
	.w2(32'h3ca89ce2),
	.w3(32'h3a0091ed),
	.w4(32'hbc18caf8),
	.w5(32'h3af87de1),
	.w6(32'hbc0ca746),
	.w7(32'h3b37d14f),
	.w8(32'h3be9a7f9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6d35),
	.w1(32'hbb8c527c),
	.w2(32'h3c4caeb9),
	.w3(32'h3a9d697a),
	.w4(32'hbc3ef964),
	.w5(32'hbc9cc64c),
	.w6(32'h3c192e14),
	.w7(32'h3c8e2cc8),
	.w8(32'h3bbc56e6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62cc86),
	.w1(32'h3c4fac8e),
	.w2(32'h3d879443),
	.w3(32'hbad6cc4d),
	.w4(32'h3c2a1c55),
	.w5(32'h3d1082e8),
	.w6(32'hbc095701),
	.w7(32'h3c595062),
	.w8(32'h3d075ade),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c112885),
	.w1(32'h3abcfbfa),
	.w2(32'h3c5d8674),
	.w3(32'h3af11729),
	.w4(32'hbb37d89e),
	.w5(32'hba8bd2d2),
	.w6(32'hb9f48667),
	.w7(32'h3b0391ab),
	.w8(32'h3bf22802),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff9058),
	.w1(32'h3ca13d1d),
	.w2(32'h3cb24b7f),
	.w3(32'h3b2868f9),
	.w4(32'h3c2db635),
	.w5(32'h3ca5842e),
	.w6(32'h3bc17379),
	.w7(32'h3bcda5f8),
	.w8(32'h3c5dd11e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e1435),
	.w1(32'hbaee6309),
	.w2(32'h3ba39a67),
	.w3(32'hbb355ff5),
	.w4(32'hbb57c874),
	.w5(32'h3c07e600),
	.w6(32'hbb97f0e7),
	.w7(32'hbbaeaa1f),
	.w8(32'h3b03e582),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e9baa),
	.w1(32'h3b577e4c),
	.w2(32'h3bb84c8f),
	.w3(32'hbc31364d),
	.w4(32'hbc30090b),
	.w5(32'hbbbfde36),
	.w6(32'h3b86a030),
	.w7(32'hbc15f559),
	.w8(32'hbb98931c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6433),
	.w1(32'h3b91f375),
	.w2(32'h3b00e236),
	.w3(32'hbbc2da38),
	.w4(32'hbc27135d),
	.w5(32'hbc22e97f),
	.w6(32'h3c02df7c),
	.w7(32'h3c0e48fa),
	.w8(32'h3c2d395d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a8b6),
	.w1(32'h3a256bab),
	.w2(32'hba683f81),
	.w3(32'hbc1b6b07),
	.w4(32'hba554d42),
	.w5(32'h39d0593c),
	.w6(32'hbc3af564),
	.w7(32'hbc242bc7),
	.w8(32'hbbaf2bb1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27865c),
	.w1(32'h3c8cb5bf),
	.w2(32'h3c8f76d6),
	.w3(32'h3b4b0301),
	.w4(32'h3cf4b424),
	.w5(32'h3d07a07f),
	.w6(32'hbc5f8925),
	.w7(32'hbcaebf7f),
	.w8(32'hbb35bacb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a240b),
	.w1(32'hbc1d596f),
	.w2(32'hbc2e1dce),
	.w3(32'h3c9e06f7),
	.w4(32'hbbc67864),
	.w5(32'hbc1589eb),
	.w6(32'hbbfccf71),
	.w7(32'hbbdeadb9),
	.w8(32'hbb18e3f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cf741),
	.w1(32'hbb764436),
	.w2(32'hbbf0ef92),
	.w3(32'hbc3923ae),
	.w4(32'h3b7a7acb),
	.w5(32'h3ba0c987),
	.w6(32'hbb9b5051),
	.w7(32'hbc18c514),
	.w8(32'hbc126f43),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e494e),
	.w1(32'h3c2cc25b),
	.w2(32'h3c4ae8af),
	.w3(32'h3b8aada8),
	.w4(32'h3b68f6e7),
	.w5(32'h3c28e274),
	.w6(32'h3b82402d),
	.w7(32'hbb4305f9),
	.w8(32'h3b2ad5c8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26417e),
	.w1(32'hbb2c848f),
	.w2(32'h389d2397),
	.w3(32'h3b54263d),
	.w4(32'h3c845d43),
	.w5(32'h3c16a3b5),
	.w6(32'hbcba9331),
	.w7(32'hbcb490cd),
	.w8(32'hbc53a39e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cb7db),
	.w1(32'h3c132803),
	.w2(32'h3d705a7d),
	.w3(32'h3c750599),
	.w4(32'hbcc6871c),
	.w5(32'hbcf2e6be),
	.w6(32'hbc134c50),
	.w7(32'h3c3322b0),
	.w8(32'h3b9593c8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4a65a),
	.w1(32'hba6abbbf),
	.w2(32'h3c2955f4),
	.w3(32'hbca74d74),
	.w4(32'hbb709300),
	.w5(32'hbc135a3e),
	.w6(32'h3aa04054),
	.w7(32'h3908a5e2),
	.w8(32'h3ba73770),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc920492),
	.w1(32'hbc23860d),
	.w2(32'h3c51a368),
	.w3(32'hbc464357),
	.w4(32'hbbf7e34e),
	.w5(32'h3c6662b2),
	.w6(32'hbc9670a7),
	.w7(32'hbc579f02),
	.w8(32'h3c2f3ea5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d01ce),
	.w1(32'h3bdde1d5),
	.w2(32'h3b44b247),
	.w3(32'hbbe0f7fb),
	.w4(32'hba342c31),
	.w5(32'hbbdee73e),
	.w6(32'hbb5a1210),
	.w7(32'hbbf3a2af),
	.w8(32'hbbfca79a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac361),
	.w1(32'h3b1f3495),
	.w2(32'h3c5d4dde),
	.w3(32'hbcb18dec),
	.w4(32'hbc4ee3e7),
	.w5(32'hbbac956c),
	.w6(32'h3a0406af),
	.w7(32'hbb9104e0),
	.w8(32'hbb604822),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba99e44),
	.w1(32'h3be39d63),
	.w2(32'h3c136e08),
	.w3(32'hbb509f03),
	.w4(32'h3b43e12a),
	.w5(32'hbb07a821),
	.w6(32'hbb8ff14e),
	.w7(32'hba14621c),
	.w8(32'h39758be7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e9ec9),
	.w1(32'h3c786824),
	.w2(32'h3d2ad20d),
	.w3(32'h3c40cdd5),
	.w4(32'h3c39f36b),
	.w5(32'h3be92f80),
	.w6(32'hbba98e32),
	.w7(32'h3b82c2ef),
	.w8(32'hb7bb19c2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f17a),
	.w1(32'h3b024000),
	.w2(32'hba86a58e),
	.w3(32'h3b933f2d),
	.w4(32'hba4205fa),
	.w5(32'hbba157b7),
	.w6(32'h3bad0694),
	.w7(32'h3bae4688),
	.w8(32'h3b01004e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a465229),
	.w1(32'h3c574569),
	.w2(32'h3c708be5),
	.w3(32'hbbeb86c1),
	.w4(32'hbbe410ea),
	.w5(32'hbbc7d4a9),
	.w6(32'h3b1d104a),
	.w7(32'h3c08b10f),
	.w8(32'h3c84248e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaac52),
	.w1(32'h3b99901d),
	.w2(32'h3c648e3c),
	.w3(32'hbc2a3d18),
	.w4(32'hbbcced5b),
	.w5(32'hbbd94743),
	.w6(32'h3a908d66),
	.w7(32'h3c04b049),
	.w8(32'hbb93c93d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ee6b),
	.w1(32'h3b115151),
	.w2(32'h3cc5f12e),
	.w3(32'hbc8a985c),
	.w4(32'hbc9f1642),
	.w5(32'hba4b95e7),
	.w6(32'hbcc3654d),
	.w7(32'hbc18f0c5),
	.w8(32'hbbf1d5dc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40b7d8),
	.w1(32'h3c82c308),
	.w2(32'h3d487ba2),
	.w3(32'hbb866e9c),
	.w4(32'h3c50cf94),
	.w5(32'h3cab5420),
	.w6(32'hbc1f41bb),
	.w7(32'h3b9df10d),
	.w8(32'h3c71019a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ab145),
	.w1(32'h3c1be210),
	.w2(32'h3c55f191),
	.w3(32'hbbae05bd),
	.w4(32'hbb2288b1),
	.w5(32'hbc217761),
	.w6(32'hb94c64a7),
	.w7(32'h3aa5e9fc),
	.w8(32'hbb595406),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa160d),
	.w1(32'h3c860528),
	.w2(32'h3cece4b2),
	.w3(32'h3b754ae6),
	.w4(32'hbbac2d5f),
	.w5(32'hbc410b5c),
	.w6(32'h3b89924a),
	.w7(32'h3bf9ce1f),
	.w8(32'h3b820624),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf2c569),
	.w1(32'h3bff7586),
	.w2(32'h3bde7a88),
	.w3(32'hbcb36999),
	.w4(32'hbc6ecc10),
	.w5(32'hbc21c0c6),
	.w6(32'h3b59904c),
	.w7(32'h3c29bd94),
	.w8(32'h3c042265),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a6ea),
	.w1(32'h3c3b8a22),
	.w2(32'h3d0103b6),
	.w3(32'hbc9712e1),
	.w4(32'hbcd6ec52),
	.w5(32'hbc441248),
	.w6(32'hbca6e868),
	.w7(32'hbc6a1aec),
	.w8(32'hba3c7a2c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30aa13),
	.w1(32'h3d20ddb8),
	.w2(32'h3d0dbbd2),
	.w3(32'h3b663fb1),
	.w4(32'h3a2e216f),
	.w5(32'hbb79bc85),
	.w6(32'hbc99cf8a),
	.w7(32'hbd26e57f),
	.w8(32'hbd2efc05),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf6eca),
	.w1(32'h3cb59af6),
	.w2(32'h3d49aa68),
	.w3(32'hbc71ae36),
	.w4(32'hbc30a29d),
	.w5(32'h3c6f1960),
	.w6(32'hbcf9e9e1),
	.w7(32'hbcc4e011),
	.w8(32'hbb92cac0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb70b19),
	.w1(32'h3cec4ce4),
	.w2(32'h3cdbd707),
	.w3(32'hbc52f581),
	.w4(32'h3c46f450),
	.w5(32'h3d0ca6aa),
	.w6(32'hbc7cec45),
	.w7(32'hbc8ba1a5),
	.w8(32'hbc32f540),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc971f),
	.w1(32'h3b805194),
	.w2(32'h3b89a697),
	.w3(32'h3b6f3211),
	.w4(32'hbb145f2e),
	.w5(32'hbb405b61),
	.w6(32'h3ab5170e),
	.w7(32'h3a2b9607),
	.w8(32'h3ad5b5be),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad8649),
	.w1(32'hbc964dec),
	.w2(32'hbce8839d),
	.w3(32'hbbc29d56),
	.w4(32'hbaf15b95),
	.w5(32'hbbfbfddf),
	.w6(32'h3c67f308),
	.w7(32'h3c90fd12),
	.w8(32'h3c006cd0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb16b64),
	.w1(32'hbb57bcff),
	.w2(32'hbad2793b),
	.w3(32'hbb7462ea),
	.w4(32'hbb531235),
	.w5(32'h3a8192a1),
	.w6(32'hbc17d269),
	.w7(32'hbc32e33b),
	.w8(32'hbbc35656),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1fa8),
	.w1(32'h3c052a2b),
	.w2(32'h3c9560b5),
	.w3(32'hbb4737f0),
	.w4(32'hbb95519a),
	.w5(32'hb8e0273f),
	.w6(32'h3b0a6857),
	.w7(32'h3b71d997),
	.w8(32'h3b343615),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd44947),
	.w1(32'h3c2a3056),
	.w2(32'h3c76c312),
	.w3(32'hb9ed47b5),
	.w4(32'h3b9b1633),
	.w5(32'hbad0c7ca),
	.w6(32'h3b180486),
	.w7(32'h3b6bc462),
	.w8(32'h3bd1672d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71674),
	.w1(32'h3b52f95e),
	.w2(32'h3b0fe093),
	.w3(32'hba9e461f),
	.w4(32'hbab5e8f5),
	.w5(32'h39ae9eff),
	.w6(32'h3a7f17e9),
	.w7(32'h3b81af29),
	.w8(32'h3c17404b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56536e),
	.w1(32'hbaa84c64),
	.w2(32'hbc608445),
	.w3(32'hbb583af6),
	.w4(32'hbbf174c5),
	.w5(32'hbc8ebecd),
	.w6(32'h3ac076d1),
	.w7(32'h39c19dda),
	.w8(32'hbafdede3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f71d84),
	.w1(32'h3b7c6294),
	.w2(32'h3c353985),
	.w3(32'hbc2535d4),
	.w4(32'hbb5cdf4e),
	.w5(32'h3b803c6e),
	.w6(32'hbc0a0685),
	.w7(32'hbb8ae6c4),
	.w8(32'h3b438a62),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab410b9),
	.w1(32'h3bea6a69),
	.w2(32'h3ce7e95c),
	.w3(32'h39fa5f1d),
	.w4(32'hbc5413ab),
	.w5(32'hbd2de636),
	.w6(32'h3b778423),
	.w7(32'h3c498ee7),
	.w8(32'h3a49359d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9806c2),
	.w1(32'h3c304141),
	.w2(32'h3cb688de),
	.w3(32'hbd08d3d2),
	.w4(32'h3bbb12fe),
	.w5(32'h3c887976),
	.w6(32'hbba93865),
	.w7(32'h3b19ee2a),
	.w8(32'h3c26057c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8269ed),
	.w1(32'h3c5043fc),
	.w2(32'h3ca50576),
	.w3(32'hbc055698),
	.w4(32'hbc7c9a3e),
	.w5(32'hbba79f33),
	.w6(32'hbc5df73b),
	.w7(32'hbc949633),
	.w8(32'h3b83ff82),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c07f3),
	.w1(32'h3badc3ce),
	.w2(32'h3c660b0c),
	.w3(32'hbc8c6156),
	.w4(32'h37d52d01),
	.w5(32'h3b9d0851),
	.w6(32'h3b9eaea5),
	.w7(32'h3c5ddedd),
	.w8(32'h3b91691d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bfac1),
	.w1(32'h3bd1f255),
	.w2(32'h3c974a8e),
	.w3(32'h3c0d74c2),
	.w4(32'h38538fa5),
	.w5(32'h3b0f9194),
	.w6(32'h3af15a9b),
	.w7(32'hba13c84c),
	.w8(32'h3b82dc90),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0e87b),
	.w1(32'h3b9dab52),
	.w2(32'hbb812589),
	.w3(32'h3c14571f),
	.w4(32'hba8eff81),
	.w5(32'h3b8f9ee6),
	.w6(32'hbafc5a14),
	.w7(32'hbb78996e),
	.w8(32'h3be061ac),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c4a4e),
	.w1(32'h3ca1e7f3),
	.w2(32'h3cb291ef),
	.w3(32'h3b34ded5),
	.w4(32'h3bc35147),
	.w5(32'h3b3e9166),
	.w6(32'hbc31510e),
	.w7(32'hbc122907),
	.w8(32'hbc193f53),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a4261),
	.w1(32'hbb28ce5e),
	.w2(32'hbc705083),
	.w3(32'h3b875986),
	.w4(32'h3ca2c83d),
	.w5(32'h3c801d4d),
	.w6(32'h3aa21a96),
	.w7(32'hbada7e68),
	.w8(32'h3b06a1fb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6dcf7),
	.w1(32'hbb844d8c),
	.w2(32'hbbb1eb5e),
	.w3(32'h3c44e3eb),
	.w4(32'hbb8c6b30),
	.w5(32'hbbf2339f),
	.w6(32'h396abcd1),
	.w7(32'h3aca753e),
	.w8(32'h3b0d2f5c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe7b3),
	.w1(32'h3c9b5b53),
	.w2(32'hba6b4843),
	.w3(32'hbc2513eb),
	.w4(32'hbc8333a3),
	.w5(32'hbceca2c5),
	.w6(32'h3c807539),
	.w7(32'h3c84d718),
	.w8(32'h3c74e5fa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c8db4),
	.w1(32'h3b80cd19),
	.w2(32'hba9c6d0d),
	.w3(32'hbc6fa3e7),
	.w4(32'hbc25fa9f),
	.w5(32'hbc3ee49c),
	.w6(32'h3b86ed85),
	.w7(32'hba9b0425),
	.w8(32'h3b0d701f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847030),
	.w1(32'h3c14d570),
	.w2(32'h3cb709ca),
	.w3(32'hbc046e9f),
	.w4(32'hbb1705f9),
	.w5(32'h3c3ecc24),
	.w6(32'hbc16c0e4),
	.w7(32'hbba52b53),
	.w8(32'h3c22b736),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5653a3),
	.w1(32'hbb87d89e),
	.w2(32'h3a5fdaad),
	.w3(32'hbafd01ad),
	.w4(32'hbb1641ee),
	.w5(32'hbb430210),
	.w6(32'hbc63a270),
	.w7(32'hbc4714f6),
	.w8(32'hbbaf997b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a003807),
	.w1(32'hbc4191f9),
	.w2(32'hbc0c85da),
	.w3(32'hbb6d41f8),
	.w4(32'hbc80c175),
	.w5(32'hbc6bd06a),
	.w6(32'h3c0954f4),
	.w7(32'h3b8b6bb6),
	.w8(32'hba82a834),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a0af),
	.w1(32'hbb771fd8),
	.w2(32'hbc707567),
	.w3(32'hbba7531b),
	.w4(32'h3bf65c7a),
	.w5(32'h3bc71c37),
	.w6(32'h3c7566fe),
	.w7(32'h3c1ba663),
	.w8(32'h3c140e23),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843383),
	.w1(32'h3b9aa098),
	.w2(32'hbb968c8b),
	.w3(32'h3c1e72f7),
	.w4(32'h3c204bd0),
	.w5(32'h3c1b77dd),
	.w6(32'h3b2d1ad9),
	.w7(32'h3af9104b),
	.w8(32'h3a9d13e2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b9a7),
	.w1(32'hbb9610b3),
	.w2(32'hbaa00f65),
	.w3(32'h3c461eb9),
	.w4(32'hbb351c34),
	.w5(32'hbac7a696),
	.w6(32'hba2d183b),
	.w7(32'h39471818),
	.w8(32'h3b8ab807),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d1520),
	.w1(32'h3b50c5da),
	.w2(32'h3b8c9f1b),
	.w3(32'hbb068e43),
	.w4(32'h38375622),
	.w5(32'h3a2bf020),
	.w6(32'h3b964949),
	.w7(32'hbb069794),
	.w8(32'h3ade7e78),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384da013),
	.w1(32'hba712f0b),
	.w2(32'hbbcac424),
	.w3(32'h3b10f134),
	.w4(32'h3c1cf74f),
	.w5(32'hbb83b771),
	.w6(32'h3ca0dd9b),
	.w7(32'h3c6aabf6),
	.w8(32'h3c261ffa),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81cde8),
	.w1(32'hbc851178),
	.w2(32'hbcb12001),
	.w3(32'h3bf66fa0),
	.w4(32'hbb6706dc),
	.w5(32'h3c207b73),
	.w6(32'hbc8b0302),
	.w7(32'hbc3a350a),
	.w8(32'hbc9019d2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca669e8),
	.w1(32'h3ac7a449),
	.w2(32'h3b844143),
	.w3(32'h3c0e4cdf),
	.w4(32'h3b86fc1d),
	.w5(32'h3c21193c),
	.w6(32'hbc543e51),
	.w7(32'hbc913e62),
	.w8(32'hbbf6af95),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b4aa3),
	.w1(32'hb8677286),
	.w2(32'hbbc926e6),
	.w3(32'h3bb8b327),
	.w4(32'h3bcf103c),
	.w5(32'h3bd57902),
	.w6(32'h39c62a02),
	.w7(32'hbb53239c),
	.w8(32'hbb4b7f2a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d627f),
	.w1(32'hbbcee5ec),
	.w2(32'hbc23c168),
	.w3(32'h3bf37b9b),
	.w4(32'h3b243736),
	.w5(32'h3b27637a),
	.w6(32'h3b84c04f),
	.w7(32'hbb214ec2),
	.w8(32'h3c01bdac),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c317b),
	.w1(32'hbba65bab),
	.w2(32'h3c178196),
	.w3(32'hba3dbd14),
	.w4(32'h3aeda777),
	.w5(32'h3c05cece),
	.w6(32'hbc1404cf),
	.w7(32'hbbcee07e),
	.w8(32'h3aa4c153),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7c6f),
	.w1(32'hbb3d10a7),
	.w2(32'hbae09ae9),
	.w3(32'h3b944e4f),
	.w4(32'h3ba89f3c),
	.w5(32'hba60af4e),
	.w6(32'hbc1c4ba4),
	.w7(32'hbc507ff7),
	.w8(32'hbc543dca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a565d),
	.w1(32'h3b2a2fb2),
	.w2(32'h3b677e56),
	.w3(32'hbbc6206a),
	.w4(32'hbb75a375),
	.w5(32'hbba1da3d),
	.w6(32'h3ba40027),
	.w7(32'h3b9d6f56),
	.w8(32'h3a8cff3f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54a78c),
	.w1(32'h3c4bfddc),
	.w2(32'h3c3d944a),
	.w3(32'hbc32f1f7),
	.w4(32'h3b9ca446),
	.w5(32'h37ae927e),
	.w6(32'h3abc328c),
	.w7(32'h3b595259),
	.w8(32'h3c283950),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4556ae),
	.w1(32'h3c3ecdda),
	.w2(32'h39c46d35),
	.w3(32'hb9190e55),
	.w4(32'hbb80adba),
	.w5(32'hbc379ab8),
	.w6(32'hbb83a423),
	.w7(32'hbac654a4),
	.w8(32'h3be8b30d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39902459),
	.w1(32'hbc217113),
	.w2(32'hbc5c328e),
	.w3(32'hbba0efe2),
	.w4(32'hbbe54b18),
	.w5(32'hbc3adddd),
	.w6(32'hbb082e87),
	.w7(32'hbb7bbf8e),
	.w8(32'hbb118f01),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7e62),
	.w1(32'h39a5493b),
	.w2(32'h3baa2b5e),
	.w3(32'hbbab83e0),
	.w4(32'h3c0e8198),
	.w5(32'h3c149d2a),
	.w6(32'h3c3852af),
	.w7(32'h3a71e097),
	.w8(32'hbb3d6a22),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccac31),
	.w1(32'hbb0b40a6),
	.w2(32'hbc30a508),
	.w3(32'h3b81f8dc),
	.w4(32'hbb084851),
	.w5(32'h3b693618),
	.w6(32'hbae33b49),
	.w7(32'hb8588555),
	.w8(32'hbbc9fd6f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e3051),
	.w1(32'h3b34c180),
	.w2(32'h3afe0206),
	.w3(32'h3c189189),
	.w4(32'hbb2a5590),
	.w5(32'hbb97227b),
	.w6(32'h3aa56805),
	.w7(32'hbb2294af),
	.w8(32'hbb83b58f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbabe74),
	.w1(32'h3a1c0f10),
	.w2(32'h3bf76605),
	.w3(32'h3b373a5d),
	.w4(32'hba89fa6c),
	.w5(32'h3aff3e66),
	.w6(32'h398bd836),
	.w7(32'h3a5289e5),
	.w8(32'h3a49759b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd5b86),
	.w1(32'hbb8e6529),
	.w2(32'h3bbd206a),
	.w3(32'hbb5ad09f),
	.w4(32'hbb0eae82),
	.w5(32'h3c137f02),
	.w6(32'hba126eb1),
	.w7(32'h3b34fb2a),
	.w8(32'h3c48dcbd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule