module layer_10_featuremap_511(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e7778),
	.w1(32'hbbe19ce7),
	.w2(32'h3b5b52a4),
	.w3(32'hbc21388a),
	.w4(32'hbb8b1cc7),
	.w5(32'hbba4942c),
	.w6(32'h3a808c3d),
	.w7(32'hbba0210b),
	.w8(32'hba325a86),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b98db),
	.w1(32'h3b98e73b),
	.w2(32'hbc292f34),
	.w3(32'hbc7ce13c),
	.w4(32'hbba76947),
	.w5(32'h3ad5ae65),
	.w6(32'hbbc42ff6),
	.w7(32'hbc2ba443),
	.w8(32'hbb665edb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac9fb8),
	.w1(32'hbb8a870d),
	.w2(32'h3b158901),
	.w3(32'h3c578f34),
	.w4(32'hbc5845eb),
	.w5(32'h3c99e54f),
	.w6(32'hba844f5c),
	.w7(32'hbbfeb2f0),
	.w8(32'hbb6832c0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49c7eb),
	.w1(32'hba2e0ec8),
	.w2(32'hbc3c1399),
	.w3(32'h3c6f1692),
	.w4(32'hbaf97a56),
	.w5(32'hbb05b980),
	.w6(32'hbca186c8),
	.w7(32'hbbe5bae6),
	.w8(32'h3cbd1c48),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836ba31),
	.w1(32'hbc2d6b44),
	.w2(32'hb935737a),
	.w3(32'hbc1fb7ef),
	.w4(32'hbbdf2380),
	.w5(32'hbad74d5b),
	.w6(32'hbb97c80a),
	.w7(32'hbc0c3a92),
	.w8(32'hbb412666),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbef7ed),
	.w1(32'hbc33fc90),
	.w2(32'hbc154391),
	.w3(32'hbc0f2dd9),
	.w4(32'hbb55a149),
	.w5(32'hbba1a08a),
	.w6(32'h3a122f3e),
	.w7(32'hbb12fa71),
	.w8(32'h3a9cec91),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae967d5),
	.w1(32'h3b963748),
	.w2(32'hbb57a4d0),
	.w3(32'hbc84010e),
	.w4(32'hbc066562),
	.w5(32'hbbf68c76),
	.w6(32'hbb9b8ece),
	.w7(32'hbc92480f),
	.w8(32'hbbb5b410),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce827b2),
	.w1(32'hbc262e72),
	.w2(32'hbc1c123e),
	.w3(32'hbc1598ba),
	.w4(32'h3bbc25fe),
	.w5(32'hb9eaa55d),
	.w6(32'h3cb7616c),
	.w7(32'hbc5cc141),
	.w8(32'h3ac16cba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b49a),
	.w1(32'h3beeb4dc),
	.w2(32'h3c030d6d),
	.w3(32'h3d111836),
	.w4(32'hbca18796),
	.w5(32'h3c6fdac1),
	.w6(32'hbb80dd87),
	.w7(32'h3b936419),
	.w8(32'hbc18ea57),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aae2fd),
	.w1(32'hbbb4c7a5),
	.w2(32'h3cc88e2b),
	.w3(32'hbc32d649),
	.w4(32'hba9de5ba),
	.w5(32'h3aa230a1),
	.w6(32'hbc2cac6c),
	.w7(32'hbc008cc8),
	.w8(32'h3c01ca77),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca560bb),
	.w1(32'hbbeb404d),
	.w2(32'h3c01383c),
	.w3(32'hbc875a26),
	.w4(32'hbbc5629e),
	.w5(32'hbbdb91ce),
	.w6(32'hbb3def28),
	.w7(32'h3c22b91a),
	.w8(32'hbc89f41c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c838380),
	.w1(32'hbc0e86b6),
	.w2(32'hbbec8868),
	.w3(32'h3c3b69bc),
	.w4(32'h3bf8daa3),
	.w5(32'hba3389d6),
	.w6(32'hbb2d94d4),
	.w7(32'h3ade92eb),
	.w8(32'hbb89b28b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc418acf),
	.w1(32'hbc2e3690),
	.w2(32'hbcd739e4),
	.w3(32'hbc403a26),
	.w4(32'h39a327b3),
	.w5(32'hbc506d59),
	.w6(32'h3b70d3f8),
	.w7(32'hbbad4568),
	.w8(32'hbc6c1830),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5e49b),
	.w1(32'hbb5e0cd1),
	.w2(32'h3c5c2983),
	.w3(32'hbb708505),
	.w4(32'hbb5218d0),
	.w5(32'hbc7094c9),
	.w6(32'h3c8186c6),
	.w7(32'hbc076774),
	.w8(32'hbc44ba92),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18efc),
	.w1(32'h3bf459d5),
	.w2(32'hbb77ecd5),
	.w3(32'h3c073bf5),
	.w4(32'h3a9f4048),
	.w5(32'h3c872067),
	.w6(32'h3b2d3281),
	.w7(32'hbcae5c38),
	.w8(32'hbbd4efcb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc169e43),
	.w1(32'hbaed3018),
	.w2(32'hbb9059bc),
	.w3(32'h3c0ae4f3),
	.w4(32'hbb8728d0),
	.w5(32'hbb3e4a7a),
	.w6(32'hbbb36357),
	.w7(32'hbc031ffb),
	.w8(32'hbc160a70),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0e664),
	.w1(32'h3c12b70f),
	.w2(32'h3c5eb556),
	.w3(32'hbbb3fb00),
	.w4(32'h3b1feec9),
	.w5(32'h3a06c5e1),
	.w6(32'hbc3b67a9),
	.w7(32'h3b45b03e),
	.w8(32'h3c886122),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be711),
	.w1(32'hb91d13dd),
	.w2(32'hbc82f312),
	.w3(32'hbc97acd6),
	.w4(32'hbc58df61),
	.w5(32'hbcb09b57),
	.w6(32'h3a2539d4),
	.w7(32'hbc1d6c76),
	.w8(32'hbbaea6e4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a1cc0),
	.w1(32'hbb1c1075),
	.w2(32'hbc84727e),
	.w3(32'hbc541022),
	.w4(32'hbb7bea29),
	.w5(32'h3b90d65d),
	.w6(32'hbc585d75),
	.w7(32'hbc56767d),
	.w8(32'hbc3aed5f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06c33),
	.w1(32'h3a4bde3e),
	.w2(32'hbb33671c),
	.w3(32'hbca1d0e8),
	.w4(32'hba8eda9e),
	.w5(32'h39a983f9),
	.w6(32'h3bf55941),
	.w7(32'h3ccfe643),
	.w8(32'h3bb099c8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf84c5),
	.w1(32'hbb91ce2c),
	.w2(32'h3b9337d2),
	.w3(32'hbb82e6af),
	.w4(32'hbb800462),
	.w5(32'hba3b35cc),
	.w6(32'hbbc619f9),
	.w7(32'h3b82d449),
	.w8(32'h3b69a2c8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083ee0),
	.w1(32'h3aad5f98),
	.w2(32'hb982b18d),
	.w3(32'hbc4ded33),
	.w4(32'hbb5e9c5e),
	.w5(32'h3bda0f6b),
	.w6(32'hba302eb0),
	.w7(32'hbb6bf10d),
	.w8(32'hbc22a605),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cdf41),
	.w1(32'hbbd5732f),
	.w2(32'h3bd92987),
	.w3(32'h3c306345),
	.w4(32'h3ba14975),
	.w5(32'hbc906da5),
	.w6(32'hbc532619),
	.w7(32'h3d323aa8),
	.w8(32'h3c051c0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061265),
	.w1(32'h3ce827ed),
	.w2(32'hbb6cba2d),
	.w3(32'h3bdee83c),
	.w4(32'h3cf20ea5),
	.w5(32'hba78d4a6),
	.w6(32'h397cb804),
	.w7(32'hbc51f7d2),
	.w8(32'hbc91d067),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77337f),
	.w1(32'hbc92fca6),
	.w2(32'h3b9d36ba),
	.w3(32'h3b3a4ab3),
	.w4(32'h3b052baa),
	.w5(32'h3c0866aa),
	.w6(32'h3b22cbfa),
	.w7(32'hbc20da92),
	.w8(32'hbb25de9f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e2f7b),
	.w1(32'h3c81033a),
	.w2(32'hbc017c5b),
	.w3(32'h3a30d519),
	.w4(32'h3d08339c),
	.w5(32'h3c3a2a14),
	.w6(32'hbc738d9d),
	.w7(32'h3b96c5c9),
	.w8(32'hbae6b666),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26cbb1),
	.w1(32'hbb569cb0),
	.w2(32'h3c4ccd2e),
	.w3(32'hbb207ddd),
	.w4(32'hbc37bf0c),
	.w5(32'h3a9f10f4),
	.w6(32'hbbcf150d),
	.w7(32'hbcbfb8ec),
	.w8(32'hbc858a89),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eae5a),
	.w1(32'hbc91a317),
	.w2(32'h3bb79bbb),
	.w3(32'hbba167af),
	.w4(32'hbbfca017),
	.w5(32'hbbb9873e),
	.w6(32'h3b50e400),
	.w7(32'h3c2099a3),
	.w8(32'hba405e36),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc717),
	.w1(32'h3c43268b),
	.w2(32'h3c11a300),
	.w3(32'h3c8bcaf1),
	.w4(32'hbc8ecf8d),
	.w5(32'hbc59ac3b),
	.w6(32'hbbd06927),
	.w7(32'hbad32b08),
	.w8(32'hbbb0221c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b4444),
	.w1(32'hba5a8221),
	.w2(32'h3c878e1e),
	.w3(32'h3c0a076c),
	.w4(32'h3b3e6d6b),
	.w5(32'h3c48e50f),
	.w6(32'hbb10281b),
	.w7(32'h3bd13dc0),
	.w8(32'hbc7d5566),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc388d6e),
	.w1(32'hbb9695a0),
	.w2(32'hbba1adb4),
	.w3(32'h3b23ac2d),
	.w4(32'h3c82cebc),
	.w5(32'hbc0ddf81),
	.w6(32'hbb62d03a),
	.w7(32'hbca5ac2b),
	.w8(32'hba103059),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcec3e9),
	.w1(32'hbbe9710c),
	.w2(32'hbd33f573),
	.w3(32'h3d247bb5),
	.w4(32'h3bb1bc5c),
	.w5(32'hbc2ec9be),
	.w6(32'h3bba1763),
	.w7(32'h3c38cf1a),
	.w8(32'hbb1a7824),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab26c0),
	.w1(32'hbc1baf2b),
	.w2(32'h3c38f552),
	.w3(32'h3b4aae4b),
	.w4(32'h3a8abbc2),
	.w5(32'h3ca130d9),
	.w6(32'h3ab6e598),
	.w7(32'hbb3ff48f),
	.w8(32'h3cfe073a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca63282),
	.w1(32'hba30d564),
	.w2(32'hbc030764),
	.w3(32'hbbe5a975),
	.w4(32'hbb7c6483),
	.w5(32'hbc022722),
	.w6(32'hbab128e0),
	.w7(32'hbb86a401),
	.w8(32'h3c96a650),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc514bbb),
	.w1(32'h3a3a1f1d),
	.w2(32'h3c7fd1ce),
	.w3(32'h3b442101),
	.w4(32'h3bee9d56),
	.w5(32'h3d1b6b82),
	.w6(32'h3b596654),
	.w7(32'h3c84dc3b),
	.w8(32'hbc8883a2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9295a7a),
	.w1(32'h3be749c6),
	.w2(32'hbc6afb79),
	.w3(32'h3ccfea43),
	.w4(32'hbc7c660e),
	.w5(32'h3afa03dd),
	.w6(32'h3ae13571),
	.w7(32'hbb47b651),
	.w8(32'hbb46c9fa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50a6f2),
	.w1(32'hbce13c6b),
	.w2(32'h3c3e99fe),
	.w3(32'h3b1d2d19),
	.w4(32'h3b82cb02),
	.w5(32'hbba8dbc5),
	.w6(32'h3c7dae7a),
	.w7(32'h3c0e96c7),
	.w8(32'hbb92d4f7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbabb4),
	.w1(32'hbc83a2f6),
	.w2(32'hbb020038),
	.w3(32'hbc129476),
	.w4(32'hbc16803c),
	.w5(32'hbb806f7f),
	.w6(32'h3c4603f5),
	.w7(32'h3ad9bee2),
	.w8(32'hbb39dea2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1365b3),
	.w1(32'h3a0ddcee),
	.w2(32'h3c81aaac),
	.w3(32'hbcde06c0),
	.w4(32'h3a95484b),
	.w5(32'h3c83918c),
	.w6(32'h39f100b1),
	.w7(32'hbbcf3f7d),
	.w8(32'h3bd8f50d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d3729),
	.w1(32'h3d144bb7),
	.w2(32'hb9225be7),
	.w3(32'hbbc08ec1),
	.w4(32'h3b053fe5),
	.w5(32'hba23ceb8),
	.w6(32'hbbde0d72),
	.w7(32'h3c25c11f),
	.w8(32'h3b5f0820),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad5a8a),
	.w1(32'hbcc5b8c9),
	.w2(32'hbc64707f),
	.w3(32'hbc4009d0),
	.w4(32'hbcb782e6),
	.w5(32'h3bd12eeb),
	.w6(32'h3932e02a),
	.w7(32'h3a7f9b5d),
	.w8(32'hbc47b5f2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc356652),
	.w1(32'h3b95a57f),
	.w2(32'h3b242eb5),
	.w3(32'hbc953f89),
	.w4(32'h3a24cd9e),
	.w5(32'h3c76dba3),
	.w6(32'hbc081b4a),
	.w7(32'h39e2e962),
	.w8(32'h3b0ad81b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05578b),
	.w1(32'h3c2bab36),
	.w2(32'h3c49fc22),
	.w3(32'h3cafc15b),
	.w4(32'hbadb8d5e),
	.w5(32'hbc213718),
	.w6(32'hbc232385),
	.w7(32'h3cb0578a),
	.w8(32'hbc867133),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9160d5),
	.w1(32'h3c479c0e),
	.w2(32'h3ba8a30a),
	.w3(32'hbbcff6f7),
	.w4(32'hbc3286a8),
	.w5(32'hbbfbe03f),
	.w6(32'hbaf1a79d),
	.w7(32'h3b91ad2b),
	.w8(32'h3bc8b58b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b985c75),
	.w1(32'hbc2176dd),
	.w2(32'h3b2196ab),
	.w3(32'h3bd94620),
	.w4(32'h384d2ee0),
	.w5(32'h3c36af99),
	.w6(32'hbc93ba8d),
	.w7(32'h3c30ae2f),
	.w8(32'hbb561667),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9f11),
	.w1(32'hbb4b981e),
	.w2(32'hbc815862),
	.w3(32'h3aca9795),
	.w4(32'h3bf52cfa),
	.w5(32'hb9a40a87),
	.w6(32'hbc5a9933),
	.w7(32'hbb29d3b6),
	.w8(32'hbb888b15),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26d5bd),
	.w1(32'hbc2472aa),
	.w2(32'hbc40b26b),
	.w3(32'hbc086188),
	.w4(32'h3b87995a),
	.w5(32'hbbac0c19),
	.w6(32'hbc0db7ea),
	.w7(32'h3c555167),
	.w8(32'hbc0d3bff),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8666dc),
	.w1(32'hbc30dfc6),
	.w2(32'h3c0ed0ee),
	.w3(32'h398a3916),
	.w4(32'hbb54c0b2),
	.w5(32'hbc1e3123),
	.w6(32'hbbcded88),
	.w7(32'h3c38e27e),
	.w8(32'h3bfb8989),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a9ff4),
	.w1(32'hbb9de685),
	.w2(32'hbb19cfa4),
	.w3(32'h3b937c38),
	.w4(32'hbb541fa3),
	.w5(32'h3af885e7),
	.w6(32'hbbc17c6a),
	.w7(32'h3c0cfa1e),
	.w8(32'h3c853a68),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89e0be),
	.w1(32'h3b9ebda6),
	.w2(32'hbb2f1a85),
	.w3(32'h3b9b1b0d),
	.w4(32'hbbd5eea3),
	.w5(32'h3b50e21f),
	.w6(32'h3cead6c6),
	.w7(32'hba25a9a2),
	.w8(32'h3c7c9999),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d06ad),
	.w1(32'h3c6b99bf),
	.w2(32'h3b58adca),
	.w3(32'h3ba816ef),
	.w4(32'h3c1cb763),
	.w5(32'hbc3be777),
	.w6(32'hba2a4c4c),
	.w7(32'hbb8b5af5),
	.w8(32'h3afda78f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e81a7),
	.w1(32'hbbf89e1f),
	.w2(32'h3ad414ec),
	.w3(32'hbbd562d2),
	.w4(32'h3cf69ee6),
	.w5(32'hbb106b00),
	.w6(32'hbb8cc190),
	.w7(32'hba8e5a6c),
	.w8(32'hbbea03d1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c185fcd),
	.w1(32'hbab89187),
	.w2(32'hbb7372de),
	.w3(32'h3c4bbd88),
	.w4(32'hbbbd901c),
	.w5(32'hbb6de9fd),
	.w6(32'h3b6bcae5),
	.w7(32'hbc1b65ad),
	.w8(32'hbba52e2c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f2fac),
	.w1(32'hbc0518cd),
	.w2(32'h39656463),
	.w3(32'h3c020867),
	.w4(32'h3b919ef3),
	.w5(32'hbcaa93b7),
	.w6(32'hbb102563),
	.w7(32'hbca18a2c),
	.w8(32'hbc3a18f8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272bec),
	.w1(32'h3b390a32),
	.w2(32'hbbd68f8a),
	.w3(32'hbc317029),
	.w4(32'hbc137b51),
	.w5(32'hbc2f9412),
	.w6(32'hbc1443c4),
	.w7(32'hbbab71cc),
	.w8(32'h3c5a7c4a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd404),
	.w1(32'hbcad1d69),
	.w2(32'hbc61898b),
	.w3(32'h3b8e7121),
	.w4(32'hbd39c0d1),
	.w5(32'hbc01035b),
	.w6(32'hba836256),
	.w7(32'hbc1e71c8),
	.w8(32'hbc577141),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1e33f),
	.w1(32'h3b21abd1),
	.w2(32'hbbfaaff6),
	.w3(32'h3c04d3b2),
	.w4(32'hbbd4c8ed),
	.w5(32'hbc59d274),
	.w6(32'h3be00fc6),
	.w7(32'h3a4e8cf3),
	.w8(32'hbc81b6ae),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f4d8),
	.w1(32'h3b03a6e8),
	.w2(32'hbb455daf),
	.w3(32'hbb4643b8),
	.w4(32'h3b4a1c95),
	.w5(32'h3c16a9ff),
	.w6(32'hbce57398),
	.w7(32'h3b9700d4),
	.w8(32'hb9b09f70),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc193156),
	.w1(32'hbbf7fc7f),
	.w2(32'hbc3551fc),
	.w3(32'h3b1997e8),
	.w4(32'hbb8d1358),
	.w5(32'hbc9c0e2c),
	.w6(32'hbb817786),
	.w7(32'h3a319aac),
	.w8(32'hbb1b78ee),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64dd50),
	.w1(32'hbc0a09e0),
	.w2(32'hbcf07176),
	.w3(32'hbaeb69c1),
	.w4(32'hbbdde4db),
	.w5(32'hbbfb8ea3),
	.w6(32'hbaf2b6e7),
	.w7(32'hbc06230b),
	.w8(32'hbc062c83),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f76a),
	.w1(32'h3c055d9b),
	.w2(32'h3c12994f),
	.w3(32'hb94f8959),
	.w4(32'hbb82439b),
	.w5(32'hbc765478),
	.w6(32'h3be17591),
	.w7(32'hbb124ab5),
	.w8(32'h3bde314b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19655e),
	.w1(32'hbb9cd8d6),
	.w2(32'hba0de841),
	.w3(32'h3c0073e9),
	.w4(32'hb953906c),
	.w5(32'h39036b89),
	.w6(32'h3bb1fad5),
	.w7(32'hbac3c045),
	.w8(32'h3b8a685f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71d77),
	.w1(32'hbbf48a86),
	.w2(32'h3b191eca),
	.w3(32'hbb63dbb5),
	.w4(32'h3936e186),
	.w5(32'h3b36f58a),
	.w6(32'hbc015d69),
	.w7(32'hbc0d3476),
	.w8(32'hbc1ae669),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbac6f),
	.w1(32'hbb6b5393),
	.w2(32'hba700fc8),
	.w3(32'h3bbf98d8),
	.w4(32'h3d4c7b4c),
	.w5(32'h3b532483),
	.w6(32'hbc0eaf2b),
	.w7(32'h3d0e039c),
	.w8(32'hbcad00f8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04c9c0),
	.w1(32'h3b82a1ce),
	.w2(32'h395c1592),
	.w3(32'h3bcf7e0d),
	.w4(32'hbca32edd),
	.w5(32'hbcba65ff),
	.w6(32'h3cdd4cf7),
	.w7(32'h3b96109a),
	.w8(32'h3ab22fb6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f40e6),
	.w1(32'hbc26e6e3),
	.w2(32'hbae5bb34),
	.w3(32'hbb96f9a9),
	.w4(32'hbc021716),
	.w5(32'h3b2aa18a),
	.w6(32'hbbd55426),
	.w7(32'h3c216605),
	.w8(32'hbc183073),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4883e9),
	.w1(32'hbbc3b7fe),
	.w2(32'hbbd9b356),
	.w3(32'h3c28f12c),
	.w4(32'h3c67e811),
	.w5(32'hbc92a314),
	.w6(32'hbc2396f2),
	.w7(32'hbbca646a),
	.w8(32'h3d133aee),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa3684),
	.w1(32'h3c4c8a3b),
	.w2(32'hbbb0aa82),
	.w3(32'h3bd7c514),
	.w4(32'hbcd3e7e4),
	.w5(32'hbba5eec1),
	.w6(32'hbbdc4e09),
	.w7(32'hbbc0f6e6),
	.w8(32'hbc3bf981),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be644b0),
	.w1(32'h3babf2a4),
	.w2(32'hbbe47929),
	.w3(32'h3bb9f395),
	.w4(32'hb919fa60),
	.w5(32'hbc898a5b),
	.w6(32'hbc6110a7),
	.w7(32'h3a2639ec),
	.w8(32'hbb6399d1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28720f),
	.w1(32'hbc0d10c0),
	.w2(32'h3c4c0555),
	.w3(32'h3c846f08),
	.w4(32'hbb87175f),
	.w5(32'hbbae8455),
	.w6(32'h3c696fa0),
	.w7(32'h3bcf2b76),
	.w8(32'hbbddeff9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dbd4e),
	.w1(32'hbb510aff),
	.w2(32'hbc243b03),
	.w3(32'h3bcac4e4),
	.w4(32'hbc1a37a5),
	.w5(32'h3b2dd6ea),
	.w6(32'h3a9b7f64),
	.w7(32'hbb1fc8eb),
	.w8(32'hbbf1ae42),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf1fa4),
	.w1(32'hbaa0cc06),
	.w2(32'hbc9adf5f),
	.w3(32'h3c502f51),
	.w4(32'h3d03321e),
	.w5(32'hb9c61d2c),
	.w6(32'hbc328ef1),
	.w7(32'hba1df9b7),
	.w8(32'hba1d99bf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13efe1),
	.w1(32'hb9858066),
	.w2(32'hbb1a6351),
	.w3(32'hbc8d9e9e),
	.w4(32'hbb09191e),
	.w5(32'h3b2d8e19),
	.w6(32'h3b969cab),
	.w7(32'hbb3370e5),
	.w8(32'hbc8e8875),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a35fb),
	.w1(32'hba5cb9e9),
	.w2(32'hbc51f5fc),
	.w3(32'h3b11df84),
	.w4(32'hbbfec5a0),
	.w5(32'hbc57e258),
	.w6(32'h3b7a8cfa),
	.w7(32'hbc8dd30a),
	.w8(32'h3c54eebf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ce2c),
	.w1(32'hbb85c722),
	.w2(32'h3b65b6f6),
	.w3(32'hbbac56fa),
	.w4(32'h3b34e9ba),
	.w5(32'hba5b3893),
	.w6(32'hbc0dcc33),
	.w7(32'h3b1d16d7),
	.w8(32'h3a5bd17b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2711ce),
	.w1(32'hbbd4c343),
	.w2(32'hbc08b3a3),
	.w3(32'h3bf1bea6),
	.w4(32'h3bc2ba51),
	.w5(32'hbc9888ae),
	.w6(32'hbb5e6681),
	.w7(32'h3b3779d8),
	.w8(32'h3b934833),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5686b1),
	.w1(32'h3c127f3c),
	.w2(32'h3857f3a8),
	.w3(32'hbbb7fd97),
	.w4(32'hbcdf9819),
	.w5(32'h3ac7905c),
	.w6(32'h3c21f85f),
	.w7(32'hba895e14),
	.w8(32'hbaf8282d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf670b6),
	.w1(32'hbacb880f),
	.w2(32'hbac847c8),
	.w3(32'hbbfe6fdb),
	.w4(32'hbb8704e7),
	.w5(32'hbb5f9ed5),
	.w6(32'hbc41e049),
	.w7(32'hbba4b7a8),
	.w8(32'h3b2a3112),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13d14b),
	.w1(32'h3c77374f),
	.w2(32'hbbf5367a),
	.w3(32'hbb432852),
	.w4(32'hb9e34739),
	.w5(32'hbbd5d86c),
	.w6(32'h3b9af916),
	.w7(32'hbc7c72cf),
	.w8(32'h3aedb09b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934248),
	.w1(32'h3bde9a3d),
	.w2(32'h3ae43c4d),
	.w3(32'h3b7ff8fb),
	.w4(32'hbcb38d3e),
	.w5(32'hbbe17102),
	.w6(32'hb7a65a2a),
	.w7(32'hbbc72c87),
	.w8(32'h3ba0b6ed),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30843a),
	.w1(32'hbd17505a),
	.w2(32'hbb744410),
	.w3(32'hbca60442),
	.w4(32'h3ae33bbf),
	.w5(32'h3bfc8df2),
	.w6(32'h3bb41785),
	.w7(32'h3babee03),
	.w8(32'hbb35cf93),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8295df),
	.w1(32'hbbabe06c),
	.w2(32'h3b5cbc17),
	.w3(32'h3a087696),
	.w4(32'h3b3e0a0b),
	.w5(32'h3a0bb646),
	.w6(32'h3865f1e7),
	.w7(32'h3b4bf1bf),
	.w8(32'hbbaf936a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc243eba),
	.w1(32'hbc70aa99),
	.w2(32'h3af8da5c),
	.w3(32'h3a803783),
	.w4(32'hbc940e1f),
	.w5(32'hbba73313),
	.w6(32'hbc64337c),
	.w7(32'h3cb8dbdb),
	.w8(32'h3c86e3d2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4be28),
	.w1(32'h3bfc73c7),
	.w2(32'hbbcb9a2a),
	.w3(32'hbc233828),
	.w4(32'hba60b589),
	.w5(32'hbbd4241f),
	.w6(32'hba873a4c),
	.w7(32'hbc756352),
	.w8(32'hbb3428a1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4309cb),
	.w1(32'h3b02d873),
	.w2(32'h3ad3cf4c),
	.w3(32'hbcb7e6b4),
	.w4(32'hb9310e08),
	.w5(32'h3a0872a6),
	.w6(32'hbd095ef8),
	.w7(32'h3c5c408a),
	.w8(32'hbbbc20cf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9080),
	.w1(32'hba909779),
	.w2(32'h3c1963bc),
	.w3(32'hbabfe83d),
	.w4(32'hba2647da),
	.w5(32'hbb11ea26),
	.w6(32'h3c6688b2),
	.w7(32'hbb615a7f),
	.w8(32'hbb69a974),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3345),
	.w1(32'hba3a38a5),
	.w2(32'h3ccd99ac),
	.w3(32'h3ca197b8),
	.w4(32'h3cefb14d),
	.w5(32'h3c0b41c6),
	.w6(32'hbc15f523),
	.w7(32'hbc96e390),
	.w8(32'hbcacffd2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130b0c),
	.w1(32'h3bee9851),
	.w2(32'h3c916243),
	.w3(32'hbaf02139),
	.w4(32'hbc4dd8e6),
	.w5(32'h3c8d0696),
	.w6(32'h3bc02eaf),
	.w7(32'h3bc7b02f),
	.w8(32'h3d054e43),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9194bd),
	.w1(32'hbbe5fbe9),
	.w2(32'h3ba7102e),
	.w3(32'hbcbb8cd9),
	.w4(32'hbb5630ae),
	.w5(32'h3c28dd4d),
	.w6(32'hbcd99eaf),
	.w7(32'hbc76a008),
	.w8(32'hbc8eb722),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f46bd),
	.w1(32'h3c03967b),
	.w2(32'hbc49a8c5),
	.w3(32'hbc220208),
	.w4(32'hbc4f1654),
	.w5(32'h3abbdab1),
	.w6(32'h3b7fee03),
	.w7(32'hbc5a3120),
	.w8(32'h3b1a6637),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2df68c),
	.w1(32'hbd3b21ed),
	.w2(32'hbd22ff1b),
	.w3(32'h3bde0e77),
	.w4(32'h3b0e14af),
	.w5(32'h3b5f081c),
	.w6(32'h3b7fe6fe),
	.w7(32'h3b955d26),
	.w8(32'hbc14ac79),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241d96),
	.w1(32'hbc449da8),
	.w2(32'hbbe16cf4),
	.w3(32'hbaaca21b),
	.w4(32'hbc0a5a24),
	.w5(32'hbc0836b8),
	.w6(32'h3a373f49),
	.w7(32'hbc53eb48),
	.w8(32'hbaf4e2ec),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c6015),
	.w1(32'h3b9160bd),
	.w2(32'hbc419f78),
	.w3(32'h39ef5bbc),
	.w4(32'hbc89f2d8),
	.w5(32'hbb3bb4df),
	.w6(32'hbbf0760f),
	.w7(32'h3bc15d12),
	.w8(32'h3ba6b5d9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a917),
	.w1(32'h3a5b341d),
	.w2(32'hbbeba29d),
	.w3(32'hbbd1cd63),
	.w4(32'hb92a64cb),
	.w5(32'hbbf3cc04),
	.w6(32'hbb1edf68),
	.w7(32'hbc1ae351),
	.w8(32'hbc6294f0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9808673),
	.w1(32'hb9bce59d),
	.w2(32'h3c8a9f1a),
	.w3(32'hbbdc191f),
	.w4(32'h3c93d082),
	.w5(32'hbd37055c),
	.w6(32'h3b3d67ab),
	.w7(32'hbc13e706),
	.w8(32'hba38af9d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe77935),
	.w1(32'hbb82cd50),
	.w2(32'h3caf3c32),
	.w3(32'hbca9131d),
	.w4(32'h3bc3f6b4),
	.w5(32'hbcd2aa3c),
	.w6(32'hba16bebd),
	.w7(32'h3ca72780),
	.w8(32'h3bc91273),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7dec3),
	.w1(32'hba8ca9e7),
	.w2(32'h3c69c44f),
	.w3(32'hbaf765b8),
	.w4(32'hba48f829),
	.w5(32'h3c55e46c),
	.w6(32'h3bf487d0),
	.w7(32'h39be9ff3),
	.w8(32'h39918c84),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca0623),
	.w1(32'hbca3041d),
	.w2(32'hb9b26c70),
	.w3(32'h3baf27a0),
	.w4(32'h396409ba),
	.w5(32'hbbb3badd),
	.w6(32'hbcd3dd53),
	.w7(32'h3c70ac5b),
	.w8(32'hbbb30451),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb42d),
	.w1(32'hbb7aaf29),
	.w2(32'h3c2b269e),
	.w3(32'h3c72aacf),
	.w4(32'hbc2f20c5),
	.w5(32'h3acc0584),
	.w6(32'h3bc3a45e),
	.w7(32'hbc98419e),
	.w8(32'h3b800c25),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c50d8),
	.w1(32'hbb59fa76),
	.w2(32'h3caa1f15),
	.w3(32'hbd24d452),
	.w4(32'h3b4722b8),
	.w5(32'hbcf05f78),
	.w6(32'hbd122da9),
	.w7(32'h3ca6de22),
	.w8(32'h3b94cdc9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc05509),
	.w1(32'hbc685122),
	.w2(32'hbbafd927),
	.w3(32'h3cecb7ea),
	.w4(32'h3c3ab5fc),
	.w5(32'h3c0bdf88),
	.w6(32'h3b18acae),
	.w7(32'h3c9701d0),
	.w8(32'hbb6b804e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefc56f),
	.w1(32'hbcb99b6e),
	.w2(32'hba9a9d8a),
	.w3(32'h3b868a19),
	.w4(32'h3b6c1d90),
	.w5(32'h3b972618),
	.w6(32'hbaf1d9d1),
	.w7(32'hb98cc29c),
	.w8(32'hbc0ebbe3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87ef8c),
	.w1(32'hbb9cf3d0),
	.w2(32'hbc5344a9),
	.w3(32'hbb469471),
	.w4(32'h3c03d739),
	.w5(32'hbbefa5e4),
	.w6(32'hbc2058ca),
	.w7(32'h39fb42a7),
	.w8(32'hbbb61b35),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19f7c),
	.w1(32'h3bce9c46),
	.w2(32'hbbe3e6b6),
	.w3(32'hbca2e632),
	.w4(32'h3c0333e4),
	.w5(32'hbbd866f2),
	.w6(32'hbb331f1a),
	.w7(32'hbbf5fc82),
	.w8(32'h3c2bf279),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95322c),
	.w1(32'h3a36ed57),
	.w2(32'hbc72e65a),
	.w3(32'h3be492ab),
	.w4(32'hbc6d158f),
	.w5(32'h3c238ace),
	.w6(32'hbad7d702),
	.w7(32'hbc627ebc),
	.w8(32'h3c096185),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93e2a2),
	.w1(32'hbb5ae567),
	.w2(32'hbb89e5cb),
	.w3(32'h3b409b0c),
	.w4(32'h3ca3cce9),
	.w5(32'h3c14f9be),
	.w6(32'hbd06cc81),
	.w7(32'hbb345a63),
	.w8(32'hba821fd0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa5b8),
	.w1(32'hbc39f252),
	.w2(32'h3c366f56),
	.w3(32'h3cff2b60),
	.w4(32'hbcdda058),
	.w5(32'h3c0a8979),
	.w6(32'hbd0f781d),
	.w7(32'hbae9e0c8),
	.w8(32'h3b498e37),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf401a4),
	.w1(32'hbc70ce0b),
	.w2(32'hbbcf4ca6),
	.w3(32'hbc33c7c5),
	.w4(32'h3bbfabf6),
	.w5(32'hbc805bf6),
	.w6(32'h3c886cab),
	.w7(32'hbb566d32),
	.w8(32'h3c070246),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c751ea2),
	.w1(32'h3d126c1a),
	.w2(32'hbc19ca20),
	.w3(32'h3ce0d6ee),
	.w4(32'hbbcb3c66),
	.w5(32'h3cac84ac),
	.w6(32'hbd7019a6),
	.w7(32'h3ca6bc26),
	.w8(32'h3cb5b938),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c5545),
	.w1(32'h3c92cbbb),
	.w2(32'hbd1d45aa),
	.w3(32'hbc4466dd),
	.w4(32'h3c24e023),
	.w5(32'hbd33768c),
	.w6(32'hbb3c03b7),
	.w7(32'h3af22e2c),
	.w8(32'hbc6b0c27),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c316380),
	.w1(32'hbc1bdd62),
	.w2(32'hbca54b17),
	.w3(32'hbb8b7d5e),
	.w4(32'h3c137c8c),
	.w5(32'hbad7de51),
	.w6(32'hbb804dcb),
	.w7(32'hbb5164cd),
	.w8(32'h3b612b9a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad34d),
	.w1(32'h3cad402c),
	.w2(32'hbc76b96a),
	.w3(32'hbc10b4b8),
	.w4(32'h3c69975a),
	.w5(32'hbcaa1a33),
	.w6(32'hbbd977db),
	.w7(32'h3d0477b5),
	.w8(32'hbbed499f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6b9b1),
	.w1(32'h3adc67b6),
	.w2(32'hbc7db336),
	.w3(32'hbbcf9ade),
	.w4(32'h3ca633b6),
	.w5(32'hbc838a1d),
	.w6(32'h3aa9f682),
	.w7(32'h3ba27644),
	.w8(32'h3b00c2a5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab9b6),
	.w1(32'h3872511d),
	.w2(32'h3b5cc77d),
	.w3(32'h3b734a4d),
	.w4(32'h3c7009de),
	.w5(32'hbc49a865),
	.w6(32'h3be78ab5),
	.w7(32'hbb33407b),
	.w8(32'hbb0eafd2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54411d),
	.w1(32'h3c1fbbc6),
	.w2(32'hbc08e0f2),
	.w3(32'h3c9bf7ca),
	.w4(32'hbb204936),
	.w5(32'hbc04c4e0),
	.w6(32'h3c9550bd),
	.w7(32'h3c0f3a8f),
	.w8(32'h3b922fc7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0e2e3),
	.w1(32'h3c6af3eb),
	.w2(32'h3b7e9fcc),
	.w3(32'hbb9541fb),
	.w4(32'h3c4ab152),
	.w5(32'hbc174a5c),
	.w6(32'hbb034f9b),
	.w7(32'h3c31aacb),
	.w8(32'h3a8a709c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb408322),
	.w1(32'hbabbf108),
	.w2(32'h3c84d7e9),
	.w3(32'h3b30cb9f),
	.w4(32'h3cd31db9),
	.w5(32'hbac2ac13),
	.w6(32'hbc528663),
	.w7(32'h3d11c3a1),
	.w8(32'h3c09143b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05141e),
	.w1(32'h3ba6c9ba),
	.w2(32'h3cace533),
	.w3(32'hbb7f9854),
	.w4(32'h3c89acf9),
	.w5(32'h3ac4f745),
	.w6(32'hbb891bff),
	.w7(32'h3b75ec79),
	.w8(32'hbc6d7f6c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01307),
	.w1(32'hbbbdd2bb),
	.w2(32'h3af549b3),
	.w3(32'hbc89379d),
	.w4(32'h3b1a5ad4),
	.w5(32'hbb75cbcd),
	.w6(32'h3b6c11ad),
	.w7(32'h3b76bd80),
	.w8(32'hbc09815b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36ff2a),
	.w1(32'hbc082256),
	.w2(32'hbbdbe957),
	.w3(32'h3c0b930f),
	.w4(32'h3c059846),
	.w5(32'h3ba8622a),
	.w6(32'hbbade7b1),
	.w7(32'h3b0ea9fa),
	.w8(32'hbc0061d4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51b627),
	.w1(32'hbc8c9438),
	.w2(32'hbbe386b9),
	.w3(32'hba922d37),
	.w4(32'hbbd1f90b),
	.w5(32'hbbe2d22c),
	.w6(32'hbc027481),
	.w7(32'h3c05b194),
	.w8(32'hbb052514),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5298f0),
	.w1(32'h3a7f60bc),
	.w2(32'h3b39552f),
	.w3(32'h3c79b473),
	.w4(32'h3bf5304b),
	.w5(32'h3c0c87e3),
	.w6(32'hbc311766),
	.w7(32'h3b4df925),
	.w8(32'h3c66babd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaa9b4),
	.w1(32'hbaaced7e),
	.w2(32'h3b216294),
	.w3(32'hbaac1577),
	.w4(32'hb993e59a),
	.w5(32'hbbee5010),
	.w6(32'hbca6b711),
	.w7(32'hbb4a0d5d),
	.w8(32'hbaf4f3e4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210465),
	.w1(32'hbb67a350),
	.w2(32'h3d18d2fa),
	.w3(32'h3bb909cc),
	.w4(32'h3c26865a),
	.w5(32'hbb8cc68f),
	.w6(32'h399b5a6c),
	.w7(32'h3a1a59cb),
	.w8(32'hbb845f31),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc65504),
	.w1(32'hbae62a1d),
	.w2(32'hbb47cf6e),
	.w3(32'h3b94be6c),
	.w4(32'hbbe962ef),
	.w5(32'h3bdf05a2),
	.w6(32'hbc0bd3e1),
	.w7(32'hbc0acfa5),
	.w8(32'h3ce7f255),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ef6aa),
	.w1(32'h38ecf068),
	.w2(32'hbcffcc1d),
	.w3(32'hbafa5f49),
	.w4(32'hbb8536e0),
	.w5(32'h3b6527e3),
	.w6(32'h3c3b91de),
	.w7(32'h3b8dcb53),
	.w8(32'h39da4d8a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4928e3),
	.w1(32'hbc6c990f),
	.w2(32'h3ad46dcb),
	.w3(32'h3c0ddfae),
	.w4(32'hbd670c43),
	.w5(32'hbb94d2eb),
	.w6(32'hbc04a522),
	.w7(32'hbac89b34),
	.w8(32'h3b0710f3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d7b25),
	.w1(32'h3b3f55ea),
	.w2(32'h3be2d0cf),
	.w3(32'h3bcae812),
	.w4(32'h3b867669),
	.w5(32'h386a3024),
	.w6(32'h3bf7de62),
	.w7(32'hbc36948f),
	.w8(32'hbbc30b5e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f957c),
	.w1(32'hbcef4f1d),
	.w2(32'h3aa717b3),
	.w3(32'hbbce851d),
	.w4(32'hbb234ef2),
	.w5(32'hbb773a70),
	.w6(32'hbc068408),
	.w7(32'h3bd865e5),
	.w8(32'hba481162),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6dfb7),
	.w1(32'hbbb45155),
	.w2(32'hb8e7e7c6),
	.w3(32'h3c20f7c7),
	.w4(32'h3c027927),
	.w5(32'hbbb9e309),
	.w6(32'h3ba5608e),
	.w7(32'hbb822848),
	.w8(32'hbb10ef97),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04892b),
	.w1(32'h3c8cf169),
	.w2(32'h3bff1c46),
	.w3(32'h3b353d6d),
	.w4(32'h3cb41a73),
	.w5(32'h3b5dee56),
	.w6(32'h37d28692),
	.w7(32'hbbca9106),
	.w8(32'hbc8b4ae7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3ca90),
	.w1(32'hbbd2456d),
	.w2(32'h3b372985),
	.w3(32'hbc15f8d3),
	.w4(32'hbb802027),
	.w5(32'h3bf80470),
	.w6(32'hbb8205e4),
	.w7(32'hbbad4fbd),
	.w8(32'h3a83a3c0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ec247),
	.w1(32'hbbf3e689),
	.w2(32'hbbdfefdd),
	.w3(32'h3b095b48),
	.w4(32'hbc53084a),
	.w5(32'h3ab7cafe),
	.w6(32'h3c4ef34a),
	.w7(32'h3bae03fa),
	.w8(32'h3c308860),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54d4ac),
	.w1(32'hbb2437b3),
	.w2(32'hbb1bc8dd),
	.w3(32'hbb1e4980),
	.w4(32'h3b396cb3),
	.w5(32'hbae995b7),
	.w6(32'h3b00138a),
	.w7(32'h3c0290c0),
	.w8(32'hbb367447),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17eef8),
	.w1(32'h3baf3266),
	.w2(32'hba60e0a5),
	.w3(32'h3c1e5ba5),
	.w4(32'h3c43757b),
	.w5(32'hbbd7d54b),
	.w6(32'hbbd3ce74),
	.w7(32'h3c86431a),
	.w8(32'hbc2b67ae),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17bb41),
	.w1(32'h39916e64),
	.w2(32'hbb705059),
	.w3(32'h3bbd10af),
	.w4(32'h3bdd0cf4),
	.w5(32'h3c1900e8),
	.w6(32'h3c04c1f0),
	.w7(32'hbad48aa0),
	.w8(32'hbb9fcfcf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09afb),
	.w1(32'hbc03d86b),
	.w2(32'h3c0d657a),
	.w3(32'hbbb11bf8),
	.w4(32'hbb91fbd7),
	.w5(32'h3c2f0d6e),
	.w6(32'h3bbf0d1c),
	.w7(32'hbc3f4a1c),
	.w8(32'hbc9be45d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4364ee),
	.w1(32'h3bdc148e),
	.w2(32'hbca2e94f),
	.w3(32'hbb89ec3b),
	.w4(32'h3c042b83),
	.w5(32'hbc05345d),
	.w6(32'hbcb87263),
	.w7(32'hbb4b820f),
	.w8(32'h3d05ef81),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9df5c),
	.w1(32'hbc0985dc),
	.w2(32'hbc0ae430),
	.w3(32'h3bd75c7c),
	.w4(32'h3bd40ab4),
	.w5(32'hba5fbf60),
	.w6(32'hbc71e884),
	.w7(32'hbc170626),
	.w8(32'h3b67f0e0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71b9d),
	.w1(32'hba0fdae7),
	.w2(32'hbae75dc2),
	.w3(32'hb9c1f128),
	.w4(32'hbb7b7c3f),
	.w5(32'hbb9865b5),
	.w6(32'hbc9dd166),
	.w7(32'hbc08662c),
	.w8(32'hbc123bb0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3155),
	.w1(32'hbc872d0b),
	.w2(32'h3b772468),
	.w3(32'h3c457ce5),
	.w4(32'h3bbc63bf),
	.w5(32'hbc16378f),
	.w6(32'h3ba093bf),
	.w7(32'hbb5727b2),
	.w8(32'hbc22442a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b202fe4),
	.w1(32'h3b9adc0e),
	.w2(32'hbb09e5d0),
	.w3(32'hbc04853b),
	.w4(32'h3bbb32f4),
	.w5(32'hbb5fe32f),
	.w6(32'hbaf220a9),
	.w7(32'hbb443497),
	.w8(32'h3ce4370d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9920),
	.w1(32'hbb0da555),
	.w2(32'h3bf1f9a0),
	.w3(32'h3baa5807),
	.w4(32'hbbc22328),
	.w5(32'hbbb210c9),
	.w6(32'h3c4e1eab),
	.w7(32'hba4b64cc),
	.w8(32'hbb87e6c1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b6d4),
	.w1(32'hbba0c528),
	.w2(32'hbbd1373d),
	.w3(32'hbbdf0803),
	.w4(32'hbc7c7d37),
	.w5(32'hbcae9b6d),
	.w6(32'hbb7cb775),
	.w7(32'hbb9e766c),
	.w8(32'hbb781b84),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d29c2),
	.w1(32'h3c066a4a),
	.w2(32'hbbebffcc),
	.w3(32'h3b76a82d),
	.w4(32'h3be0107d),
	.w5(32'hbbf125f1),
	.w6(32'h3bd43bb2),
	.w7(32'hb9eee0f4),
	.w8(32'h3c772d8f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6aa361),
	.w1(32'h3bbfe46d),
	.w2(32'hbbe05a13),
	.w3(32'hbb1034b2),
	.w4(32'hbcaef572),
	.w5(32'hbb1e4219),
	.w6(32'h3c6be143),
	.w7(32'h3c191259),
	.w8(32'h3a448d64),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5749b2),
	.w1(32'hbb4f6a1c),
	.w2(32'h3ae088e0),
	.w3(32'hba7c4bfd),
	.w4(32'h3c31faf6),
	.w5(32'h3b435cc8),
	.w6(32'h3a8d90be),
	.w7(32'hbc2d2a31),
	.w8(32'hbb9d4fd9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ed2eb6),
	.w1(32'hbc54114c),
	.w2(32'hbb697c29),
	.w3(32'hbb7e57c0),
	.w4(32'hbc0556a6),
	.w5(32'h3c200f19),
	.w6(32'h3b7e0059),
	.w7(32'hbb89b590),
	.w8(32'hbb0890d9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7aba92),
	.w1(32'hbb8adddf),
	.w2(32'h38946a81),
	.w3(32'hbc29bfcb),
	.w4(32'hbc916cec),
	.w5(32'h3ca37e7f),
	.w6(32'hbc36ce86),
	.w7(32'h3c06549a),
	.w8(32'hbaf410cc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf68ce),
	.w1(32'hbba73576),
	.w2(32'h3bd0bf27),
	.w3(32'hbbb71204),
	.w4(32'hba342daf),
	.w5(32'hbb458f3a),
	.w6(32'hbc678fac),
	.w7(32'h3c0759a9),
	.w8(32'hbab2e764),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e26691),
	.w1(32'h3c4fc590),
	.w2(32'h3ca882e3),
	.w3(32'h3b457ffa),
	.w4(32'h3af6c277),
	.w5(32'hbb51c9ee),
	.w6(32'hbbd840e5),
	.w7(32'h3ab27d88),
	.w8(32'hbc3aaa35),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ec57a),
	.w1(32'hbc55e494),
	.w2(32'hbc4b62d6),
	.w3(32'hbbde5031),
	.w4(32'hbc2dc49b),
	.w5(32'hbbda00cf),
	.w6(32'h3bebb483),
	.w7(32'hbbd1b893),
	.w8(32'hbbbe128d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d61a),
	.w1(32'h3cdf5646),
	.w2(32'hb9c94aac),
	.w3(32'hbb965d43),
	.w4(32'hbbddc6a6),
	.w5(32'h3a63862e),
	.w6(32'hbb35cd72),
	.w7(32'hbbed8963),
	.w8(32'h3b616b43),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76d105),
	.w1(32'h3beddb8a),
	.w2(32'hbc68913d),
	.w3(32'hbb96c86f),
	.w4(32'h3c0e9ca3),
	.w5(32'h3a29cb8e),
	.w6(32'h3b9803d7),
	.w7(32'h3ba30852),
	.w8(32'h3bb3baaf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4b5d8),
	.w1(32'h3c458377),
	.w2(32'h3c527760),
	.w3(32'hbb9a8bdd),
	.w4(32'hb944bfaa),
	.w5(32'h3c81e72b),
	.w6(32'hbcb305f6),
	.w7(32'hbb9d11d2),
	.w8(32'h3bc9683e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e68b1),
	.w1(32'hbb0c242c),
	.w2(32'h3bafd036),
	.w3(32'hbb86f674),
	.w4(32'hbb81c646),
	.w5(32'h3b2ce9f4),
	.w6(32'hbc1a6728),
	.w7(32'hbbf79e5d),
	.w8(32'hbaf09f4d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba421d30),
	.w1(32'hbb6a76e2),
	.w2(32'hbba17f92),
	.w3(32'hbb5f1de7),
	.w4(32'hbb1de2c9),
	.w5(32'hbb43816f),
	.w6(32'hbc24a095),
	.w7(32'h3bed2364),
	.w8(32'hbbc831de),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2e2f),
	.w1(32'hbb4361c6),
	.w2(32'h39aa3c48),
	.w3(32'h3b3e0b9c),
	.w4(32'hbc0b40f2),
	.w5(32'h3b230cdf),
	.w6(32'h3b9f8d87),
	.w7(32'h3c086df9),
	.w8(32'hbbbcc0a1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50017f),
	.w1(32'h3bb2ad9a),
	.w2(32'hba489fb3),
	.w3(32'hbb7d3f69),
	.w4(32'hbbeace69),
	.w5(32'hba662036),
	.w6(32'hbb192972),
	.w7(32'hbb2e19b5),
	.w8(32'hbba71d6c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5e326),
	.w1(32'h3a56fd7d),
	.w2(32'h3c0a440a),
	.w3(32'h3b4cf2a8),
	.w4(32'h3cb8e907),
	.w5(32'h3b36c6ca),
	.w6(32'hbc5ccf9b),
	.w7(32'hbc7f5466),
	.w8(32'hbc471313),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0cfc1),
	.w1(32'h3bb9f84c),
	.w2(32'hbb9a6d73),
	.w3(32'h3ba00cf1),
	.w4(32'hbaab48fa),
	.w5(32'hbbf5faf9),
	.w6(32'h3b16825d),
	.w7(32'h3b80ce16),
	.w8(32'hbb13926f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad57baf),
	.w1(32'h3bb6ac29),
	.w2(32'hba885664),
	.w3(32'hbc1f698a),
	.w4(32'hb969ab36),
	.w5(32'h3bbdd984),
	.w6(32'hbbd95079),
	.w7(32'h3c99cb22),
	.w8(32'h3abb6efa),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafed454),
	.w1(32'hbb74bea8),
	.w2(32'h3ceaab9a),
	.w3(32'hbbff78a8),
	.w4(32'hbb517204),
	.w5(32'hba69a2d3),
	.w6(32'h3c4cd549),
	.w7(32'h3bb2435d),
	.w8(32'h3bc8729e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc522be1),
	.w1(32'h3b766cde),
	.w2(32'h3acab2ec),
	.w3(32'h3c3961a5),
	.w4(32'hbb7e82e0),
	.w5(32'h3a690ac8),
	.w6(32'h3aa6c142),
	.w7(32'h3c0d504e),
	.w8(32'hbaae4251),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c014c67),
	.w1(32'hba06c72d),
	.w2(32'h3b0b9160),
	.w3(32'h3b83541b),
	.w4(32'h3a5d9b35),
	.w5(32'h3bb9cefb),
	.w6(32'h3ccb67f9),
	.w7(32'hbaa3a6df),
	.w8(32'hbbef7709),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058eba),
	.w1(32'hb9bd7ff7),
	.w2(32'hbc39c5d2),
	.w3(32'hba447ecf),
	.w4(32'h3ba7f7e9),
	.w5(32'h3bc7cca3),
	.w6(32'hbb8ab570),
	.w7(32'h3c12a9d1),
	.w8(32'hbc86c0af),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba5f6),
	.w1(32'hbc670e06),
	.w2(32'hba8727df),
	.w3(32'h3b897f6f),
	.w4(32'hbbb013fb),
	.w5(32'h3c11a882),
	.w6(32'h39c2ea4a),
	.w7(32'hbc27444f),
	.w8(32'hbb7e6ddf),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13a261),
	.w1(32'hbcde3e26),
	.w2(32'h3bd22c02),
	.w3(32'hbc4a9062),
	.w4(32'h3be6bc1a),
	.w5(32'hbc24f21c),
	.w6(32'hbb9bdcfb),
	.w7(32'h3b781f67),
	.w8(32'h3cbff3b8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45a31b),
	.w1(32'hbba7ed6d),
	.w2(32'hbae1f4e5),
	.w3(32'h3be5903b),
	.w4(32'h3bd0d155),
	.w5(32'h3c619783),
	.w6(32'hbbc36ee1),
	.w7(32'hbaf2f29b),
	.w8(32'hb914656c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf36ca),
	.w1(32'h3b0a3628),
	.w2(32'h3ba7d841),
	.w3(32'hbc37f209),
	.w4(32'hbb630025),
	.w5(32'hbc1aeb04),
	.w6(32'hbccc6f3a),
	.w7(32'h3c2a249e),
	.w8(32'h3b6ed72a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ca975),
	.w1(32'hbca12c36),
	.w2(32'hbc773e09),
	.w3(32'h3b11807a),
	.w4(32'hbc373b58),
	.w5(32'hb926ab54),
	.w6(32'h3b6e4a28),
	.w7(32'h3b035de4),
	.w8(32'hbbe7af9d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3d3c),
	.w1(32'hbc515fe9),
	.w2(32'h3b0504b2),
	.w3(32'h38506a69),
	.w4(32'h3c295a96),
	.w5(32'hbbb65027),
	.w6(32'hbc6d37da),
	.w7(32'hbbd3a9ae),
	.w8(32'h39de780b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3399c2),
	.w1(32'h3b74fafc),
	.w2(32'hbc80ed60),
	.w3(32'h3bcf1761),
	.w4(32'h3b57f253),
	.w5(32'hbcb31ef0),
	.w6(32'h3abf3a43),
	.w7(32'h3b3c5c79),
	.w8(32'h3bb022ca),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b58c5),
	.w1(32'h3c0e8fc4),
	.w2(32'h3b829e41),
	.w3(32'h3c7ab42f),
	.w4(32'h3b94436a),
	.w5(32'hbc75e20a),
	.w6(32'h3c019b6f),
	.w7(32'hbb53fe3b),
	.w8(32'hbc88dd51),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547f12),
	.w1(32'h3a08211f),
	.w2(32'h3cb9dacc),
	.w3(32'hbb3ad9c7),
	.w4(32'h3c0461ac),
	.w5(32'h3c174da5),
	.w6(32'h3a695ffb),
	.w7(32'h3c509c53),
	.w8(32'hbb83d4a4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059a87),
	.w1(32'h3a28ff11),
	.w2(32'h3ac64188),
	.w3(32'hbba6d203),
	.w4(32'h3b6b1979),
	.w5(32'h3b22df1d),
	.w6(32'hbc69a617),
	.w7(32'h3a853c5c),
	.w8(32'h3a6b0fb2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cb018),
	.w1(32'h3c7e5e9c),
	.w2(32'hbaaa5cd2),
	.w3(32'h3bc55b52),
	.w4(32'h3b1ca615),
	.w5(32'h3c480705),
	.w6(32'hbb465757),
	.w7(32'h39fd24c3),
	.w8(32'h3b0dde73),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab6fb),
	.w1(32'h3bbd8b27),
	.w2(32'h3c27feeb),
	.w3(32'hbb81dd05),
	.w4(32'h3b9aa105),
	.w5(32'hbbadd5df),
	.w6(32'hbc2158c5),
	.w7(32'hbbe71d63),
	.w8(32'hbbfdcefb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb085c27),
	.w1(32'hba6a5a41),
	.w2(32'hbb83f4ad),
	.w3(32'hbc524372),
	.w4(32'h3aa9d220),
	.w5(32'h3c785539),
	.w6(32'h3c2067ce),
	.w7(32'hbbeb468a),
	.w8(32'h3c304e1f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87192),
	.w1(32'h3b62c764),
	.w2(32'h3c10cc2b),
	.w3(32'hbcb65664),
	.w4(32'hbb8b23d0),
	.w5(32'h3bf1acf1),
	.w6(32'h3b98c9a5),
	.w7(32'hba39aa0b),
	.w8(32'h3b8bed47),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9b5bd),
	.w1(32'hbd08a588),
	.w2(32'h3b73c8f3),
	.w3(32'h3b9b6599),
	.w4(32'hba621526),
	.w5(32'h3b3328e4),
	.w6(32'hbc0dbbaa),
	.w7(32'hbc8c3c18),
	.w8(32'hbc755f5e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c509),
	.w1(32'h3b74b5c3),
	.w2(32'h3c2bcd3e),
	.w3(32'hbbb81d13),
	.w4(32'h3b435683),
	.w5(32'h3c1c05e8),
	.w6(32'hba87fe0b),
	.w7(32'hbcd5e9cc),
	.w8(32'h3bcb634b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc530da4),
	.w1(32'hbae1d826),
	.w2(32'h3c87c33d),
	.w3(32'hbbba2f31),
	.w4(32'hbb26c94e),
	.w5(32'hbc54962b),
	.w6(32'h38c74d3f),
	.w7(32'hbc4f112d),
	.w8(32'h3abfe3f0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd113ee),
	.w1(32'h3c7c1c28),
	.w2(32'hbbb3ec12),
	.w3(32'h3b412bb9),
	.w4(32'hbc8ff3e5),
	.w5(32'hbbee9fde),
	.w6(32'h3bfaeefd),
	.w7(32'hbc578746),
	.w8(32'hbc709132),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed25f),
	.w1(32'hbba07cde),
	.w2(32'h3abc0f15),
	.w3(32'h3b1f7c66),
	.w4(32'hb9fb17ec),
	.w5(32'hbc436a74),
	.w6(32'h3bbfebd1),
	.w7(32'hbc008ba1),
	.w8(32'hbc95dcf2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c177),
	.w1(32'hba96ac36),
	.w2(32'hbbe7b790),
	.w3(32'hba297850),
	.w4(32'h3c2fdeea),
	.w5(32'h3b0b3b45),
	.w6(32'hbbb79f97),
	.w7(32'hbb230238),
	.w8(32'hba87b212),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bdf8b),
	.w1(32'h3ad4e573),
	.w2(32'h3b6a54c1),
	.w3(32'hba8738cb),
	.w4(32'hbc25bddc),
	.w5(32'h3c58ece4),
	.w6(32'h3b82630b),
	.w7(32'h3900cd94),
	.w8(32'h3b5ffaf7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12911b),
	.w1(32'h3ab2e7e4),
	.w2(32'h3bcc58db),
	.w3(32'h3b8ef529),
	.w4(32'hba02a467),
	.w5(32'hbb06d072),
	.w6(32'h39071b04),
	.w7(32'h3b75dcc0),
	.w8(32'hbc8db9af),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11bfbd),
	.w1(32'hbc31a6f6),
	.w2(32'h3b0f5ac6),
	.w3(32'hbc5660a8),
	.w4(32'hbb20c7d8),
	.w5(32'hbb84657e),
	.w6(32'h3a4be4cc),
	.w7(32'hbab3c586),
	.w8(32'hbb04af19),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55a53),
	.w1(32'hbbc74c5e),
	.w2(32'hb9d66dfe),
	.w3(32'h3be67abe),
	.w4(32'h3c1fddbc),
	.w5(32'hba291238),
	.w6(32'h3b06b9eb),
	.w7(32'hbbbc9a4d),
	.w8(32'hbc8c43f2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575c67),
	.w1(32'hbb5de193),
	.w2(32'h3babc248),
	.w3(32'h3baf8640),
	.w4(32'h3bad6712),
	.w5(32'hbb470fea),
	.w6(32'h3bc3a1a2),
	.w7(32'h3c07c8c2),
	.w8(32'hbbba9a0f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3211fe),
	.w1(32'hbb7218d9),
	.w2(32'hbc40471b),
	.w3(32'hbbb6f9c8),
	.w4(32'h3c876919),
	.w5(32'hbb939e8c),
	.w6(32'hbb81b0e5),
	.w7(32'hbc1f2f7e),
	.w8(32'hbb035da3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12f2be),
	.w1(32'h3c11c8de),
	.w2(32'hbb8eba30),
	.w3(32'hba84c006),
	.w4(32'hbbb83bb4),
	.w5(32'h3b8e7b29),
	.w6(32'hbb1ef19f),
	.w7(32'hbc235e6b),
	.w8(32'hba6756b1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1495de),
	.w1(32'h3c46b540),
	.w2(32'hbc5d8f68),
	.w3(32'hbbac1d68),
	.w4(32'h3c2a2ba5),
	.w5(32'h3c7ff29a),
	.w6(32'hbba88a98),
	.w7(32'hbcacdb8c),
	.w8(32'h3c34b719),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f8861),
	.w1(32'hbb7e4b69),
	.w2(32'h3c05ad8f),
	.w3(32'hba95e620),
	.w4(32'hbaa555db),
	.w5(32'hbce1cec4),
	.w6(32'h3b8cbfdb),
	.w7(32'hbc036406),
	.w8(32'hbbc1e977),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c62fd),
	.w1(32'h3ab7bacd),
	.w2(32'hbc0d658c),
	.w3(32'h3ca298d2),
	.w4(32'hbbfa0348),
	.w5(32'h3897cdf2),
	.w6(32'h3ba22051),
	.w7(32'hbb501832),
	.w8(32'hbad6cbfe),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c517f6e),
	.w1(32'hbcb378ff),
	.w2(32'hbba18d29),
	.w3(32'hbc0de138),
	.w4(32'h3c3eb8c6),
	.w5(32'hba9f8f39),
	.w6(32'h3c874983),
	.w7(32'hbba78001),
	.w8(32'h3bf009a5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d82e7),
	.w1(32'hbd0117d3),
	.w2(32'h39daaee8),
	.w3(32'hb94d7971),
	.w4(32'hbb6eb54e),
	.w5(32'h393e4727),
	.w6(32'hbb315dae),
	.w7(32'hbcf94f6d),
	.w8(32'hbb83fa5f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cf7c4),
	.w1(32'h3b320614),
	.w2(32'hbbf9b578),
	.w3(32'h3b3a3c2d),
	.w4(32'h3bb5cf8d),
	.w5(32'hb8e9de0c),
	.w6(32'h3bab63f6),
	.w7(32'hbb863568),
	.w8(32'hbb5b1453),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5e416),
	.w1(32'hbb04b3ed),
	.w2(32'hbc464802),
	.w3(32'hbc24fed9),
	.w4(32'hb9f09dc8),
	.w5(32'h3abe7bae),
	.w6(32'hbb845130),
	.w7(32'h3c23dda7),
	.w8(32'h3cd415c5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5399de),
	.w1(32'hba13704d),
	.w2(32'h3c3f8e8c),
	.w3(32'hbbcc8650),
	.w4(32'hbc93e55a),
	.w5(32'hbbb35b84),
	.w6(32'h3babfff2),
	.w7(32'h3bb4e755),
	.w8(32'h3c1be48b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7be1aa),
	.w1(32'h3b9290b3),
	.w2(32'h39f0ffbb),
	.w3(32'hbcd412e1),
	.w4(32'h3ab65e82),
	.w5(32'hba4b8369),
	.w6(32'h3c418a16),
	.w7(32'h3bbbca7d),
	.w8(32'h3ae18db7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f1b4),
	.w1(32'hbb2c2bf8),
	.w2(32'h3b3da008),
	.w3(32'h3bfd4ca5),
	.w4(32'hbb91d4c9),
	.w5(32'hbba130f3),
	.w6(32'h3d24655c),
	.w7(32'h3cb36383),
	.w8(32'h3c029646),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4acf13),
	.w1(32'h3c5d6c0d),
	.w2(32'h3bab5597),
	.w3(32'h3cfa8f7f),
	.w4(32'hbaeb5eac),
	.w5(32'hbb04b493),
	.w6(32'h3baa500e),
	.w7(32'h3b922a01),
	.w8(32'h3b7c644f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a307880),
	.w1(32'hbbf14e92),
	.w2(32'hbc30c1f4),
	.w3(32'hbce464b2),
	.w4(32'h3b2c1f27),
	.w5(32'hbae231f5),
	.w6(32'hbc0d43b0),
	.w7(32'h3967ce07),
	.w8(32'h3bbc74c7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96822d),
	.w1(32'h3c3c7dcc),
	.w2(32'h3a5e41d0),
	.w3(32'hbcacf530),
	.w4(32'hbbe63b3b),
	.w5(32'h3c32cfeb),
	.w6(32'h3c2ffaa6),
	.w7(32'hbb300bab),
	.w8(32'hb9fa4fe5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c68f6e),
	.w1(32'hbc549396),
	.w2(32'h3afecb80),
	.w3(32'h3bd40fdd),
	.w4(32'h3bd6e9b8),
	.w5(32'h3c2e03d3),
	.w6(32'hbc3fc41d),
	.w7(32'h39d73266),
	.w8(32'h3ac46866),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022ba7),
	.w1(32'h3a97b052),
	.w2(32'h3b05a612),
	.w3(32'h3bcbadac),
	.w4(32'h3abbc63d),
	.w5(32'h3a1ba836),
	.w6(32'hbba20226),
	.w7(32'h39ff0969),
	.w8(32'h3cf7bfab),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a831b),
	.w1(32'h3bc25e8f),
	.w2(32'h3c043b41),
	.w3(32'hbb03e254),
	.w4(32'hbb86c586),
	.w5(32'hbc4b13b5),
	.w6(32'h3bc29212),
	.w7(32'hbbba7480),
	.w8(32'hbbc34178),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc48cb8),
	.w1(32'h3c5687e2),
	.w2(32'h3b698dc0),
	.w3(32'h3c3ba473),
	.w4(32'hbc71a941),
	.w5(32'hbb7c0610),
	.w6(32'hbc01a01f),
	.w7(32'hbc442b33),
	.w8(32'h3c1be68e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1bf09),
	.w1(32'hbb9c38f7),
	.w2(32'hb90c9eef),
	.w3(32'hba8fcfa0),
	.w4(32'hbb7eda1e),
	.w5(32'h3b8e94c8),
	.w6(32'hbc32fcf4),
	.w7(32'hbc714451),
	.w8(32'h3af90e14),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c178ca6),
	.w1(32'h3bc7ef50),
	.w2(32'hbc1951da),
	.w3(32'hbca9195f),
	.w4(32'h3c030b20),
	.w5(32'hbc44a914),
	.w6(32'hbb3e30fd),
	.w7(32'h3b5c5dd5),
	.w8(32'h3ba02a72),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec60d9),
	.w1(32'h3ccbc40f),
	.w2(32'h3b7c0364),
	.w3(32'hbca2317f),
	.w4(32'h3cd55c18),
	.w5(32'h3c3042a5),
	.w6(32'hbab836c4),
	.w7(32'h3bc4775c),
	.w8(32'hbc8c657b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63228d),
	.w1(32'hbc3054e0),
	.w2(32'h3c238dcf),
	.w3(32'hbc146a30),
	.w4(32'hbc0c6998),
	.w5(32'h3c082369),
	.w6(32'h3a63eff0),
	.w7(32'h3af1fe0e),
	.w8(32'hbbd0f5ab),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc441951),
	.w1(32'h3c1cf748),
	.w2(32'h3b4a99b5),
	.w3(32'h3bde5edb),
	.w4(32'h3bf35225),
	.w5(32'h3c5c20aa),
	.w6(32'h3c46175e),
	.w7(32'hbb143f28),
	.w8(32'h3c428c21),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bd643),
	.w1(32'h3c783f93),
	.w2(32'h3b631424),
	.w3(32'h3b469d4b),
	.w4(32'h3c27c7b8),
	.w5(32'hbc9e50dc),
	.w6(32'h3b835d67),
	.w7(32'h3a0662d7),
	.w8(32'h3b7846a9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ae49),
	.w1(32'hbbc0d491),
	.w2(32'hbb1925a3),
	.w3(32'h3c3005f5),
	.w4(32'hbbab8577),
	.w5(32'h3a1bc560),
	.w6(32'h3bbd35f4),
	.w7(32'hbb86e763),
	.w8(32'hbbb5bbf1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb730e),
	.w1(32'hba575e60),
	.w2(32'h3c1f87d7),
	.w3(32'h3bdcf0eb),
	.w4(32'h3a50b379),
	.w5(32'h3acc48b5),
	.w6(32'hbb6c7622),
	.w7(32'h3bd91ef6),
	.w8(32'hbd880c0c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ab26),
	.w1(32'h3d344323),
	.w2(32'hbbe535a1),
	.w3(32'h3bd1db89),
	.w4(32'hbc6ee1a3),
	.w5(32'h3b86df68),
	.w6(32'hbbd123df),
	.w7(32'hbba76cf4),
	.w8(32'h3b2e50c1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3d02),
	.w1(32'h3b05d5ea),
	.w2(32'hbc07e292),
	.w3(32'hbb5ce2e3),
	.w4(32'hbb5e7e2d),
	.w5(32'h3a3fbfaa),
	.w6(32'hbb485c83),
	.w7(32'h3c088618),
	.w8(32'hbb5bab65),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780f8f),
	.w1(32'hbb8053c4),
	.w2(32'h3baacff2),
	.w3(32'h3c54cf84),
	.w4(32'h3ca9383c),
	.w5(32'hbb29e5e7),
	.w6(32'hbb24ca55),
	.w7(32'h3a6d651a),
	.w8(32'hbb14d675),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e6a0),
	.w1(32'h3b448aeb),
	.w2(32'hbce67a24),
	.w3(32'hbae84fd1),
	.w4(32'h3c3a7bc8),
	.w5(32'h3bd44734),
	.w6(32'hbb6903eb),
	.w7(32'h37ba04e6),
	.w8(32'hbc53e2f6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85d509),
	.w1(32'h3b57087f),
	.w2(32'hbc19a0ba),
	.w3(32'hbb505521),
	.w4(32'h3bc6e822),
	.w5(32'hbcc49501),
	.w6(32'h3b7b7243),
	.w7(32'h3a892cc5),
	.w8(32'hbc2f309c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39438d),
	.w1(32'h3c79a97e),
	.w2(32'hbbc24a01),
	.w3(32'hbacdee11),
	.w4(32'h3c62f018),
	.w5(32'hb8bd101a),
	.w6(32'h3b6d5ddd),
	.w7(32'hbd2e17be),
	.w8(32'hbc3f7cb7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6dd4),
	.w1(32'h39bc7b9a),
	.w2(32'h3bac37c3),
	.w3(32'hbbea15d0),
	.w4(32'h3abe2937),
	.w5(32'hbb67779e),
	.w6(32'h3b0fae6a),
	.w7(32'hb98d1655),
	.w8(32'h3b4fb3c4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb30db),
	.w1(32'h3c4294b3),
	.w2(32'h3b38f4ae),
	.w3(32'h3b46477a),
	.w4(32'hbb67161e),
	.w5(32'h3bac26d1),
	.w6(32'hba73ee28),
	.w7(32'hbcc5895c),
	.w8(32'h3b35d320),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59fd06),
	.w1(32'h3c5958c4),
	.w2(32'hbc49b8b2),
	.w3(32'h3994678a),
	.w4(32'hbc0d681a),
	.w5(32'h3d01bc26),
	.w6(32'h3c2de5ca),
	.w7(32'hba6502af),
	.w8(32'h3bc0b1f2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7145f1),
	.w1(32'h3bc2d54c),
	.w2(32'hbb49d498),
	.w3(32'h3b862b85),
	.w4(32'h3b97f1d1),
	.w5(32'hba675c7b),
	.w6(32'hbc738739),
	.w7(32'h39fd0f61),
	.w8(32'hbc25649a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe11987),
	.w1(32'h3c9dd3e2),
	.w2(32'h3b350b08),
	.w3(32'h3c3000bc),
	.w4(32'h3a78c35d),
	.w5(32'hba4e5d01),
	.w6(32'h3b1e7453),
	.w7(32'h3bb9f07a),
	.w8(32'hbbaeba8d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bf744),
	.w1(32'h39339e25),
	.w2(32'hba971e5e),
	.w3(32'h3bf2186a),
	.w4(32'hbbb67bc7),
	.w5(32'h3a53d5a4),
	.w6(32'h3b33ebed),
	.w7(32'h3b3d0473),
	.w8(32'h3b0c18f5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c542e44),
	.w1(32'hbb6323c9),
	.w2(32'hbcc29c80),
	.w3(32'h3c0ad2ab),
	.w4(32'h3cb9a4bb),
	.w5(32'hbc6d1203),
	.w6(32'hb915c8fa),
	.w7(32'h3aa14f07),
	.w8(32'hbcf1d4d3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06ee74),
	.w1(32'hbb30e591),
	.w2(32'hbc458736),
	.w3(32'h3bff73c0),
	.w4(32'hbc223996),
	.w5(32'hbccb9923),
	.w6(32'hba89c5f7),
	.w7(32'h3c00edad),
	.w8(32'hbc8b1757),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc08f65),
	.w1(32'hb92aa701),
	.w2(32'h3bd98051),
	.w3(32'hbc1f966c),
	.w4(32'hbc5cd631),
	.w5(32'hbc514aeb),
	.w6(32'hba600a32),
	.w7(32'h3c339102),
	.w8(32'hbbeaf88d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c00bb),
	.w1(32'h3c11bf0f),
	.w2(32'h39c9bf30),
	.w3(32'hbc038c2d),
	.w4(32'hbb6a5a38),
	.w5(32'h3a085b82),
	.w6(32'hbc02f326),
	.w7(32'h3bdae17f),
	.w8(32'hbc3dd5c6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857a9d),
	.w1(32'hb9b781fe),
	.w2(32'hbaa4163d),
	.w3(32'h3babb575),
	.w4(32'hbb86b577),
	.w5(32'hbc2553b7),
	.w6(32'h3a0bcc4f),
	.w7(32'hbbdba8a4),
	.w8(32'h3ad11487),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac01e64),
	.w1(32'h3b7960cf),
	.w2(32'h3bb4c4f7),
	.w3(32'hbbd1bc4e),
	.w4(32'h3ae354b0),
	.w5(32'h3ba57dd1),
	.w6(32'hbb1c7eb9),
	.w7(32'h398f3f3f),
	.w8(32'hbb294dca),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8d652),
	.w1(32'h3ba3a7ac),
	.w2(32'h3ad53fe5),
	.w3(32'h3ba5ecd0),
	.w4(32'hba58e106),
	.w5(32'h3987f01a),
	.w6(32'h3c901921),
	.w7(32'h3b5d7c31),
	.w8(32'h3be4232a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f850),
	.w1(32'h3b355f66),
	.w2(32'hbb1bce50),
	.w3(32'hbb2b6c12),
	.w4(32'hbb3cf4b9),
	.w5(32'hbbecbcdd),
	.w6(32'h3c6c56df),
	.w7(32'hbb46bf05),
	.w8(32'hbb0f0404),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4745),
	.w1(32'hba9fc97d),
	.w2(32'h3b1d65bc),
	.w3(32'hbc182d02),
	.w4(32'hbc84c29e),
	.w5(32'hbb8f8fbc),
	.w6(32'hbb7fb5e0),
	.w7(32'h3bb68d1a),
	.w8(32'h3b4fd747),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa49451),
	.w1(32'h3b6a0144),
	.w2(32'hbb19ace3),
	.w3(32'h3b916533),
	.w4(32'h3ce31cb2),
	.w5(32'h3c0df22e),
	.w6(32'hbba61cd2),
	.w7(32'hbc5e6eb4),
	.w8(32'h3b9f043b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36e032),
	.w1(32'hbbfbc151),
	.w2(32'hbbc809d6),
	.w3(32'hbc1cbd1e),
	.w4(32'hbbb8d1a1),
	.w5(32'hbd1be818),
	.w6(32'h3be7ba71),
	.w7(32'hbbd3a903),
	.w8(32'hbb5496a8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd0172),
	.w1(32'hbc01842a),
	.w2(32'h3b96750c),
	.w3(32'h3c1cf220),
	.w4(32'hbb9915e8),
	.w5(32'hbcdb0467),
	.w6(32'h3b9208ba),
	.w7(32'h3b166746),
	.w8(32'hbc460904),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12307e),
	.w1(32'hbb2d1ad3),
	.w2(32'hbb9524b8),
	.w3(32'h393ce66e),
	.w4(32'h3bb312b1),
	.w5(32'hbbaa0a0d),
	.w6(32'hbbd98c98),
	.w7(32'hbc9f64fd),
	.w8(32'h3bba3fb1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b9532),
	.w1(32'hbc83f830),
	.w2(32'hbc767b9b),
	.w3(32'h3a68b81c),
	.w4(32'hbbcbe4be),
	.w5(32'h3c0b6676),
	.w6(32'hbbd75ee5),
	.w7(32'hbc85b936),
	.w8(32'h3a4ad9ec),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7928240),
	.w1(32'h3b7dd23b),
	.w2(32'h3c05eb2c),
	.w3(32'hbb75346d),
	.w4(32'h3b4d69c1),
	.w5(32'hbc645041),
	.w6(32'h3c8a0114),
	.w7(32'h3c1afd8f),
	.w8(32'h39ff201a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eaa73),
	.w1(32'h3bd591d3),
	.w2(32'h3a1e0b4e),
	.w3(32'h3c32d64a),
	.w4(32'hbc420a37),
	.w5(32'h3c3d951f),
	.w6(32'h3be7fd59),
	.w7(32'h399009c0),
	.w8(32'h3a19c910),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba200b3),
	.w1(32'hbb341b7d),
	.w2(32'hbc7fabb1),
	.w3(32'h3d2421f5),
	.w4(32'h3b2b5eed),
	.w5(32'hbcda750e),
	.w6(32'h3bdc528e),
	.w7(32'h3ad47a39),
	.w8(32'hbc68c43a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb69c1c),
	.w1(32'hbbbf9461),
	.w2(32'h3b4bda09),
	.w3(32'hbad6dbf8),
	.w4(32'hbba6745c),
	.w5(32'h3c1c06b6),
	.w6(32'h39fcd33e),
	.w7(32'h3b2bf45d),
	.w8(32'hba6d8ed1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1486),
	.w1(32'h3a95d784),
	.w2(32'hbb253c02),
	.w3(32'h3b0a5bb8),
	.w4(32'hbc0006c1),
	.w5(32'hbb8051b8),
	.w6(32'h3bb4e87f),
	.w7(32'h3aa3df5a),
	.w8(32'h3b84b7bf),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f794),
	.w1(32'h3b8d6b45),
	.w2(32'hbbbec5fd),
	.w3(32'h3a619daf),
	.w4(32'hbc3e4331),
	.w5(32'h3bb03777),
	.w6(32'hbc079ed9),
	.w7(32'hb9a3a4bf),
	.w8(32'h3c1f31f3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc120afd),
	.w1(32'h3bc44825),
	.w2(32'hbb084afa),
	.w3(32'hba193fda),
	.w4(32'hbbf46311),
	.w5(32'h3b65a39f),
	.w6(32'hb956d808),
	.w7(32'h3b30b023),
	.w8(32'hbbad1bc6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db4b2c),
	.w1(32'hba8d1a82),
	.w2(32'h3b83c9af),
	.w3(32'h3bd4fc28),
	.w4(32'hbbbab5f2),
	.w5(32'hbb4da858),
	.w6(32'h3c04e01c),
	.w7(32'hbc4f2ffe),
	.w8(32'hbcbebdb0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe306f),
	.w1(32'hbc141684),
	.w2(32'hbc826911),
	.w3(32'hbb97b413),
	.w4(32'hbb890050),
	.w5(32'h3a518140),
	.w6(32'hbc052a0e),
	.w7(32'hbc36b7fb),
	.w8(32'h3b7d98ff),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c4d36),
	.w1(32'hbb539ee7),
	.w2(32'hbc2fe3ec),
	.w3(32'h3c0d44b6),
	.w4(32'h3aa0b823),
	.w5(32'h3be59241),
	.w6(32'hbb4aacf4),
	.w7(32'hbc0b6d6f),
	.w8(32'hbb89e8e5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe8370),
	.w1(32'hbbe2196f),
	.w2(32'hbc3ed905),
	.w3(32'h3ad06c18),
	.w4(32'hbc8939af),
	.w5(32'h3cd4fd84),
	.w6(32'h3c5f357d),
	.w7(32'h3a0a0cc7),
	.w8(32'h3c755dc6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e72e6),
	.w1(32'h3aa2eb3d),
	.w2(32'hbba8f68b),
	.w3(32'hbc27512d),
	.w4(32'hba681076),
	.w5(32'hbc3d5d9b),
	.w6(32'h3c4aae34),
	.w7(32'hba9d66f1),
	.w8(32'hbcdf7e50),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule