module layer_10_featuremap_160(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcae6b),
	.w1(32'h3977e8a8),
	.w2(32'hb91aaf06),
	.w3(32'h3a018b5c),
	.w4(32'hb8a43764),
	.w5(32'hb9a7a7e5),
	.w6(32'h3a0f40fe),
	.w7(32'h3a0cac1c),
	.w8(32'h3a6e7639),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8ad79),
	.w1(32'h3a78fd5b),
	.w2(32'hb9e1fd4c),
	.w3(32'h3ae94b7a),
	.w4(32'h3ab9faeb),
	.w5(32'h374c1402),
	.w6(32'h3b26d401),
	.w7(32'h3ab6192a),
	.w8(32'h3aa6a621),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f225bf),
	.w1(32'h3a056bb2),
	.w2(32'h39d92140),
	.w3(32'h39dc16cb),
	.w4(32'h3a0e80bb),
	.w5(32'h39f9ab9e),
	.w6(32'h3a13f61a),
	.w7(32'h39d53883),
	.w8(32'h39ed95cf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29142d),
	.w1(32'h3a0f8b5c),
	.w2(32'h3997ce79),
	.w3(32'h3a0780a9),
	.w4(32'h39903934),
	.w5(32'h37409cba),
	.w6(32'hb90f909e),
	.w7(32'hba027a2c),
	.w8(32'hb9b14d35),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874520),
	.w1(32'hb9f7be67),
	.w2(32'hba22c94b),
	.w3(32'h39968ab8),
	.w4(32'hb964c337),
	.w5(32'hb989f3be),
	.w6(32'hb95a4796),
	.w7(32'hb83100cc),
	.w8(32'hb9a6644a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21f20b),
	.w1(32'h39dcfc76),
	.w2(32'h38e0135b),
	.w3(32'h39019bcf),
	.w4(32'h3a1faf6e),
	.w5(32'h3a09cfe9),
	.w6(32'h39fa45ce),
	.w7(32'h39dd08b6),
	.w8(32'h3a19bd05),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a61209),
	.w1(32'h3a84019b),
	.w2(32'h3b4b4625),
	.w3(32'h39408d19),
	.w4(32'h39b47a88),
	.w5(32'h3b17fae3),
	.w6(32'h39e61c1f),
	.w7(32'h3a4c86c6),
	.w8(32'h3b1b26dd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99795df),
	.w1(32'h39dc46c3),
	.w2(32'h3bbe0b2b),
	.w3(32'h3848d213),
	.w4(32'hba6373a6),
	.w5(32'h3a228897),
	.w6(32'h3a82724f),
	.w7(32'h39d3f496),
	.w8(32'h3994540f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b01e87),
	.w1(32'hb9d70863),
	.w2(32'hba4e7674),
	.w3(32'h3a214a5b),
	.w4(32'h380d75d6),
	.w5(32'hb9ed1f0d),
	.w6(32'h3a501f2d),
	.w7(32'h39d3214a),
	.w8(32'hb9416cf3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb7433),
	.w1(32'h3b46399f),
	.w2(32'h3b97c6f4),
	.w3(32'h3b879ac2),
	.w4(32'h39a54fad),
	.w5(32'h3b32f45d),
	.w6(32'h3ba2cfd9),
	.w7(32'hb93a9071),
	.w8(32'h3a124ae8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14f3f3),
	.w1(32'h38095e88),
	.w2(32'hb99cbbfd),
	.w3(32'hb9c61abe),
	.w4(32'h3a132fa3),
	.w5(32'hba1490c1),
	.w6(32'h395cb1bd),
	.w7(32'h3946d542),
	.w8(32'hba0d54b4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a882cf3),
	.w1(32'hbb54a23b),
	.w2(32'hb8aaa2ff),
	.w3(32'h3a58cabe),
	.w4(32'hbb6cae47),
	.w5(32'hba906301),
	.w6(32'h3af424f4),
	.w7(32'hbaf055ff),
	.w8(32'h3a32a1bd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54dd7c),
	.w1(32'h3af5f771),
	.w2(32'h3bb53136),
	.w3(32'h3a9b55a1),
	.w4(32'hba8e5740),
	.w5(32'h3b7b8ad6),
	.w6(32'h3ac660af),
	.w7(32'hbb11d343),
	.w8(32'h3a6c38d3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab472e0),
	.w1(32'hb9c3dc96),
	.w2(32'hba8ba017),
	.w3(32'h3aaf26e7),
	.w4(32'hb88a6862),
	.w5(32'hba840c61),
	.w6(32'h3b561a69),
	.w7(32'h38a4bccb),
	.w8(32'hb9279477),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398c81),
	.w1(32'h3a8f5658),
	.w2(32'h3ae51076),
	.w3(32'h3b11482d),
	.w4(32'h38bb894d),
	.w5(32'h39a6d00c),
	.w6(32'h3b16c134),
	.w7(32'h38840779),
	.w8(32'h38aef11f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a84c9),
	.w1(32'h3b3302b1),
	.w2(32'h3acb1edf),
	.w3(32'h3b3ddb9d),
	.w4(32'h3a636459),
	.w5(32'h3a40bd94),
	.w6(32'h3b69010d),
	.w7(32'h39cfc6ab),
	.w8(32'hb9647345),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2907b6),
	.w1(32'h39735f27),
	.w2(32'hb9247ec2),
	.w3(32'h3a726a1c),
	.w4(32'h3a80d60b),
	.w5(32'h39629810),
	.w6(32'h3935eee8),
	.w7(32'h3a5bd064),
	.w8(32'h39f8ac24),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253e96),
	.w1(32'h3b2a42fa),
	.w2(32'h3bc71dd1),
	.w3(32'h3a839d6a),
	.w4(32'h39f621ad),
	.w5(32'h3b50d769),
	.w6(32'h3b3175b3),
	.w7(32'hb7051613),
	.w8(32'h3aac89be),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00f88),
	.w1(32'h3a8bc515),
	.w2(32'h3b67e122),
	.w3(32'h3a594a4d),
	.w4(32'hba1566d2),
	.w5(32'h3b1aa8d4),
	.w6(32'h3af321e7),
	.w7(32'hba7e9861),
	.w8(32'h39fa6f81),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393930b7),
	.w1(32'h39245730),
	.w2(32'h391e7853),
	.w3(32'h3849dc03),
	.w4(32'h39618a80),
	.w5(32'h393caf70),
	.w6(32'h39643018),
	.w7(32'h39a216f6),
	.w8(32'h393dc6ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39314a2d),
	.w1(32'hb8a0828d),
	.w2(32'hb9b659f5),
	.w3(32'h38d7ab3a),
	.w4(32'hb8ba1caf),
	.w5(32'hb995b653),
	.w6(32'hb9949739),
	.w7(32'hb9c45b87),
	.w8(32'hb9781146),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9948f74),
	.w1(32'hb89e4503),
	.w2(32'h3a91080d),
	.w3(32'hb9f4e379),
	.w4(32'hb9bc4ca5),
	.w5(32'hba124506),
	.w6(32'h3a484052),
	.w7(32'h396c7af5),
	.w8(32'h3abe3e35),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aab52),
	.w1(32'h3b2515c6),
	.w2(32'hb9ea5f19),
	.w3(32'h3c07fbe8),
	.w4(32'h3b327328),
	.w5(32'h3b0e8087),
	.w6(32'h3c2c4220),
	.w7(32'h3b677aec),
	.w8(32'h3b58846e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35512c),
	.w1(32'h3b007cee),
	.w2(32'h3b4339e6),
	.w3(32'h3afc71c9),
	.w4(32'h39ab5e7e),
	.w5(32'h3a9c9124),
	.w6(32'h3b92c469),
	.w7(32'h39d8cb3c),
	.w8(32'h3a49c186),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7591e0),
	.w1(32'hba99e978),
	.w2(32'hbad1543c),
	.w3(32'h3b4eac58),
	.w4(32'hbb012d4b),
	.w5(32'hbb3dd214),
	.w6(32'h3b8032c9),
	.w7(32'hbad39ece),
	.w8(32'hbb03a7df),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cb031),
	.w1(32'hb87c238a),
	.w2(32'h399e89eb),
	.w3(32'h3a194f4b),
	.w4(32'h391f2e1e),
	.w5(32'h3a2cdf1e),
	.w6(32'hb9755282),
	.w7(32'h37ace34b),
	.w8(32'h391e48fa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dc748),
	.w1(32'h392240b9),
	.w2(32'h38f544e0),
	.w3(32'hb9d81266),
	.w4(32'h390134ef),
	.w5(32'h38af7f07),
	.w6(32'h383f238a),
	.w7(32'h39634437),
	.w8(32'h38fb766c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063613),
	.w1(32'h3a5c875a),
	.w2(32'hba0d50c6),
	.w3(32'h3af7e417),
	.w4(32'hba178823),
	.w5(32'hbafae385),
	.w6(32'h3b1ca9b5),
	.w7(32'hb9376a15),
	.w8(32'hbabda84f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07aed9),
	.w1(32'hba99778b),
	.w2(32'hba78f4ff),
	.w3(32'h3b0ac2ff),
	.w4(32'hba7de517),
	.w5(32'hbaa1c560),
	.w6(32'h3b1d725f),
	.w7(32'hb93a59c1),
	.w8(32'h38e930a8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba247e6),
	.w1(32'h3b3324a6),
	.w2(32'h3a768c8c),
	.w3(32'h3b81b7a7),
	.w4(32'h3a55c6fc),
	.w5(32'h3912aefc),
	.w6(32'h3b790ae4),
	.w7(32'h393c8d51),
	.w8(32'hba59070e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d49ea),
	.w1(32'h396b0a6e),
	.w2(32'h35d4f412),
	.w3(32'hb9d2fd33),
	.w4(32'h39770cf7),
	.w5(32'h38aff9bd),
	.w6(32'h3914f7b5),
	.w7(32'h38bf6381),
	.w8(32'h3895f9a0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901213d),
	.w1(32'hb918aefe),
	.w2(32'hb9818e62),
	.w3(32'h37e2c2c8),
	.w4(32'h38d0244c),
	.w5(32'hb82db2a4),
	.w6(32'hb6b75d99),
	.w7(32'h38cf6266),
	.w8(32'hb7c9e299),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a88a32),
	.w1(32'h3a6a727f),
	.w2(32'h3af97db1),
	.w3(32'h39817f60),
	.w4(32'h3948eb76),
	.w5(32'h3a2087fe),
	.w6(32'h3ad04f85),
	.w7(32'h3a1cf772),
	.w8(32'h39a8a1ff),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fac97),
	.w1(32'hba32c4f7),
	.w2(32'hba5efa76),
	.w3(32'h3a75b158),
	.w4(32'hba2cc821),
	.w5(32'hbaa49c1d),
	.w6(32'h38f150ad),
	.w7(32'h38081b36),
	.w8(32'hb9199657),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391154e9),
	.w1(32'h39e605b0),
	.w2(32'h39e05f7d),
	.w3(32'h39c3fe6c),
	.w4(32'h39792f5f),
	.w5(32'h39663dba),
	.w6(32'h399de717),
	.w7(32'h393160f6),
	.w8(32'h38e4e0c1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e5de8),
	.w1(32'hb8532379),
	.w2(32'h3afe1aff),
	.w3(32'hba1f6f6a),
	.w4(32'hba33ce28),
	.w5(32'h3a9652fd),
	.w6(32'hb89d0372),
	.w7(32'hba7fc895),
	.w8(32'h3a6cd112),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76c06d),
	.w1(32'h3ac05e2e),
	.w2(32'h3b5c9ee2),
	.w3(32'h3a7550cc),
	.w4(32'hba296ba6),
	.w5(32'h3a8f80b1),
	.w6(32'h3adedba7),
	.w7(32'h3984f272),
	.w8(32'h3a74992a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3040a5),
	.w1(32'hbb867f61),
	.w2(32'hbbed04f3),
	.w3(32'h3c438913),
	.w4(32'h3994f624),
	.w5(32'hbb716f93),
	.w6(32'h3c767597),
	.w7(32'h3b4e7cce),
	.w8(32'h3b296b3a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e42a5),
	.w1(32'hba2211c7),
	.w2(32'hbbd01b31),
	.w3(32'h3c18fb8b),
	.w4(32'h3a8a6097),
	.w5(32'hbb1407d4),
	.w6(32'h3c31dfd1),
	.w7(32'h3b6ff72f),
	.w8(32'h3b6c3dda),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfe96a),
	.w1(32'hb99440f3),
	.w2(32'hba510e26),
	.w3(32'h3aec0867),
	.w4(32'hb884454e),
	.w5(32'hba4273df),
	.w6(32'h3b0eba74),
	.w7(32'h3a0a4854),
	.w8(32'h388f2529),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cceb41),
	.w1(32'hb9035db9),
	.w2(32'hb89b2390),
	.w3(32'h390002ec),
	.w4(32'hb9804d35),
	.w5(32'hb961660f),
	.w6(32'hb9922a6e),
	.w7(32'hb921498a),
	.w8(32'hb8e3f3c0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85829e8),
	.w1(32'h3a38d192),
	.w2(32'h3a008846),
	.w3(32'hb98920f9),
	.w4(32'h3a5744c1),
	.w5(32'h3a1c700b),
	.w6(32'h39fbdc3d),
	.w7(32'h3976f983),
	.w8(32'h39a4096e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b887f58),
	.w1(32'hb90054af),
	.w2(32'hba4e602a),
	.w3(32'h3babe0d2),
	.w4(32'h3abdccdc),
	.w5(32'h3a663a51),
	.w6(32'h3b568c28),
	.w7(32'h3ab100f5),
	.w8(32'h3984c4ee),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be501c7),
	.w1(32'h3ba01e1c),
	.w2(32'h3b2b6601),
	.w3(32'h3bb25b5a),
	.w4(32'h3b3a41e8),
	.w5(32'h3a8e0fba),
	.w6(32'h3bf381bd),
	.w7(32'h3ae506ec),
	.w8(32'hb8bb98ec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b656946),
	.w1(32'h3aa70327),
	.w2(32'h3afcbe86),
	.w3(32'h3b15eeab),
	.w4(32'hba2e2017),
	.w5(32'hb822410d),
	.w6(32'h3b8d33ba),
	.w7(32'hb999ec82),
	.w8(32'hb83a225d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932737),
	.w1(32'h3b2419c6),
	.w2(32'h3b779ed7),
	.w3(32'h3b286109),
	.w4(32'hba2a873b),
	.w5(32'h3a33e9b7),
	.w6(32'h3ba36fc1),
	.w7(32'hb9b13935),
	.w8(32'h39e9a91a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67e463),
	.w1(32'hba13e554),
	.w2(32'hb8cd02b8),
	.w3(32'h3b786f76),
	.w4(32'hb9d9fe3c),
	.w5(32'hb9a78419),
	.w6(32'h3b896dd3),
	.w7(32'hb896307f),
	.w8(32'hb71c6f79),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec04a),
	.w1(32'h3aa753da),
	.w2(32'h3b9dd0e2),
	.w3(32'h3ab7dd82),
	.w4(32'h3a0fc012),
	.w5(32'h3b581cbe),
	.w6(32'h3a823ae6),
	.w7(32'hb91f8512),
	.w8(32'h3a672c43),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a79a53),
	.w1(32'hb885db3c),
	.w2(32'hb871acd9),
	.w3(32'h38ad2db6),
	.w4(32'hb6854388),
	.w5(32'hb90690b6),
	.w6(32'hb9782a55),
	.w7(32'hb8dda1b1),
	.w8(32'hb9b55ab2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91af084),
	.w1(32'h39749ec9),
	.w2(32'hb99a015b),
	.w3(32'hb97bafd3),
	.w4(32'h392cd2da),
	.w5(32'hb8957bf1),
	.w6(32'h396ae90b),
	.w7(32'hb91c3bd8),
	.w8(32'hb9ad298d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8c8b4),
	.w1(32'h3a3b068c),
	.w2(32'h39be469e),
	.w3(32'h3a1d027c),
	.w4(32'h3a082b50),
	.w5(32'h393059a7),
	.w6(32'h3a134cff),
	.w7(32'h38703ac9),
	.w8(32'hb89bc710),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26622f),
	.w1(32'h3aaeffa3),
	.w2(32'h3b700242),
	.w3(32'h3a93f857),
	.w4(32'hb98f0f97),
	.w5(32'h3a322166),
	.w6(32'h3a7b1e47),
	.w7(32'hb9fba337),
	.w8(32'hba018bd1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4edb2),
	.w1(32'h3a63e42e),
	.w2(32'h3a1feef0),
	.w3(32'h3a70aaab),
	.w4(32'h3a4c984c),
	.w5(32'h3a44632d),
	.w6(32'h3a8986cc),
	.w7(32'h3a163adc),
	.w8(32'h3a541b66),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b711897),
	.w1(32'h3b1243b6),
	.w2(32'h3bb882d9),
	.w3(32'h3ada68b8),
	.w4(32'hba071d35),
	.w5(32'h3b3e836f),
	.w6(32'h3b14b54e),
	.w7(32'hba529701),
	.w8(32'h3aa974be),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862a7b2),
	.w1(32'hb9ab7a7a),
	.w2(32'hba360d71),
	.w3(32'h3a1826cf),
	.w4(32'hb9c63cc5),
	.w5(32'hb99d199b),
	.w6(32'h3a985c4a),
	.w7(32'h3a2bc59b),
	.w8(32'h39bc9f4b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399943f8),
	.w1(32'h38f3045e),
	.w2(32'h391a68d4),
	.w3(32'hb88c5eb1),
	.w4(32'h398e0a33),
	.w5(32'h39512e01),
	.w6(32'hb903050f),
	.w7(32'hb9596c0d),
	.w8(32'h3768e5c4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c09cf9),
	.w1(32'h3a2a2480),
	.w2(32'h39c8c87e),
	.w3(32'hb69660c5),
	.w4(32'h3a456247),
	.w5(32'h3a01d32b),
	.w6(32'h3a26b5d6),
	.w7(32'h3a53481a),
	.w8(32'h3a5b7ef3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6bfb),
	.w1(32'hb875eee3),
	.w2(32'hb96c4332),
	.w3(32'h3a2b626b),
	.w4(32'hb83e8777),
	.w5(32'h38a26e4a),
	.w6(32'hb8678b27),
	.w7(32'h38818e9f),
	.w8(32'h3981447e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2661c6),
	.w1(32'h39bb8c01),
	.w2(32'h39c1b6c3),
	.w3(32'h3abb14ef),
	.w4(32'h3a389fd4),
	.w5(32'h39cdade2),
	.w6(32'h3ada62f8),
	.w7(32'h3a72153c),
	.w8(32'h3a33c97a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c2137),
	.w1(32'h3a130da6),
	.w2(32'h39a73dd1),
	.w3(32'h3a1d7751),
	.w4(32'h3a65a05d),
	.w5(32'h3a35ab4a),
	.w6(32'h3a2797eb),
	.w7(32'h3a6dfb4d),
	.w8(32'h3a121e26),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf9791),
	.w1(32'h39774c41),
	.w2(32'h3b138394),
	.w3(32'h3a86e8b9),
	.w4(32'hba3f0274),
	.w5(32'h39c83a72),
	.w6(32'h3ab7ed66),
	.w7(32'hbab85479),
	.w8(32'hb9fa1c83),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264a87),
	.w1(32'h3aea60cd),
	.w2(32'h3aaf6232),
	.w3(32'h3af57299),
	.w4(32'h3a7d445e),
	.w5(32'h3ada3ce3),
	.w6(32'h3af3baa0),
	.w7(32'h3a857e2f),
	.w8(32'h3a5276cf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a5d76),
	.w1(32'h3910fc1b),
	.w2(32'h39bcce94),
	.w3(32'h3991a1a5),
	.w4(32'h37ee5fd2),
	.w5(32'h38c5d49f),
	.w6(32'h39ae50b0),
	.w7(32'h39d40f4e),
	.w8(32'h3a448317),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a171f82),
	.w1(32'h39af7208),
	.w2(32'h38cd2cfc),
	.w3(32'h39c2b9ca),
	.w4(32'h3909ad9d),
	.w5(32'hb926f5a8),
	.w6(32'h390caaf9),
	.w7(32'h37432a79),
	.w8(32'hb880f047),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915d368),
	.w1(32'h38be9e49),
	.w2(32'h38eadfc0),
	.w3(32'hb9a76b0b),
	.w4(32'h379b7a5e),
	.w5(32'h3739797b),
	.w6(32'h37c0682a),
	.w7(32'h397104f1),
	.w8(32'h386764d7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8906d32),
	.w1(32'hb9ab51fc),
	.w2(32'hb880b844),
	.w3(32'hb8b6fd6c),
	.w4(32'hb93891dc),
	.w5(32'hb93010fd),
	.w6(32'hba1b4967),
	.w7(32'hb928f026),
	.w8(32'h3a0a00f2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f36cfd),
	.w1(32'h3a86e7d1),
	.w2(32'h3b3cda21),
	.w3(32'h3a073082),
	.w4(32'hba860082),
	.w5(32'h3a429310),
	.w6(32'h3a7d57fb),
	.w7(32'h39f2bbd3),
	.w8(32'h3a94aa1a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd2ba),
	.w1(32'hbae3a549),
	.w2(32'h39c84ef5),
	.w3(32'h3a499be1),
	.w4(32'hbb2949b7),
	.w5(32'hb7ef4b0b),
	.w6(32'h3b5bc495),
	.w7(32'hb9e9261a),
	.w8(32'h3a357c9e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e2c41),
	.w1(32'hbab08028),
	.w2(32'hbb03e291),
	.w3(32'h3a5ed112),
	.w4(32'hbb266e01),
	.w5(32'hbb4f3266),
	.w6(32'h3b7a44d9),
	.w7(32'h399eeeff),
	.w8(32'hba2bf1cb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55abae),
	.w1(32'hbbe714b6),
	.w2(32'hbb3d8377),
	.w3(32'h3b266df4),
	.w4(32'hbbe762c5),
	.w5(32'hbc0d8b0f),
	.w6(32'h3b9b1b87),
	.w7(32'hbb7c2678),
	.w8(32'hbb788d0a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2a5a9),
	.w1(32'h3a38db16),
	.w2(32'h39ded5fd),
	.w3(32'hb8ad9677),
	.w4(32'h39f1eecd),
	.w5(32'h3992ec90),
	.w6(32'h3a0ea862),
	.w7(32'h3a188575),
	.w8(32'h39acf6a7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39504af5),
	.w1(32'h38f68fd8),
	.w2(32'h385217a4),
	.w3(32'h38365e84),
	.w4(32'h39a2e672),
	.w5(32'h3992d91c),
	.w6(32'hb822131f),
	.w7(32'h3862ab86),
	.w8(32'h39a14ed9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390faf05),
	.w1(32'h39c12eea),
	.w2(32'h398d0602),
	.w3(32'h38efebbe),
	.w4(32'h39e9379d),
	.w5(32'h39e47ca6),
	.w6(32'h392b440b),
	.w7(32'h3971355a),
	.w8(32'h39a8383d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a29147),
	.w1(32'hb91a2652),
	.w2(32'hb86a0500),
	.w3(32'h39aee4d5),
	.w4(32'hba01513f),
	.w5(32'h392855c7),
	.w6(32'h3a0bc632),
	.w7(32'hb8e1085c),
	.w8(32'h382a947b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978c978),
	.w1(32'h39e8046f),
	.w2(32'h39d3f27a),
	.w3(32'hb90fdc68),
	.w4(32'h3a1a7644),
	.w5(32'h3a0b3a4f),
	.w6(32'h39c6abe2),
	.w7(32'h39a92162),
	.w8(32'h396c3225),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7640),
	.w1(32'h399ca9c1),
	.w2(32'h3b7ca499),
	.w3(32'h3a11ae72),
	.w4(32'hb9ae1d01),
	.w5(32'h3acfe105),
	.w6(32'h39e0baba),
	.w7(32'hba56c657),
	.w8(32'hba0fe4d4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3938),
	.w1(32'hb97bf70f),
	.w2(32'h3a7818b4),
	.w3(32'h3b3c649b),
	.w4(32'hb9f60c30),
	.w5(32'hbb1f0ab5),
	.w6(32'h3b7bb543),
	.w7(32'hb9e6d4a1),
	.w8(32'hba896648),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77a386),
	.w1(32'h3ad9c6e5),
	.w2(32'h3b431a9f),
	.w3(32'h3b094335),
	.w4(32'hb99040bd),
	.w5(32'h3a2753e5),
	.w6(32'h3b18b93f),
	.w7(32'hba2b355e),
	.w8(32'hb9f5f2a8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6ee80),
	.w1(32'hba275791),
	.w2(32'h394d0b22),
	.w3(32'h3a7287fc),
	.w4(32'hba946adc),
	.w5(32'hb71c261d),
	.w6(32'h3af19c46),
	.w7(32'hb7f25269),
	.w8(32'hb863661f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0653d),
	.w1(32'h397840d2),
	.w2(32'h3aed44e4),
	.w3(32'hba46cbbf),
	.w4(32'hba5b6385),
	.w5(32'h3aa4c00b),
	.w6(32'h390122fe),
	.w7(32'hba4c2f39),
	.w8(32'h3a4f587c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace0708),
	.w1(32'h3a34ef5c),
	.w2(32'h38d1859f),
	.w3(32'h3a8f2548),
	.w4(32'hb8d08ba6),
	.w5(32'hb904dfd1),
	.w6(32'h3a8fb340),
	.w7(32'hb8ffd5d0),
	.w8(32'hba3c271a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a313669),
	.w1(32'h3b1d5aac),
	.w2(32'h3b8301fc),
	.w3(32'h3901131f),
	.w4(32'h3aaaf3f5),
	.w5(32'h3b738a8b),
	.w6(32'h3aa8c170),
	.w7(32'h3a266231),
	.w8(32'h3ae05933),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de6c34),
	.w1(32'h3783f986),
	.w2(32'hb94b426f),
	.w3(32'h3a133fc2),
	.w4(32'h3923db04),
	.w5(32'h389c7460),
	.w6(32'h38df5aa9),
	.w7(32'hb8d5934c),
	.w8(32'hb8942258),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d216f6),
	.w1(32'h39e00d08),
	.w2(32'h399ee2c4),
	.w3(32'h378f0b6f),
	.w4(32'h39a35b52),
	.w5(32'h39313398),
	.w6(32'h3a08cf68),
	.w7(32'h39f56dc6),
	.w8(32'h39c50c02),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396074b9),
	.w1(32'hb9bbdf7b),
	.w2(32'hb9821c47),
	.w3(32'h390f2e4f),
	.w4(32'hb9f67cc2),
	.w5(32'hb9ae6be9),
	.w6(32'hb9a5e254),
	.w7(32'hb9303e94),
	.w8(32'hb804832e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ac5cb),
	.w1(32'h3999c874),
	.w2(32'h38cc422a),
	.w3(32'hb94745ec),
	.w4(32'h3945bf74),
	.w5(32'h3907865c),
	.w6(32'h399dc5e5),
	.w7(32'h399416e6),
	.w8(32'h39915508),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cf441),
	.w1(32'hba01e72a),
	.w2(32'hbad367d1),
	.w3(32'h3b52cc7a),
	.w4(32'h3a657b84),
	.w5(32'hba5214b5),
	.w6(32'h3b5f2b5e),
	.w7(32'h3a0db0a4),
	.w8(32'h3a815de6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd3eb4),
	.w1(32'h385ab816),
	.w2(32'hb944ead3),
	.w3(32'hb992ffb1),
	.w4(32'hb9f9f0b1),
	.w5(32'hb9d26ba7),
	.w6(32'h38940315),
	.w7(32'h39800946),
	.w8(32'h3a026981),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc281e),
	.w1(32'h3afe99f4),
	.w2(32'h3b597022),
	.w3(32'h3a3a3ab3),
	.w4(32'h3abe8055),
	.w5(32'h3b113912),
	.w6(32'h3ac857f9),
	.w7(32'h3a859129),
	.w8(32'h3abf84d0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b988af1),
	.w1(32'h3b287ba2),
	.w2(32'h3a9f6b45),
	.w3(32'h3baff293),
	.w4(32'h3aff7929),
	.w5(32'hba8a0cd6),
	.w6(32'h3bb6b858),
	.w7(32'h3b5876b8),
	.w8(32'h3938cd01),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5726bc),
	.w1(32'hba39eec6),
	.w2(32'hbb18cb9f),
	.w3(32'h3b329280),
	.w4(32'hba1888b7),
	.w5(32'hbaf84715),
	.w6(32'h3b6a471f),
	.w7(32'h3a5c6f40),
	.w8(32'h3956eba2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf734a),
	.w1(32'hb885eae9),
	.w2(32'hba97f591),
	.w3(32'h3aa9eaad),
	.w4(32'hbadeb5f7),
	.w5(32'hbac23eda),
	.w6(32'h3b688dbc),
	.w7(32'h3b543a4a),
	.w8(32'h3b31b31e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b04b77),
	.w1(32'hba468107),
	.w2(32'hbadd1ae0),
	.w3(32'hbac10b4b),
	.w4(32'hbac8884c),
	.w5(32'hbb08e6c4),
	.w6(32'h3a3a79e6),
	.w7(32'hba93105f),
	.w8(32'hbaa3f160),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b045a2c),
	.w1(32'hbb2aecde),
	.w2(32'hbb365794),
	.w3(32'h3aaed958),
	.w4(32'hbb28e62d),
	.w5(32'hbb4558dd),
	.w6(32'h3b7af38b),
	.w7(32'hba16d120),
	.w8(32'hbad2f2d6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b168ad6),
	.w1(32'h3b047479),
	.w2(32'h3af6bed3),
	.w3(32'h3ac8a1ea),
	.w4(32'h3b0297e1),
	.w5(32'h3a83bf84),
	.w6(32'h3b21fed2),
	.w7(32'h3aba6a17),
	.w8(32'h3a7a61e3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b765455),
	.w1(32'h386c6f39),
	.w2(32'h3a521a43),
	.w3(32'h3b275895),
	.w4(32'hba8c82fa),
	.w5(32'hb8a2e04d),
	.w6(32'h3b968f16),
	.w7(32'h39adffe2),
	.w8(32'h3a2c7be7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9113318),
	.w1(32'hb9cf2518),
	.w2(32'hb773630a),
	.w3(32'hb920c2ea),
	.w4(32'hb9d02c51),
	.w5(32'hb8d36695),
	.w6(32'hba31b28b),
	.w7(32'hba2b1a92),
	.w8(32'hba082c66),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e3e9),
	.w1(32'h3b144079),
	.w2(32'h3b748eb2),
	.w3(32'h3b288a71),
	.w4(32'h38ccb9b9),
	.w5(32'h3a461e39),
	.w6(32'h3b7a09fa),
	.w7(32'hb9bde3c3),
	.w8(32'h39c532a9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87eb32),
	.w1(32'hb9149f99),
	.w2(32'h3a9447fa),
	.w3(32'h3a2058f0),
	.w4(32'hba76d816),
	.w5(32'hba1442f0),
	.w6(32'h3aff2c2c),
	.w7(32'h3a622b2d),
	.w8(32'h3a6b0c45),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c76c1b),
	.w1(32'h395caa68),
	.w2(32'h3b38d6a8),
	.w3(32'hba6a8980),
	.w4(32'hba99cbf7),
	.w5(32'h3a4bea87),
	.w6(32'hb95f5045),
	.w7(32'hba2f3377),
	.w8(32'h3b229bad),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7037f3),
	.w1(32'hbb92d0e9),
	.w2(32'hbbab8038),
	.w3(32'h3c8257a0),
	.w4(32'h3acd8340),
	.w5(32'hba06edee),
	.w6(32'h3c6cc258),
	.w7(32'h3b805b28),
	.w8(32'h3b849ccf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1836e),
	.w1(32'h3b7f8865),
	.w2(32'h3b971b9d),
	.w3(32'h3b714f9c),
	.w4(32'h3adb02be),
	.w5(32'h3afb24ab),
	.w6(32'h3b8789d5),
	.w7(32'h3a01372f),
	.w8(32'h3949de02),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa644eb),
	.w1(32'hba830fa2),
	.w2(32'hb9d97237),
	.w3(32'h3ad9b238),
	.w4(32'hbab17c8e),
	.w5(32'hb94cd6fe),
	.w6(32'h3aed3b36),
	.w7(32'hba080e02),
	.w8(32'h3a2ec4ab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606b8d),
	.w1(32'h3a4276c2),
	.w2(32'h39f2d3f3),
	.w3(32'h3a93ba82),
	.w4(32'h3a3031e3),
	.w5(32'h3a3cc6ab),
	.w6(32'hb8e8fea0),
	.w7(32'hb937daf7),
	.w8(32'hb9913456),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f1de3),
	.w1(32'hb908a9ff),
	.w2(32'h3bb48a34),
	.w3(32'hba12ac87),
	.w4(32'hbb2a35ce),
	.w5(32'h3b1c6ccc),
	.w6(32'h38eb6315),
	.w7(32'hbac559c8),
	.w8(32'h3a86ed56),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15bd6e),
	.w1(32'hba192191),
	.w2(32'hbb12ba08),
	.w3(32'h3a7c97d0),
	.w4(32'hba7c8fa4),
	.w5(32'hbb5e6f8c),
	.w6(32'h38da0dd1),
	.w7(32'hba260c84),
	.w8(32'hbb6276da),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a194b1),
	.w1(32'h39ce9102),
	.w2(32'h39ae761d),
	.w3(32'hb7173dda),
	.w4(32'h39ccfb4b),
	.w5(32'h39291ce3),
	.w6(32'h3a19b619),
	.w7(32'h3a042287),
	.w8(32'h399cddb6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a172306),
	.w1(32'h389c981e),
	.w2(32'h397bbb7f),
	.w3(32'h39e8935d),
	.w4(32'h396765a9),
	.w5(32'h39e2746d),
	.w6(32'h39796226),
	.w7(32'hb7ca62e8),
	.w8(32'h39ac5172),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b984cf1),
	.w1(32'h3b2f7c8d),
	.w2(32'h3ac5a9ee),
	.w3(32'h3b6f703d),
	.w4(32'h3ae34c34),
	.w5(32'h3a493f10),
	.w6(32'h3b86a0d8),
	.w7(32'h3a9be7b9),
	.w8(32'hba3917e7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a373),
	.w1(32'h3b0f70f1),
	.w2(32'h3b217a64),
	.w3(32'h3a9caa46),
	.w4(32'hb980041f),
	.w5(32'h39afd4bb),
	.w6(32'h3af2b1bc),
	.w7(32'hbaae7bad),
	.w8(32'hba9cd387),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59c5a8),
	.w1(32'h3aff6626),
	.w2(32'hb9cd6336),
	.w3(32'h3b6c8219),
	.w4(32'h3ae526a2),
	.w5(32'h3a331200),
	.w6(32'h3b8a391e),
	.w7(32'h3b48ba01),
	.w8(32'h3b068ca2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fd27f),
	.w1(32'hb8b79807),
	.w2(32'hb9deae4c),
	.w3(32'h3af280ee),
	.w4(32'h39c73bbe),
	.w5(32'hb8dacf75),
	.w6(32'h3ad63cd6),
	.w7(32'h3adade38),
	.w8(32'h3a30f32a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adef470),
	.w1(32'hbaced4de),
	.w2(32'hba8205eb),
	.w3(32'h3ac02ece),
	.w4(32'hba0e43aa),
	.w5(32'hb8b40f08),
	.w6(32'h3b57be08),
	.w7(32'h3a2019c4),
	.w8(32'h3a9c5ad1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac531c8),
	.w1(32'h3b1c5e03),
	.w2(32'h3b1a90ce),
	.w3(32'h39eda700),
	.w4(32'h3b0f867c),
	.w5(32'h3b26530e),
	.w6(32'h3a9a58ac),
	.w7(32'h3abb1841),
	.w8(32'h3a4f6a14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b475a50),
	.w1(32'h3a474aad),
	.w2(32'h38d9f248),
	.w3(32'h3b1f79cf),
	.w4(32'h392ed156),
	.w5(32'hb98ee6cf),
	.w6(32'h3b1d834d),
	.w7(32'h3a00bd33),
	.w8(32'hb9ce893a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba0511),
	.w1(32'h3881c9fb),
	.w2(32'hb8e03186),
	.w3(32'h398d17c0),
	.w4(32'h397d30d2),
	.w5(32'h389ab00f),
	.w6(32'h39406983),
	.w7(32'hb82493cc),
	.w8(32'h39a8d27c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395093c5),
	.w1(32'h39831256),
	.w2(32'h39099029),
	.w3(32'h39b1ab1b),
	.w4(32'h39a41d28),
	.w5(32'h39a11156),
	.w6(32'h398db90a),
	.w7(32'h3924f855),
	.w8(32'h39af5771),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39712d52),
	.w1(32'h38fe9d95),
	.w2(32'h389be4b1),
	.w3(32'h39e26a82),
	.w4(32'h39a8a682),
	.w5(32'h39ab1de2),
	.w6(32'h3985e7f5),
	.w7(32'h392c4b6a),
	.w8(32'h39b6aac5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381640bf),
	.w1(32'h39b3261b),
	.w2(32'hb62e0569),
	.w3(32'h3995acf9),
	.w4(32'h3823e4dc),
	.w5(32'hba112d47),
	.w6(32'h3a4623d6),
	.w7(32'h39cd8700),
	.w8(32'h39d5b727),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35c0d0),
	.w1(32'h3adc0ad9),
	.w2(32'h3b04c86c),
	.w3(32'h3ad1f4c0),
	.w4(32'h3996689b),
	.w5(32'h3a880363),
	.w6(32'h3b2990fa),
	.w7(32'h3916ebec),
	.w8(32'h387ce0c1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396018a1),
	.w1(32'hb85e78a0),
	.w2(32'hba26d1a5),
	.w3(32'h392fd3f8),
	.w4(32'h392bd34a),
	.w5(32'hb9d08800),
	.w6(32'h39f40113),
	.w7(32'h3985e5c8),
	.w8(32'hb9928689),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9d200),
	.w1(32'h396aa7c7),
	.w2(32'h3a9f79b4),
	.w3(32'h3900ae25),
	.w4(32'hb90060d8),
	.w5(32'hb883be16),
	.w6(32'h398d539d),
	.w7(32'h39195a2f),
	.w8(32'hb859126c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d7349),
	.w1(32'h3b2fb985),
	.w2(32'hbaa983e6),
	.w3(32'h3b534d50),
	.w4(32'h3b215589),
	.w5(32'hba4e788f),
	.w6(32'h3b90e7bb),
	.w7(32'h3b461e2c),
	.w8(32'h3af7804c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a720c2),
	.w1(32'h399d543c),
	.w2(32'h3a00c225),
	.w3(32'h39d25413),
	.w4(32'hb99d7d25),
	.w5(32'hba06d727),
	.w6(32'h390c5206),
	.w7(32'hb8ab1fec),
	.w8(32'h3947da7f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a21fb),
	.w1(32'h3a2a7a5c),
	.w2(32'h393295b5),
	.w3(32'hba163121),
	.w4(32'h3a53bb95),
	.w5(32'h3a1ae4c4),
	.w6(32'h3a6174eb),
	.w7(32'h3a843a5d),
	.w8(32'h3a918fdb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a26c9f),
	.w1(32'h391ea7f5),
	.w2(32'hb9468e8f),
	.w3(32'h3a288580),
	.w4(32'h390ff4f7),
	.w5(32'hb900d5de),
	.w6(32'h3919e03a),
	.w7(32'hb7376c86),
	.w8(32'hb85dda28),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa23df8),
	.w1(32'h3b06273c),
	.w2(32'hbbcb2ba4),
	.w3(32'h3a964191),
	.w4(32'h3b19249a),
	.w5(32'hbbe9ed2f),
	.w6(32'h3b635c4e),
	.w7(32'hbb0f44e1),
	.w8(32'hb9e3a74d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e9955b),
	.w1(32'h3ac4cd52),
	.w2(32'h3af5404f),
	.w3(32'h3a69f490),
	.w4(32'hba24bf30),
	.w5(32'hba074300),
	.w6(32'h39e399a1),
	.w7(32'h390ed5c3),
	.w8(32'hba771f86),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27fb7a),
	.w1(32'h3c297cc0),
	.w2(32'h3b834ddc),
	.w3(32'h38cf6858),
	.w4(32'hb9fbe6e3),
	.w5(32'h38019b3f),
	.w6(32'h3b3b6f83),
	.w7(32'hbb55e5ea),
	.w8(32'hbbc4ddeb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0614b),
	.w1(32'h3a7f2077),
	.w2(32'h3927d67c),
	.w3(32'hbbd8417f),
	.w4(32'h3b483a8b),
	.w5(32'h3b2ac46f),
	.w6(32'h3b09735d),
	.w7(32'h3a3d280a),
	.w8(32'h39d7adfd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af426b5),
	.w1(32'h39b810ec),
	.w2(32'h3b64a180),
	.w3(32'h3b39c628),
	.w4(32'h3afde7b2),
	.w5(32'h3ada80e3),
	.w6(32'h3b80c7fd),
	.w7(32'h3b1e8604),
	.w8(32'h3b5a0de1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45d5ed),
	.w1(32'h3b8f997f),
	.w2(32'h3c6621e8),
	.w3(32'h3a5281ef),
	.w4(32'hbadbf6e1),
	.w5(32'hbbc5d3b5),
	.w6(32'h3b679ec3),
	.w7(32'h3ae64fc3),
	.w8(32'h3b65c9e6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01f14d),
	.w1(32'hbb067506),
	.w2(32'h3b1ae148),
	.w3(32'hbc003e94),
	.w4(32'hbb89bcbb),
	.w5(32'hba0a68d2),
	.w6(32'hb9478396),
	.w7(32'h3bbdf282),
	.w8(32'hba38c066),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163601),
	.w1(32'h3a5118d8),
	.w2(32'hb9ca9f1f),
	.w3(32'hbb5af74c),
	.w4(32'h3aa141d0),
	.w5(32'h3ae82d64),
	.w6(32'hbb5ffc4b),
	.w7(32'hba50a23e),
	.w8(32'hbb040587),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab81c66),
	.w1(32'h3b0a4620),
	.w2(32'h3bd012ef),
	.w3(32'h3ab35090),
	.w4(32'h3ab4ba9d),
	.w5(32'h3b7f34e2),
	.w6(32'h3b65ea44),
	.w7(32'h3b12e002),
	.w8(32'h3b5155f6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce6d1),
	.w1(32'h3aa16962),
	.w2(32'hbacbdf15),
	.w3(32'h3b8de377),
	.w4(32'hba046626),
	.w5(32'hbb7b2ce0),
	.w6(32'h3a8c35ac),
	.w7(32'hba90187c),
	.w8(32'hbb2daed6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8686bd),
	.w1(32'h3ac5ea01),
	.w2(32'h3b01698a),
	.w3(32'hb8cec61a),
	.w4(32'h39d51510),
	.w5(32'hb9042b69),
	.w6(32'h3b89e9b2),
	.w7(32'hb9ef969f),
	.w8(32'h3aea72ae),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160ca8),
	.w1(32'hbb8d0cb6),
	.w2(32'h3b846b30),
	.w3(32'h3a6cf2e6),
	.w4(32'hbab1511c),
	.w5(32'h3bd78fd8),
	.w6(32'hbbf98e73),
	.w7(32'hbbc7d8b0),
	.w8(32'hbaad1e30),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9e92),
	.w1(32'hb9bbdbe3),
	.w2(32'hbbef1763),
	.w3(32'h3b94ccd3),
	.w4(32'hbb8004c7),
	.w5(32'hbc02835d),
	.w6(32'h3a8685f0),
	.w7(32'hba6fa991),
	.w8(32'h3b16a4e0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1c81),
	.w1(32'h3b62bfba),
	.w2(32'h3ae9905a),
	.w3(32'hbb2b3969),
	.w4(32'h3b009f15),
	.w5(32'hbb190ebd),
	.w6(32'h3ac5ffe3),
	.w7(32'hbb5fe3ca),
	.w8(32'hbaf62a54),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72c27c),
	.w1(32'h3b077b02),
	.w2(32'hbb5eb7e6),
	.w3(32'hba53a9f6),
	.w4(32'h3ac6185e),
	.w5(32'hba2ffdaa),
	.w6(32'h3b36129a),
	.w7(32'h38e56822),
	.w8(32'h3a93a5fd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb867c2),
	.w1(32'h3af72346),
	.w2(32'h3a0f5428),
	.w3(32'h3be2e2c1),
	.w4(32'hbaa46791),
	.w5(32'hb9d084e4),
	.w6(32'hbab86c3d),
	.w7(32'hbb14ed92),
	.w8(32'h3a368870),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae150),
	.w1(32'h3b33fa46),
	.w2(32'hbbe35a20),
	.w3(32'h3bf44188),
	.w4(32'hbb866f86),
	.w5(32'hbc1a4a1c),
	.w6(32'h3b5723fb),
	.w7(32'hbb41c783),
	.w8(32'hbba424a8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034323),
	.w1(32'h3b59b65c),
	.w2(32'h3ac833c8),
	.w3(32'hbb91d311),
	.w4(32'h3b402fb3),
	.w5(32'h39a7ea2f),
	.w6(32'h3b3cb503),
	.w7(32'h3aa4049a),
	.w8(32'h3aafa9c4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cb6c7),
	.w1(32'h3b1ad0e9),
	.w2(32'h3b7c2821),
	.w3(32'hb9244e8b),
	.w4(32'h3a2ab043),
	.w5(32'h3bc7a31b),
	.w6(32'hba8a1492),
	.w7(32'h3ab8425f),
	.w8(32'h3b875b0a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd64e7c),
	.w1(32'hbb78d5b5),
	.w2(32'hba7d80ba),
	.w3(32'h3c13801d),
	.w4(32'hb9c08e1b),
	.w5(32'hba5295eb),
	.w6(32'hb9aae7c8),
	.w7(32'hbac102f8),
	.w8(32'hbacc717c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05b249),
	.w1(32'hbb82e5bb),
	.w2(32'hbb468d3d),
	.w3(32'hbabe618d),
	.w4(32'hbb309ace),
	.w5(32'hbb7f9a16),
	.w6(32'h3b00796c),
	.w7(32'hba92454b),
	.w8(32'hbae5ba04),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34e67a),
	.w1(32'hbaa41d96),
	.w2(32'h3b2996bb),
	.w3(32'hbaac29c5),
	.w4(32'hbb2baa4c),
	.w5(32'h3a2e2713),
	.w6(32'h3b297f70),
	.w7(32'hbb843078),
	.w8(32'hba260ebc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a178501),
	.w1(32'h3a0b1426),
	.w2(32'hbb775754),
	.w3(32'hb9b6a544),
	.w4(32'h3a841109),
	.w5(32'hbbb89af7),
	.w6(32'h3aab8653),
	.w7(32'hbb12d982),
	.w8(32'h392050e4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60dad0),
	.w1(32'h3b96f536),
	.w2(32'h3b84825a),
	.w3(32'h39e4ce5e),
	.w4(32'hbb31a273),
	.w5(32'h39b37133),
	.w6(32'h3b95c3a9),
	.w7(32'hbb3d9c23),
	.w8(32'hbae23bd3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc4a73),
	.w1(32'hba88153a),
	.w2(32'h3c83e1c4),
	.w3(32'h3a05d79d),
	.w4(32'hb90369da),
	.w5(32'h3c5c5969),
	.w6(32'h3b09176e),
	.w7(32'h3c137775),
	.w8(32'hbbb0193e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba951316),
	.w1(32'h3a94b484),
	.w2(32'h3ade9fc7),
	.w3(32'hbbb2804b),
	.w4(32'hbad3736f),
	.w5(32'hb9863981),
	.w6(32'h39ea5afe),
	.w7(32'hba8c748a),
	.w8(32'h38b45aba),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810952),
	.w1(32'h3bb1716f),
	.w2(32'h3c3a7694),
	.w3(32'hba4fd4ff),
	.w4(32'h3b75895f),
	.w5(32'h3be4761e),
	.w6(32'h3b8a1cd4),
	.w7(32'h3b3b3bf1),
	.w8(32'h3b3139f9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77dcc),
	.w1(32'h3c01d56a),
	.w2(32'h3cb75b9e),
	.w3(32'h3bced120),
	.w4(32'h3c51905c),
	.w5(32'h3c772bf0),
	.w6(32'h39ab959e),
	.w7(32'hbbaeaa6c),
	.w8(32'h3b984629),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce065f6),
	.w1(32'hbb1aca81),
	.w2(32'hba92e603),
	.w3(32'h3c85149a),
	.w4(32'hba10bce4),
	.w5(32'h38c4818e),
	.w6(32'hbac82fb1),
	.w7(32'hbb3a3361),
	.w8(32'h39cb138a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804ea4),
	.w1(32'hbb06fa84),
	.w2(32'h3ab12727),
	.w3(32'h3b5266b5),
	.w4(32'h3a25b5b4),
	.w5(32'hba77c22b),
	.w6(32'h3b1f741c),
	.w7(32'hbb3a450c),
	.w8(32'hbaafbdaf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a4277),
	.w1(32'h3c0493a7),
	.w2(32'h3cb2b412),
	.w3(32'h3b1038cb),
	.w4(32'h3bec3a45),
	.w5(32'h3cca4584),
	.w6(32'h3c1bad61),
	.w7(32'h3c5d348d),
	.w8(32'h3be115df),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d77b2),
	.w1(32'h3be63428),
	.w2(32'h3a8939aa),
	.w3(32'h3bc51229),
	.w4(32'h3b93b1d2),
	.w5(32'hbb3c95e7),
	.w6(32'h3c0a4e3f),
	.w7(32'h3b93c400),
	.w8(32'h3bfa7810),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baea01d),
	.w1(32'h3a2c2f93),
	.w2(32'hbb34346c),
	.w3(32'h3b67f117),
	.w4(32'h3adf774d),
	.w5(32'hbb1f30f5),
	.w6(32'h3a3e5d41),
	.w7(32'hbac49997),
	.w8(32'h3a2bd9c2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f01ff),
	.w1(32'h3b33f87a),
	.w2(32'hbaec0042),
	.w3(32'hb949184d),
	.w4(32'h3b3a942b),
	.w5(32'hb9ccb23d),
	.w6(32'h3b583fff),
	.w7(32'h3ac24cd9),
	.w8(32'h3b28418c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64fc48),
	.w1(32'hba27d33b),
	.w2(32'h3c0ca425),
	.w3(32'h3b937ad3),
	.w4(32'h3b2d7c83),
	.w5(32'h3c5202cf),
	.w6(32'h3b4d3133),
	.w7(32'h3bec26a4),
	.w8(32'h3bbaafe4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9719),
	.w1(32'hbbb1dbe9),
	.w2(32'hbc66a00e),
	.w3(32'h3ba50a19),
	.w4(32'hbbdab075),
	.w5(32'hbc9bd170),
	.w6(32'hbb9f5482),
	.w7(32'hbc4c17e8),
	.w8(32'hbabdaa83),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf03b5),
	.w1(32'hba9d1e64),
	.w2(32'h3a0c8ae6),
	.w3(32'h3bf0d203),
	.w4(32'h3ac1dec0),
	.w5(32'h3886f495),
	.w6(32'hba8926cb),
	.w7(32'hbbba5bf3),
	.w8(32'hbb2237a5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b226e23),
	.w1(32'hb9126a02),
	.w2(32'hbb1a43fb),
	.w3(32'h3979202f),
	.w4(32'h3b120207),
	.w5(32'hba57289e),
	.w6(32'h3b08cfce),
	.w7(32'hba3e3ae4),
	.w8(32'h3ab9098a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d2377),
	.w1(32'hbb545b39),
	.w2(32'hb9a2fecc),
	.w3(32'hba4e2bb3),
	.w4(32'hbae01a9f),
	.w5(32'h38ba3663),
	.w6(32'h388143ad),
	.w7(32'hbb4aa79d),
	.w8(32'hbb1e2afd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a6fd),
	.w1(32'h3b0771f6),
	.w2(32'h3b1b2f25),
	.w3(32'hbacecd1a),
	.w4(32'h3b3f9a8c),
	.w5(32'h3b507812),
	.w6(32'h3b03bf78),
	.w7(32'h3b1a6a90),
	.w8(32'h3adde52b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf3aee),
	.w1(32'h3b10a75e),
	.w2(32'h3a115c56),
	.w3(32'h3b69b9b0),
	.w4(32'h3aa06476),
	.w5(32'hba8b21a7),
	.w6(32'h3ab0c619),
	.w7(32'h3b0d3596),
	.w8(32'h3a26d145),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dd217),
	.w1(32'h3a5afeeb),
	.w2(32'hbb46108c),
	.w3(32'h3b418c7e),
	.w4(32'h3a626667),
	.w5(32'hbb1a6545),
	.w6(32'h3baadfb6),
	.w7(32'h3b0c0372),
	.w8(32'hba651549),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82d632),
	.w1(32'h3c484a41),
	.w2(32'h3af5ce3d),
	.w3(32'h3b074dbf),
	.w4(32'h3be18712),
	.w5(32'hb9e8077e),
	.w6(32'h3c30c4d5),
	.w7(32'h3bcd0500),
	.w8(32'h3c0ebdc2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba79641),
	.w1(32'hb9b9bbfd),
	.w2(32'h3a1204bd),
	.w3(32'h3b2e3740),
	.w4(32'h3a012f49),
	.w5(32'hbb753f01),
	.w6(32'h3b316fdb),
	.w7(32'h392ed89f),
	.w8(32'h3b08d149),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817617),
	.w1(32'h3b41a9c6),
	.w2(32'h3aea73ad),
	.w3(32'hbb0bb64e),
	.w4(32'h3b659e59),
	.w5(32'h3b92f026),
	.w6(32'h3ba38649),
	.w7(32'h3b0fa219),
	.w8(32'h3b23a11b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819fe4),
	.w1(32'hbc196383),
	.w2(32'hbb42a3c7),
	.w3(32'h3bca6a07),
	.w4(32'hbbb0e292),
	.w5(32'h394f81f0),
	.w6(32'hbc9d6a5b),
	.w7(32'hbc4cf9b1),
	.w8(32'hbc0a0e6f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e493),
	.w1(32'h3a2ff3dd),
	.w2(32'h3b651290),
	.w3(32'h3bec2534),
	.w4(32'hbb62ec3e),
	.w5(32'h3adccc6c),
	.w6(32'h3b86a4f2),
	.w7(32'hba2d6f01),
	.w8(32'h3b1d76d1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05a000),
	.w1(32'h3a0c7977),
	.w2(32'h3b92d058),
	.w3(32'h3b01491c),
	.w4(32'hba060a08),
	.w5(32'h3a9173e9),
	.w6(32'h3b9190c2),
	.w7(32'h3aedf73f),
	.w8(32'h3af2fa64),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7e61),
	.w1(32'h3c38c420),
	.w2(32'h3c193a8a),
	.w3(32'h3a9a4823),
	.w4(32'h3b251980),
	.w5(32'hbaa8d373),
	.w6(32'h3ba3cda8),
	.w7(32'h3adb70c1),
	.w8(32'h3b13dc3c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2898f),
	.w1(32'h3bc311d7),
	.w2(32'h3a05c0b4),
	.w3(32'hbb75f366),
	.w4(32'h3bc4a600),
	.w5(32'h3b290e76),
	.w6(32'h3b8f27fe),
	.w7(32'hbb458ea4),
	.w8(32'h39f1689a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80d32),
	.w1(32'h3b0734fa),
	.w2(32'h3b52507b),
	.w3(32'hb9d643d1),
	.w4(32'h3b005566),
	.w5(32'h3b992ade),
	.w6(32'h3b3634c3),
	.w7(32'h3a5caa97),
	.w8(32'h3b5959bf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b468d89),
	.w1(32'h3a907c3d),
	.w2(32'h3ac4f0aa),
	.w3(32'h3b7895d4),
	.w4(32'hbaa63559),
	.w5(32'hb9b1076f),
	.w6(32'hbb0b83f0),
	.w7(32'hb9b267fb),
	.w8(32'hba70f52a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90473f),
	.w1(32'h3b8716ad),
	.w2(32'h3b9e6832),
	.w3(32'h3a0eb481),
	.w4(32'h3b5cc9bf),
	.w5(32'h3b68a79a),
	.w6(32'h3a515d35),
	.w7(32'h3afad9bc),
	.w8(32'h3b16d893),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9004ad),
	.w1(32'h3b7f5453),
	.w2(32'hbb1e7925),
	.w3(32'h3ba1c00f),
	.w4(32'hbb0ae8ba),
	.w5(32'hbb9e3e77),
	.w6(32'h3b880110),
	.w7(32'h3845375f),
	.w8(32'hbb3b7dd7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13f5e),
	.w1(32'h3b52b743),
	.w2(32'h3b9f23d2),
	.w3(32'hbb01fffd),
	.w4(32'h3b67f2c5),
	.w5(32'h3ba4b8c9),
	.w6(32'h3aa4bf94),
	.w7(32'h3a41c4e1),
	.w8(32'h39a94f27),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18f9b),
	.w1(32'hbb495fbd),
	.w2(32'hba86752d),
	.w3(32'h3b5ba147),
	.w4(32'hbafaff72),
	.w5(32'hba03e2a4),
	.w6(32'hbb332100),
	.w7(32'hba614735),
	.w8(32'hb95edd6d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24a410),
	.w1(32'h3b318f83),
	.w2(32'h3c1cee4b),
	.w3(32'h39eed278),
	.w4(32'h3be1e633),
	.w5(32'h3c57f39f),
	.w6(32'h3b61a8bb),
	.w7(32'h3bd6910f),
	.w8(32'h3c413a08),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4463),
	.w1(32'h3bf40b1f),
	.w2(32'h3bb737e4),
	.w3(32'h3c42ac69),
	.w4(32'hb9c20705),
	.w5(32'hbb75ca7e),
	.w6(32'h3bddea02),
	.w7(32'h3c5993ae),
	.w8(32'h3c2ae9f1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb3bc4),
	.w1(32'h3a6851cc),
	.w2(32'h39e3626f),
	.w3(32'hbb643ccd),
	.w4(32'h3ab98cbf),
	.w5(32'h3ad043d1),
	.w6(32'h3b806591),
	.w7(32'h399cb29b),
	.w8(32'h3b524ce9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c85d2),
	.w1(32'h3aa94aef),
	.w2(32'hbb1e89ca),
	.w3(32'h3bb1a061),
	.w4(32'h38a19d29),
	.w5(32'h3a6e7084),
	.w6(32'h38476655),
	.w7(32'hbb179be9),
	.w8(32'hbb92f23c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b28d),
	.w1(32'h3b198d44),
	.w2(32'h39536867),
	.w3(32'hb9b881c2),
	.w4(32'h3b4bf765),
	.w5(32'h39a43961),
	.w6(32'h3b3c0d82),
	.w7(32'h3931c860),
	.w8(32'hb9255b16),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb66d10),
	.w1(32'h3abc4af8),
	.w2(32'h3c2b2452),
	.w3(32'h3b939b94),
	.w4(32'hbb4498ce),
	.w5(32'h3b2afd8e),
	.w6(32'h3b76fdb8),
	.w7(32'hbbf71aef),
	.w8(32'hbb58c546),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d727),
	.w1(32'h3b04b3e5),
	.w2(32'hbad39da8),
	.w3(32'h3bbf310a),
	.w4(32'h3b6d4f32),
	.w5(32'hba87a38b),
	.w6(32'h3c1bdee8),
	.w7(32'h3ba15f1b),
	.w8(32'h3a9dda85),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d6ccb),
	.w1(32'h3ab17f75),
	.w2(32'hb963a4b2),
	.w3(32'hbb298fdb),
	.w4(32'hbaf5d0f3),
	.w5(32'hb9743346),
	.w6(32'hb9c85af7),
	.w7(32'h39905b4b),
	.w8(32'hb8fc0918),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e5679),
	.w1(32'hbb8899ec),
	.w2(32'h3a6615a0),
	.w3(32'h3a0057dc),
	.w4(32'hbb970810),
	.w5(32'h3a9cd0d2),
	.w6(32'h3a1a28d0),
	.w7(32'h3b276f96),
	.w8(32'hbb1f282e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d03a),
	.w1(32'hbbc7eb63),
	.w2(32'hbb27a3bd),
	.w3(32'hbb4db582),
	.w4(32'hbb424573),
	.w5(32'h398f3378),
	.w6(32'hbc49a324),
	.w7(32'hbc068a19),
	.w8(32'hbbb0f7d6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0a90),
	.w1(32'hbb9751a5),
	.w2(32'h399ec329),
	.w3(32'h3b2b1970),
	.w4(32'hba8ba978),
	.w5(32'h3b958033),
	.w6(32'hba6dda3f),
	.w7(32'h3b126e20),
	.w8(32'hba2af36c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb220eea),
	.w1(32'h3bca9056),
	.w2(32'h3b083c0e),
	.w3(32'hbaac21fd),
	.w4(32'h3ad5d609),
	.w5(32'hbb2f1811),
	.w6(32'h3b82ce13),
	.w7(32'h3b843ec0),
	.w8(32'hb88cad10),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8c97),
	.w1(32'h3bf46bfa),
	.w2(32'h3ab0d3a7),
	.w3(32'h3ba29f7d),
	.w4(32'h3bfcd529),
	.w5(32'h371f2796),
	.w6(32'h3c14d759),
	.w7(32'h3c022c16),
	.w8(32'h3bfdedeb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a359b),
	.w1(32'h3b621f7f),
	.w2(32'h3a30da77),
	.w3(32'hb928fdaa),
	.w4(32'h3ac7bc6a),
	.w5(32'hbb4c0b45),
	.w6(32'h3af2febc),
	.w7(32'hbb8314a6),
	.w8(32'h3a097218),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c181),
	.w1(32'h3ada3a7e),
	.w2(32'h3a6e6214),
	.w3(32'h3a183389),
	.w4(32'h3ae99133),
	.w5(32'h39e413f0),
	.w6(32'h3b2cd9a7),
	.w7(32'h3aab082b),
	.w8(32'h3a23628a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88be17),
	.w1(32'h39ba68a6),
	.w2(32'h3c14148e),
	.w3(32'h3b08f744),
	.w4(32'hbb0f3298),
	.w5(32'h3baef914),
	.w6(32'h3a2ae9c7),
	.w7(32'h3b351027),
	.w8(32'hbb175d80),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e4a9),
	.w1(32'hbb06512d),
	.w2(32'hbaed5886),
	.w3(32'h3b3eca74),
	.w4(32'h3a274d3b),
	.w5(32'hbaef3676),
	.w6(32'h39fa1ac6),
	.w7(32'hbb096745),
	.w8(32'hba933882),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4fd2),
	.w1(32'h3a860cd7),
	.w2(32'hba31909a),
	.w3(32'hba9261f4),
	.w4(32'h3ad1407a),
	.w5(32'hbae771d8),
	.w6(32'h3ab826a3),
	.w7(32'h3a850f0c),
	.w8(32'h3ac6d4b3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3d896),
	.w1(32'h3b047106),
	.w2(32'h3a4a4a1c),
	.w3(32'hba8d30b8),
	.w4(32'h3a3ce881),
	.w5(32'hba8db290),
	.w6(32'h3a742abe),
	.w7(32'h3ad79063),
	.w8(32'h3a29b0d3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91af2d2),
	.w1(32'h3a740578),
	.w2(32'hbac01c6a),
	.w3(32'hba9f7091),
	.w4(32'h3b4c91a6),
	.w5(32'h3aafec52),
	.w6(32'h3b117785),
	.w7(32'h3a86d2a1),
	.w8(32'h3b2c1835),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858f1d),
	.w1(32'hbaa63d67),
	.w2(32'hbba01702),
	.w3(32'h3b8e8e4f),
	.w4(32'hbac20864),
	.w5(32'hbb97924a),
	.w6(32'h3b6b07df),
	.w7(32'hbaace917),
	.w8(32'hbb48a512),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd7a3),
	.w1(32'h380aa96b),
	.w2(32'h3c5e7ef9),
	.w3(32'h3ae0aef6),
	.w4(32'h3bd8f1f5),
	.w5(32'hba9ad9f3),
	.w6(32'h3b04d544),
	.w7(32'hbb9d475f),
	.w8(32'h3be7c464),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc0f31),
	.w1(32'hbb3239f1),
	.w2(32'h3a02a87c),
	.w3(32'h3b18b399),
	.w4(32'hbb64fca7),
	.w5(32'hbabb8f1f),
	.w6(32'hbbb47044),
	.w7(32'hbb24674c),
	.w8(32'hbb809cea),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b937d5a),
	.w1(32'hbaf92d58),
	.w2(32'hbace0aed),
	.w3(32'h3b199a6c),
	.w4(32'hba9e199f),
	.w5(32'hbabc902d),
	.w6(32'h3b52f5a0),
	.w7(32'h3b208d54),
	.w8(32'hba0016c2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3758d),
	.w1(32'hba9850e3),
	.w2(32'h3ca3fba0),
	.w3(32'hba616a85),
	.w4(32'h3c1c7ef3),
	.w5(32'h3cc4ba67),
	.w6(32'h3af1a0d0),
	.w7(32'h3ba9ce0c),
	.w8(32'h3c4b0085),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9644f7),
	.w1(32'h3afc3dee),
	.w2(32'hbb44892f),
	.w3(32'h3c7ecc93),
	.w4(32'h3a9adaa4),
	.w5(32'hbb85931c),
	.w6(32'h3b3c1398),
	.w7(32'hbb3f84fc),
	.w8(32'hba5fe786),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6bd5a),
	.w1(32'h3a143731),
	.w2(32'hba3628b2),
	.w3(32'hba1bfbd7),
	.w4(32'h38c2d176),
	.w5(32'hbb886c20),
	.w6(32'h3a9fc5a8),
	.w7(32'hba91f411),
	.w8(32'h3b4353be),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad805a7),
	.w1(32'hb9d9273a),
	.w2(32'hbb4b0b1e),
	.w3(32'hbabc8edc),
	.w4(32'hb9f9f8e1),
	.w5(32'hba73ffba),
	.w6(32'h3b3456a0),
	.w7(32'hba734f30),
	.w8(32'hba563a11),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa23a21),
	.w1(32'h3b7d471e),
	.w2(32'h3b9ba463),
	.w3(32'hb904e266),
	.w4(32'h3b8d1bd6),
	.w5(32'h3b226f84),
	.w6(32'h3b34c97a),
	.w7(32'h3ad22126),
	.w8(32'h3b53d642),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78debd),
	.w1(32'hbb2be797),
	.w2(32'hbb8428d4),
	.w3(32'h3b2e3190),
	.w4(32'hbadb3c7a),
	.w5(32'hbb3f279b),
	.w6(32'h3b60c938),
	.w7(32'h398f64f8),
	.w8(32'hba938a8b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9543dae),
	.w1(32'hbaae3b54),
	.w2(32'hbbdcb042),
	.w3(32'hba2cddb7),
	.w4(32'h3c18e509),
	.w5(32'h3b2fff72),
	.w6(32'h3c08c547),
	.w7(32'h3b1876df),
	.w8(32'h3b4c7304),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b1389),
	.w1(32'h3a8c8020),
	.w2(32'hbae47e23),
	.w3(32'h3baa39d7),
	.w4(32'hb9876714),
	.w5(32'hbaf8f2b6),
	.w6(32'h3bd24f31),
	.w7(32'h396ca8b3),
	.w8(32'hbb3127ea),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de396),
	.w1(32'h3a6dc488),
	.w2(32'hbab19d04),
	.w3(32'hbb32963c),
	.w4(32'h3ab9df32),
	.w5(32'hbb9ead5b),
	.w6(32'hbaebc4d5),
	.w7(32'hbbc85ae9),
	.w8(32'hba4d1b5a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61baf9),
	.w1(32'h3946404c),
	.w2(32'hbb6bb3cb),
	.w3(32'hba33375d),
	.w4(32'h3a153325),
	.w5(32'hbb4e1c25),
	.w6(32'h3a29fa28),
	.w7(32'hba83a8b0),
	.w8(32'h3935f20f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab121eb),
	.w1(32'h3baad9db),
	.w2(32'h3bf667ae),
	.w3(32'hba47087a),
	.w4(32'h3c040916),
	.w5(32'h3c40891f),
	.w6(32'h3ba7032d),
	.w7(32'h3bc68ec2),
	.w8(32'h3c22cbd7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23620d),
	.w1(32'hb8f41041),
	.w2(32'hbb10293b),
	.w3(32'h3c466565),
	.w4(32'h39d8a8d1),
	.w5(32'hbb622b75),
	.w6(32'h3ae56ab6),
	.w7(32'hbaf08e59),
	.w8(32'h3aa42065),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a45a6),
	.w1(32'h39d49972),
	.w2(32'h3bbbc1c0),
	.w3(32'h3b1dc706),
	.w4(32'hbabedaa3),
	.w5(32'h3b225613),
	.w6(32'h3b8f63fc),
	.w7(32'hbb4ae79c),
	.w8(32'h3b27695e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dcb55),
	.w1(32'hbb7d811d),
	.w2(32'h39c4ce82),
	.w3(32'h39415083),
	.w4(32'hba10ad6b),
	.w5(32'h3b0de367),
	.w6(32'hbb3ebcfe),
	.w7(32'hba872b70),
	.w8(32'h3a831cda),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c47c8),
	.w1(32'hbb78a8e8),
	.w2(32'hbbbb00d2),
	.w3(32'h3b82f543),
	.w4(32'h3a29e4c8),
	.w5(32'h3a646546),
	.w6(32'h3ac811d2),
	.w7(32'hbb030a42),
	.w8(32'hbaf6ec15),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2583a),
	.w1(32'h3bb6c573),
	.w2(32'h3c02ee87),
	.w3(32'h3b49bd34),
	.w4(32'h3b2ce993),
	.w5(32'h3b75beb8),
	.w6(32'h3b3c105c),
	.w7(32'h3c443ba7),
	.w8(32'h3b64ff95),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37f505),
	.w1(32'h3b0bdc47),
	.w2(32'h3b1264c6),
	.w3(32'h3b2fb1b8),
	.w4(32'h3aeab9d4),
	.w5(32'hbabea5e2),
	.w6(32'h3b4825c5),
	.w7(32'h3a90c09d),
	.w8(32'h39908a4e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa54184),
	.w1(32'h3ad47d9e),
	.w2(32'hbaec55c2),
	.w3(32'hbb3da5b9),
	.w4(32'h3b87e3ce),
	.w5(32'h3ab91dc1),
	.w6(32'hbb0702c4),
	.w7(32'hba5c1761),
	.w8(32'hbade69dd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802d56),
	.w1(32'hb747a560),
	.w2(32'h3c42ecb9),
	.w3(32'h3ac9e0ab),
	.w4(32'h3a10dbae),
	.w5(32'h3c41bbda),
	.w6(32'h3a53bc07),
	.w7(32'h3bc4a91a),
	.w8(32'hbad2cb58),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b57c32),
	.w1(32'hbadcae78),
	.w2(32'hbb8b9d6a),
	.w3(32'hbbb4f379),
	.w4(32'hbb2df524),
	.w5(32'hbb41eccf),
	.w6(32'h38eb305e),
	.w7(32'hbb8b6bff),
	.w8(32'hbb1f81b8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04231),
	.w1(32'hbb678ebc),
	.w2(32'hbbb481a1),
	.w3(32'hbb41ed0c),
	.w4(32'hbb66a796),
	.w5(32'hbb8415ee),
	.w6(32'h3aeb90b9),
	.w7(32'hbaece5ec),
	.w8(32'hbb38703d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1ff0a),
	.w1(32'h3a11a17d),
	.w2(32'h3b5b3d52),
	.w3(32'hbacc5d3a),
	.w4(32'h3b4b7d0a),
	.w5(32'h3baa7fa3),
	.w6(32'h3b268b5b),
	.w7(32'hba35264a),
	.w8(32'hbaf0c9fc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6d7a1),
	.w1(32'hbb327127),
	.w2(32'hbbc9848a),
	.w3(32'h3b8adb46),
	.w4(32'hbac31d5d),
	.w5(32'hbb435b4b),
	.w6(32'h3b18c2e7),
	.w7(32'hbb761f2d),
	.w8(32'hbb11472e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31318f),
	.w1(32'hbb346307),
	.w2(32'hbb7ae774),
	.w3(32'h3b5dd44f),
	.w4(32'hbb7ae4e3),
	.w5(32'hba483b2f),
	.w6(32'hbb4070fd),
	.w7(32'hbaa14b92),
	.w8(32'hbbab5910),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f1e00),
	.w1(32'hbb4cbc38),
	.w2(32'h3bdbec8c),
	.w3(32'h3b3ee461),
	.w4(32'hbbc0b13c),
	.w5(32'h3ac80c78),
	.w6(32'hbc55df59),
	.w7(32'hbbb939ee),
	.w8(32'hbb927031),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84f37f),
	.w1(32'h3b2305a9),
	.w2(32'h3b21e39e),
	.w3(32'h395802ff),
	.w4(32'h3aade2a3),
	.w5(32'h38265e0f),
	.w6(32'h3a5a8246),
	.w7(32'h39c134e2),
	.w8(32'h39a5cad9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab06f26),
	.w1(32'hbaf14229),
	.w2(32'h3a8a7bcc),
	.w3(32'hb9920605),
	.w4(32'hbb1b5b2a),
	.w5(32'hb9a6ef08),
	.w6(32'hbbdcfd7d),
	.w7(32'hbb149126),
	.w8(32'hbb2356c1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b9a02),
	.w1(32'hbaf18e77),
	.w2(32'h3b14d6c0),
	.w3(32'h3a3a909a),
	.w4(32'h39f66ebe),
	.w5(32'h3b0ab613),
	.w6(32'h392bb7a4),
	.w7(32'hbb22be89),
	.w8(32'h3aa62107),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e360b),
	.w1(32'hba967aed),
	.w2(32'hbb280cd2),
	.w3(32'h399f7ca2),
	.w4(32'hb9c4a87b),
	.w5(32'hbb20e0ad),
	.w6(32'h3b122613),
	.w7(32'h3a516305),
	.w8(32'h383cb319),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b318),
	.w1(32'h3918e906),
	.w2(32'hba95405b),
	.w3(32'hbb6b81f8),
	.w4(32'h3a8fb160),
	.w5(32'hbb106246),
	.w6(32'h3aa9fbb0),
	.w7(32'h3a34c2d3),
	.w8(32'h3a0f075c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fdae9),
	.w1(32'hbac60b32),
	.w2(32'h3aefc485),
	.w3(32'hbb14bf61),
	.w4(32'hbb1ef171),
	.w5(32'hb89a0158),
	.w6(32'hbbe6ac10),
	.w7(32'hbb2119bc),
	.w8(32'hbb423a7e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd36e),
	.w1(32'hba92ae55),
	.w2(32'h3b3e5588),
	.w3(32'h39ad8f56),
	.w4(32'hba3f7e82),
	.w5(32'h3b1b89cc),
	.w6(32'h3b23eb16),
	.w7(32'h3b52a69c),
	.w8(32'h3b33fbe5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae88c76),
	.w1(32'h3b155f7a),
	.w2(32'h3af3ee41),
	.w3(32'hb9bf66f4),
	.w4(32'h3ad92871),
	.w5(32'hbac9ec9b),
	.w6(32'h3b38edf5),
	.w7(32'h3ae45d96),
	.w8(32'h3a03942a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40eb1e),
	.w1(32'hbad8ef85),
	.w2(32'h3a1611d4),
	.w3(32'hb99dedd2),
	.w4(32'hbbdfae86),
	.w5(32'h3a7e9fa8),
	.w6(32'h3af7e087),
	.w7(32'h3af60d48),
	.w8(32'h3b88d99f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0709d0),
	.w1(32'h3b98abb2),
	.w2(32'h3b8efd5a),
	.w3(32'hba87f26e),
	.w4(32'h3abe98f5),
	.w5(32'h3a672732),
	.w6(32'h3b83740d),
	.w7(32'h3abf39d6),
	.w8(32'h3a3917de),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53e738),
	.w1(32'h3bb0967a),
	.w2(32'h3b91666c),
	.w3(32'h3ae84881),
	.w4(32'h3b38edee),
	.w5(32'h396842f9),
	.w6(32'h3bd56eb8),
	.w7(32'h3afcc106),
	.w8(32'h3b070925),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62bbf0),
	.w1(32'hbbef1d14),
	.w2(32'hbb51af6d),
	.w3(32'hbb2ade93),
	.w4(32'hbb9e7939),
	.w5(32'h39d0ddfc),
	.w6(32'hbba97075),
	.w7(32'hbbd9e709),
	.w8(32'h399c831c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001f18),
	.w1(32'hbb23b4c6),
	.w2(32'h3b15a710),
	.w3(32'h3b624c9f),
	.w4(32'hbb6ce039),
	.w5(32'hb8e062a1),
	.w6(32'hbc2a1aa6),
	.w7(32'hbb668b02),
	.w8(32'hbb86bb91),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374f7b),
	.w1(32'hbb05f45d),
	.w2(32'hbb042caa),
	.w3(32'h39f88058),
	.w4(32'hbb03a5aa),
	.w5(32'hbb133529),
	.w6(32'hbb486dfa),
	.w7(32'hba83ce72),
	.w8(32'hbb263306),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602d1b),
	.w1(32'hbb2ac664),
	.w2(32'hbb3dcda3),
	.w3(32'hbb65ac2a),
	.w4(32'hbb297e8d),
	.w5(32'hbb24f991),
	.w6(32'hbb96b76d),
	.w7(32'hbb183228),
	.w8(32'hbb66131e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6008b8),
	.w1(32'h3b9c7769),
	.w2(32'h3acda67e),
	.w3(32'hbb5c927e),
	.w4(32'hbac0a137),
	.w5(32'h3b35b3c2),
	.w6(32'h3bb7b81b),
	.w7(32'h3b6c8ca5),
	.w8(32'hb9c0f88f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6f508),
	.w1(32'hba3216a2),
	.w2(32'hb9810938),
	.w3(32'h3a62ef20),
	.w4(32'hb96e002f),
	.w5(32'h3a8bde40),
	.w6(32'h3ab542c0),
	.w7(32'h3a5f721b),
	.w8(32'hba60ad95),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcc35d),
	.w1(32'hba957d49),
	.w2(32'hbb5d312e),
	.w3(32'h3a33755d),
	.w4(32'h39bc78e2),
	.w5(32'hbbd22432),
	.w6(32'h3947120d),
	.w7(32'hbb0e47c3),
	.w8(32'h39aed817),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0afe8f),
	.w1(32'hbb018be8),
	.w2(32'hbb61f4b6),
	.w3(32'hbaae700c),
	.w4(32'hba207fac),
	.w5(32'hbb5a5cee),
	.w6(32'hb9c3ab96),
	.w7(32'hbb773f34),
	.w8(32'hbae90021),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac86fa6),
	.w1(32'h3abc2a47),
	.w2(32'hb9cea3bc),
	.w3(32'hbb57c8da),
	.w4(32'h38e44e8c),
	.w5(32'hbac254ef),
	.w6(32'hb934531c),
	.w7(32'h39b60d47),
	.w8(32'hba0b0c7a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3b988),
	.w1(32'h3abc7137),
	.w2(32'h3b430bb0),
	.w3(32'h398932ed),
	.w4(32'h3a38c70d),
	.w5(32'h3a062525),
	.w6(32'hb9e0077b),
	.w7(32'hbae32c79),
	.w8(32'hbc0ecfab),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b9ce),
	.w1(32'h39934fc6),
	.w2(32'hba8ba254),
	.w3(32'hbb3396d4),
	.w4(32'h3a7b92e2),
	.w5(32'h3b059f7e),
	.w6(32'hbb547aaa),
	.w7(32'hba90deab),
	.w8(32'hbb40f182),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb884a),
	.w1(32'hba6314cc),
	.w2(32'hbba290d8),
	.w3(32'h3b86851b),
	.w4(32'hb69f4c02),
	.w5(32'hbb3237d6),
	.w6(32'h3b457079),
	.w7(32'hbb25886b),
	.w8(32'h3abf761a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18591a),
	.w1(32'hba4658b6),
	.w2(32'hbb24a75e),
	.w3(32'hbaa2c826),
	.w4(32'hbb23d255),
	.w5(32'hbb2de141),
	.w6(32'h3ab1c1aa),
	.w7(32'hb90c7634),
	.w8(32'hba934351),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a567c77),
	.w1(32'hbadec034),
	.w2(32'hbabcc982),
	.w3(32'h3aa412aa),
	.w4(32'hbb8ad8bc),
	.w5(32'hbbb01fe6),
	.w6(32'h3bcb8b07),
	.w7(32'h3a968d20),
	.w8(32'hbb78c837),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule