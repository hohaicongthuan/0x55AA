module layer_10_featuremap_315(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3e185),
	.w1(32'h38995668),
	.w2(32'h3a26ae6a),
	.w3(32'h391ab44c),
	.w4(32'h3aefb197),
	.w5(32'h3a02b45c),
	.w6(32'h3904fc60),
	.w7(32'h3a1e8baa),
	.w8(32'h3a4a6e38),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698690),
	.w1(32'h3b94fb49),
	.w2(32'h3bb0f2bb),
	.w3(32'h3b2ec9a7),
	.w4(32'h3b382de8),
	.w5(32'h3b28218d),
	.w6(32'h3b48725a),
	.w7(32'h3aec5ede),
	.w8(32'h3b42b65b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b7514),
	.w1(32'h3ab0358a),
	.w2(32'h3ab1abf4),
	.w3(32'h39c39150),
	.w4(32'hb7a492bf),
	.w5(32'h396b8f39),
	.w6(32'h3a136010),
	.w7(32'hb89a9ce7),
	.w8(32'h38f97218),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3e70a),
	.w1(32'h39816b67),
	.w2(32'h39cc2724),
	.w3(32'h3958e88c),
	.w4(32'h3a09032a),
	.w5(32'hba957244),
	.w6(32'hb9be55a4),
	.w7(32'h3a44bb72),
	.w8(32'hba4ffbd3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d739a),
	.w1(32'hbab4e98e),
	.w2(32'hb992cd77),
	.w3(32'hbaca1980),
	.w4(32'hb8d279cd),
	.w5(32'hba1031e6),
	.w6(32'hbb06b8e4),
	.w7(32'h38a00465),
	.w8(32'hb995ba42),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c4cfc),
	.w1(32'hba2c8796),
	.w2(32'h399952e0),
	.w3(32'hb9f88ad5),
	.w4(32'h39aa65f2),
	.w5(32'h39d94bd4),
	.w6(32'hba67596c),
	.w7(32'hb84112a9),
	.w8(32'h3932694e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a332205),
	.w1(32'h3857af5d),
	.w2(32'hb9c76240),
	.w3(32'h3af596bf),
	.w4(32'h3a8561bc),
	.w5(32'h390dc8a6),
	.w6(32'h3a1e1ece),
	.w7(32'hb9ab149c),
	.w8(32'hbad08a4d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98706d),
	.w1(32'hbbb9b029),
	.w2(32'hbc0b02f4),
	.w3(32'hbbdcb76d),
	.w4(32'hbb6d5a5e),
	.w5(32'hbadcbbb9),
	.w6(32'hbbd3b60d),
	.w7(32'hbbffcad8),
	.w8(32'hbbf61339),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808e55),
	.w1(32'h388d7242),
	.w2(32'h3a020248),
	.w3(32'h3a72b6d6),
	.w4(32'h3ab90d56),
	.w5(32'hba991e29),
	.w6(32'h3a51bc80),
	.w7(32'h3a5c956d),
	.w8(32'hbaa58dd9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85c678),
	.w1(32'h3a661d73),
	.w2(32'h3aff74c3),
	.w3(32'hbb3fecc2),
	.w4(32'hb8b9ff2d),
	.w5(32'h39e84430),
	.w6(32'hbb175d42),
	.w7(32'hbb1e573e),
	.w8(32'hba768ecc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bd15e),
	.w1(32'hb8dc0f22),
	.w2(32'hb84d6ed2),
	.w3(32'hb994e446),
	.w4(32'h39760973),
	.w5(32'hb9ef736f),
	.w6(32'h38dc3203),
	.w7(32'h39ad96c5),
	.w8(32'hb971f997),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8256b2),
	.w1(32'h39fe978d),
	.w2(32'hbb2c5fd6),
	.w3(32'h3aa410b3),
	.w4(32'h3ac40f0a),
	.w5(32'hbadc990b),
	.w6(32'h3a89e23a),
	.w7(32'h368e02cf),
	.w8(32'hbbb33179),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868c2d),
	.w1(32'hb9a38067),
	.w2(32'hbb0d64a2),
	.w3(32'hba29e050),
	.w4(32'hbb517c08),
	.w5(32'h38a35f56),
	.w6(32'hb5a9052c),
	.w7(32'hbb5a64c4),
	.w8(32'hb9b75e50),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69f19),
	.w1(32'hb83aaa59),
	.w2(32'h38db0ef4),
	.w3(32'hba3f1baf),
	.w4(32'h380dd113),
	.w5(32'hba383115),
	.w6(32'h39b2e275),
	.w7(32'hb9d71bf2),
	.w8(32'hba008dcf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a658039),
	.w1(32'h3b1671a4),
	.w2(32'h3acfcb6f),
	.w3(32'h3a85c598),
	.w4(32'h39cc2356),
	.w5(32'hb9372987),
	.w6(32'h3ab6cb5f),
	.w7(32'h3ad7cb0a),
	.w8(32'h3b271910),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae72533),
	.w1(32'hb9d2660d),
	.w2(32'h3a7bb0dc),
	.w3(32'hba90b64f),
	.w4(32'hba8c9aa1),
	.w5(32'h3a4967f4),
	.w6(32'hbb136494),
	.w7(32'hbae60a5f),
	.w8(32'hba159411),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a553efe),
	.w1(32'hb9e86a5e),
	.w2(32'h3982e268),
	.w3(32'h3a137900),
	.w4(32'h39e3b109),
	.w5(32'hb869b433),
	.w6(32'hba8ba6fc),
	.w7(32'hba4c1063),
	.w8(32'hba5b5d1c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a3f48),
	.w1(32'hbc908037),
	.w2(32'hbc9656ba),
	.w3(32'hbc7a8478),
	.w4(32'hbc461e56),
	.w5(32'hbc816f3b),
	.w6(32'hbc40624e),
	.w7(32'hbc54f1aa),
	.w8(32'hbc61a487),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83aaf5),
	.w1(32'hbbbed45c),
	.w2(32'hbb878fb7),
	.w3(32'hbbc92a38),
	.w4(32'hbba10677),
	.w5(32'hbbb29c0a),
	.w6(32'hbb812a1e),
	.w7(32'hbb485fd9),
	.w8(32'hbb94a46a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921a36),
	.w1(32'hbade1cdd),
	.w2(32'hb991a023),
	.w3(32'hba610666),
	.w4(32'hb88ccb0b),
	.w5(32'hb904818b),
	.w6(32'hbac243a5),
	.w7(32'hb98c7838),
	.w8(32'h39df63e0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8948b0),
	.w1(32'h390afd27),
	.w2(32'h3a440eef),
	.w3(32'hb95f510a),
	.w4(32'h39e4c766),
	.w5(32'h3ab94799),
	.w6(32'h38f2a4d7),
	.w7(32'h3aef23fc),
	.w8(32'h3ac7c78e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302d20),
	.w1(32'h3b5990f6),
	.w2(32'h3b0dedec),
	.w3(32'h3b68b045),
	.w4(32'h3b8c4498),
	.w5(32'h3a735072),
	.w6(32'h3b509769),
	.w7(32'h3b5e4b83),
	.w8(32'h3a69889c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8607b5),
	.w1(32'hbc8bbc4c),
	.w2(32'hbc7f7a42),
	.w3(32'hbc85291c),
	.w4(32'hbc2086c1),
	.w5(32'hbca22608),
	.w6(32'hbcb889e7),
	.w7(32'hbc0dba87),
	.w8(32'hbc9f33a0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6a9d5),
	.w1(32'h3abf72b5),
	.w2(32'h3b53503b),
	.w3(32'h39538ac1),
	.w4(32'h3ad11e5f),
	.w5(32'h3b3388b6),
	.w6(32'h3a0c7aca),
	.w7(32'h38485df3),
	.w8(32'h3ac14ace),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f3345),
	.w1(32'h3bbcfcf3),
	.w2(32'h3bc5c9fe),
	.w3(32'h3b49d2c6),
	.w4(32'h3bb02eb2),
	.w5(32'h3bab645a),
	.w6(32'h3a93e92b),
	.w7(32'h3a9dfbca),
	.w8(32'h3a81d434),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31cd13),
	.w1(32'h3ac8f2d5),
	.w2(32'h3a378566),
	.w3(32'hb8707884),
	.w4(32'h3a3c8b2b),
	.w5(32'hbad0b1de),
	.w6(32'h3a4f57dc),
	.w7(32'h3a70ebc4),
	.w8(32'hba52541c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a196b5),
	.w1(32'hb706b70e),
	.w2(32'hba529932),
	.w3(32'hb9a8d163),
	.w4(32'hba23abe9),
	.w5(32'h3a3fb400),
	.w6(32'h3931c881),
	.w7(32'hba00d7e5),
	.w8(32'h3a467cb5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3faccd),
	.w1(32'h3b97c9fe),
	.w2(32'h3b916e71),
	.w3(32'h3b830ce9),
	.w4(32'h3bab2322),
	.w5(32'h3a993f24),
	.w6(32'h3b899e4b),
	.w7(32'h3b8e4c65),
	.w8(32'h3b3e2651),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6d272),
	.w1(32'h3ad28f11),
	.w2(32'h3ad4dc6b),
	.w3(32'h39ae53d5),
	.w4(32'h3aec999e),
	.w5(32'h39e29fdb),
	.w6(32'h3a959a14),
	.w7(32'h3ae174df),
	.w8(32'h393b7297),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd1625),
	.w1(32'h3b3bf7e8),
	.w2(32'h3b775d70),
	.w3(32'h3a12794d),
	.w4(32'h3b397583),
	.w5(32'h3b1c9a3b),
	.w6(32'h3b0bf1d8),
	.w7(32'h3b2658a8),
	.w8(32'h3b5ab1db),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaea500),
	.w1(32'hba3c2e30),
	.w2(32'hb9f2156c),
	.w3(32'hba5ff01b),
	.w4(32'hbaaec335),
	.w5(32'h3ad04079),
	.w6(32'h39540f54),
	.w7(32'hb99cad3c),
	.w8(32'h3a25c247),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca7c8f),
	.w1(32'h3a999e75),
	.w2(32'h3a877882),
	.w3(32'h3abc4eea),
	.w4(32'h39a78983),
	.w5(32'h395453a9),
	.w6(32'h3a5fad28),
	.w7(32'h3a856bb2),
	.w8(32'hb9dcdce1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab37b69),
	.w1(32'h39edfd50),
	.w2(32'h387400e1),
	.w3(32'hbac6e9c2),
	.w4(32'h3a06a48c),
	.w5(32'h3a02a624),
	.w6(32'h3a89aaa0),
	.w7(32'h3ab16f5d),
	.w8(32'hb8df84da),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1240ba),
	.w1(32'hba2b3d3f),
	.w2(32'h3a8ce2f2),
	.w3(32'hb92d66cf),
	.w4(32'hb9d7c552),
	.w5(32'h3acfde89),
	.w6(32'hba9cf62f),
	.w7(32'hbabb453a),
	.w8(32'h3aaecb4e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7e72),
	.w1(32'h3a01e5fe),
	.w2(32'h38b3c235),
	.w3(32'hba1319eb),
	.w4(32'hb9ae0037),
	.w5(32'hb9c28d87),
	.w6(32'hba380dad),
	.w7(32'hba7cb0d7),
	.w8(32'hbb027e42),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5733d),
	.w1(32'hba38038c),
	.w2(32'hbaaa6575),
	.w3(32'hbac96816),
	.w4(32'hba4a187c),
	.w5(32'h38c66bfb),
	.w6(32'hbad048a0),
	.w7(32'hbb22a8b3),
	.w8(32'hba41353f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5fe8a),
	.w1(32'hbb9738e2),
	.w2(32'hbb50fdd8),
	.w3(32'hbb980b28),
	.w4(32'hbb1fa2d2),
	.w5(32'hbb41e00a),
	.w6(32'hbbb803c6),
	.w7(32'hbaac049d),
	.w8(32'hbba8c392),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbe4f6),
	.w1(32'h3c335549),
	.w2(32'h3bda27a7),
	.w3(32'h3c02900c),
	.w4(32'h3c5080cf),
	.w5(32'h3c0dc391),
	.w6(32'h3bf913e3),
	.w7(32'h3c1a6e4a),
	.w8(32'h3c103493),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d9a4),
	.w1(32'h3c762ba8),
	.w2(32'h3c11c0f5),
	.w3(32'h3c6a384c),
	.w4(32'h3c5ccd43),
	.w5(32'h3bf0f404),
	.w6(32'h3c476414),
	.w7(32'h3c022b14),
	.w8(32'h3bf1889a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac529e1),
	.w1(32'h39971484),
	.w2(32'h37ee245f),
	.w3(32'h3b28b45a),
	.w4(32'h3b3a5427),
	.w5(32'h3ab87dd1),
	.w6(32'h3a451c86),
	.w7(32'h3a81ab4b),
	.w8(32'h3a62bcb9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3a481),
	.w1(32'hbaa0f845),
	.w2(32'hba16a63b),
	.w3(32'hbb064a74),
	.w4(32'hb96baab6),
	.w5(32'h394148d8),
	.w6(32'hba81b4fc),
	.w7(32'hba5fddf9),
	.w8(32'h39c9695d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f821c),
	.w1(32'h3a95cf5b),
	.w2(32'h3a68014f),
	.w3(32'h3a7ff401),
	.w4(32'h3ac473b6),
	.w5(32'h3a87e1e3),
	.w6(32'h3aad87e6),
	.w7(32'h3a56d881),
	.w8(32'h3a6967a5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30f385),
	.w1(32'h3b007e63),
	.w2(32'h3b003136),
	.w3(32'h383ec08c),
	.w4(32'h3b342502),
	.w5(32'hbb53f136),
	.w6(32'hb9ca3433),
	.w7(32'h3b1f0b64),
	.w8(32'hbb84624b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9012aa),
	.w1(32'hbb9e99c5),
	.w2(32'hba8c2e91),
	.w3(32'hbc0f8258),
	.w4(32'hbbd00bd0),
	.w5(32'hbb2ead6c),
	.w6(32'hbc064358),
	.w7(32'hbb9a1bc2),
	.w8(32'hbb0d3b78),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c56a),
	.w1(32'h3a4ea052),
	.w2(32'h398e9552),
	.w3(32'hbb0f6cd9),
	.w4(32'h3a7d4aff),
	.w5(32'h3a9e8027),
	.w6(32'hbaaada88),
	.w7(32'hb989ad40),
	.w8(32'h3aee484d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fda5d),
	.w1(32'h3b15ff9a),
	.w2(32'h3b3e435c),
	.w3(32'hba688b7b),
	.w4(32'h3a5b547c),
	.w5(32'h3ade340b),
	.w6(32'hbaad12d0),
	.w7(32'hba88beb0),
	.w8(32'h3a2a30bb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482f43),
	.w1(32'hbb5e6b04),
	.w2(32'hbb0d2ef6),
	.w3(32'hbb89b334),
	.w4(32'hbb334cce),
	.w5(32'h3bb1c62c),
	.w6(32'hbc02d10e),
	.w7(32'hbb507f06),
	.w8(32'h3b24d1da),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d7e62),
	.w1(32'hbc4a8461),
	.w2(32'hbc730966),
	.w3(32'hbc4250ba),
	.w4(32'hbc04fd30),
	.w5(32'hbc99817f),
	.w6(32'hbc1d2dbb),
	.w7(32'hbbe95d5c),
	.w8(32'hbc965b09),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4ba4),
	.w1(32'hba9b98ea),
	.w2(32'hbaf90c24),
	.w3(32'hbaa8973f),
	.w4(32'hbac61ee2),
	.w5(32'h3ae4d088),
	.w6(32'hba46cada),
	.w7(32'hbb03a747),
	.w8(32'h3af0fbe6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d0ce),
	.w1(32'h3b0b11a7),
	.w2(32'h3ae809c9),
	.w3(32'h3ab99e5f),
	.w4(32'h3aeb06a2),
	.w5(32'hb9597375),
	.w6(32'h3a772bc2),
	.w7(32'h39d49cb9),
	.w8(32'hbb2595b5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f584b5),
	.w1(32'hbae2e32b),
	.w2(32'hb8539699),
	.w3(32'hb95931e1),
	.w4(32'hb77cb63b),
	.w5(32'h39f22a84),
	.w6(32'hbaca979a),
	.w7(32'h37a7faff),
	.w8(32'h3a290be2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a61974),
	.w1(32'hb902143f),
	.w2(32'hbaa3ca7d),
	.w3(32'hba8f7850),
	.w4(32'h39d86bce),
	.w5(32'hbb0a0266),
	.w6(32'hba0b06f4),
	.w7(32'hba30c935),
	.w8(32'hbb78d8cd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb187c61),
	.w1(32'hbb0c94bd),
	.w2(32'hbad7587a),
	.w3(32'hbb0bb6ba),
	.w4(32'hbac61bd0),
	.w5(32'hba3d078a),
	.w6(32'hbb369775),
	.w7(32'hbb1be511),
	.w8(32'hba5ddf2b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc45172),
	.w1(32'hbc435aae),
	.w2(32'hbc18b1f0),
	.w3(32'hbc4a3b95),
	.w4(32'hbc11be89),
	.w5(32'hbc06a075),
	.w6(32'hbbfc1a8d),
	.w7(32'hbc02d0ea),
	.w8(32'hbbc6c9aa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed70f6),
	.w1(32'hbb0f420b),
	.w2(32'hbb49f49d),
	.w3(32'hb98a2566),
	.w4(32'h39c87cd1),
	.w5(32'hbabdcd15),
	.w6(32'hba8ac58a),
	.w7(32'hba6e3c8e),
	.w8(32'hbabb0747),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9a83),
	.w1(32'hb91bc9c8),
	.w2(32'hb9eb9a6b),
	.w3(32'hb9cdad83),
	.w4(32'hb9863062),
	.w5(32'h383ab645),
	.w6(32'hba8215dc),
	.w7(32'hba7d1d3c),
	.w8(32'h39878308),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17c59d),
	.w1(32'hb8564174),
	.w2(32'hb98063b0),
	.w3(32'hba16079c),
	.w4(32'h3a06e6c0),
	.w5(32'hb9110419),
	.w6(32'hb7813c1e),
	.w7(32'h34db42bb),
	.w8(32'hb98a3984),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f540d),
	.w1(32'hbae233b4),
	.w2(32'hb88d6770),
	.w3(32'hba748832),
	.w4(32'h39020832),
	.w5(32'h3b0a9bbd),
	.w6(32'hbab3f8cf),
	.w7(32'hb9b4db21),
	.w8(32'h3b08e3a8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0f16),
	.w1(32'h3b3f1d02),
	.w2(32'h3b0ae641),
	.w3(32'h3b32d548),
	.w4(32'h3b7396ed),
	.w5(32'h3aa177ac),
	.w6(32'h3b251e8e),
	.w7(32'h3b226d36),
	.w8(32'h3980bcbe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94c2d3),
	.w1(32'h3a8175b9),
	.w2(32'h3b03a1df),
	.w3(32'h3afbac12),
	.w4(32'h3b00f2c2),
	.w5(32'hb948fa35),
	.w6(32'hba41e6e7),
	.w7(32'h39e9ce8a),
	.w8(32'hb964a5f4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edb77),
	.w1(32'hbb5ecb18),
	.w2(32'hbb6f6c0a),
	.w3(32'hbb92ad19),
	.w4(32'hbb55ac55),
	.w5(32'hbb73666a),
	.w6(32'hbb536ddf),
	.w7(32'hbb4e6b30),
	.w8(32'hbb86bfc1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd457d8),
	.w1(32'hbb6ea736),
	.w2(32'hbbaf4c96),
	.w3(32'hbbc1dbf8),
	.w4(32'hbb44af5b),
	.w5(32'hbbf95d2a),
	.w6(32'hbb9ff24a),
	.w7(32'hbb58b14e),
	.w8(32'hbbdcffce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775e20),
	.w1(32'hba09808a),
	.w2(32'hb9be6df1),
	.w3(32'hba808db7),
	.w4(32'hba1181b7),
	.w5(32'hba341f12),
	.w6(32'hbad8c2dd),
	.w7(32'hbab06989),
	.w8(32'hba1d9967),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cf088),
	.w1(32'hba4a6cd5),
	.w2(32'hba5c6194),
	.w3(32'hbae684f2),
	.w4(32'hb9816f2f),
	.w5(32'hb9be42fa),
	.w6(32'hba61b9e6),
	.w7(32'hba872cb3),
	.w8(32'h39231659),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e43a4),
	.w1(32'hba8c8b98),
	.w2(32'hba9782f3),
	.w3(32'hbabe1fdc),
	.w4(32'hba51cc62),
	.w5(32'hba79bffe),
	.w6(32'hbb004c2b),
	.w7(32'hbb033479),
	.w8(32'hbaf436dd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada841b),
	.w1(32'hba3797de),
	.w2(32'hba239e1f),
	.w3(32'hba317c9c),
	.w4(32'hb9a07692),
	.w5(32'h39b4f964),
	.w6(32'hbaf228ae),
	.w7(32'hbaa3d304),
	.w8(32'hb6008328),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585f91),
	.w1(32'hba8cc582),
	.w2(32'hba073167),
	.w3(32'hba2cde63),
	.w4(32'hb9533a23),
	.w5(32'hbb6e1763),
	.w6(32'hbac9dabc),
	.w7(32'hbad6ff1c),
	.w8(32'hbb662f92),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ad54),
	.w1(32'h3a91d04c),
	.w2(32'hb9d85ebc),
	.w3(32'hba950221),
	.w4(32'h3aaa3cbf),
	.w5(32'h3b8f5a62),
	.w6(32'hbb52b6dc),
	.w7(32'hbb18c44b),
	.w8(32'hbb040cb3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03363),
	.w1(32'hbbd64de7),
	.w2(32'hbc2e5d0b),
	.w3(32'hbbc8cf33),
	.w4(32'hb9f4f4a2),
	.w5(32'hbc166594),
	.w6(32'hbc0a77ff),
	.w7(32'hbbb79f27),
	.w8(32'hbc61f6d2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf51174),
	.w1(32'h3b707e5d),
	.w2(32'h3bc479e4),
	.w3(32'h39d6467a),
	.w4(32'h3b87659a),
	.w5(32'h3bfbf5a2),
	.w6(32'hba15a091),
	.w7(32'h3b3736b2),
	.w8(32'h3bed1be5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e6ad),
	.w1(32'h3a302a5a),
	.w2(32'h39db77f5),
	.w3(32'h39cab483),
	.w4(32'h3a66441d),
	.w5(32'hb79e4658),
	.w6(32'h3a55ac84),
	.w7(32'h3a5525a2),
	.w8(32'hba3727ee),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1534b7),
	.w1(32'hb9bb2831),
	.w2(32'h39d1e593),
	.w3(32'h3980c547),
	.w4(32'h39e3f248),
	.w5(32'h3b12b59f),
	.w6(32'h38e3f969),
	.w7(32'h39a12aad),
	.w8(32'h3a999e6d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58e1f7),
	.w1(32'h3af9f9b1),
	.w2(32'h3a97e4d6),
	.w3(32'h3b07dea3),
	.w4(32'h3ad48506),
	.w5(32'hba804819),
	.w6(32'h3accb8ee),
	.w7(32'hb9a9cfbe),
	.w8(32'hba8a50c6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dffd9),
	.w1(32'hbb884df0),
	.w2(32'hbb565876),
	.w3(32'hbaecc50b),
	.w4(32'hba8cb133),
	.w5(32'hba91b3f4),
	.w6(32'hbb43c6db),
	.w7(32'hbb1b63b7),
	.w8(32'hbaf2be42),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8697a38),
	.w1(32'h3a488f74),
	.w2(32'h3a13c3e1),
	.w3(32'h39951508),
	.w4(32'h392b87f2),
	.w5(32'hba9747af),
	.w6(32'h38ac8f2c),
	.w7(32'h38815faf),
	.w8(32'hbb02703f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba690e4),
	.w1(32'hbc479402),
	.w2(32'hbbfaaee3),
	.w3(32'hbc2756ca),
	.w4(32'hbc1b3dd7),
	.w5(32'hbba5c3ba),
	.w6(32'hbc0218e2),
	.w7(32'hbb972690),
	.w8(32'hbb95d0a9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700564),
	.w1(32'hbc711227),
	.w2(32'hbc2e895a),
	.w3(32'hbc5a1503),
	.w4(32'hbc5cd621),
	.w5(32'hbc1fa3f4),
	.w6(32'hbc3a5ff0),
	.w7(32'hbc266f1c),
	.w8(32'hbc3826c4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39143864),
	.w1(32'h3a901cac),
	.w2(32'hba74698f),
	.w3(32'h3acbaa11),
	.w4(32'hb8d8b8e3),
	.w5(32'hbb28ffc9),
	.w6(32'h3a94bfb6),
	.w7(32'hbab868bb),
	.w8(32'hbac4687d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f044),
	.w1(32'hbb8607df),
	.w2(32'hbb6b326a),
	.w3(32'hbb86fe8e),
	.w4(32'hbaf79483),
	.w5(32'hbaad3e5e),
	.w6(32'hbb816439),
	.w7(32'hbb5aab87),
	.w8(32'hbb0fe96a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811d8a),
	.w1(32'hbab7eb53),
	.w2(32'hb9ef5fa4),
	.w3(32'hb9a3d904),
	.w4(32'h3a9ac3ef),
	.w5(32'h3a651866),
	.w6(32'hbad5fe59),
	.w7(32'hbadbaf50),
	.w8(32'hba3ef7df),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a224c74),
	.w1(32'h3aa66fd9),
	.w2(32'h3a28d4d1),
	.w3(32'h393f4930),
	.w4(32'h39cc88d1),
	.w5(32'hbaa8e15d),
	.w6(32'h3a7cc768),
	.w7(32'h3a8db42d),
	.w8(32'hbac83100),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd713be),
	.w1(32'hbc21f640),
	.w2(32'hbc0489a2),
	.w3(32'hbbd2e1cc),
	.w4(32'hbbb25313),
	.w5(32'hbb8642ed),
	.w6(32'hbbd50e28),
	.w7(32'hbbacbcf9),
	.w8(32'hbb7f2de3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c2cd),
	.w1(32'h3a0ccab0),
	.w2(32'h3a29eb8a),
	.w3(32'h3a2514c7),
	.w4(32'h39550da6),
	.w5(32'hbac7be6e),
	.w6(32'h3a425df5),
	.w7(32'h3a2df551),
	.w8(32'hba91759f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8005f),
	.w1(32'h39dd89e7),
	.w2(32'h3a9ee0f9),
	.w3(32'hb9986830),
	.w4(32'hb9565e6d),
	.w5(32'hb8d11d9e),
	.w6(32'h3a60e77f),
	.w7(32'h3a4d3df9),
	.w8(32'hb8a3e1b7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ba108),
	.w1(32'h3abb6dd4),
	.w2(32'h3a80c203),
	.w3(32'h3973d7ef),
	.w4(32'hb92b687c),
	.w5(32'hb856dce4),
	.w6(32'h3a3117a6),
	.w7(32'h395f5f9a),
	.w8(32'hba390036),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d06af),
	.w1(32'h3a2aca80),
	.w2(32'h3a091d45),
	.w3(32'h390115dc),
	.w4(32'hba21359e),
	.w5(32'h396c5144),
	.w6(32'h3907dabf),
	.w7(32'h3980c0fc),
	.w8(32'h3a59f4a5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72240f),
	.w1(32'h3aaf6311),
	.w2(32'h3b362c55),
	.w3(32'h3a95f0a1),
	.w4(32'h3b003248),
	.w5(32'h3b1981b2),
	.w6(32'h3aa38465),
	.w7(32'hba5395d8),
	.w8(32'h3abec36b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba130055),
	.w1(32'h397454de),
	.w2(32'h3a632af1),
	.w3(32'hbab1c80c),
	.w4(32'hbaa4d857),
	.w5(32'h39fb47b3),
	.w6(32'hba785b6f),
	.w7(32'h392a3f58),
	.w8(32'h399e0a3e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6effb9),
	.w1(32'hbab8d7d6),
	.w2(32'h3919800c),
	.w3(32'hba8369a0),
	.w4(32'hba98ae5f),
	.w5(32'hb9a274b2),
	.w6(32'hbadf62e5),
	.w7(32'hbaa3a62b),
	.w8(32'h3a22be33),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc526360),
	.w1(32'hbc580281),
	.w2(32'hbc157cba),
	.w3(32'hbca70147),
	.w4(32'hbc2d97df),
	.w5(32'hbc1dc306),
	.w6(32'hbc726463),
	.w7(32'hbc33751f),
	.w8(32'hbc574655),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bbf25),
	.w1(32'h3b2d1e8f),
	.w2(32'h3a1e16b1),
	.w3(32'h3b38fbff),
	.w4(32'h3b716d66),
	.w5(32'h3ab87c0b),
	.w6(32'h3b0ce15a),
	.w7(32'h3adddf51),
	.w8(32'h3a1cb274),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ad340),
	.w1(32'hba61aa02),
	.w2(32'h3aa798f9),
	.w3(32'hbb0fc04a),
	.w4(32'h3abacec2),
	.w5(32'hbacbd286),
	.w6(32'hbaca2ee0),
	.w7(32'h3b54b038),
	.w8(32'hbac6470a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a0ea7),
	.w1(32'h3b44fe91),
	.w2(32'h3b122152),
	.w3(32'h3afee485),
	.w4(32'h3b82cf31),
	.w5(32'h3b5d151d),
	.w6(32'h3b42dd29),
	.w7(32'h3b55c305),
	.w8(32'h3b6b2b35),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba847184),
	.w1(32'hbae5a1ca),
	.w2(32'hb962c2e4),
	.w3(32'hbb5cf369),
	.w4(32'hba9c3e7d),
	.w5(32'hb8702c44),
	.w6(32'hbaec0521),
	.w7(32'hbb08a566),
	.w8(32'hbb228aff),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f081a),
	.w1(32'h3a29f174),
	.w2(32'h3b4e0a35),
	.w3(32'h3ab49ec4),
	.w4(32'h3b590349),
	.w5(32'h3b64dd6a),
	.w6(32'h3a64f1f8),
	.w7(32'h3a2f4a7f),
	.w8(32'h3b005028),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd1890),
	.w1(32'h3b994bdd),
	.w2(32'h3b0fd892),
	.w3(32'h3b597d7f),
	.w4(32'h3b4809ea),
	.w5(32'h3adb34ea),
	.w6(32'h3b89bad4),
	.w7(32'h3bacbbbf),
	.w8(32'h3b031ad4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92b98c),
	.w1(32'hbb0a6cbd),
	.w2(32'hbb101a28),
	.w3(32'hb840b8b8),
	.w4(32'h399341cc),
	.w5(32'h3b320028),
	.w6(32'hbb45e1d7),
	.w7(32'hbafeaebd),
	.w8(32'h3aa5a931),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a570444),
	.w1(32'h3a0a4668),
	.w2(32'hba87902d),
	.w3(32'hbae69117),
	.w4(32'hba218d1c),
	.w5(32'hbba5179f),
	.w6(32'hb9975559),
	.w7(32'hb94347d0),
	.w8(32'hbbeb5ca5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7bfa),
	.w1(32'h39a4d2d3),
	.w2(32'hbbb03e99),
	.w3(32'h3b341721),
	.w4(32'h39106e13),
	.w5(32'hbc2ac5b6),
	.w6(32'hb814f130),
	.w7(32'hbbbc9bb3),
	.w8(32'hbbdec580),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0176fe),
	.w1(32'hbc25a6a2),
	.w2(32'h3a960e08),
	.w3(32'hbbbcd439),
	.w4(32'hbc0f0772),
	.w5(32'hbc55dbd2),
	.w6(32'hba40c330),
	.w7(32'h3a1cf28a),
	.w8(32'hbc8d2ba9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169c0b),
	.w1(32'h3b76397c),
	.w2(32'h3b967aa0),
	.w3(32'h3be8ee11),
	.w4(32'h3c472b70),
	.w5(32'hbcce7c78),
	.w6(32'hbb308628),
	.w7(32'h3b94e8f0),
	.w8(32'hbcbf45c2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a142b),
	.w1(32'hbc6e606b),
	.w2(32'hbc6d8572),
	.w3(32'hbc1a1000),
	.w4(32'hbbb9dc42),
	.w5(32'hb9398750),
	.w6(32'hbbdce6c8),
	.w7(32'hbc48b2a8),
	.w8(32'hbc481753),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68e58c),
	.w1(32'hbc9dc41a),
	.w2(32'h3b9d2cea),
	.w3(32'hbcab5544),
	.w4(32'hbb4c6460),
	.w5(32'hbb794297),
	.w6(32'hbc82c481),
	.w7(32'hbbcf0723),
	.w8(32'hbc20d711),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba109ac8),
	.w1(32'hbb97a45b),
	.w2(32'h3b93c7a0),
	.w3(32'h3b383f2b),
	.w4(32'h3bcf40db),
	.w5(32'h3afc794b),
	.w6(32'h39e82605),
	.w7(32'h3bc777ef),
	.w8(32'hb9de07ab),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92eaeb),
	.w1(32'hbceb77ec),
	.w2(32'hbcc951cd),
	.w3(32'hbc8bf92e),
	.w4(32'hbce46eef),
	.w5(32'hbc651758),
	.w6(32'hbc8fcbf8),
	.w7(32'hbc819a7c),
	.w8(32'hbc753ded),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfe713),
	.w1(32'h3b875b0b),
	.w2(32'h3c193138),
	.w3(32'h39a767c5),
	.w4(32'h3bc141af),
	.w5(32'h3ad03751),
	.w6(32'hbae17475),
	.w7(32'h3b53a018),
	.w8(32'hba038065),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a437ce0),
	.w1(32'h3b8d21fc),
	.w2(32'h3b937563),
	.w3(32'h3b269e2b),
	.w4(32'hbb15f60e),
	.w5(32'hbb34ae8e),
	.w6(32'h3c19ac93),
	.w7(32'hbbe0beb6),
	.w8(32'hbac117ae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68fe14),
	.w1(32'h3a5b49fa),
	.w2(32'h389bbf78),
	.w3(32'hb9c46d4a),
	.w4(32'hbae062f6),
	.w5(32'h3ae06176),
	.w6(32'h3a7b65b2),
	.w7(32'hbb44efca),
	.w8(32'hba02a25f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedfc14),
	.w1(32'h3ae0f65c),
	.w2(32'hbb1ab752),
	.w3(32'h3b17d8ac),
	.w4(32'hbb55b92d),
	.w5(32'h3a89a227),
	.w6(32'hbbd43d81),
	.w7(32'hbb12d3be),
	.w8(32'hbaa3ea78),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5856da),
	.w1(32'h3bb37181),
	.w2(32'h3a84c4d5),
	.w3(32'h3b9e0be6),
	.w4(32'h398b77a9),
	.w5(32'h3bc5b0ed),
	.w6(32'h3b560d2c),
	.w7(32'h399532c4),
	.w8(32'h3bd50dea),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12dec2),
	.w1(32'h3b61ac63),
	.w2(32'hba8ad148),
	.w3(32'h3bdcfad0),
	.w4(32'hb8143d4f),
	.w5(32'h3b9ef187),
	.w6(32'h3b34f7ab),
	.w7(32'h3a382df5),
	.w8(32'h3d0218a8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca43614),
	.w1(32'h3cc464bc),
	.w2(32'h3c9e3b0e),
	.w3(32'h3c9ed1c3),
	.w4(32'h3cb1bf42),
	.w5(32'h3af45437),
	.w6(32'h3ccd4321),
	.w7(32'h3cc22b5f),
	.w8(32'hbae1b93b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a76a0),
	.w1(32'h3a20414a),
	.w2(32'hbb9ba484),
	.w3(32'hbb4009bc),
	.w4(32'h3a72b2c5),
	.w5(32'h3d00ab2d),
	.w6(32'hba01ab6c),
	.w7(32'hbb818b74),
	.w8(32'h3cc44fa5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc863ba),
	.w1(32'hbc433c67),
	.w2(32'h3b918c8f),
	.w3(32'hbbb48c3a),
	.w4(32'hbc0d85ae),
	.w5(32'hba8067db),
	.w6(32'hbc9091e6),
	.w7(32'hbc1305f8),
	.w8(32'h3bcea191),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbac6d9),
	.w1(32'h3be00b31),
	.w2(32'hb9d04005),
	.w3(32'h39ce2fb2),
	.w4(32'h3bf339e3),
	.w5(32'hba932cb5),
	.w6(32'h3acaaba1),
	.w7(32'h39960320),
	.w8(32'h3c6b168f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c926b33),
	.w1(32'h3c585d60),
	.w2(32'hbbf2c826),
	.w3(32'h3ca5061f),
	.w4(32'h3c162f8b),
	.w5(32'hbbaf648e),
	.w6(32'h3d24726e),
	.w7(32'h3c0b583f),
	.w8(32'hbba8e447),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae6b3),
	.w1(32'hba1c31e4),
	.w2(32'hba52ebac),
	.w3(32'hbb497188),
	.w4(32'hb9bb19a3),
	.w5(32'hbb5602c0),
	.w6(32'hbaf3ad61),
	.w7(32'h38e17333),
	.w8(32'hbb355462),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd189a),
	.w1(32'h3bce822e),
	.w2(32'h38840ec4),
	.w3(32'h3adfe4eb),
	.w4(32'h3ba90b06),
	.w5(32'hbbc085fd),
	.w6(32'h3c08b7ac),
	.w7(32'hbb78852f),
	.w8(32'hbc0a496a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0786f3),
	.w1(32'hbb022d0d),
	.w2(32'h39a1825a),
	.w3(32'hba7f81aa),
	.w4(32'hbb1c168e),
	.w5(32'h3c1f4885),
	.w6(32'hb9812c19),
	.w7(32'hbb8ecd51),
	.w8(32'h3ba7c355),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04f2a6),
	.w1(32'hba35aaaf),
	.w2(32'hbbdd7067),
	.w3(32'h3a4a7f51),
	.w4(32'hbbbd3031),
	.w5(32'h3b069ee3),
	.w6(32'hba9033c1),
	.w7(32'hbc0e5ade),
	.w8(32'h3ce00118),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0c509),
	.w1(32'h3cdb2b92),
	.w2(32'h3d0a9193),
	.w3(32'h3bc36a33),
	.w4(32'h3af5f0e8),
	.w5(32'hbbe3873b),
	.w6(32'hbbd2e2d2),
	.w7(32'h3cdc1452),
	.w8(32'hbc1bfd73),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61ab86),
	.w1(32'h3c375f11),
	.w2(32'hbbf897a2),
	.w3(32'h3bde80f2),
	.w4(32'hbb6dc908),
	.w5(32'hbbf36ce5),
	.w6(32'h3c92f56d),
	.w7(32'hbbcd465d),
	.w8(32'hbc16c64a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07db4a),
	.w1(32'h3b2f78ce),
	.w2(32'h3c0384eb),
	.w3(32'h3b90792a),
	.w4(32'h3bfea6dc),
	.w5(32'hb9b62fb8),
	.w6(32'hba418533),
	.w7(32'h3a115608),
	.w8(32'hbbfea5cf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0c63),
	.w1(32'h3b02af88),
	.w2(32'hbb930f55),
	.w3(32'hbb809e28),
	.w4(32'h3b7bd0f2),
	.w5(32'hbba29e3c),
	.w6(32'h3973b9e2),
	.w7(32'h3a8e1dbe),
	.w8(32'hbaa381de),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb211ce2),
	.w1(32'h3b260f84),
	.w2(32'h3aa83791),
	.w3(32'h3b1b01f9),
	.w4(32'h38cbda0f),
	.w5(32'h3ca979d9),
	.w6(32'hbb1e7d89),
	.w7(32'hbac46740),
	.w8(32'h3d309be2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bac00),
	.w1(32'h3bca7afa),
	.w2(32'h3c218311),
	.w3(32'h3b848783),
	.w4(32'h3be9a518),
	.w5(32'hba8f8ef1),
	.w6(32'hbaf2e1dd),
	.w7(32'h3c50feb3),
	.w8(32'hbb7734ae),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa84b),
	.w1(32'hba699288),
	.w2(32'hbb8c2cd5),
	.w3(32'hba3ff69d),
	.w4(32'h3a27de45),
	.w5(32'h3c8e1cf2),
	.w6(32'hbb3e4f1a),
	.w7(32'hbbb0b5a5),
	.w8(32'h3d089da1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbf140),
	.w1(32'h3b91655c),
	.w2(32'hbb8dfa54),
	.w3(32'h3aa10215),
	.w4(32'hbb6aba9e),
	.w5(32'hbb708d93),
	.w6(32'hbc351358),
	.w7(32'hbbd03dba),
	.w8(32'hbc139cbc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f537e),
	.w1(32'hbc486829),
	.w2(32'hbbfd8510),
	.w3(32'hbc36e566),
	.w4(32'hbbdeb78a),
	.w5(32'hbab31bf8),
	.w6(32'hbc61596d),
	.w7(32'hbc0df3d1),
	.w8(32'hbaf0dea9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f508),
	.w1(32'hba75c92a),
	.w2(32'hbad0c92e),
	.w3(32'h3af1e05d),
	.w4(32'hbab6a177),
	.w5(32'hbc057a63),
	.w6(32'hb9b25573),
	.w7(32'hbb4cd586),
	.w8(32'hbc43c91a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34526),
	.w1(32'h3b0b52bb),
	.w2(32'hbbbb684d),
	.w3(32'hb8643753),
	.w4(32'hba89b700),
	.w5(32'hbba1365e),
	.w6(32'h3c36ff17),
	.w7(32'hba3fe637),
	.w8(32'hbbfd79c0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91282d0),
	.w1(32'hbb31a1e1),
	.w2(32'hbb925cb7),
	.w3(32'hbb287b62),
	.w4(32'hbac76ffa),
	.w5(32'h3c60a441),
	.w6(32'h37b9a74f),
	.w7(32'hbb02862d),
	.w8(32'h3c420beb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05f661),
	.w1(32'hbbe77cbd),
	.w2(32'hbb85034c),
	.w3(32'hbbea6d61),
	.w4(32'hbb2d245d),
	.w5(32'h3ab4f0b4),
	.w6(32'hbb06e8a3),
	.w7(32'hbbe0ea70),
	.w8(32'h3acd6943),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3b089),
	.w1(32'h3b7f779a),
	.w2(32'h3b956fd7),
	.w3(32'hbb270c84),
	.w4(32'h397731a5),
	.w5(32'h3b9253d6),
	.w6(32'h372a6c4e),
	.w7(32'hbb19d841),
	.w8(32'h3b607686),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b3aa),
	.w1(32'hbbf190fb),
	.w2(32'hbc1724c1),
	.w3(32'hbc2fec90),
	.w4(32'hbc04465e),
	.w5(32'hbc0af581),
	.w6(32'hbbdf293a),
	.w7(32'hbc12f45d),
	.w8(32'hbc3fd35f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3af521),
	.w1(32'hb8c62567),
	.w2(32'h3b4666c3),
	.w3(32'h3bbae721),
	.w4(32'h3b148100),
	.w5(32'h3b884251),
	.w6(32'hba03393b),
	.w7(32'h3afb681e),
	.w8(32'h3b7f7f32),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3236ee),
	.w1(32'h3a3765d9),
	.w2(32'hbb5a44fd),
	.w3(32'hbaafc8e9),
	.w4(32'hb9fa5961),
	.w5(32'hbb73a534),
	.w6(32'hbb99f1d1),
	.w7(32'hbbb2a7ba),
	.w8(32'hbb1afe51),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59f8b2),
	.w1(32'hbbcc6179),
	.w2(32'hbc1b0f28),
	.w3(32'hbc359749),
	.w4(32'hbbf107db),
	.w5(32'hbb9255f3),
	.w6(32'hbbc7a23a),
	.w7(32'hbbc53551),
	.w8(32'hbb06e2be),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6b73),
	.w1(32'h3b4148f4),
	.w2(32'hbaba585f),
	.w3(32'hbb97e5f5),
	.w4(32'hbba90820),
	.w5(32'h3c11934b),
	.w6(32'h3b823acd),
	.w7(32'hbb7a2c31),
	.w8(32'hbab24c36),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bac0c),
	.w1(32'hbac08a16),
	.w2(32'h3b4bcff1),
	.w3(32'hba6819c0),
	.w4(32'hbbe52b2f),
	.w5(32'h3b88d4a6),
	.w6(32'hbc1a5aff),
	.w7(32'hba286160),
	.w8(32'hbb4de348),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9294e2a),
	.w1(32'hbb45eeb5),
	.w2(32'h3b855d51),
	.w3(32'hbb5a460f),
	.w4(32'h3b443cca),
	.w5(32'h3caff94b),
	.w6(32'hbb68ab8d),
	.w7(32'h3b12fbef),
	.w8(32'h3d02243b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98e718),
	.w1(32'h3c81810a),
	.w2(32'hbb98a4d8),
	.w3(32'h3cb933fe),
	.w4(32'hbbbb4eb9),
	.w5(32'h3bbd3201),
	.w6(32'h3c955c0b),
	.w7(32'hbb2c405a),
	.w8(32'h3bf05e14),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86957f),
	.w1(32'h3b14ea02),
	.w2(32'h39bec6ef),
	.w3(32'hbb27d672),
	.w4(32'hbb0f9210),
	.w5(32'hbb84316f),
	.w6(32'hbab3a23c),
	.w7(32'h3ad3bd7f),
	.w8(32'hbb176532),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f524d),
	.w1(32'hbb10ba32),
	.w2(32'hbaa0f3b3),
	.w3(32'hbb895426),
	.w4(32'h3b8657fb),
	.w5(32'h3b8ed359),
	.w6(32'h3a53ffac),
	.w7(32'h3b88050c),
	.w8(32'hba92a733),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab83a),
	.w1(32'hba4546a3),
	.w2(32'h3b9084ae),
	.w3(32'hbaadbd6e),
	.w4(32'hba0de98f),
	.w5(32'hbb192670),
	.w6(32'hbbb77cbe),
	.w7(32'hba7853e7),
	.w8(32'hbb17b73a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace98a2),
	.w1(32'h3b51c62b),
	.w2(32'h39ed777d),
	.w3(32'hbb086464),
	.w4(32'hbacd5e1b),
	.w5(32'hbaba75dc),
	.w6(32'hb9abb3d6),
	.w7(32'hbb1eaf89),
	.w8(32'h3bacc97d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b31d5),
	.w1(32'h39897c79),
	.w2(32'h3a6d4414),
	.w3(32'h3a6ed041),
	.w4(32'h3b6d1a97),
	.w5(32'h3ca38032),
	.w6(32'h39b3cbbe),
	.w7(32'hb9fdda99),
	.w8(32'h3cb67d6a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe689),
	.w1(32'h3c9cc9ae),
	.w2(32'h3c24ba24),
	.w3(32'h3c6e2741),
	.w4(32'h3b02e21f),
	.w5(32'hbb89d652),
	.w6(32'h3cc36995),
	.w7(32'h3c091409),
	.w8(32'hbb2de1aa),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa6fc),
	.w1(32'h3bd4baa3),
	.w2(32'h3bef0b62),
	.w3(32'hb9828cde),
	.w4(32'h3bb1a78c),
	.w5(32'h3a2c16f8),
	.w6(32'h3c464637),
	.w7(32'h3c0ed12b),
	.w8(32'hbae95d77),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fda6e),
	.w1(32'hbae06f53),
	.w2(32'h3b0a99f2),
	.w3(32'hbb98c537),
	.w4(32'h3a3c1744),
	.w5(32'h3c806928),
	.w6(32'hbbe743e4),
	.w7(32'hb9205d66),
	.w8(32'hbb297ea0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c418a59),
	.w1(32'hbc2ab68e),
	.w2(32'h3b8bddef),
	.w3(32'hbc5b4c97),
	.w4(32'hbc80eccb),
	.w5(32'h3ac6543e),
	.w6(32'hbc2a0963),
	.w7(32'hbcc7b0f4),
	.w8(32'h3c059588),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c746f),
	.w1(32'hbbb1cbf0),
	.w2(32'hbb95cc7d),
	.w3(32'hbc4a08a8),
	.w4(32'hbb8f8db2),
	.w5(32'hbc8e3e4d),
	.w6(32'hbb55b62d),
	.w7(32'h3a6f4946),
	.w8(32'hbc4ae8b5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc82fc),
	.w1(32'hbc318783),
	.w2(32'hbc9e4cca),
	.w3(32'h3ab4350f),
	.w4(32'h3bc09c28),
	.w5(32'h3a969fa1),
	.w6(32'h3bceb35a),
	.w7(32'h3b512a0f),
	.w8(32'h3b4b13ff),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9549b3b),
	.w1(32'h3b5db5cd),
	.w2(32'h3ad0cc85),
	.w3(32'h398c3290),
	.w4(32'h3b5a891c),
	.w5(32'h3bb169f7),
	.w6(32'hbae1d895),
	.w7(32'h3a367ebd),
	.w8(32'h3b272471),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3539cc),
	.w1(32'hba1d71f0),
	.w2(32'hbb735ea0),
	.w3(32'h39f81a15),
	.w4(32'hbbe96b6b),
	.w5(32'h3b33f48d),
	.w6(32'h3b652e60),
	.w7(32'hbbb4202d),
	.w8(32'hbadffbc7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f4c72),
	.w1(32'h36f4ad1e),
	.w2(32'hbbab7a39),
	.w3(32'hbb68f2c0),
	.w4(32'hbb6b6777),
	.w5(32'hbbd363b5),
	.w6(32'hbb851405),
	.w7(32'hbbbea830),
	.w8(32'h3c0ceccd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ea9df),
	.w1(32'h3c395d0b),
	.w2(32'hbb860e78),
	.w3(32'hb7cf3b70),
	.w4(32'hbaa6d3c6),
	.w5(32'h3c0da758),
	.w6(32'h3c1366dd),
	.w7(32'h3ad0e099),
	.w8(32'h3bfce53d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0aeed),
	.w1(32'h3be9a37d),
	.w2(32'hbb8d0589),
	.w3(32'h3be3fb1d),
	.w4(32'hbb6e73fd),
	.w5(32'h3abe4c0a),
	.w6(32'h3c96a674),
	.w7(32'hbc0afe6c),
	.w8(32'hbbb79f34),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92ff77),
	.w1(32'hbc195b93),
	.w2(32'hbba35d5c),
	.w3(32'h3b3b3a0d),
	.w4(32'hbaa9527f),
	.w5(32'hbc719c95),
	.w6(32'h3b11d8bc),
	.w7(32'h3c007f58),
	.w8(32'hbba238b4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de50d),
	.w1(32'h3bfe5009),
	.w2(32'h3bac619a),
	.w3(32'hba8b87eb),
	.w4(32'hbb1d7fcd),
	.w5(32'hbb0223d9),
	.w6(32'h3ba06e4d),
	.w7(32'h3b287882),
	.w8(32'h3c5e6bc9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40ca51),
	.w1(32'hb9af551c),
	.w2(32'hbc065f05),
	.w3(32'h3b67ef67),
	.w4(32'hb9cdc3eb),
	.w5(32'hbbdacc9b),
	.w6(32'h3aea82b1),
	.w7(32'hbb6faa83),
	.w8(32'hbb885e75),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b8f5),
	.w1(32'h3aed3980),
	.w2(32'hba787213),
	.w3(32'hbb853507),
	.w4(32'h3a711f84),
	.w5(32'hbaa1495c),
	.w6(32'hb92057e0),
	.w7(32'h3ac2ab1e),
	.w8(32'hbb6dd2a4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b1d67),
	.w1(32'hbbd72e92),
	.w2(32'hbbcf7146),
	.w3(32'hbc70cc18),
	.w4(32'h3bda064f),
	.w5(32'hbc1bf2b6),
	.w6(32'hbc64486b),
	.w7(32'hbbdb51d8),
	.w8(32'hbc0a8266),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ef08),
	.w1(32'h3a279e15),
	.w2(32'hbac0cd89),
	.w3(32'h3b5a4aa5),
	.w4(32'h3bbe1581),
	.w5(32'hbb22c646),
	.w6(32'h3c637fd7),
	.w7(32'h3b61a2b1),
	.w8(32'h3b371d95),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a4f2),
	.w1(32'h3b816a42),
	.w2(32'hbbc1f9a8),
	.w3(32'h3990bcf5),
	.w4(32'hb9b618f4),
	.w5(32'h3b0a5935),
	.w6(32'h3b6b1bba),
	.w7(32'hba96ce12),
	.w8(32'hb6d54e9d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e070c),
	.w1(32'hbb00dc0d),
	.w2(32'hbadd0a8e),
	.w3(32'hbba145f9),
	.w4(32'hbb604f8f),
	.w5(32'hbbc88951),
	.w6(32'hbb568d6c),
	.w7(32'hbb86466f),
	.w8(32'hbc297787),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5fd49),
	.w1(32'hbad2cd75),
	.w2(32'hbb8d7b0d),
	.w3(32'hbb5a2ea8),
	.w4(32'hbb23fc67),
	.w5(32'h3bcdc757),
	.w6(32'hbb8f5a83),
	.w7(32'hba9a4346),
	.w8(32'hbaabd6ea),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396ac7),
	.w1(32'hbbba2031),
	.w2(32'hbadd66f9),
	.w3(32'h3b97be9c),
	.w4(32'h3bb5a584),
	.w5(32'hbc2af8ae),
	.w6(32'hbad7b336),
	.w7(32'h3bc4db71),
	.w8(32'hbafd7b87),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb589fff),
	.w1(32'hbc5264b8),
	.w2(32'hbc21ed6f),
	.w3(32'hbc5cabc9),
	.w4(32'hbc670e62),
	.w5(32'hbb43c358),
	.w6(32'hbc9737d7),
	.w7(32'hbc141a38),
	.w8(32'hbc28e155),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b4591),
	.w1(32'hba609e05),
	.w2(32'h3b3abfcc),
	.w3(32'hbb8c9944),
	.w4(32'h3b15320f),
	.w5(32'h38338370),
	.w6(32'hbbe00750),
	.w7(32'hbaace959),
	.w8(32'hbb2eb45c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64257d),
	.w1(32'h3ba7aef6),
	.w2(32'hbaf5039c),
	.w3(32'hba3ebf85),
	.w4(32'h3b3f5c91),
	.w5(32'h3b089cd6),
	.w6(32'h3b826138),
	.w7(32'hbaf30a8a),
	.w8(32'h3bf129e7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16ecdf),
	.w1(32'h3affd178),
	.w2(32'hb903a328),
	.w3(32'h38f202bc),
	.w4(32'hbc1175e9),
	.w5(32'hbc12c339),
	.w6(32'h3bb36fd8),
	.w7(32'hbb1cd818),
	.w8(32'hbb6328da),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc348aa5),
	.w1(32'hbc1d7fe6),
	.w2(32'hbbcfeda2),
	.w3(32'hbc25c95a),
	.w4(32'hbbc42642),
	.w5(32'h3b5d79bb),
	.w6(32'hbbc59c2b),
	.w7(32'hbc170069),
	.w8(32'hbae3911a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33202e),
	.w1(32'hbb12dcd6),
	.w2(32'hba1c3b24),
	.w3(32'h3b96b449),
	.w4(32'hb909bb3e),
	.w5(32'h3b25d87a),
	.w6(32'hbae89c46),
	.w7(32'h3ad77bc8),
	.w8(32'hb81eefa9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06e70),
	.w1(32'hbb27c6b4),
	.w2(32'hbb49681a),
	.w3(32'hb96c7e88),
	.w4(32'hbb9ae3c7),
	.w5(32'hbb682c47),
	.w6(32'hbb8eff2e),
	.w7(32'hbbca6203),
	.w8(32'hbc05eef7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a9a7),
	.w1(32'h3b20971e),
	.w2(32'h39a7c75f),
	.w3(32'hbaa4f8bb),
	.w4(32'h3b66b49d),
	.w5(32'hbb919d99),
	.w6(32'hbba1a76d),
	.w7(32'h3a9cdade),
	.w8(32'hbbc76f1b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641f85),
	.w1(32'hbbc34bec),
	.w2(32'hbc015cf5),
	.w3(32'hbc1057f1),
	.w4(32'hbb7bc411),
	.w5(32'hba6a93ee),
	.w6(32'hbbc353f6),
	.w7(32'hbbd71def),
	.w8(32'hbbb68d43),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab817f5),
	.w1(32'hbb5ccad6),
	.w2(32'h3954cfe6),
	.w3(32'hbb5f59a2),
	.w4(32'h3b2536f6),
	.w5(32'h3d069156),
	.w6(32'hbbc93d31),
	.w7(32'hbab4151e),
	.w8(32'h3d4206a8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29329e),
	.w1(32'h3c5c4ad1),
	.w2(32'hbb16b421),
	.w3(32'h3c3935f2),
	.w4(32'hbbb82c5b),
	.w5(32'h3c074953),
	.w6(32'h3b940c18),
	.w7(32'hbbe1346b),
	.w8(32'h3bac006f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eccf3),
	.w1(32'h3bf29fb8),
	.w2(32'h3aeb3cea),
	.w3(32'hbaf59250),
	.w4(32'h3b170489),
	.w5(32'hbcda6dd6),
	.w6(32'h3bc39ecc),
	.w7(32'hbaf7ff44),
	.w8(32'hba10427b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92eee0),
	.w1(32'h3bc98774),
	.w2(32'hbc047ddb),
	.w3(32'h3b388a03),
	.w4(32'hbc759b0a),
	.w5(32'hbbea5270),
	.w6(32'h3c1de258),
	.w7(32'hbab1b776),
	.w8(32'hbc1bf570),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c66a3),
	.w1(32'h3bd31d4a),
	.w2(32'hbb03ab83),
	.w3(32'hb9e55d40),
	.w4(32'hb98b5612),
	.w5(32'h3b4c775d),
	.w6(32'h3c144793),
	.w7(32'h3b80b3df),
	.w8(32'h39a21634),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91aefb),
	.w1(32'h3c2dff5e),
	.w2(32'hba45d0c9),
	.w3(32'h3a98e5c5),
	.w4(32'hbc44f954),
	.w5(32'hbbfdaa3d),
	.w6(32'h3c1ad97c),
	.w7(32'hbc1ac5a4),
	.w8(32'hbbda6a20),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f5de7),
	.w1(32'hbb00a5c1),
	.w2(32'hbba7c058),
	.w3(32'hbc3f76d8),
	.w4(32'hbb9d0906),
	.w5(32'hbaa2b67f),
	.w6(32'hbc042a71),
	.w7(32'hbb191580),
	.w8(32'hb9fd9f3e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3155e8),
	.w1(32'hbbfb4144),
	.w2(32'hba002869),
	.w3(32'hbb942430),
	.w4(32'h3bd1d20a),
	.w5(32'hbb28f821),
	.w6(32'hbc38dade),
	.w7(32'h3b639a4a),
	.w8(32'hbb9f313a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97b3b),
	.w1(32'h3c67a157),
	.w2(32'hbb3dbc7d),
	.w3(32'h3bb03a28),
	.w4(32'hbb8d394e),
	.w5(32'h3aa8aa7c),
	.w6(32'h3cd255c4),
	.w7(32'hbae98f87),
	.w8(32'hbb94ccb1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3654e),
	.w1(32'hbb9b600d),
	.w2(32'hbba3ed9f),
	.w3(32'hbb8b709d),
	.w4(32'hb9d31293),
	.w5(32'hbc22f4b1),
	.w6(32'hbbc6d8cc),
	.w7(32'hbb883e77),
	.w8(32'hbc0a2db7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe97de),
	.w1(32'hbc144b35),
	.w2(32'hbaf66c48),
	.w3(32'hbc1add8c),
	.w4(32'hbc4d4587),
	.w5(32'hbb7055fe),
	.w6(32'hbc5adf54),
	.w7(32'hbc4dc91f),
	.w8(32'hbc077db3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaa2db),
	.w1(32'h3be1edaf),
	.w2(32'h3b6dbd54),
	.w3(32'h3bf85593),
	.w4(32'h3bf4f293),
	.w5(32'h391ced59),
	.w6(32'h3bd6c0c0),
	.w7(32'h3b83aa3b),
	.w8(32'hb9998b6b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fcd2),
	.w1(32'hbb6f612c),
	.w2(32'hbb9585f8),
	.w3(32'h3a8b6eb9),
	.w4(32'h38874c98),
	.w5(32'h3a415163),
	.w6(32'hbb7bfecc),
	.w7(32'hbb3606e9),
	.w8(32'h3bcd0b90),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b4129),
	.w1(32'hbb995a7a),
	.w2(32'hbbbbe227),
	.w3(32'hbb7021da),
	.w4(32'h3a97146f),
	.w5(32'h3ba53d22),
	.w6(32'hbc39110a),
	.w7(32'hbc08c2fa),
	.w8(32'hba0dd4e9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15ff9c),
	.w1(32'hbb0a0766),
	.w2(32'h3b89c249),
	.w3(32'hbbd8032b),
	.w4(32'h3c4008c0),
	.w5(32'hbc9b8fd2),
	.w6(32'hb90c21ef),
	.w7(32'hbb44b9fe),
	.w8(32'hbcaa2b61),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dbf1b),
	.w1(32'hbc84ea6a),
	.w2(32'hbba639e2),
	.w3(32'hbcbacf84),
	.w4(32'h3b4ee413),
	.w5(32'hbc380e5c),
	.w6(32'hbc54914e),
	.w7(32'hbc61ff89),
	.w8(32'hbc57d0dd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1f7eb),
	.w1(32'hbb850deb),
	.w2(32'hbb985c1a),
	.w3(32'hbc24f75f),
	.w4(32'hbc6f59bd),
	.w5(32'hbb88b1db),
	.w6(32'hbc5fe841),
	.w7(32'hbc2eef2e),
	.w8(32'hbba60999),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7af6af),
	.w1(32'h3afbea91),
	.w2(32'h3b9953b4),
	.w3(32'h3bc0ce0e),
	.w4(32'h3bee95b1),
	.w5(32'h3c6b17e9),
	.w6(32'h3b7ebde9),
	.w7(32'h3a519ae1),
	.w8(32'h3c1283be),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e1376),
	.w1(32'h38c86ff5),
	.w2(32'h3a1a856a),
	.w3(32'h3b98bced),
	.w4(32'h3ad29ee4),
	.w5(32'h3ba39415),
	.w6(32'h3b642fe4),
	.w7(32'h39a40d98),
	.w8(32'h3c10df0f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85b621),
	.w1(32'hbc22c6ef),
	.w2(32'hbc10b79b),
	.w3(32'hbbb11a7a),
	.w4(32'hbbe6b42a),
	.w5(32'h3bc82856),
	.w6(32'h3b8a08ba),
	.w7(32'hbc3a5743),
	.w8(32'hbb7d06b1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b7cfd),
	.w1(32'hba1001aa),
	.w2(32'h3bc6c40b),
	.w3(32'h3b642223),
	.w4(32'h3ba8cb67),
	.w5(32'hba9c2c94),
	.w6(32'hbbcb316c),
	.w7(32'h3b52890e),
	.w8(32'hbb9e4c6b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7243ed),
	.w1(32'hbb0f7b6d),
	.w2(32'hba260d28),
	.w3(32'hbbbfbb01),
	.w4(32'hba91332f),
	.w5(32'h3ad1b900),
	.w6(32'hbbeb1dfb),
	.w7(32'h3aba66a4),
	.w8(32'hbb3aabf1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87050e),
	.w1(32'h3b5e310c),
	.w2(32'h3bd398eb),
	.w3(32'h3bb97e21),
	.w4(32'h3b1ec268),
	.w5(32'hb8dc198e),
	.w6(32'hbaaad4b2),
	.w7(32'h3b9d22ee),
	.w8(32'hbbf54ba6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3f3d),
	.w1(32'h39b6ff62),
	.w2(32'hbad31df1),
	.w3(32'hbb811e7b),
	.w4(32'hbb6a4801),
	.w5(32'h3b10f9db),
	.w6(32'hbb34d62b),
	.w7(32'hbb54afd0),
	.w8(32'hbbc39288),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3588cc),
	.w1(32'hbac8017a),
	.w2(32'hbac7500e),
	.w3(32'hbb57fb59),
	.w4(32'hba6d65f6),
	.w5(32'hbbc38d7e),
	.w6(32'h39b63957),
	.w7(32'hbb9603b2),
	.w8(32'hbbf7beae),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d8ec),
	.w1(32'hbb4cc63c),
	.w2(32'h398582c0),
	.w3(32'hbabdc95b),
	.w4(32'h3b0be43b),
	.w5(32'hb98daa5d),
	.w6(32'h3999e47b),
	.w7(32'hb88d4da0),
	.w8(32'hbb2aa8fd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a07386),
	.w1(32'hbb8fc3e6),
	.w2(32'h3b457336),
	.w3(32'hbbd93bcb),
	.w4(32'h3b83ff91),
	.w5(32'h3c1e3c70),
	.w6(32'hbb29f80d),
	.w7(32'h3adc413b),
	.w8(32'hbb95a0d6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbf6a),
	.w1(32'hbc060dbb),
	.w2(32'h3c01516f),
	.w3(32'hbc225920),
	.w4(32'hbbabcc5e),
	.w5(32'h3b9b8e83),
	.w6(32'hbbea7332),
	.w7(32'hbaf73b3a),
	.w8(32'h3b02a3c2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8030c3),
	.w1(32'h398b2a37),
	.w2(32'h3baba6b8),
	.w3(32'h3b858dfa),
	.w4(32'h3b9ab2dc),
	.w5(32'h3a0f8eb9),
	.w6(32'h3b4aa6c5),
	.w7(32'h3bd84633),
	.w8(32'hbb401fda),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11a2e2),
	.w1(32'h3adb583e),
	.w2(32'h3bff207d),
	.w3(32'h3b3561e8),
	.w4(32'h3ba8b1ed),
	.w5(32'h3b1cc117),
	.w6(32'hbae5df0c),
	.w7(32'h3c2dd075),
	.w8(32'h3b234d97),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b0a41),
	.w1(32'hba145a2a),
	.w2(32'h3a0a4688),
	.w3(32'hbb370f36),
	.w4(32'hbaadca71),
	.w5(32'hbb9a4cd7),
	.w6(32'hbb41097f),
	.w7(32'hbb6d7df5),
	.w8(32'hbbebf7f9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa428a3),
	.w1(32'hbbcd3d8c),
	.w2(32'hbaf83c94),
	.w3(32'hbad976ca),
	.w4(32'hb8913f64),
	.w5(32'hbb75c494),
	.w6(32'hbbdf63b7),
	.w7(32'hbb75aceb),
	.w8(32'hbbf74c4f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba873f7),
	.w1(32'hbbb0b5c7),
	.w2(32'h3a4b68e9),
	.w3(32'hbb9ea0d6),
	.w4(32'h3b37c32b),
	.w5(32'hbb5c51a9),
	.w6(32'hbb1ebabc),
	.w7(32'h3b418308),
	.w8(32'hbca56cfe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e1a4),
	.w1(32'hbcc43623),
	.w2(32'hbab3c255),
	.w3(32'hbc86471f),
	.w4(32'hbc1cd8a2),
	.w5(32'hbb94748b),
	.w6(32'hbc10b508),
	.w7(32'hbc6f56ec),
	.w8(32'hba915cab),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f680b),
	.w1(32'hbaa8ef25),
	.w2(32'hbb267d8a),
	.w3(32'hbaa60a94),
	.w4(32'h397f5a4a),
	.w5(32'h3c3ce792),
	.w6(32'h3a87e897),
	.w7(32'hbb81fbba),
	.w8(32'hbb1fdee1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e5c5a),
	.w1(32'hbcbb6794),
	.w2(32'hbc797263),
	.w3(32'hbc93f96e),
	.w4(32'hbc6b2068),
	.w5(32'hbb8b48b4),
	.w6(32'hbcc75c6d),
	.w7(32'hbcb768f1),
	.w8(32'hbc331a06),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e8ec),
	.w1(32'h3b894911),
	.w2(32'hbb793a58),
	.w3(32'h3b113a73),
	.w4(32'hbc15bc28),
	.w5(32'h3c0e51ea),
	.w6(32'h3c0d1718),
	.w7(32'hbbdf99dd),
	.w8(32'h3b9268d3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c38a),
	.w1(32'h3bb3ae30),
	.w2(32'h3b1b4dc5),
	.w3(32'h3bda7a4e),
	.w4(32'h3adb948c),
	.w5(32'h3b7d53d6),
	.w6(32'h3bf6e768),
	.w7(32'hb8e8d88e),
	.w8(32'h3c20722d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f631c),
	.w1(32'hba9a8ed7),
	.w2(32'h3ae312a0),
	.w3(32'hbba476cc),
	.w4(32'hbc13992c),
	.w5(32'h3a050f8c),
	.w6(32'h3b7bc5a5),
	.w7(32'hba7e13bd),
	.w8(32'hb9432115),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa51c90),
	.w1(32'hba10ccbc),
	.w2(32'h3ac7970f),
	.w3(32'hbad78081),
	.w4(32'h39b76369),
	.w5(32'hbb2164af),
	.w6(32'hbb944aa3),
	.w7(32'h39c543d5),
	.w8(32'h3af21e51),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0cea),
	.w1(32'hbb9c6526),
	.w2(32'hbb393a7c),
	.w3(32'hba9d6f3b),
	.w4(32'h3971a627),
	.w5(32'hbb97cae8),
	.w6(32'hbb8609fc),
	.w7(32'hbaac48f7),
	.w8(32'hbb34b05f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2a68),
	.w1(32'hbbb7ba1d),
	.w2(32'hba255ac3),
	.w3(32'hbc1303c1),
	.w4(32'hbae591d9),
	.w5(32'hbc868a68),
	.w6(32'hbbeb9607),
	.w7(32'hba492bad),
	.w8(32'hbb31e498),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbac9a5),
	.w1(32'hbbef40e8),
	.w2(32'hbc3e8c35),
	.w3(32'hbc12bb3e),
	.w4(32'hbbf129d9),
	.w5(32'hbc208d50),
	.w6(32'h3b29df06),
	.w7(32'hbc316ee5),
	.w8(32'hbb4d1007),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f861b),
	.w1(32'h3932d07d),
	.w2(32'h3b0d741d),
	.w3(32'hbb87a2b9),
	.w4(32'h3b281391),
	.w5(32'h3bcbe305),
	.w6(32'hbb8fa7c4),
	.w7(32'h3a375816),
	.w8(32'h3ba9ec24),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24c3c7),
	.w1(32'h3bb3652e),
	.w2(32'h3aabf564),
	.w3(32'h3ac1171e),
	.w4(32'h3b877779),
	.w5(32'hbb743e95),
	.w6(32'h3c1c7314),
	.w7(32'h3a9886c6),
	.w8(32'hbad3346c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86192d),
	.w1(32'hba662d63),
	.w2(32'h3a14785d),
	.w3(32'hbb2fd849),
	.w4(32'hbb458dc7),
	.w5(32'hbb113fc6),
	.w6(32'hb9c2ea18),
	.w7(32'h3a76aefb),
	.w8(32'hbb691aff),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ee36),
	.w1(32'hbb1c68f6),
	.w2(32'h3b92e80d),
	.w3(32'hbbbfe331),
	.w4(32'hbbf894d3),
	.w5(32'h3a084c65),
	.w6(32'hbbafc715),
	.w7(32'hbbca2156),
	.w8(32'hbc212f5a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd2f7f),
	.w1(32'hba8bfe25),
	.w2(32'h3c025e7a),
	.w3(32'hbaaf4eec),
	.w4(32'h3be96353),
	.w5(32'h3b7bb2a4),
	.w6(32'hbbb038c6),
	.w7(32'h3c3b658a),
	.w8(32'h3b10277a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eecff),
	.w1(32'hbc258957),
	.w2(32'hbc0787be),
	.w3(32'hbbf49c71),
	.w4(32'hbb377b1e),
	.w5(32'hbb841835),
	.w6(32'hbb64a1b4),
	.w7(32'h3a611fd1),
	.w8(32'hbb96b460),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e1ec),
	.w1(32'hbbb1f184),
	.w2(32'hba21f5b3),
	.w3(32'hbba9750d),
	.w4(32'hba32d7af),
	.w5(32'hbb966d6d),
	.w6(32'hbbc86c81),
	.w7(32'hbaa66103),
	.w8(32'hbb5fde2d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b889f),
	.w1(32'hbbafef85),
	.w2(32'hbb6c36f3),
	.w3(32'hbbe57957),
	.w4(32'hbb42cdcc),
	.w5(32'hbaf82a80),
	.w6(32'hbbc1ab50),
	.w7(32'hbb1cafad),
	.w8(32'hbbef0110),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2fba),
	.w1(32'hbb7cd990),
	.w2(32'hbb54b765),
	.w3(32'hbb40f7ce),
	.w4(32'hb9d760b7),
	.w5(32'h3b1d67c8),
	.w6(32'hbbaf57e0),
	.w7(32'hbb9256a9),
	.w8(32'hb991c24b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9bf3),
	.w1(32'hbb0338d0),
	.w2(32'hbb189bb0),
	.w3(32'hbb0dd906),
	.w4(32'hba8c373d),
	.w5(32'h3a52b9b0),
	.w6(32'hbb3f71a0),
	.w7(32'hbabd9b82),
	.w8(32'h3a03f82f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce7225),
	.w1(32'hbc445bf6),
	.w2(32'hbc2d3514),
	.w3(32'hbc3a8370),
	.w4(32'hbbd1034c),
	.w5(32'hbb8a829f),
	.w6(32'hbc304bf3),
	.w7(32'hbbaed363),
	.w8(32'hbbc13a67),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b35d3),
	.w1(32'h3aa3c6b6),
	.w2(32'h3b2811bb),
	.w3(32'h3abe2654),
	.w4(32'h39ce6d9c),
	.w5(32'hba1b2f42),
	.w6(32'h3a26b1ab),
	.w7(32'h3a4fafb6),
	.w8(32'hb9e6de17),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aa0a0),
	.w1(32'h3a9dfb9d),
	.w2(32'h3a266309),
	.w3(32'h3a12dd99),
	.w4(32'h3a9c872c),
	.w5(32'h3b0b0163),
	.w6(32'h3a6f1ef2),
	.w7(32'hb9cf8c7a),
	.w8(32'h3b3980a4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a712aec),
	.w1(32'hb9c8275f),
	.w2(32'hbaf409a8),
	.w3(32'hbb577dfc),
	.w4(32'hbad25c57),
	.w5(32'hbb81e9cf),
	.w6(32'hbb42df35),
	.w7(32'hbb8be956),
	.w8(32'hbb3e3cd5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccca8f),
	.w1(32'hba7ef906),
	.w2(32'hbb0be7e4),
	.w3(32'hbac647cb),
	.w4(32'hbb2b0e34),
	.w5(32'h3a3653e7),
	.w6(32'hba811209),
	.w7(32'hbb7f390c),
	.w8(32'hbb020793),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8451b),
	.w1(32'h39cefee1),
	.w2(32'h3b368574),
	.w3(32'h3a16cc89),
	.w4(32'h3b1bd1ff),
	.w5(32'hbbc973b3),
	.w6(32'hbb16ed8b),
	.w7(32'h395195af),
	.w8(32'hbbc37de8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860b68),
	.w1(32'hbbfe16b9),
	.w2(32'hba7b5990),
	.w3(32'hbbf70ce6),
	.w4(32'hbb29ab2f),
	.w5(32'h3c07b922),
	.w6(32'hbc014756),
	.w7(32'hbb0b439b),
	.w8(32'h3c087c96),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c257665),
	.w1(32'h3c0cfd0b),
	.w2(32'h3c171894),
	.w3(32'h3bed77b6),
	.w4(32'h3c51f65f),
	.w5(32'hba1b6af8),
	.w6(32'h3c0c997c),
	.w7(32'h3c1f92ae),
	.w8(32'hbaf93bca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf72cb),
	.w1(32'h3ad5ade1),
	.w2(32'h3b09060f),
	.w3(32'h39605916),
	.w4(32'h3baa11f4),
	.w5(32'h3baad274),
	.w6(32'h3b0bd905),
	.w7(32'h3b9fd430),
	.w8(32'h3b0efa9f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacca2fa),
	.w1(32'h3bc59ea0),
	.w2(32'h3b7e0d11),
	.w3(32'h3bab71f8),
	.w4(32'hb98f0cee),
	.w5(32'hbb2a85fc),
	.w6(32'h3b84495d),
	.w7(32'hbad10c85),
	.w8(32'hbb198af1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb597c5f),
	.w1(32'hba023c9e),
	.w2(32'hba30a115),
	.w3(32'h3abaa61e),
	.w4(32'h3a650bed),
	.w5(32'hbb188ab8),
	.w6(32'h3b8bd1b3),
	.w7(32'hb8dc18d4),
	.w8(32'hbb0374fb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70b462),
	.w1(32'hbb6e61e4),
	.w2(32'hbb4cd8d6),
	.w3(32'hbb5c476e),
	.w4(32'hbb474f1a),
	.w5(32'hbb85e309),
	.w6(32'hbbbbd763),
	.w7(32'hbbaed073),
	.w8(32'hbb78b036),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0591),
	.w1(32'hbb80bf99),
	.w2(32'hbab8636b),
	.w3(32'hbb319ea5),
	.w4(32'h3a90433a),
	.w5(32'hb9aab076),
	.w6(32'hbba66dba),
	.w7(32'hba68bfc2),
	.w8(32'hbb42aaae),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb916154),
	.w1(32'hb900de88),
	.w2(32'h3ab8f16b),
	.w3(32'h3924dbe4),
	.w4(32'hbb3e1a5f),
	.w5(32'hbaa96559),
	.w6(32'hb9c8b454),
	.w7(32'hbab9d3a6),
	.w8(32'hbb0c01f2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f2556),
	.w1(32'hba33c05f),
	.w2(32'hba7a12d4),
	.w3(32'hb98f6f5c),
	.w4(32'h3a4bdcbd),
	.w5(32'h3a8bf084),
	.w6(32'h3a0a6351),
	.w7(32'h37b4436b),
	.w8(32'h3aabea6b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ef8b),
	.w1(32'hbb4ef3cd),
	.w2(32'hbb373562),
	.w3(32'hbb5eea82),
	.w4(32'hbb92c12d),
	.w5(32'hbb308450),
	.w6(32'hbacc428a),
	.w7(32'hbb690a44),
	.w8(32'hbb7f5fe1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2738e),
	.w1(32'hbc1cf5b4),
	.w2(32'hbb9519d2),
	.w3(32'hbc22ccbb),
	.w4(32'hbb8df88a),
	.w5(32'hbc0e7d53),
	.w6(32'hbc2458f4),
	.w7(32'hbb8380ce),
	.w8(32'hbc0b8afb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a67bf),
	.w1(32'hbbdfb2bb),
	.w2(32'hbbb9a8d5),
	.w3(32'hbbf68f0d),
	.w4(32'hbbf115c4),
	.w5(32'hbb444114),
	.w6(32'hbc20db22),
	.w7(32'hbbee7219),
	.w8(32'hbb620316),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399847bf),
	.w1(32'h3b7f18c0),
	.w2(32'h3af83b2a),
	.w3(32'h3b84d14c),
	.w4(32'h3b6e5767),
	.w5(32'hbaf330f0),
	.w6(32'h3aba88d8),
	.w7(32'h3ae40b74),
	.w8(32'h3aacc800),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ae58c),
	.w1(32'hbc1d9a19),
	.w2(32'hbb1f70c5),
	.w3(32'hbbb33e8f),
	.w4(32'h3a9fa0a5),
	.w5(32'h3b3d95b2),
	.w6(32'hbbd2b8b8),
	.w7(32'h3ac30780),
	.w8(32'h3b92f245),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a890865),
	.w1(32'h3a847318),
	.w2(32'hbabfa3c1),
	.w3(32'h3ab844b1),
	.w4(32'hba474d76),
	.w5(32'hbb01149a),
	.w6(32'h3b817cb1),
	.w7(32'hba646f32),
	.w8(32'h3a3e79ac),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc43036),
	.w1(32'hbb3750c4),
	.w2(32'hbb79b588),
	.w3(32'h3b5f258b),
	.w4(32'h3b4f48ff),
	.w5(32'h3bd70462),
	.w6(32'hba79beae),
	.w7(32'h3ad226ba),
	.w8(32'h3b031938),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5f16c),
	.w1(32'h3b2970ef),
	.w2(32'hbb4d49b1),
	.w3(32'h3b371aee),
	.w4(32'h3b12a447),
	.w5(32'hbb4cb033),
	.w6(32'hb8d56249),
	.w7(32'hbae7e840),
	.w8(32'hba932b1c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc21c89),
	.w1(32'hba851215),
	.w2(32'hbbcf7f09),
	.w3(32'hbb32cee4),
	.w4(32'hbb6aa95c),
	.w5(32'hbc20503e),
	.w6(32'hbb6a69f6),
	.w7(32'hbbfd229e),
	.w8(32'hbc128062),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aaf1f),
	.w1(32'hbb47d1b9),
	.w2(32'hbb3423bd),
	.w3(32'hba987045),
	.w4(32'hb92f4feb),
	.w5(32'h3a6eac87),
	.w6(32'hbb1f0e1a),
	.w7(32'hbaf1fba2),
	.w8(32'h38769ee1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a249),
	.w1(32'hbba9051e),
	.w2(32'hbb65b7ed),
	.w3(32'hbbbe173c),
	.w4(32'hb8bd7778),
	.w5(32'h3bdc4781),
	.w6(32'hbba57728),
	.w7(32'hba96b914),
	.w8(32'hbb966ba5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule