module layer_8_featuremap_234(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080262),
	.w1(32'h3b52e3d3),
	.w2(32'h3cc1db9b),
	.w3(32'hbb08f6da),
	.w4(32'hb984de03),
	.w5(32'h3c8ce321),
	.w6(32'h3c08b0ee),
	.w7(32'h3c31cdf1),
	.w8(32'hbba9d807),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0b8df),
	.w1(32'hba57f6e7),
	.w2(32'hb8e71da5),
	.w3(32'h3859ff72),
	.w4(32'h3b30e975),
	.w5(32'h3ab7a50e),
	.w6(32'hbb5922f3),
	.w7(32'hbb64853d),
	.w8(32'hbbb6ccbd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56932),
	.w1(32'h3c3d552c),
	.w2(32'hbc402453),
	.w3(32'h3b360797),
	.w4(32'h3c89c6b1),
	.w5(32'hbb6b9a56),
	.w6(32'h3c31faa8),
	.w7(32'hba82b90a),
	.w8(32'hbbd93b60),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7d3b9),
	.w1(32'hbbdd08f2),
	.w2(32'hbc2c39b1),
	.w3(32'hbc098cd6),
	.w4(32'h3b4b5104),
	.w5(32'hbc5f285c),
	.w6(32'hbbd48318),
	.w7(32'h3b4a4cc1),
	.w8(32'h3b218312),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0781ce),
	.w1(32'h3bea5832),
	.w2(32'hbafed072),
	.w3(32'hbc483995),
	.w4(32'h3c147855),
	.w5(32'h3a5d41d5),
	.w6(32'h3b60608a),
	.w7(32'hbbbf0a1b),
	.w8(32'hbc60fdbf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b0bbf),
	.w1(32'h3b8adc5c),
	.w2(32'h3be6cfeb),
	.w3(32'hbc00bee1),
	.w4(32'h3ba50f40),
	.w5(32'h3bacb0b4),
	.w6(32'h3b393669),
	.w7(32'hb9bad087),
	.w8(32'h3b84a4bc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5d9b),
	.w1(32'h386cae7f),
	.w2(32'hbbb49dc8),
	.w3(32'h3a6895e0),
	.w4(32'h3a8975e1),
	.w5(32'hbb81e715),
	.w6(32'h3adcce06),
	.w7(32'hbb322c5d),
	.w8(32'hbb7e7ef1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf669),
	.w1(32'hbcf3bd4c),
	.w2(32'hbcd41dd2),
	.w3(32'hbbf0384f),
	.w4(32'hbc9df403),
	.w5(32'hbccee67a),
	.w6(32'hbcc816e4),
	.w7(32'hbc924625),
	.w8(32'h3b6bb181),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e73df),
	.w1(32'h3c18300c),
	.w2(32'h3b90e691),
	.w3(32'h3b7bbd17),
	.w4(32'h3c094622),
	.w5(32'h3bc3bdd8),
	.w6(32'h3c176d59),
	.w7(32'hba299ecf),
	.w8(32'hbbcd49e8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac48502),
	.w1(32'h3c94a59c),
	.w2(32'hba89f1e0),
	.w3(32'h3b6a1f63),
	.w4(32'hbbf5b0a0),
	.w5(32'h3bd6abe6),
	.w6(32'h3bf77e88),
	.w7(32'h3ba62ebe),
	.w8(32'h3c1f57d4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf42c),
	.w1(32'hbc91599f),
	.w2(32'hbc87aaa1),
	.w3(32'hba16b083),
	.w4(32'hbc395151),
	.w5(32'hbcaed2d4),
	.w6(32'hbcb8c976),
	.w7(32'hbc595804),
	.w8(32'hbb8686a3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8056b4),
	.w1(32'h3baf80c0),
	.w2(32'hbbbbaea6),
	.w3(32'hba400afa),
	.w4(32'h3c009642),
	.w5(32'hbba878ac),
	.w6(32'h3bbf1e82),
	.w7(32'hbba0b3ef),
	.w8(32'h3b85b72d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0894cd),
	.w1(32'hbc1dd0ef),
	.w2(32'h3b17d55e),
	.w3(32'hb85508e4),
	.w4(32'hbbceae01),
	.w5(32'h3a90ffc1),
	.w6(32'hbb0b9ca6),
	.w7(32'h3ae14c24),
	.w8(32'h3bbc02d3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b1fe6),
	.w1(32'h3c722260),
	.w2(32'hbb712703),
	.w3(32'hbafc640c),
	.w4(32'h3c1cdfc8),
	.w5(32'hbba6f350),
	.w6(32'h3b917f6e),
	.w7(32'h3b50ecfa),
	.w8(32'hba2b1bf8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696da3),
	.w1(32'h3be25fc8),
	.w2(32'hbade2afa),
	.w3(32'hbc40224b),
	.w4(32'h3bb084ff),
	.w5(32'h3a296004),
	.w6(32'h3bf8d218),
	.w7(32'h39fc51fb),
	.w8(32'h3b3f8a63),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615fdc),
	.w1(32'h3d2055cb),
	.w2(32'h3d361de3),
	.w3(32'h3b19355b),
	.w4(32'h3d14c6ff),
	.w5(32'h3d34bb15),
	.w6(32'h3cd66734),
	.w7(32'h3c96803b),
	.w8(32'hbb21a25c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc2649),
	.w1(32'h3be565f8),
	.w2(32'h3bb59371),
	.w3(32'h3cb696e0),
	.w4(32'h3c08e7dc),
	.w5(32'h3ad0206e),
	.w6(32'hbc224bdd),
	.w7(32'hba4449b7),
	.w8(32'hbc07cdbf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c4ef1),
	.w1(32'h3b2157fe),
	.w2(32'hbb025504),
	.w3(32'hba853a10),
	.w4(32'hbbcabb07),
	.w5(32'h3b67aca3),
	.w6(32'h3bbf47c2),
	.w7(32'hb9ba8f66),
	.w8(32'hbbb1a31a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab31ce),
	.w1(32'h3c5c62e8),
	.w2(32'h3c4fd84c),
	.w3(32'hbbdcfafb),
	.w4(32'h3c866ea9),
	.w5(32'h3c855a0f),
	.w6(32'h3c310178),
	.w7(32'h399e0c1e),
	.w8(32'hbbf83190),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0715ef),
	.w1(32'hbb80869b),
	.w2(32'hba417c40),
	.w3(32'hbbcabcf7),
	.w4(32'hbc06230f),
	.w5(32'hbb0d7657),
	.w6(32'hbb0f49c3),
	.w7(32'h3ab02343),
	.w8(32'h3b14f02b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5e96d),
	.w1(32'hbbab8241),
	.w2(32'hbb1afba6),
	.w3(32'hb92278b7),
	.w4(32'hbc7c39a1),
	.w5(32'h3b596762),
	.w6(32'h39de61f1),
	.w7(32'h3be0e569),
	.w8(32'hbbf44119),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69248d),
	.w1(32'h3ba1e5a8),
	.w2(32'hbb3057bf),
	.w3(32'hbc5ffa66),
	.w4(32'h3b8cb8d5),
	.w5(32'hbab9a54b),
	.w6(32'hba2c6316),
	.w7(32'hbc08ac04),
	.w8(32'hbbb32300),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20eb42),
	.w1(32'hbc7adf36),
	.w2(32'hbc95e6ce),
	.w3(32'hbc00d339),
	.w4(32'hbae7ae84),
	.w5(32'hbc54ab49),
	.w6(32'hbc95d579),
	.w7(32'hbcbb6828),
	.w8(32'hbb61baa3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923e3c7),
	.w1(32'h3b6a3106),
	.w2(32'hbb87667a),
	.w3(32'h3b584250),
	.w4(32'h3bc5f7ff),
	.w5(32'h3a8f7cac),
	.w6(32'h3c057e55),
	.w7(32'hbc0bc1ce),
	.w8(32'hbc5836c7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51e420),
	.w1(32'hbc1585bc),
	.w2(32'hba9d1e06),
	.w3(32'hbad0cf74),
	.w4(32'hbc794fdb),
	.w5(32'h390889f4),
	.w6(32'hbb56836e),
	.w7(32'h3ac55b90),
	.w8(32'h38ed44a7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba271ee),
	.w1(32'h3c996ee9),
	.w2(32'h3cc1d022),
	.w3(32'h3bb525d3),
	.w4(32'h3b2e977b),
	.w5(32'h3c796278),
	.w6(32'h3c99cd71),
	.w7(32'h3c2c3efb),
	.w8(32'hbc906a7f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02a5da),
	.w1(32'h3b5d519d),
	.w2(32'h3a9118fc),
	.w3(32'h3b85c0b6),
	.w4(32'h3c96e1c2),
	.w5(32'hbb8117f7),
	.w6(32'hbb75c39a),
	.w7(32'h3b63db43),
	.w8(32'h3b80ddba),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ace3b),
	.w1(32'h3b1e56c1),
	.w2(32'hbc437037),
	.w3(32'hbc5c830f),
	.w4(32'hbc010dd2),
	.w5(32'hbb9782d9),
	.w6(32'h3ba4a4bc),
	.w7(32'hbc460ffd),
	.w8(32'hbb975a94),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9016),
	.w1(32'hb9aaafda),
	.w2(32'hbb4a801f),
	.w3(32'hbb9c8577),
	.w4(32'hbb83663d),
	.w5(32'hbbe6703e),
	.w6(32'h3ae605eb),
	.w7(32'hbbc083e4),
	.w8(32'h38b2afa1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b313b9d),
	.w1(32'h3b185772),
	.w2(32'hbb99880f),
	.w3(32'h3b97f176),
	.w4(32'h3b3d7fd8),
	.w5(32'hbb8e4ba6),
	.w6(32'h3b35177f),
	.w7(32'hbb53433c),
	.w8(32'h3b8e7200),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd87ec),
	.w1(32'hbba04d10),
	.w2(32'hbc104574),
	.w3(32'h3bbe90a9),
	.w4(32'hbb4a0d4d),
	.w5(32'hbb7f371c),
	.w6(32'hba56b66e),
	.w7(32'hba82dd76),
	.w8(32'h39ac92a0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd2c7),
	.w1(32'h3c90efbe),
	.w2(32'h3c441c8f),
	.w3(32'hba5c7c97),
	.w4(32'h3c7fc508),
	.w5(32'h3bf647dc),
	.w6(32'h3c1f1614),
	.w7(32'h3b72d03a),
	.w8(32'hbbe4237e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39703698),
	.w1(32'hbc3d35a5),
	.w2(32'h39c4acc3),
	.w3(32'hb768c962),
	.w4(32'hbcc73aca),
	.w5(32'hbc2b182e),
	.w6(32'hbbb08e33),
	.w7(32'hba848a2a),
	.w8(32'hb7bf6e60),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8185ce),
	.w1(32'h3c1ae627),
	.w2(32'hbaf47430),
	.w3(32'hbb89e2de),
	.w4(32'h3bb07b99),
	.w5(32'h381c09bf),
	.w6(32'h3ba1377a),
	.w7(32'h3b96f01f),
	.w8(32'hbb70086f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a260ef3),
	.w1(32'hbb6dca20),
	.w2(32'h3b922eb9),
	.w3(32'hba2ed28c),
	.w4(32'hbbf719de),
	.w5(32'hbba350b5),
	.w6(32'hbba19093),
	.w7(32'h3a851534),
	.w8(32'h3ba2a5b3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c514e85),
	.w1(32'h3c627f56),
	.w2(32'hbc18cc4b),
	.w3(32'h3aa9d124),
	.w4(32'h3c9b55e2),
	.w5(32'hbb4b49df),
	.w6(32'h3bf9e1db),
	.w7(32'hbb56faea),
	.w8(32'hbc12283b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70a9e1),
	.w1(32'hbbeb73a2),
	.w2(32'hbadac7f6),
	.w3(32'hbc8f2529),
	.w4(32'h3988093c),
	.w5(32'h3a65fb37),
	.w6(32'hbbac8055),
	.w7(32'h3b2ac11e),
	.w8(32'h3c2d79d7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22c4e7),
	.w1(32'h3bb26982),
	.w2(32'h3ae8df6d),
	.w3(32'h3c0a74f2),
	.w4(32'h3b869c15),
	.w5(32'h3b8beea9),
	.w6(32'h3ba1c384),
	.w7(32'hba82dafe),
	.w8(32'h3a279015),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c4af),
	.w1(32'h3bd8fe48),
	.w2(32'hbbd0d8c2),
	.w3(32'h3bce8eab),
	.w4(32'hba579ca1),
	.w5(32'hbb2f8612),
	.w6(32'hbb5aa198),
	.w7(32'hbc24a151),
	.w8(32'hbb7d64dc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5d2d7),
	.w1(32'h3c0570ce),
	.w2(32'hbc3178e1),
	.w3(32'hbb836456),
	.w4(32'h3c0f09d6),
	.w5(32'hbb840b60),
	.w6(32'h3b6ab53f),
	.w7(32'hbc063600),
	.w8(32'hbb7c90c8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ba347),
	.w1(32'hbbca4453),
	.w2(32'h3b1314cd),
	.w3(32'hbc17faa7),
	.w4(32'hbc11636c),
	.w5(32'hbadcf197),
	.w6(32'hbb7acae6),
	.w7(32'h3b8bb32e),
	.w8(32'h3c0baa5f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001360),
	.w1(32'h3bbb9290),
	.w2(32'h386386ab),
	.w3(32'h3ba6c7a0),
	.w4(32'h3c72f423),
	.w5(32'h3b106a9c),
	.w6(32'h395bdd51),
	.w7(32'hb9b1c8cc),
	.w8(32'h3bbc1c11),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc27059),
	.w1(32'hbbf9ec4d),
	.w2(32'hbb8e8c8f),
	.w3(32'h3b4ff953),
	.w4(32'hba890137),
	.w5(32'hbb7a2818),
	.w6(32'hbb0fec44),
	.w7(32'h3ac236c7),
	.w8(32'h3b357d74),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e72e),
	.w1(32'hbbd817dd),
	.w2(32'hbbf76e84),
	.w3(32'hba0a5728),
	.w4(32'h3a9050f7),
	.w5(32'hbb02d708),
	.w6(32'hb9df5b85),
	.w7(32'hbc10a02f),
	.w8(32'hbc02be24),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ac9f),
	.w1(32'h3c35fb66),
	.w2(32'hbc2bd031),
	.w3(32'hbacf6bf7),
	.w4(32'h3c1c48ba),
	.w5(32'hbc06a887),
	.w6(32'hba8ecb6d),
	.w7(32'hbc517d62),
	.w8(32'h3b7ff4b7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c561653),
	.w1(32'h39c060be),
	.w2(32'h3af57ff7),
	.w3(32'h3ad900f4),
	.w4(32'h39dc5ca7),
	.w5(32'h3af4fbb1),
	.w6(32'h3b2fa10c),
	.w7(32'h3b751eac),
	.w8(32'h3b97929f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3a1a),
	.w1(32'h3ca82088),
	.w2(32'hbc141b0a),
	.w3(32'h3bab4eb3),
	.w4(32'h3cafff6f),
	.w5(32'h3b4d4f4d),
	.w6(32'h3bc274aa),
	.w7(32'hbc538ed7),
	.w8(32'hbc7693b0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2acbf),
	.w1(32'h3c90fb1b),
	.w2(32'hbbb97c55),
	.w3(32'hbc5f4247),
	.w4(32'h3c91554c),
	.w5(32'h3c80d46d),
	.w6(32'h3c38b172),
	.w7(32'hbb8004fd),
	.w8(32'hbc58acea),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8aba31),
	.w1(32'h3c7237ef),
	.w2(32'hbc12c559),
	.w3(32'hbc0ec5a9),
	.w4(32'h3cb3888f),
	.w5(32'h3c412ca4),
	.w6(32'h3b9f8617),
	.w7(32'hbc561f09),
	.w8(32'hbc5be0bb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d6059),
	.w1(32'h3a17e396),
	.w2(32'h3c9b74e1),
	.w3(32'hbc09408a),
	.w4(32'hbb653dd8),
	.w5(32'h3c084fb9),
	.w6(32'h388b8c28),
	.w7(32'h3b6d9c0e),
	.w8(32'hbb04f2c8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfb418),
	.w1(32'hb9e9b8cd),
	.w2(32'hbb2ec4a2),
	.w3(32'h3abab2e7),
	.w4(32'h3930b26f),
	.w5(32'hbb20fd3c),
	.w6(32'hb83a8ac6),
	.w7(32'hbb29e781),
	.w8(32'h3adf3f88),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b386efe),
	.w1(32'h3b43574c),
	.w2(32'hbc51951e),
	.w3(32'h3aa63031),
	.w4(32'h3bd7152a),
	.w5(32'hbc465380),
	.w6(32'hbabdcaee),
	.w7(32'hbc2c55ce),
	.w8(32'hba4ec509),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259d73),
	.w1(32'h3b4dfefb),
	.w2(32'hbb9f694f),
	.w3(32'hbbef6699),
	.w4(32'h3b8c3c82),
	.w5(32'hbb2d8d29),
	.w6(32'hba380f3b),
	.w7(32'hbc1166a5),
	.w8(32'hbbebecb1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f41a1),
	.w1(32'hbc93fd1e),
	.w2(32'hbc800939),
	.w3(32'hbaf4d97f),
	.w4(32'hbb69c7fb),
	.w5(32'hbbf58eea),
	.w6(32'hbb4ecd3c),
	.w7(32'hbb02d358),
	.w8(32'h3c398eae),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f0a93),
	.w1(32'hba310098),
	.w2(32'h3be441ff),
	.w3(32'h3be17314),
	.w4(32'hbb81f2e6),
	.w5(32'h3bb8a653),
	.w6(32'h3bc67253),
	.w7(32'h3ba8ecbe),
	.w8(32'h3b6b79a1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ef103),
	.w1(32'hbbd45df9),
	.w2(32'h3b6feed4),
	.w3(32'h3b1301e2),
	.w4(32'hbb895a10),
	.w5(32'hbb4ceee5),
	.w6(32'h3b8cbf3b),
	.w7(32'hbc1be4d3),
	.w8(32'hba76fc42),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46ba3),
	.w1(32'h3b61a90b),
	.w2(32'hbc1419aa),
	.w3(32'h380c357e),
	.w4(32'h3b884ece),
	.w5(32'hbbc2f523),
	.w6(32'hbb66b317),
	.w7(32'hbc49e3c9),
	.w8(32'h3855e70c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24732c),
	.w1(32'hbb3a41f6),
	.w2(32'hbc1d2bfa),
	.w3(32'h3b2fc4fc),
	.w4(32'h3b431180),
	.w5(32'hbc105668),
	.w6(32'hba81734f),
	.w7(32'hbb9094c3),
	.w8(32'h3bb6b4d1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6a367),
	.w1(32'hba90e6f3),
	.w2(32'hbb1a7e34),
	.w3(32'h3b24402c),
	.w4(32'hba31e732),
	.w5(32'hbb84fc61),
	.w6(32'hba9e0679),
	.w7(32'hbaf60617),
	.w8(32'h3a82b7a2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d8d88e),
	.w1(32'h3b8bb29a),
	.w2(32'hbbdd9ca4),
	.w3(32'hba0a35a8),
	.w4(32'h3c153ba6),
	.w5(32'hbabc65c9),
	.w6(32'hbb010678),
	.w7(32'hbc613836),
	.w8(32'hbb966a54),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11e26f),
	.w1(32'hbc5bb774),
	.w2(32'hbbc990c3),
	.w3(32'hbc037087),
	.w4(32'hbb8f60c0),
	.w5(32'hba4c902e),
	.w6(32'h399d6696),
	.w7(32'h3ad57db2),
	.w8(32'h3c5c99c4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98bc79),
	.w1(32'hbb477a7d),
	.w2(32'hbaa93dc1),
	.w3(32'h3b3284da),
	.w4(32'hbbebe023),
	.w5(32'h3bac4c5a),
	.w6(32'h3b7885a1),
	.w7(32'h3a5dc672),
	.w8(32'hbb13838b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827534),
	.w1(32'h3b6a143a),
	.w2(32'h3c5f35b8),
	.w3(32'h3bec2255),
	.w4(32'h3b4e8d4f),
	.w5(32'h3c0789fe),
	.w6(32'h3c0f0aca),
	.w7(32'h3c0be251),
	.w8(32'h3b83fd2b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a83aa),
	.w1(32'hbb046db4),
	.w2(32'hbbbd4bb5),
	.w3(32'h3b9aeadf),
	.w4(32'hbad3e7ea),
	.w5(32'hbbf3d049),
	.w6(32'hbaa228f9),
	.w7(32'hbbc4c65d),
	.w8(32'hbc019eec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08515),
	.w1(32'hbb0ec5ee),
	.w2(32'hbabb08f8),
	.w3(32'hbbfc70fe),
	.w4(32'hba50e47c),
	.w5(32'hba480ce7),
	.w6(32'hbb56ea2c),
	.w7(32'hbb837fc1),
	.w8(32'h39ef5845),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba7a8),
	.w1(32'h3beaca59),
	.w2(32'hbac23153),
	.w3(32'h3ba9d825),
	.w4(32'h3be22e37),
	.w5(32'h3b2da7f0),
	.w6(32'h3b97db14),
	.w7(32'hbbe21ab7),
	.w8(32'hbc060708),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c3e02),
	.w1(32'hbc812b08),
	.w2(32'h3bf79089),
	.w3(32'hbbb888f4),
	.w4(32'hbc15d70c),
	.w5(32'h3c06ab0f),
	.w6(32'hbb0e3fab),
	.w7(32'h3c0e7bb6),
	.w8(32'h3ba6fb9a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb9d10),
	.w1(32'h3b46c20c),
	.w2(32'hbbdb4e32),
	.w3(32'hbb3aa86c),
	.w4(32'hbb010b08),
	.w5(32'hbc0f1e36),
	.w6(32'hbb1ca3e1),
	.w7(32'hbb85768c),
	.w8(32'hbc0ebe6b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9220a),
	.w1(32'hbafa65c3),
	.w2(32'hbc30b0c4),
	.w3(32'hbae17c4f),
	.w4(32'hbc058831),
	.w5(32'hbc293834),
	.w6(32'h3bd9a350),
	.w7(32'hbc01217d),
	.w8(32'hbb96a945),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83fdd3),
	.w1(32'h3b94ef5b),
	.w2(32'hbbc9e1ab),
	.w3(32'hbbe8a9a2),
	.w4(32'h3cbe1e40),
	.w5(32'h3b3768ae),
	.w6(32'h3a806235),
	.w7(32'hbb4075cc),
	.w8(32'hbba54a42),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39eea7),
	.w1(32'h3a8de9ff),
	.w2(32'hbbb315bf),
	.w3(32'hbbafb058),
	.w4(32'h3bcdb4b5),
	.w5(32'hbb1515b4),
	.w6(32'h3a3492bc),
	.w7(32'hbc0fc993),
	.w8(32'hbc009ce2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab45c6d),
	.w1(32'h3ca7545f),
	.w2(32'hbbd4e0a8),
	.w3(32'hbab9ff5c),
	.w4(32'h3c61c2bb),
	.w5(32'hbbaa05a8),
	.w6(32'h3c14209b),
	.w7(32'hbba2d2d7),
	.w8(32'hbc7ac292),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd06df9),
	.w1(32'h3c8aaddb),
	.w2(32'hbc8aeed6),
	.w3(32'hbcaa2855),
	.w4(32'h3cbc6357),
	.w5(32'hbb7aa441),
	.w6(32'h3c13b50d),
	.w7(32'h39f73ae7),
	.w8(32'hbbe3d79f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5e852),
	.w1(32'hbba751ad),
	.w2(32'hbc86a4dc),
	.w3(32'hbcd1e5c8),
	.w4(32'hba9a3089),
	.w5(32'hbc3d7803),
	.w6(32'h3a05ba11),
	.w7(32'hbb89318a),
	.w8(32'h3bb3f6f6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba9076),
	.w1(32'hbb12432a),
	.w2(32'hbc6723b1),
	.w3(32'h3ad437fd),
	.w4(32'hbc064eb1),
	.w5(32'hbc6940c2),
	.w6(32'h3be88621),
	.w7(32'hbb815d91),
	.w8(32'h3aadbb50),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b06974),
	.w1(32'hbbb3b296),
	.w2(32'h3c1b1110),
	.w3(32'h3b9803b8),
	.w4(32'hbb40a7f6),
	.w5(32'h3c2e3ce7),
	.w6(32'hbbab322b),
	.w7(32'h3b654ef4),
	.w8(32'h3b70dd60),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a835),
	.w1(32'hbbc16d8c),
	.w2(32'hbc07e06f),
	.w3(32'h3ba77b22),
	.w4(32'h3a26d152),
	.w5(32'hbc23673d),
	.w6(32'hbb041db9),
	.w7(32'hbb2e3b5d),
	.w8(32'h3b76ae66),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3501d),
	.w1(32'hbbc2e5cc),
	.w2(32'hbc033168),
	.w3(32'h3b4ea8b8),
	.w4(32'hbac2898c),
	.w5(32'hbc324d83),
	.w6(32'hbb8868cf),
	.w7(32'hbb14f3e0),
	.w8(32'h3b03d642),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a5b39),
	.w1(32'hbbe33c08),
	.w2(32'hbc8ebb15),
	.w3(32'hbb07f5ab),
	.w4(32'h3bb25e86),
	.w5(32'hbbf3a562),
	.w6(32'hbbf361c1),
	.w7(32'hbbcb8419),
	.w8(32'h3c358fdd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44d3d5),
	.w1(32'h3b7710c4),
	.w2(32'hbb27dd27),
	.w3(32'hba8aec7a),
	.w4(32'hbaa01c15),
	.w5(32'hba635b68),
	.w6(32'h3c0f95ce),
	.w7(32'hbb81908a),
	.w8(32'hbb67250a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06095a),
	.w1(32'h3c511fd3),
	.w2(32'hbafccda2),
	.w3(32'hbb7ff3d1),
	.w4(32'h3c48eaa4),
	.w5(32'hbbdc197f),
	.w6(32'h3c152b47),
	.w7(32'h3a110858),
	.w8(32'hbbaaadac),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58fe02),
	.w1(32'h3c33a631),
	.w2(32'h3b8700eb),
	.w3(32'hbc4eed5c),
	.w4(32'h3b3cab66),
	.w5(32'hbbc96ea5),
	.w6(32'hbb2affbf),
	.w7(32'hbb87a5e9),
	.w8(32'hbb0fbf74),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e1640),
	.w1(32'hbb063dff),
	.w2(32'hbae33204),
	.w3(32'hbb8f540a),
	.w4(32'hbaa7d84f),
	.w5(32'h39cd58cf),
	.w6(32'hbbb4032a),
	.w7(32'hbbdc0ccc),
	.w8(32'hbb11aae7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4663d),
	.w1(32'hbc2c31d1),
	.w2(32'hbc1bb3e8),
	.w3(32'h3b95485b),
	.w4(32'hbc4efa6b),
	.w5(32'hbc250ead),
	.w6(32'h3a9dd14a),
	.w7(32'hbbf4cec4),
	.w8(32'hbc135920),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d2954),
	.w1(32'h3be92299),
	.w2(32'hbbde4faa),
	.w3(32'hbb148833),
	.w4(32'h3b1ea510),
	.w5(32'hbc5dcb3f),
	.w6(32'h3bdb721a),
	.w7(32'hb96224b8),
	.w8(32'h39ee1db8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7974),
	.w1(32'h3ca08fae),
	.w2(32'h3c47f09c),
	.w3(32'hbc1b895b),
	.w4(32'h3c96b5fb),
	.w5(32'h3bb18f42),
	.w6(32'h3c333fe8),
	.w7(32'h39c79f4f),
	.w8(32'hba0707c7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ad848),
	.w1(32'hbbd3ee1a),
	.w2(32'hba40dd23),
	.w3(32'hbc423cd2),
	.w4(32'hbb7e27a5),
	.w5(32'hb91d0306),
	.w6(32'hbbbd9f7d),
	.w7(32'h3b52c835),
	.w8(32'h3c0f86ae),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba66934),
	.w1(32'hbb9c738b),
	.w2(32'h3a462b4b),
	.w3(32'h3b34a963),
	.w4(32'h38ef60c2),
	.w5(32'h3aa4725b),
	.w6(32'hbb19f626),
	.w7(32'h3b801a71),
	.w8(32'h3bcd0bc4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d0d55),
	.w1(32'hbafe56b1),
	.w2(32'hbb598f9c),
	.w3(32'h3c044778),
	.w4(32'hbbca8618),
	.w5(32'hbb68540f),
	.w6(32'h3b19284d),
	.w7(32'h3bc96875),
	.w8(32'h3bccd20c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bda91),
	.w1(32'h3c9cfbfc),
	.w2(32'hbc3c3c4c),
	.w3(32'hbba6d0c7),
	.w4(32'h3cbe0fe7),
	.w5(32'h3b99f8fa),
	.w6(32'hbba8ad7d),
	.w7(32'hbc5d9d63),
	.w8(32'h3b31f539),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2d24),
	.w1(32'h3c803c4c),
	.w2(32'hbc362f14),
	.w3(32'hbb42dc7a),
	.w4(32'h3cbb3467),
	.w5(32'hbbdb633d),
	.w6(32'h3bd6fb36),
	.w7(32'hbb71840e),
	.w8(32'hbc2ce261),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9652e7),
	.w1(32'h3c96befc),
	.w2(32'h3b20d33f),
	.w3(32'hbca16f9a),
	.w4(32'h3b4c01c7),
	.w5(32'h3a236eb3),
	.w6(32'h3bfdc120),
	.w7(32'h3a00389a),
	.w8(32'hbb786178),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9491f0),
	.w1(32'hbaec76e3),
	.w2(32'hba898142),
	.w3(32'hbb6d4fb2),
	.w4(32'hbae5c278),
	.w5(32'hbb2d079e),
	.w6(32'h3a0a0ad7),
	.w7(32'h39444526),
	.w8(32'hbad5703f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3353b5),
	.w1(32'h3b840c26),
	.w2(32'h3a0489e6),
	.w3(32'hbb2db130),
	.w4(32'h3b71b5ee),
	.w5(32'h3a7abf30),
	.w6(32'hbb5a51a9),
	.w7(32'hbb626d3a),
	.w8(32'hbba523d1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c745),
	.w1(32'h3c91fdec),
	.w2(32'h3bc73bbe),
	.w3(32'hb9e5d315),
	.w4(32'h3c6b5e88),
	.w5(32'h3c8f0b30),
	.w6(32'h3c915c1b),
	.w7(32'hb9795d8c),
	.w8(32'hbc853c10),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dff1a),
	.w1(32'hbb269b54),
	.w2(32'h39eaa2b4),
	.w3(32'hbb988632),
	.w4(32'hbbe67eeb),
	.w5(32'hbb639092),
	.w6(32'h3ad27595),
	.w7(32'h3b508561),
	.w8(32'h3bb56469),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba97cc8),
	.w1(32'h3bba94a0),
	.w2(32'hbb0de107),
	.w3(32'h3b65af83),
	.w4(32'h3c2813a6),
	.w5(32'h3b35dcf1),
	.w6(32'hbbac3128),
	.w7(32'hbbcaa8e9),
	.w8(32'hbbbc0a4d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dd430),
	.w1(32'hbc69e54d),
	.w2(32'h3b769961),
	.w3(32'h3b7c8abc),
	.w4(32'h3a875327),
	.w5(32'h3b072f70),
	.w6(32'hbc2a831d),
	.w7(32'hbc0358c2),
	.w8(32'hbb88e1f4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc165155),
	.w1(32'hbbc91d64),
	.w2(32'hbbb18d59),
	.w3(32'hbb02d616),
	.w4(32'h3b833406),
	.w5(32'hbb8df955),
	.w6(32'hbb0e4791),
	.w7(32'hbbce1ecd),
	.w8(32'hbbd9f4be),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08eeb7),
	.w1(32'hbc933644),
	.w2(32'hbc8887ca),
	.w3(32'hbb81f9ef),
	.w4(32'hbcbf1b9c),
	.w5(32'hbc90028c),
	.w6(32'hbbba5793),
	.w7(32'h3ae1fede),
	.w8(32'h3b74a3da),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3817),
	.w1(32'hbd382e92),
	.w2(32'hbcec7f5e),
	.w3(32'h3aa43ff3),
	.w4(32'hbd1abd94),
	.w5(32'hbd11ab84),
	.w6(32'hbc57e322),
	.w7(32'hbaabdfca),
	.w8(32'h3bd6f988),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44b33c),
	.w1(32'hbc3232f0),
	.w2(32'h3ba88974),
	.w3(32'hba96686f),
	.w4(32'hbc43e458),
	.w5(32'h3b1bf5c6),
	.w6(32'hbad08995),
	.w7(32'h3c127258),
	.w8(32'h3c04131d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c7f2f),
	.w1(32'h3c1dd8e2),
	.w2(32'h3c0e3182),
	.w3(32'h3c2410cf),
	.w4(32'h3b70dda1),
	.w5(32'h3b160964),
	.w6(32'h3ba2cf07),
	.w7(32'h3b7ddf06),
	.w8(32'hb87042cb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc137a1e),
	.w1(32'h3bdb95cf),
	.w2(32'hbc308bd6),
	.w3(32'hbc668b68),
	.w4(32'h3c4da503),
	.w5(32'h3aa945f1),
	.w6(32'hbb375c74),
	.w7(32'hbca30723),
	.w8(32'hbbd8dbc0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027e6f),
	.w1(32'h3c58a32d),
	.w2(32'hbbe39626),
	.w3(32'hbb9698fb),
	.w4(32'h3c7a1830),
	.w5(32'hbb01aa36),
	.w6(32'h398413f1),
	.w7(32'hbc1e1a28),
	.w8(32'hbc31eda5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c324a),
	.w1(32'h3a107c19),
	.w2(32'hbc15af5f),
	.w3(32'hbbeb83e0),
	.w4(32'h3b0b98d6),
	.w5(32'hbb953d30),
	.w6(32'hb86e25e1),
	.w7(32'hbbb57947),
	.w8(32'hbb72e092),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad3f52),
	.w1(32'hbbb19da7),
	.w2(32'hbb9f506c),
	.w3(32'hba8f77eb),
	.w4(32'hbb8c7fa1),
	.w5(32'hbbb202c4),
	.w6(32'hbbbe1ccd),
	.w7(32'h3b569b5a),
	.w8(32'h3b40635a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e03d1),
	.w1(32'hbc6590d4),
	.w2(32'hbc2af3b3),
	.w3(32'hbb39a896),
	.w4(32'hbc0fbd68),
	.w5(32'hbb5029c5),
	.w6(32'hbc19d903),
	.w7(32'hbb8e1eb4),
	.w8(32'h3abd8ffa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5571),
	.w1(32'h3bfb9f55),
	.w2(32'h3b61b270),
	.w3(32'hb9d8be5d),
	.w4(32'h3bd3c041),
	.w5(32'h3b656f11),
	.w6(32'h3c124893),
	.w7(32'hb9a54edd),
	.w8(32'hba8b4313),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85b0e2),
	.w1(32'h3af3f959),
	.w2(32'hba160074),
	.w3(32'h3a5c3125),
	.w4(32'h3b5ee13f),
	.w5(32'h3853a9c1),
	.w6(32'hba6ac9c7),
	.w7(32'hbb932545),
	.w8(32'hbbabc42b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb116be2),
	.w1(32'h3c4e4686),
	.w2(32'h3b22e205),
	.w3(32'hbaf97643),
	.w4(32'h3bf8ede3),
	.w5(32'hbb20fa55),
	.w6(32'hbb7bd283),
	.w7(32'h3bd9f51e),
	.w8(32'hbc5ad81c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2df9ee),
	.w1(32'hbb3adf8e),
	.w2(32'h3ae93e8f),
	.w3(32'hbc6e8335),
	.w4(32'hba6c8aa1),
	.w5(32'h3a3fe624),
	.w6(32'hbb9123d9),
	.w7(32'hbadd63d2),
	.w8(32'h37543fa5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b166541),
	.w1(32'hbb761e50),
	.w2(32'hbc0a52fb),
	.w3(32'h3b915799),
	.w4(32'hbb812598),
	.w5(32'hbc2839d7),
	.w6(32'h3968dd72),
	.w7(32'hbc260608),
	.w8(32'hbc651aba),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88deba),
	.w1(32'h3b69e088),
	.w2(32'hbb450172),
	.w3(32'hbb94ec39),
	.w4(32'h3b6228f6),
	.w5(32'h3b765f4b),
	.w6(32'h3c2e7eaf),
	.w7(32'hbc26d239),
	.w8(32'hbc1ffe93),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944a7f),
	.w1(32'hbb253465),
	.w2(32'hbb6053f4),
	.w3(32'hbbfd0eef),
	.w4(32'h3afbf100),
	.w5(32'hbabfdf9c),
	.w6(32'h3a96d48d),
	.w7(32'h3b4eb4ab),
	.w8(32'h3c47c917),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2c88),
	.w1(32'hb9c72886),
	.w2(32'h3a6d8acd),
	.w3(32'h3ab51470),
	.w4(32'h3b2c3849),
	.w5(32'h3a3b97bc),
	.w6(32'hbada99cb),
	.w7(32'hbadf523d),
	.w8(32'h39eced58),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f310c),
	.w1(32'h3b8711cb),
	.w2(32'h3bb04ec1),
	.w3(32'h3b67afc7),
	.w4(32'hbb33c804),
	.w5(32'h3a64d31c),
	.w6(32'h3aa89ef1),
	.w7(32'h3b54c068),
	.w8(32'h3c25de12),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56d873),
	.w1(32'hbb1a2adf),
	.w2(32'hbb90c1b4),
	.w3(32'h3c29d5d8),
	.w4(32'h3a223c67),
	.w5(32'hbba1d7ad),
	.w6(32'hbb44a110),
	.w7(32'hbc0542bc),
	.w8(32'h395a7a44),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9290eb),
	.w1(32'hbbd3562d),
	.w2(32'h3b79b2be),
	.w3(32'h371439e0),
	.w4(32'hbb9ed907),
	.w5(32'hbb5cb810),
	.w6(32'hb929eaa0),
	.w7(32'hbaed2771),
	.w8(32'h3b18a271),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae58cb3),
	.w1(32'h3bb2862a),
	.w2(32'hbb3f869d),
	.w3(32'hbc1ef7a0),
	.w4(32'h3b9755df),
	.w5(32'hbbba707d),
	.w6(32'h3b5d1de9),
	.w7(32'hb862bbf7),
	.w8(32'h3b4c07a3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1514f3),
	.w1(32'h3b734d8a),
	.w2(32'hbbcbfb34),
	.w3(32'h3af69ae5),
	.w4(32'h3aff313e),
	.w5(32'hbbe98534),
	.w6(32'h3c0171a9),
	.w7(32'hbc2129eb),
	.w8(32'hbab1e30a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05a37),
	.w1(32'hbc0076d7),
	.w2(32'hbc270013),
	.w3(32'hba93c3a7),
	.w4(32'h3b94878e),
	.w5(32'hbc27ad7f),
	.w6(32'hbb796fe1),
	.w7(32'hbb70ba73),
	.w8(32'h3ad1d933),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27a516),
	.w1(32'h3b02eb6f),
	.w2(32'h39ba29b4),
	.w3(32'hbbdb68db),
	.w4(32'h3b376c91),
	.w5(32'hba295b92),
	.w6(32'hbb1474b4),
	.w7(32'hbb78674e),
	.w8(32'hbc1486a2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e32a5),
	.w1(32'hbb1d535f),
	.w2(32'hbc133938),
	.w3(32'hbaea72db),
	.w4(32'h39577f83),
	.w5(32'hbba52aa3),
	.w6(32'hbb80f6af),
	.w7(32'hbc2531cd),
	.w8(32'hbb020028),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3435c8),
	.w1(32'h3c19974b),
	.w2(32'hbc455464),
	.w3(32'hbb9728b2),
	.w4(32'h3b24326d),
	.w5(32'hbc692c03),
	.w6(32'h3b04a9c9),
	.w7(32'hbb0443aa),
	.w8(32'hbb9d3a43),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f09a3),
	.w1(32'h3c877a6b),
	.w2(32'hbc11c099),
	.w3(32'hbbb861b6),
	.w4(32'h3c7126ca),
	.w5(32'h3bbd55c6),
	.w6(32'h3b59f1f6),
	.w7(32'hbc1b5f71),
	.w8(32'hbc773a0b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81bf8f),
	.w1(32'h3b5a35e5),
	.w2(32'h3d17c1cf),
	.w3(32'h39b3affa),
	.w4(32'hbb24386a),
	.w5(32'h3c8417e2),
	.w6(32'hbb7e55c1),
	.w7(32'h3c236a63),
	.w8(32'hb588de7a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30b697),
	.w1(32'hbb08d7c5),
	.w2(32'h3b23c138),
	.w3(32'h3a095889),
	.w4(32'hbb4a42a6),
	.w5(32'hba0f6191),
	.w6(32'hbae0d97c),
	.w7(32'hba4e7a50),
	.w8(32'hbbf0d66f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule