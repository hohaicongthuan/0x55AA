module layer_10_featuremap_75(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc985581),
	.w1(32'hbb4668f8),
	.w2(32'h38374f99),
	.w3(32'h3a1e3f02),
	.w4(32'hbc5e540f),
	.w5(32'hb98ff64a),
	.w6(32'h3bee06a5),
	.w7(32'hbca08ed2),
	.w8(32'hbb3e23d6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c595620),
	.w1(32'h3b4b20aa),
	.w2(32'h3a96b1ea),
	.w3(32'h3c7b1c39),
	.w4(32'hbbfe0969),
	.w5(32'h3c0e7a14),
	.w6(32'h3c015c0c),
	.w7(32'h3c277578),
	.w8(32'hbb3616c5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd94abe),
	.w1(32'h3ca784b5),
	.w2(32'hbb74a044),
	.w3(32'hbcde6820),
	.w4(32'h3c3fff92),
	.w5(32'hbbb085fa),
	.w6(32'h3aa711b8),
	.w7(32'hbca60ae8),
	.w8(32'h39ec6607),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9a0f),
	.w1(32'hbb8eae9a),
	.w2(32'h3b83f702),
	.w3(32'hbbc66e63),
	.w4(32'hbc4786fa),
	.w5(32'h3c1a587d),
	.w6(32'hbc4465b4),
	.w7(32'hbbb8b1e1),
	.w8(32'h3c19422a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4aea1),
	.w1(32'h3c494ef2),
	.w2(32'h3ccc0920),
	.w3(32'hbac99558),
	.w4(32'h3c723785),
	.w5(32'h3ce1541a),
	.w6(32'h3c168625),
	.w7(32'h39d47220),
	.w8(32'h3c0de2f2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c9a88),
	.w1(32'h3c93cdf4),
	.w2(32'hbba7f175),
	.w3(32'h3d525542),
	.w4(32'hb9a7bb98),
	.w5(32'hba45bf5d),
	.w6(32'h3d8edb47),
	.w7(32'hbbb56ec5),
	.w8(32'hba908369),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251be7),
	.w1(32'hbb224084),
	.w2(32'h3b6a4a62),
	.w3(32'h3b176f55),
	.w4(32'hbab8a19b),
	.w5(32'h3b2ad413),
	.w6(32'h3b7a7430),
	.w7(32'hb9349e84),
	.w8(32'h3b455b9b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7507de),
	.w1(32'hbc1124af),
	.w2(32'hbc6b04bd),
	.w3(32'hbb961c5f),
	.w4(32'hbbd7d397),
	.w5(32'hbbf2c907),
	.w6(32'h3a38eed5),
	.w7(32'h3a2131b0),
	.w8(32'hbb7668ec),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97fdb8),
	.w1(32'h3ba10204),
	.w2(32'h3ac87d8b),
	.w3(32'hbbd887ef),
	.w4(32'h3c261181),
	.w5(32'hba5ce788),
	.w6(32'hbcaf2be1),
	.w7(32'h3bf38306),
	.w8(32'hb881c678),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a9f7),
	.w1(32'hba440818),
	.w2(32'h3becf6dd),
	.w3(32'h3bb8b182),
	.w4(32'h3b7e357f),
	.w5(32'hbaee91e7),
	.w6(32'hbbd0a5cb),
	.w7(32'h3bf84353),
	.w8(32'hbafe9045),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae1bfe),
	.w1(32'hba953b48),
	.w2(32'h3b96002a),
	.w3(32'hbad0269c),
	.w4(32'hbb682e97),
	.w5(32'h3c3264d8),
	.w6(32'h3b2c78da),
	.w7(32'hbb5f03bd),
	.w8(32'h3b7a7729),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16ef2b),
	.w1(32'hbb9b6e46),
	.w2(32'hbba62b80),
	.w3(32'hbc6af27b),
	.w4(32'hbc3b5def),
	.w5(32'hbafede28),
	.w6(32'hbb29bab0),
	.w7(32'hbc121c2e),
	.w8(32'hbbb21a6a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f38a5),
	.w1(32'h3b8910a6),
	.w2(32'h3b75644e),
	.w3(32'h3b11f5ff),
	.w4(32'hba144d64),
	.w5(32'hbb7f04c1),
	.w6(32'hbaf8279f),
	.w7(32'hbb368640),
	.w8(32'hbb0b27ad),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c441bf4),
	.w1(32'h3b4e4e51),
	.w2(32'hbb367cab),
	.w3(32'h3ba49e1e),
	.w4(32'h3b53ffb1),
	.w5(32'h3ba5257a),
	.w6(32'h3c3dffc0),
	.w7(32'h3c09345e),
	.w8(32'h39b6056d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ebcc3),
	.w1(32'h3c093f06),
	.w2(32'h3b6438cf),
	.w3(32'h3b9bfb66),
	.w4(32'hbb8567a7),
	.w5(32'hbbfe079e),
	.w6(32'h3aab74fa),
	.w7(32'hbc26e729),
	.w8(32'hbbf34aa0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf3a0),
	.w1(32'hbbcfad0a),
	.w2(32'hba7134bb),
	.w3(32'h3b3ec524),
	.w4(32'hbc680220),
	.w5(32'h3901e2aa),
	.w6(32'h3ab15be4),
	.w7(32'hbc07573c),
	.w8(32'hbad28f96),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2454ae),
	.w1(32'hba903b44),
	.w2(32'h3a57e71f),
	.w3(32'hbae8f9f2),
	.w4(32'hbb07dce2),
	.w5(32'h3bbfd5af),
	.w6(32'h3aa51b86),
	.w7(32'hbb7aeaf2),
	.w8(32'hb9080bde),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce63b93),
	.w1(32'hbd071906),
	.w2(32'hbbd3b9c7),
	.w3(32'hbcaf9f2b),
	.w4(32'hbcd91340),
	.w5(32'hbb06341e),
	.w6(32'hbc08cdcd),
	.w7(32'hbbdeb936),
	.w8(32'hbb7e3369),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dad0a),
	.w1(32'hbb7cdbc9),
	.w2(32'hbc428021),
	.w3(32'hbb327a7b),
	.w4(32'hbbbfd37f),
	.w5(32'hbc4025f7),
	.w6(32'hbb88f025),
	.w7(32'h3b23d13f),
	.w8(32'hbc0bf591),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba724831),
	.w1(32'hbacf69f7),
	.w2(32'hba63858c),
	.w3(32'hbc498a5a),
	.w4(32'hbc4617c5),
	.w5(32'hbaf6872a),
	.w6(32'hbcb80705),
	.w7(32'hbb2d7a0c),
	.w8(32'hba825ff0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bc71e),
	.w1(32'hbb6fe50f),
	.w2(32'hbb603af3),
	.w3(32'h3b0ed728),
	.w4(32'hbb5378f3),
	.w5(32'hbca834e1),
	.w6(32'h3b8e42ab),
	.w7(32'hb9ddb3e5),
	.w8(32'hbb8b21a5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98458b),
	.w1(32'hbc1ba5a3),
	.w2(32'h3bc0e50c),
	.w3(32'h3b9ec9ce),
	.w4(32'hbbb38d88),
	.w5(32'h3ad0eaec),
	.w6(32'hbc808509),
	.w7(32'h3c469f4d),
	.w8(32'hbc433b24),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf1faae),
	.w1(32'hbcd9542d),
	.w2(32'hbabc3e92),
	.w3(32'hbcbb2659),
	.w4(32'hbcc643a6),
	.w5(32'h3c13a994),
	.w6(32'hbc7d508e),
	.w7(32'hbc85c0d1),
	.w8(32'h3c4c0c77),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911f63),
	.w1(32'hb9e8b04d),
	.w2(32'h3c5f4413),
	.w3(32'hba0ac07f),
	.w4(32'hba2ab1ea),
	.w5(32'h3b7b64f1),
	.w6(32'hbbda5f9f),
	.w7(32'hbbfbd58d),
	.w8(32'h3b35685a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d474a),
	.w1(32'h3bfe8a77),
	.w2(32'h3c4f7f14),
	.w3(32'h3c1d2bde),
	.w4(32'h3b57e972),
	.w5(32'h3c85e3e1),
	.w6(32'h3b923c2c),
	.w7(32'hbadd4275),
	.w8(32'h3c1ca021),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba7bf5),
	.w1(32'h3bf11d4b),
	.w2(32'h3b6768d2),
	.w3(32'h3a547b6c),
	.w4(32'h3d121534),
	.w5(32'hb9ea777c),
	.w6(32'h3a545cd9),
	.w7(32'h3c9219f4),
	.w8(32'hbbed66fa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf77c14),
	.w1(32'h3a1ee835),
	.w2(32'h3b46063e),
	.w3(32'hbc0ed864),
	.w4(32'hbb041746),
	.w5(32'h3b65358d),
	.w6(32'hbb8a66ef),
	.w7(32'hbc4bc30c),
	.w8(32'h3b2b4340),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c6c8),
	.w1(32'h3be17d76),
	.w2(32'hbb6405b2),
	.w3(32'h3c03edad),
	.w4(32'h3b9d9ac8),
	.w5(32'hbc187191),
	.w6(32'h3b9e7965),
	.w7(32'h3a8bfad6),
	.w8(32'hbbfd5dad),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffd298),
	.w1(32'h388ba308),
	.w2(32'hbb525917),
	.w3(32'hbc1ee334),
	.w4(32'hbb3387d2),
	.w5(32'h3b16a4ee),
	.w6(32'hbabb006a),
	.w7(32'hb910ef96),
	.w8(32'hbb0b3358),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3ed68),
	.w1(32'h3bc046bd),
	.w2(32'h3c159699),
	.w3(32'h3c7992fc),
	.w4(32'h3c6d8064),
	.w5(32'h3bb1758d),
	.w6(32'h3bb01227),
	.w7(32'h3c5210c5),
	.w8(32'h3bf1bc03),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf163d6),
	.w1(32'h3bcf57e4),
	.w2(32'hbafe01d5),
	.w3(32'h3c6129fe),
	.w4(32'h3c474df2),
	.w5(32'h3bb810ff),
	.w6(32'h3c7e5d95),
	.w7(32'h3c08ab53),
	.w8(32'h3c176f9a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed7df),
	.w1(32'h3c83630f),
	.w2(32'hba7c3eb3),
	.w3(32'h3c81caa0),
	.w4(32'h3c893a8e),
	.w5(32'hbbc77f75),
	.w6(32'h3c77588f),
	.w7(32'h3c2388e0),
	.w8(32'hbab39efe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f4d0a),
	.w1(32'h3c0ed149),
	.w2(32'h3be3d968),
	.w3(32'h3c18af2a),
	.w4(32'h3c5101e7),
	.w5(32'hbb867c9a),
	.w6(32'hbb9f8ebe),
	.w7(32'h3c0434cd),
	.w8(32'hbbd3a85b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4adb0),
	.w1(32'hba30dced),
	.w2(32'hbad21848),
	.w3(32'hbbfdcfd9),
	.w4(32'hbb62f6b9),
	.w5(32'h3aa55d9b),
	.w6(32'hbc363ae3),
	.w7(32'hbb783cbd),
	.w8(32'hbb229ad3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5e30),
	.w1(32'hba2443c3),
	.w2(32'hbba3b59d),
	.w3(32'h3c09788a),
	.w4(32'h3acc0cf8),
	.w5(32'hbc5b8f3c),
	.w6(32'h3c1a7537),
	.w7(32'h3b87c0d3),
	.w8(32'hbc814224),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65da04),
	.w1(32'hbc624dea),
	.w2(32'hbca155de),
	.w3(32'hbc9a34e5),
	.w4(32'hbcb35f4f),
	.w5(32'hbc3d159a),
	.w6(32'hbca7ea3e),
	.w7(32'hbc898ebf),
	.w8(32'h3a5cc39d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f69e0),
	.w1(32'hbbaf8bd1),
	.w2(32'hbba8bde3),
	.w3(32'h3aa429df),
	.w4(32'h3b52f58a),
	.w5(32'h3ae833ae),
	.w6(32'h3c9b0069),
	.w7(32'h3cab2b9b),
	.w8(32'hbb4785f1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc23e18),
	.w1(32'h3c7522bc),
	.w2(32'hbb751876),
	.w3(32'h3cd17c07),
	.w4(32'h3c4caa2a),
	.w5(32'hbcc85890),
	.w6(32'h3c8efed6),
	.w7(32'h3ba09429),
	.w8(32'hbc9106a4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc002aa9),
	.w1(32'h3afeff43),
	.w2(32'h3ac603ca),
	.w3(32'h3c260101),
	.w4(32'h3c17e410),
	.w5(32'hbca451c4),
	.w6(32'h3b9a9b24),
	.w7(32'h3b515c5c),
	.w8(32'hbcaad142),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d2785),
	.w1(32'h3c37b898),
	.w2(32'hbbe1c08e),
	.w3(32'h3c057a31),
	.w4(32'h3c8a6967),
	.w5(32'hbc8dd927),
	.w6(32'h3a03f9d8),
	.w7(32'h3b9f2dae),
	.w8(32'hbc272d62),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f870c),
	.w1(32'hba19e3a6),
	.w2(32'hbbc1e06b),
	.w3(32'hbc9e6993),
	.w4(32'hbbd2c35d),
	.w5(32'h3a8f6d64),
	.w6(32'hbbc9bc81),
	.w7(32'h3bdbfab1),
	.w8(32'hbab13e69),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e6f0),
	.w1(32'hbbfc774d),
	.w2(32'hba1b6959),
	.w3(32'h3bf99c3d),
	.w4(32'h3c051992),
	.w5(32'hbb5a0a49),
	.w6(32'hb88effaf),
	.w7(32'hbb8f9e32),
	.w8(32'h3af2b55d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85d3b9),
	.w1(32'h3bdb714d),
	.w2(32'hbb419899),
	.w3(32'hbc5ce416),
	.w4(32'hb97ca652),
	.w5(32'hb9dfc07e),
	.w6(32'hbbef1e2f),
	.w7(32'hbb4b0f2f),
	.w8(32'hb9ad7a87),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a37694),
	.w1(32'h3b63db73),
	.w2(32'h3c8951b3),
	.w3(32'hba94c19e),
	.w4(32'h3a5c00b5),
	.w5(32'h3ce8500d),
	.w6(32'hbb7dc27b),
	.w7(32'hb9ec6f3d),
	.w8(32'h3c29dbec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c536cad),
	.w1(32'h3c3913b5),
	.w2(32'h3c499818),
	.w3(32'h3ceccb1d),
	.w4(32'hba6af3c0),
	.w5(32'hbb7056c0),
	.w6(32'h3c015b59),
	.w7(32'hbb8b5ce3),
	.w8(32'hbc419aae),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe204),
	.w1(32'hbc221f12),
	.w2(32'h3c550ffb),
	.w3(32'hbb802c84),
	.w4(32'hbc84b77a),
	.w5(32'h3c317d74),
	.w6(32'hbc84c5bc),
	.w7(32'hbc229a5e),
	.w8(32'h3b433551),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019423),
	.w1(32'h3b8f7cf9),
	.w2(32'h394a5dfa),
	.w3(32'h3bdcf640),
	.w4(32'hbc006b50),
	.w5(32'h3bda5336),
	.w6(32'hbbf50b3d),
	.w7(32'hbc31bb6b),
	.w8(32'h3c76685d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95a6e6),
	.w1(32'hbcd5d639),
	.w2(32'hbc4f842c),
	.w3(32'hbc0ff7bb),
	.w4(32'hbcb4bd15),
	.w5(32'h3bd80bd6),
	.w6(32'hbb6dab12),
	.w7(32'h39d2bd18),
	.w8(32'h3b230e4f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9f03),
	.w1(32'h3bd927c9),
	.w2(32'h3a8a695c),
	.w3(32'h3c29c047),
	.w4(32'h3c083416),
	.w5(32'h3b7b6eed),
	.w6(32'h3bd2600b),
	.w7(32'h3bea9d18),
	.w8(32'h3c1cf8ea),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77e06f),
	.w1(32'h3c5e9da6),
	.w2(32'h396c1236),
	.w3(32'hbb1dcdda),
	.w4(32'h3be9eb4e),
	.w5(32'h3bb70606),
	.w6(32'hbc10f5cc),
	.w7(32'hb97348ce),
	.w8(32'h3b40e803),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4757b0),
	.w1(32'h3c05855c),
	.w2(32'hbb9b8228),
	.w3(32'h3c705022),
	.w4(32'h3c8a76a0),
	.w5(32'h3baecc95),
	.w6(32'h3c39ea63),
	.w7(32'h3b8c6691),
	.w8(32'hbacc39d5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc5509),
	.w1(32'h3a2efa4e),
	.w2(32'hbbede987),
	.w3(32'h3b9e8746),
	.w4(32'h3c0cffe2),
	.w5(32'hbb053798),
	.w6(32'h3b398b7d),
	.w7(32'hba957b91),
	.w8(32'hbb3ffa33),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0855),
	.w1(32'hb9effef0),
	.w2(32'hbc8f79d6),
	.w3(32'h3c025c81),
	.w4(32'hbae5e73d),
	.w5(32'hbbd8d769),
	.w6(32'hba51b510),
	.w7(32'hbc222732),
	.w8(32'hbb86d607),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c980f),
	.w1(32'hbcd5f3bc),
	.w2(32'hbc623b35),
	.w3(32'hbcb54f0a),
	.w4(32'hbcb98c39),
	.w5(32'hbc0b1ca7),
	.w6(32'hbc63e468),
	.w7(32'hbc256038),
	.w8(32'h39fc0c5c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca40843),
	.w1(32'hbb2fa06a),
	.w2(32'hbbd7f999),
	.w3(32'hbba3b634),
	.w4(32'h3ba84bfd),
	.w5(32'h3c3aa6df),
	.w6(32'h3cbb2d21),
	.w7(32'h3ca3d778),
	.w8(32'h3c11f18d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb87d50),
	.w1(32'h3ad13034),
	.w2(32'h3b950e30),
	.w3(32'h3c98bc3c),
	.w4(32'h3c320ce8),
	.w5(32'hbba4a840),
	.w6(32'h3c822493),
	.w7(32'h3c43e497),
	.w8(32'h3b089634),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97f9fd),
	.w1(32'h3c8941f6),
	.w2(32'hbbb6455a),
	.w3(32'h3b550712),
	.w4(32'h3c37ecca),
	.w5(32'hbabaf999),
	.w6(32'hbba47ff8),
	.w7(32'h3c1b8b9f),
	.w8(32'hbbb6984f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6126c),
	.w1(32'hbacbf130),
	.w2(32'hbb8c3a01),
	.w3(32'hb78643be),
	.w4(32'h3abf6178),
	.w5(32'hbbc30152),
	.w6(32'hbab5c8a3),
	.w7(32'hbb04d355),
	.w8(32'hbc199b14),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e984),
	.w1(32'hbbce87b6),
	.w2(32'hbb51f6b1),
	.w3(32'hbba49055),
	.w4(32'hbbb92261),
	.w5(32'hbb896c22),
	.w6(32'hbbe23615),
	.w7(32'hbbe9f48e),
	.w8(32'hbbd96f6f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc218570),
	.w1(32'hbb91d32f),
	.w2(32'hbaaf6518),
	.w3(32'hbc21a241),
	.w4(32'hbbfb09de),
	.w5(32'h3c0614bb),
	.w6(32'hbaadfb74),
	.w7(32'hbc047f90),
	.w8(32'h3b523526),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc91a0),
	.w1(32'hbc0c112a),
	.w2(32'h3b6fcf04),
	.w3(32'h3bd2a59b),
	.w4(32'hbbc557a7),
	.w5(32'h3c9156c4),
	.w6(32'h3ae1401c),
	.w7(32'h3b2c5f0e),
	.w8(32'h3c6229f6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167f1a),
	.w1(32'h3c74353a),
	.w2(32'hbc9258a7),
	.w3(32'h3caf8a90),
	.w4(32'h3d073884),
	.w5(32'hbd300002),
	.w6(32'h3cc728bd),
	.w7(32'h3ce1ccb8),
	.w8(32'hbd02ee52),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b352e),
	.w1(32'hbd047a8a),
	.w2(32'hbb68beed),
	.w3(32'hbd9d8e7c),
	.w4(32'hbd5626ce),
	.w5(32'h3aef9842),
	.w6(32'hbd4f4ed6),
	.w7(32'hbd26918d),
	.w8(32'hbb66a6e9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c08dd1),
	.w1(32'hbbad7800),
	.w2(32'h3aa73b0e),
	.w3(32'h3bffcdaa),
	.w4(32'h3b4c8d6c),
	.w5(32'h3b15eed9),
	.w6(32'h3c1fc643),
	.w7(32'h3a9e46ca),
	.w8(32'hbad72051),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39200a5b),
	.w1(32'hbb20e0b7),
	.w2(32'hbb140c10),
	.w3(32'hba5f7eb8),
	.w4(32'hbb50074f),
	.w5(32'h3bccfb50),
	.w6(32'hbab88a99),
	.w7(32'hbb116a0b),
	.w8(32'h3b2b6180),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48631),
	.w1(32'hbab3459e),
	.w2(32'hbbcfb124),
	.w3(32'h3c7e3a6a),
	.w4(32'h3bbf978a),
	.w5(32'hbb4bca2f),
	.w6(32'h3be7775e),
	.w7(32'h37d1e8a0),
	.w8(32'hbb34682c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dafef3),
	.w1(32'hba578c66),
	.w2(32'hbba1d994),
	.w3(32'hba6a9544),
	.w4(32'h3b22579c),
	.w5(32'h3c0f5ab5),
	.w6(32'hba2f418c),
	.w7(32'hb8c66e9c),
	.w8(32'h3c259f13),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be83f87),
	.w1(32'h3bef7531),
	.w2(32'hbbbb45b0),
	.w3(32'h3c71b74b),
	.w4(32'h3bf373c7),
	.w5(32'hbcbaf20e),
	.w6(32'h3b9201eb),
	.w7(32'hbb8e6673),
	.w8(32'hbcda35bf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c08c5),
	.w1(32'hbd15bf8a),
	.w2(32'h3b835648),
	.w3(32'hbd2ede3d),
	.w4(32'hbcb0b31b),
	.w5(32'h3c22321e),
	.w6(32'hbce73d1b),
	.w7(32'hbcc42da9),
	.w8(32'h3c06d8d3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f8608),
	.w1(32'h3c47bf67),
	.w2(32'hbbefec6e),
	.w3(32'h3d02d04c),
	.w4(32'h3c915ea0),
	.w5(32'hbc4a294d),
	.w6(32'h3c9972cf),
	.w7(32'h3c0792aa),
	.w8(32'hbc37ca39),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68a915),
	.w1(32'h3beb42f8),
	.w2(32'hbb09830a),
	.w3(32'h3aeb365d),
	.w4(32'h3b016e92),
	.w5(32'h3b7158ab),
	.w6(32'h3bdd3438),
	.w7(32'h3b96cfe2),
	.w8(32'h3b049c02),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94a2e0),
	.w1(32'h3b9040f5),
	.w2(32'h3ab676cb),
	.w3(32'hbb5c7211),
	.w4(32'hba905e5c),
	.w5(32'hbb3d6624),
	.w6(32'hbbced2ad),
	.w7(32'hbc3a9b53),
	.w8(32'hbb32d877),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38cc7a),
	.w1(32'hbb261f88),
	.w2(32'hb9b0d756),
	.w3(32'hbc6852a5),
	.w4(32'hbc8e7018),
	.w5(32'h3c5c3b5b),
	.w6(32'hbca0be77),
	.w7(32'hbc490bf3),
	.w8(32'h3c475b5d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca31991),
	.w1(32'h3c8aea28),
	.w2(32'hba0dc55b),
	.w3(32'h3d31ab1a),
	.w4(32'h3d48496f),
	.w5(32'hbabffd2d),
	.w6(32'h3d2b5143),
	.w7(32'h3d04f8a4),
	.w8(32'h391137a4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77bf7c),
	.w1(32'h3a9b6235),
	.w2(32'hbc89e8a4),
	.w3(32'h3bd2a0ea),
	.w4(32'hbb31634d),
	.w5(32'hbd019324),
	.w6(32'h3b7b0f9f),
	.w7(32'hbb6fc9f6),
	.w8(32'hbcaabd01),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0358e1),
	.w1(32'hbd01d457),
	.w2(32'hbc0671f3),
	.w3(32'hbd6ae40f),
	.w4(32'hbd39851c),
	.w5(32'h3c0d84fd),
	.w6(32'hbd41f45a),
	.w7(32'hbcdf0ce2),
	.w8(32'h3bb3aca9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a8bd0),
	.w1(32'hbc09adca),
	.w2(32'hbc39b5c9),
	.w3(32'hba944c8d),
	.w4(32'hbca08095),
	.w5(32'h3ca43690),
	.w6(32'hbb5a8732),
	.w7(32'hbb9e1d3d),
	.w8(32'h3bfd06f8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbd080),
	.w1(32'h3c813679),
	.w2(32'h3b8ab46c),
	.w3(32'h3cb7b93f),
	.w4(32'h3c9c69c5),
	.w5(32'h3bbd1ec1),
	.w6(32'h3cef76c5),
	.w7(32'h3c073c25),
	.w8(32'h3c059b35),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3f720),
	.w1(32'h3c734d3f),
	.w2(32'h3b8d75b7),
	.w3(32'h3c7452ce),
	.w4(32'h3bbcea38),
	.w5(32'h3a6d839b),
	.w6(32'h3c20f202),
	.w7(32'h3c2fd358),
	.w8(32'h3b967227),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c1a0b),
	.w1(32'h3b034c77),
	.w2(32'hbb78f113),
	.w3(32'hbbaa799b),
	.w4(32'hbb3d6156),
	.w5(32'hbb5e33f2),
	.w6(32'hba761e6c),
	.w7(32'hbb2837a7),
	.w8(32'hbbd2a50b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8b16a),
	.w1(32'hbb3853bd),
	.w2(32'h3a938b77),
	.w3(32'h3bad5438),
	.w4(32'h3b891b6b),
	.w5(32'hbb81ce08),
	.w6(32'h3b98e839),
	.w7(32'hbaedbfcc),
	.w8(32'hbb575af3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba584b0a),
	.w1(32'hbc5f6946),
	.w2(32'hbbfef360),
	.w3(32'hbbef9799),
	.w4(32'hbc62371c),
	.w5(32'hbb647766),
	.w6(32'hbbbc44e4),
	.w7(32'hbc48bed0),
	.w8(32'hbb11b4b4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba90c8c),
	.w1(32'h3c423a25),
	.w2(32'h3b0aecab),
	.w3(32'h3c9087f3),
	.w4(32'h3ca5fb98),
	.w5(32'h3c0e0e61),
	.w6(32'h3c1ed53c),
	.w7(32'h3c491d2f),
	.w8(32'h3ca5ba78),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf79d),
	.w1(32'h3bf30594),
	.w2(32'hbc44c55a),
	.w3(32'h3c0c2b5d),
	.w4(32'hbb318140),
	.w5(32'hbcb87f5a),
	.w6(32'h3c78947f),
	.w7(32'hbb643dfa),
	.w8(32'hbc9f8396),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5b0e0),
	.w1(32'hbc59ad5d),
	.w2(32'h3afab093),
	.w3(32'hbd5de06b),
	.w4(32'hbd0bb552),
	.w5(32'hbc1c2a0f),
	.w6(32'hbce7ac42),
	.w7(32'hbca06f71),
	.w8(32'hbb3021c4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3928d),
	.w1(32'hbaf970a6),
	.w2(32'h3b6d2f0b),
	.w3(32'h3c1c74df),
	.w4(32'h3be55f69),
	.w5(32'h3b81ace6),
	.w6(32'h3c235bfe),
	.w7(32'hbb669307),
	.w8(32'h3b8db684),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa1db),
	.w1(32'h3b827ae2),
	.w2(32'hbb85d233),
	.w3(32'h3bc14926),
	.w4(32'hbb5bb4be),
	.w5(32'hbc1c5bcc),
	.w6(32'hba896db3),
	.w7(32'hbc4b8b29),
	.w8(32'hbab3a08b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667107),
	.w1(32'hba5fc721),
	.w2(32'hbaf17e5f),
	.w3(32'hbbe47b04),
	.w4(32'hbb04caa6),
	.w5(32'h3bf30437),
	.w6(32'hbb133cb2),
	.w7(32'h3b2fc9b1),
	.w8(32'h3abe4cfd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac8dd0),
	.w1(32'h3bb84b61),
	.w2(32'h39b48a93),
	.w3(32'h3c4ab0e5),
	.w4(32'h3c3be20a),
	.w5(32'hb98cf295),
	.w6(32'h3ba2050f),
	.w7(32'hbb9c50a6),
	.w8(32'hbb178883),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae99a6),
	.w1(32'hbc8bfb09),
	.w2(32'h3b8f4e0a),
	.w3(32'hbd0a97b0),
	.w4(32'hbc317c24),
	.w5(32'h3c865534),
	.w6(32'hbc2ad60d),
	.w7(32'h3a9a7ecf),
	.w8(32'hbb176c53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270181),
	.w1(32'hbc0e8cd0),
	.w2(32'hbbf88e34),
	.w3(32'hbb42d7b4),
	.w4(32'hbc5d0346),
	.w5(32'h3a67cc2c),
	.w6(32'hbc962cc1),
	.w7(32'hbc57d807),
	.w8(32'hbbdf54ba),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79f83b),
	.w1(32'hbcb55309),
	.w2(32'hbc065da0),
	.w3(32'hbc06b05b),
	.w4(32'hbcd6075a),
	.w5(32'hbc5fab73),
	.w6(32'hbc6354bd),
	.w7(32'hbcbaa4f6),
	.w8(32'hbaa76f97),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e1926),
	.w1(32'h3a9d7101),
	.w2(32'hbb842609),
	.w3(32'hbc20dd67),
	.w4(32'hbaa119e5),
	.w5(32'hbb1f75a4),
	.w6(32'hbbb328dc),
	.w7(32'hba3ef802),
	.w8(32'hbb5caa4a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864fe9),
	.w1(32'hba99952a),
	.w2(32'hbb974821),
	.w3(32'hbb3bdae8),
	.w4(32'h3a63cba0),
	.w5(32'hbc34bcb2),
	.w6(32'hb977b8d4),
	.w7(32'h3b8d66e2),
	.w8(32'hbc8e14f3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8009e9),
	.w1(32'hbc817adb),
	.w2(32'h3c1b58ba),
	.w3(32'hbce3c543),
	.w4(32'hbc8ea085),
	.w5(32'h3c798fa1),
	.w6(32'hbcae9fb8),
	.w7(32'hbc996019),
	.w8(32'h3c12bb30),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4faa04),
	.w1(32'h3c237693),
	.w2(32'hbbad2ea2),
	.w3(32'h3c402886),
	.w4(32'hbab122db),
	.w5(32'hbc058717),
	.w6(32'hbc13528c),
	.w7(32'hbc96d0eb),
	.w8(32'hbc1abe7a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f5e11),
	.w1(32'hb9b84e60),
	.w2(32'hbc693b25),
	.w3(32'hbccb1df6),
	.w4(32'hbbb6404a),
	.w5(32'hbc90cb38),
	.w6(32'hbc85e9f6),
	.w7(32'hb9ec2d35),
	.w8(32'hbc287a1f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce61c68),
	.w1(32'hbc0b5988),
	.w2(32'hbb60f3cf),
	.w3(32'hbd557efe),
	.w4(32'hbce8be9f),
	.w5(32'hbb341ab4),
	.w6(32'hbd0177b6),
	.w7(32'hbc87031f),
	.w8(32'h3b9a9ce4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd69fa),
	.w1(32'hbc22798e),
	.w2(32'hbb822820),
	.w3(32'h3b828a46),
	.w4(32'h3c18961c),
	.w5(32'hbbf3fab9),
	.w6(32'h3bc47725),
	.w7(32'hba1c2a1d),
	.w8(32'hbbe95ead),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904e9f),
	.w1(32'hbcde74b1),
	.w2(32'hbba5e5a0),
	.w3(32'hbcba5e24),
	.w4(32'hbcc568e0),
	.w5(32'h3b81c73f),
	.w6(32'hbcc1aa3a),
	.w7(32'hbbfa70df),
	.w8(32'hba158684),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be991b0),
	.w1(32'h3c58394b),
	.w2(32'h3b36894c),
	.w3(32'hbacc8145),
	.w4(32'h3b7ee0d9),
	.w5(32'hba3f1d2b),
	.w6(32'hbbb2672a),
	.w7(32'hbc08210c),
	.w8(32'hbb2ec94b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb7f1b),
	.w1(32'h3bcebac2),
	.w2(32'h3c3e0c72),
	.w3(32'h3c6a55b9),
	.w4(32'h3c261ff8),
	.w5(32'hbaa7f2ff),
	.w6(32'hba04ec51),
	.w7(32'hbb794e47),
	.w8(32'hbbe4851c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a3302),
	.w1(32'hbc575e6e),
	.w2(32'hbb1ad941),
	.w3(32'hbc0fd471),
	.w4(32'hbb94341a),
	.w5(32'h39267147),
	.w6(32'hbc052262),
	.w7(32'hbc1f65af),
	.w8(32'hbbdfb915),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042648),
	.w1(32'hbc1d9b88),
	.w2(32'hba397c18),
	.w3(32'hbc0819bf),
	.w4(32'hbb89ee07),
	.w5(32'hbb0858a9),
	.w6(32'hbbbab051),
	.w7(32'hbbed038a),
	.w8(32'h3bea44ee),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d3f7b),
	.w1(32'hbcb6d19b),
	.w2(32'hbca73a6a),
	.w3(32'hb9f3f3c8),
	.w4(32'hbc7b369f),
	.w5(32'hbbc1bc4c),
	.w6(32'hbbbfb932),
	.w7(32'hbc2cec07),
	.w8(32'hbbcd5efa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870e39),
	.w1(32'h3a018b05),
	.w2(32'hbc17f5db),
	.w3(32'hbb38a27c),
	.w4(32'h3b6c22ff),
	.w5(32'hbc49bc52),
	.w6(32'hbba8d378),
	.w7(32'hbb42d8e6),
	.w8(32'hbbae89b7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bddb0),
	.w1(32'h3af847c7),
	.w2(32'hba192826),
	.w3(32'h3c0bdfcc),
	.w4(32'h3bd54436),
	.w5(32'hbab8f000),
	.w6(32'h3b49262a),
	.w7(32'h3a128e62),
	.w8(32'h3b4e75a8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb726502f),
	.w1(32'h3c026237),
	.w2(32'hbb90a50b),
	.w3(32'h3bf20676),
	.w4(32'h3c86a7e7),
	.w5(32'hbc958fb6),
	.w6(32'h3bbc1d57),
	.w7(32'h3c021d60),
	.w8(32'hbc2d26bd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcc4d6),
	.w1(32'h3b8cfede),
	.w2(32'h3bad627a),
	.w3(32'hbcea2014),
	.w4(32'h3c0e596b),
	.w5(32'h3bba8316),
	.w6(32'hbc547cf4),
	.w7(32'hb97b79b4),
	.w8(32'h3b87d308),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f58f3),
	.w1(32'h3c60213f),
	.w2(32'hbc99c54b),
	.w3(32'h3c805ee2),
	.w4(32'h3c480141),
	.w5(32'hbd1487b6),
	.w6(32'h3c10eec2),
	.w7(32'h3bd680ad),
	.w8(32'hbc960e90),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd021629),
	.w1(32'hbc1e8977),
	.w2(32'hbb217ea0),
	.w3(32'hbd6eb7ed),
	.w4(32'hbca7c119),
	.w5(32'h3c475dd1),
	.w6(32'hbcec3f6a),
	.w7(32'hbc918642),
	.w8(32'h3c3c568c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d5965),
	.w1(32'h3c8c451a),
	.w2(32'hbbf7040e),
	.w3(32'h3d131498),
	.w4(32'h3cd95ae9),
	.w5(32'hbc0fb7b7),
	.w6(32'h3cd6d4bb),
	.w7(32'h3c33af1e),
	.w8(32'hbb30e2b0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21ea21),
	.w1(32'hbb1880ca),
	.w2(32'h3c513003),
	.w3(32'h3982fe8c),
	.w4(32'h3bf2b70a),
	.w5(32'h3c7d0edb),
	.w6(32'hbb078d14),
	.w7(32'h3af18cc8),
	.w8(32'h3c3b22de),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd2f8c),
	.w1(32'h3cb5156d),
	.w2(32'h3ba3c5f3),
	.w3(32'h3cc90b60),
	.w4(32'h3cc319bf),
	.w5(32'h3bd80292),
	.w6(32'h3c43edd9),
	.w7(32'h3c559adc),
	.w8(32'h3bbd9c0b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287a5b),
	.w1(32'h3b9d3093),
	.w2(32'hbb3edb5e),
	.w3(32'h3ae6fe95),
	.w4(32'hbb84e788),
	.w5(32'hbb50c819),
	.w6(32'hbbcdc7b0),
	.w7(32'h3b681d53),
	.w8(32'hbbfbb6ec),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956fd5a),
	.w1(32'hbb482a77),
	.w2(32'hbc1b2b7e),
	.w3(32'h3ad0f252),
	.w4(32'hba8cddcb),
	.w5(32'hbc3fef16),
	.w6(32'hbaa31785),
	.w7(32'hbb614b53),
	.w8(32'hbbc82bc3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0235a),
	.w1(32'h3b116ad7),
	.w2(32'h3a3a7d34),
	.w3(32'h3ad3f8e8),
	.w4(32'h3bc253b7),
	.w5(32'h3aa5d21f),
	.w6(32'h3a5f25ab),
	.w7(32'h3c559300),
	.w8(32'hbaba3191),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab23da5),
	.w1(32'hbad16432),
	.w2(32'hbabb6e50),
	.w3(32'hbb2c2cff),
	.w4(32'hbb2f61bf),
	.w5(32'hbadd0269),
	.w6(32'h3a97c386),
	.w7(32'hbb037a97),
	.w8(32'h3baf7d3b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eb43b),
	.w1(32'hbb898d71),
	.w2(32'h3bce1b71),
	.w3(32'h3b9458f3),
	.w4(32'h3bfafa41),
	.w5(32'hba663095),
	.w6(32'h3c314fe8),
	.w7(32'hbb4ab74e),
	.w8(32'hbb780b59),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440e26),
	.w1(32'h3c2eb280),
	.w2(32'hbccc92ad),
	.w3(32'hbbd4e000),
	.w4(32'hbbad977e),
	.w5(32'hbd4c8d89),
	.w6(32'hbb7a3ca6),
	.w7(32'hbc2de2db),
	.w8(32'hbd2e00cc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36e475),
	.w1(32'hbd0fe6c4),
	.w2(32'h39e89c0b),
	.w3(32'hbda87e08),
	.w4(32'hbd91dcce),
	.w5(32'h38cb825b),
	.w6(32'hbd8395e5),
	.w7(32'hbd5f2e4f),
	.w8(32'h3a85ae71),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe382b1),
	.w1(32'hbc27e2fb),
	.w2(32'hb88e491c),
	.w3(32'hbb773085),
	.w4(32'hbbc2a268),
	.w5(32'h3a86c2f4),
	.w6(32'hbade3d76),
	.w7(32'h3b1224bc),
	.w8(32'h3ae32b61),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ec4d),
	.w1(32'h3bd06da5),
	.w2(32'h3bf977f9),
	.w3(32'h3b5219ab),
	.w4(32'h3a439634),
	.w5(32'h3b8861d7),
	.w6(32'h3a948dd1),
	.w7(32'hbac57f86),
	.w8(32'h3b643f12),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f52c),
	.w1(32'hbab2f647),
	.w2(32'h3b2ee47c),
	.w3(32'h3aeb86d5),
	.w4(32'hbbb0db93),
	.w5(32'hbb296686),
	.w6(32'h3b586c5b),
	.w7(32'hbbb468f0),
	.w8(32'hbbd3e2dc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a913ec),
	.w1(32'hbb413a4b),
	.w2(32'h3acc6aed),
	.w3(32'hbbc63757),
	.w4(32'hbc03ccd1),
	.w5(32'h3c7e64fe),
	.w6(32'hbbc504cb),
	.w7(32'hbc28d79f),
	.w8(32'h3c8b57ac),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c506893),
	.w1(32'h3be5bde1),
	.w2(32'h3b817597),
	.w3(32'h3ca9e5c5),
	.w4(32'h3c19a521),
	.w5(32'h3c9005ff),
	.w6(32'h3c2bdbb4),
	.w7(32'h3a0f0f38),
	.w8(32'h3c30ef9d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c855e07),
	.w1(32'h3c5b329e),
	.w2(32'hbab39f72),
	.w3(32'h3cf3b4db),
	.w4(32'h3c1c4b19),
	.w5(32'hbbb2af9c),
	.w6(32'h3c4d6f66),
	.w7(32'h3b6517dd),
	.w8(32'hbbe0771b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61b809),
	.w1(32'hbac93839),
	.w2(32'hb89957c2),
	.w3(32'h3b1e1548),
	.w4(32'h3afb7333),
	.w5(32'h3ac147e8),
	.w6(32'hbbfefd25),
	.w7(32'hbc1bf459),
	.w8(32'hbae4c9cb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38445d),
	.w1(32'h3c67714b),
	.w2(32'h3c3a1c7e),
	.w3(32'h3bab673a),
	.w4(32'h3c67d09f),
	.w5(32'h3c07d045),
	.w6(32'h3a245317),
	.w7(32'h3c1d5a19),
	.w8(32'h3c8b3657),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a13cc),
	.w1(32'h3ce02f08),
	.w2(32'hbc496b1a),
	.w3(32'h3c52030f),
	.w4(32'h3c787a3f),
	.w5(32'h3b8b3a64),
	.w6(32'h3c905b18),
	.w7(32'h3c7a22b3),
	.w8(32'h3c021e53),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd805),
	.w1(32'hb941e226),
	.w2(32'hbb8edf0c),
	.w3(32'h3c8eb661),
	.w4(32'h3bfccc2d),
	.w5(32'hbcdd1efb),
	.w6(32'h3bcc3579),
	.w7(32'h3ba6e284),
	.w8(32'hbc8cce74),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87d351),
	.w1(32'hbb893225),
	.w2(32'h3c78d267),
	.w3(32'hbd2ed5ad),
	.w4(32'hbcea5c5b),
	.w5(32'h3bf4e4a7),
	.w6(32'hbd2d1e50),
	.w7(32'hbce524fe),
	.w8(32'h3ab15e9a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f3353),
	.w1(32'h3b988e6d),
	.w2(32'h3c23b8be),
	.w3(32'h3c3de644),
	.w4(32'h3bbaa5b0),
	.w5(32'h3c3c6ced),
	.w6(32'h3bf29f2a),
	.w7(32'hba8a571a),
	.w8(32'h3c415484),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59a74b),
	.w1(32'h3c4fce62),
	.w2(32'h3c5f8672),
	.w3(32'h3ca2994d),
	.w4(32'h3c62e98d),
	.w5(32'h3c1c33ad),
	.w6(32'h3c8c4184),
	.w7(32'h3bc59ce2),
	.w8(32'h3c0b111e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8193b7),
	.w1(32'hbc9ac889),
	.w2(32'hbb618f55),
	.w3(32'hbc6d9e36),
	.w4(32'hbc8ef5b8),
	.w5(32'h3b6fed46),
	.w6(32'hbc18130d),
	.w7(32'hbc67872f),
	.w8(32'h3b0a9358),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38647897),
	.w1(32'hbb843f28),
	.w2(32'hbb6ed17c),
	.w3(32'hbaa8e3d3),
	.w4(32'hbbe001f4),
	.w5(32'h3bd86d07),
	.w6(32'h3bc55aa2),
	.w7(32'hbc82a47c),
	.w8(32'h3c279b01),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0603b),
	.w1(32'h3c1fb96a),
	.w2(32'hbbca6d09),
	.w3(32'h3c5790f7),
	.w4(32'h3b86c292),
	.w5(32'hbcb766ad),
	.w6(32'h3bf2a52c),
	.w7(32'h3b073b5b),
	.w8(32'hbcf4635a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd176ab4),
	.w1(32'hbd15a783),
	.w2(32'hbbbdba28),
	.w3(32'hbd839555),
	.w4(32'hbd5d0f22),
	.w5(32'hbb363ff4),
	.w6(32'hbd5f6661),
	.w7(32'hbd12fc5e),
	.w8(32'hbba196ff),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3a18),
	.w1(32'hbb8abb23),
	.w2(32'h3bab0893),
	.w3(32'hbc1e2d65),
	.w4(32'hbc06d1ff),
	.w5(32'hbc68ebcb),
	.w6(32'hbc52f88a),
	.w7(32'hbbf8052e),
	.w8(32'hbc8a510c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acab2de),
	.w1(32'h3a21419f),
	.w2(32'h3c2334aa),
	.w3(32'hbcd86b8e),
	.w4(32'hbc56f58a),
	.w5(32'h3bd59e3a),
	.w6(32'hbd2a1f24),
	.w7(32'hbcd048e4),
	.w8(32'h3b88982e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd57834),
	.w1(32'h3ba881e5),
	.w2(32'h3b8b2c87),
	.w3(32'h3c12a75e),
	.w4(32'h3bb39fdb),
	.w5(32'h3bfdc422),
	.w6(32'h3c118a86),
	.w7(32'h3c5d0895),
	.w8(32'h3b7a649e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5c0f5),
	.w1(32'h3c32c53e),
	.w2(32'hbb243a75),
	.w3(32'h3b73bc62),
	.w4(32'h3c18a3ef),
	.w5(32'hba5e835e),
	.w6(32'h3ba64b08),
	.w7(32'h3bb2338e),
	.w8(32'hbb49fef4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7194e9),
	.w1(32'hbb276a50),
	.w2(32'hbbd88990),
	.w3(32'h3c3351c4),
	.w4(32'h3c00e02e),
	.w5(32'hbaa1c7b1),
	.w6(32'h39ac1798),
	.w7(32'h3b79c486),
	.w8(32'hbac1d058),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa6af3),
	.w1(32'hbb6e4178),
	.w2(32'hbb5dba32),
	.w3(32'hbb49d75c),
	.w4(32'hbb6763cb),
	.w5(32'hb8dc2f4c),
	.w6(32'h3b150990),
	.w7(32'hbad95749),
	.w8(32'h3b466d7e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7856f4),
	.w1(32'hbab945e8),
	.w2(32'hbbbe29a4),
	.w3(32'h3b013605),
	.w4(32'hb8ea07de),
	.w5(32'hbaef0751),
	.w6(32'h3b7f33ac),
	.w7(32'h3a06e1c3),
	.w8(32'h3a368965),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19cd5d),
	.w1(32'hbbd4f00e),
	.w2(32'hba1d46cf),
	.w3(32'h3bf3eb46),
	.w4(32'h3b82bd66),
	.w5(32'hbc0cad09),
	.w6(32'h3ba1f142),
	.w7(32'h3b691d3c),
	.w8(32'hbb25775c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00187a),
	.w1(32'h3b84f71a),
	.w2(32'hbc16918f),
	.w3(32'hbbd7fa1d),
	.w4(32'hbb753eff),
	.w5(32'hb9fc05f1),
	.w6(32'hbbe2bacf),
	.w7(32'hbb42bc7c),
	.w8(32'h3c498514),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04912b),
	.w1(32'h3c1408ab),
	.w2(32'h399105af),
	.w3(32'h3ab7c975),
	.w4(32'h3b09c1b1),
	.w5(32'hba7b1b0e),
	.w6(32'h3c5e0b19),
	.w7(32'h3a85b82d),
	.w8(32'hbb9745f0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b6295),
	.w1(32'hbbb819b3),
	.w2(32'hbc6a9948),
	.w3(32'hbadc11a6),
	.w4(32'hbbc9a68f),
	.w5(32'hbcf5e7de),
	.w6(32'hbbef2f0b),
	.w7(32'hbc764ac6),
	.w8(32'hbca1f4e6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14296a),
	.w1(32'hbc7891ba),
	.w2(32'h3a3277f9),
	.w3(32'hbd80aecc),
	.w4(32'hbd188792),
	.w5(32'h3b01ef36),
	.w6(32'hbd2f0ab1),
	.w7(32'hbd02c5f4),
	.w8(32'h3c259fed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c352d3c),
	.w1(32'h3ca2955e),
	.w2(32'h3bf5935c),
	.w3(32'h3c988ca6),
	.w4(32'h3cc86624),
	.w5(32'hbb21b120),
	.w6(32'h3c74bee6),
	.w7(32'h3c659624),
	.w8(32'hbb47250f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d922f),
	.w1(32'hbc3fa0a9),
	.w2(32'hbaa7d26e),
	.w3(32'hbc408d27),
	.w4(32'hbc438b78),
	.w5(32'h3a993724),
	.w6(32'hbbc84d59),
	.w7(32'hbb9288a7),
	.w8(32'h3b21c604),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91cdd5),
	.w1(32'h3b96a137),
	.w2(32'h3b9f3825),
	.w3(32'hbafeadbf),
	.w4(32'h3b38551a),
	.w5(32'h3b9b6ff2),
	.w6(32'h3bc0f427),
	.w7(32'h39eb1615),
	.w8(32'hba5494a1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aca54),
	.w1(32'h3c562d6a),
	.w2(32'hb8b80287),
	.w3(32'hbb96f40c),
	.w4(32'hbbd3837e),
	.w5(32'hbb138aba),
	.w6(32'h3bbfce79),
	.w7(32'hbba8ff55),
	.w8(32'h3addab18),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b490a),
	.w1(32'h3a2d1c4b),
	.w2(32'hba20042a),
	.w3(32'h3c07f91e),
	.w4(32'h3c7f3808),
	.w5(32'h39b0bdd0),
	.w6(32'h3c453257),
	.w7(32'h3abcbd79),
	.w8(32'hba55fd28),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6f7ab),
	.w1(32'h3aad192c),
	.w2(32'h3bdbdb3a),
	.w3(32'h3a0eb564),
	.w4(32'h3b1b166d),
	.w5(32'h3b6618aa),
	.w6(32'hbb228458),
	.w7(32'h38fa6ecc),
	.w8(32'h3b4dc503),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcc81),
	.w1(32'h3bda077f),
	.w2(32'h3af9097a),
	.w3(32'h3c1f1e17),
	.w4(32'h3c82d512),
	.w5(32'hbc4c85f1),
	.w6(32'hb99cd678),
	.w7(32'h3c0f5be5),
	.w8(32'hbbafd514),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5618f2),
	.w1(32'hbc143bd7),
	.w2(32'hbb01fbf3),
	.w3(32'hbc6e69eb),
	.w4(32'h3a69ecdf),
	.w5(32'h3afcac8d),
	.w6(32'hbc2dff0d),
	.w7(32'hbc83cf94),
	.w8(32'h3b2aa061),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32197),
	.w1(32'hbc198502),
	.w2(32'h3b416c77),
	.w3(32'hbb8e35a8),
	.w4(32'hbc06ccf4),
	.w5(32'hb91a79f8),
	.w6(32'h3b08344d),
	.w7(32'h3abcdccf),
	.w8(32'hbbe86a0f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fa2c2),
	.w1(32'h3aa1f856),
	.w2(32'h3c90a672),
	.w3(32'h3c6936aa),
	.w4(32'h3ce6d457),
	.w5(32'h3d02d2e9),
	.w6(32'hbc483641),
	.w7(32'h3c127f86),
	.w8(32'hbc3b5648),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6273a2),
	.w1(32'hbc9e05ea),
	.w2(32'h3ac6a0b5),
	.w3(32'h3d83b4fd),
	.w4(32'h3d1f1059),
	.w5(32'hba4b354d),
	.w6(32'h3c42bcf8),
	.w7(32'h3d1b033b),
	.w8(32'hbb81e93d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f06c2),
	.w1(32'hbb8f9399),
	.w2(32'h3c28e0a2),
	.w3(32'h3b992cdb),
	.w4(32'h3a988ea5),
	.w5(32'hba453bf3),
	.w6(32'h3a2e4055),
	.w7(32'h3b38785f),
	.w8(32'h3bda3b8f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21946e),
	.w1(32'h3bac5418),
	.w2(32'h3b4770ff),
	.w3(32'hb8c0a781),
	.w4(32'hba6e1de5),
	.w5(32'h39d4f2c8),
	.w6(32'h3bdebbfe),
	.w7(32'h3b72d475),
	.w8(32'hbafa6e67),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16677d),
	.w1(32'hbb63d3a4),
	.w2(32'h3b64d28d),
	.w3(32'h3b8063da),
	.w4(32'h3b2ae948),
	.w5(32'hbb1a9311),
	.w6(32'hba60d199),
	.w7(32'h3b164c1e),
	.w8(32'h3a0e2a7a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af130b),
	.w1(32'hbc819eae),
	.w2(32'hbb66b156),
	.w3(32'h39b0600b),
	.w4(32'h3ba8bebf),
	.w5(32'hba9bb474),
	.w6(32'hbbcff921),
	.w7(32'hbbaf9d75),
	.w8(32'hbc177aa2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1418ac),
	.w1(32'hbc5fa291),
	.w2(32'hbc88a425),
	.w3(32'h3b5ae8cd),
	.w4(32'hbb8c9ddb),
	.w5(32'h3c3c0048),
	.w6(32'hbbbd8763),
	.w7(32'hb9a31e34),
	.w8(32'h3b38bf49),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb00fa7),
	.w1(32'hbbf06faa),
	.w2(32'hbc44e7d7),
	.w3(32'hbc51abf8),
	.w4(32'hbcf8977b),
	.w5(32'h3b05eb8b),
	.w6(32'h3c1ec586),
	.w7(32'hbb9ae7c0),
	.w8(32'hbbb8dd86),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fbcd3),
	.w1(32'h3c33223b),
	.w2(32'h3b8df75d),
	.w3(32'hbb939941),
	.w4(32'hbbefb742),
	.w5(32'h39f1fae6),
	.w6(32'hbbe78390),
	.w7(32'hbba54104),
	.w8(32'h3b0494e2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b3b8),
	.w1(32'hbb8aa64a),
	.w2(32'h39da865c),
	.w3(32'hbc16db80),
	.w4(32'hbc02e7cd),
	.w5(32'h3c9406dd),
	.w6(32'hbc48591e),
	.w7(32'hbbda31f2),
	.w8(32'h3c8c1009),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4311ba),
	.w1(32'hbb63b5ec),
	.w2(32'h3bcbae0d),
	.w3(32'h3c88e2d9),
	.w4(32'hbbfab8e0),
	.w5(32'hbc4bb832),
	.w6(32'h3cecd61f),
	.w7(32'h3cb3b302),
	.w8(32'h3b845530),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c41a2),
	.w1(32'h3c3726ce),
	.w2(32'h3aecc01e),
	.w3(32'h39b85749),
	.w4(32'h3cbefca3),
	.w5(32'hbb7e20a1),
	.w6(32'hbbce1a45),
	.w7(32'hbc4264dd),
	.w8(32'hbb894a68),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3d4d3),
	.w1(32'hb77cb771),
	.w2(32'h3b651ca9),
	.w3(32'hbaaf1d42),
	.w4(32'h3af13aa8),
	.w5(32'h3a8a02ce),
	.w6(32'hbc07e5cc),
	.w7(32'hb952f30e),
	.w8(32'h3c4401f3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cb1de),
	.w1(32'hbbb8afc8),
	.w2(32'hbb86e8aa),
	.w3(32'hbc80075e),
	.w4(32'hbc7323fe),
	.w5(32'h3b5f23ff),
	.w6(32'hbb946c8e),
	.w7(32'hbca55cf9),
	.w8(32'hbc47e3ee),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a40f8),
	.w1(32'hbb8b10e3),
	.w2(32'h3bb884f9),
	.w3(32'h3bacee39),
	.w4(32'hbc09c9bf),
	.w5(32'h3b7dc1be),
	.w6(32'hb91d5b8a),
	.w7(32'h3bd087c3),
	.w8(32'hbb74e7fa),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ceaea1),
	.w1(32'h3baa7687),
	.w2(32'hbc34d738),
	.w3(32'hbb329523),
	.w4(32'h3974ef3b),
	.w5(32'h3c8adb89),
	.w6(32'hbb9da85a),
	.w7(32'hbb8a4c52),
	.w8(32'h3c587be4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0051e8),
	.w1(32'h3bac3c5f),
	.w2(32'h3999379e),
	.w3(32'hbc730ec8),
	.w4(32'hbcae9f2b),
	.w5(32'hbb137e77),
	.w6(32'h3c60ea00),
	.w7(32'hbbdd8fea),
	.w8(32'hbb889d27),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1836a),
	.w1(32'hbb921a1f),
	.w2(32'hbb1cae45),
	.w3(32'hbb9b8cbd),
	.w4(32'hb9b708ae),
	.w5(32'hbc3e4d0f),
	.w6(32'hbc1ad845),
	.w7(32'hbbccca71),
	.w8(32'hbc4a5589),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f5569),
	.w1(32'h39dc5076),
	.w2(32'hbb23a74f),
	.w3(32'hbc72dfba),
	.w4(32'h3b80a351),
	.w5(32'h3b231629),
	.w6(32'hbca92105),
	.w7(32'hbc5fb5b3),
	.w8(32'hbad71795),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb866bcf3),
	.w1(32'hbaa0904e),
	.w2(32'h3b809c07),
	.w3(32'hbbb86eab),
	.w4(32'h3aa6af2a),
	.w5(32'hbbd383de),
	.w6(32'hba99c11f),
	.w7(32'h3b8feedf),
	.w8(32'hba574886),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257382),
	.w1(32'hba1e2cc0),
	.w2(32'h3b8d9b10),
	.w3(32'hbb910e5f),
	.w4(32'hbb1b54b7),
	.w5(32'h3ba01344),
	.w6(32'hba681a62),
	.w7(32'hbbe44361),
	.w8(32'h3c229086),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8621913),
	.w1(32'h3b02616f),
	.w2(32'hbb874143),
	.w3(32'h3c0dcbef),
	.w4(32'h3b948b58),
	.w5(32'hbc5059c9),
	.w6(32'h3c217b86),
	.w7(32'hbaa0c192),
	.w8(32'hbbd5570f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c3937),
	.w1(32'h3bc632bc),
	.w2(32'hbc3917fb),
	.w3(32'hbbad649f),
	.w4(32'h3c2ea7fd),
	.w5(32'hbb23dc44),
	.w6(32'hbc69212f),
	.w7(32'hbbd81e57),
	.w8(32'h3b5632e6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0854c9),
	.w1(32'h3b3e3953),
	.w2(32'h3b2f3305),
	.w3(32'hbcb28ae6),
	.w4(32'h3b8e087f),
	.w5(32'hbc7c66fa),
	.w6(32'h3b1f1879),
	.w7(32'hbc3ccd85),
	.w8(32'hbc0ef726),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56341a),
	.w1(32'h3b7e32c8),
	.w2(32'h3ce8eb58),
	.w3(32'h3b4a19bf),
	.w4(32'h3c582e82),
	.w5(32'h3c0dfbe3),
	.w6(32'hbc9abdb3),
	.w7(32'hbb11b6ad),
	.w8(32'hbc5b38c7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff4d4d),
	.w1(32'hbca51bfa),
	.w2(32'hbb6d7a9f),
	.w3(32'h3d434d12),
	.w4(32'h3cbe2f2a),
	.w5(32'hbbb824eb),
	.w6(32'hbb1adc3f),
	.w7(32'h3c832f6b),
	.w8(32'hbb11862c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922be3),
	.w1(32'hbb7119bd),
	.w2(32'hba5ee98d),
	.w3(32'hbc2a7614),
	.w4(32'hbba32f47),
	.w5(32'hba4c4442),
	.w6(32'hbb3d613f),
	.w7(32'hbb8b5a82),
	.w8(32'hba25ad69),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3957),
	.w1(32'hbbaeb3bf),
	.w2(32'h3b1b6060),
	.w3(32'hbb98b7fc),
	.w4(32'h3ba3da06),
	.w5(32'h3aa17ac0),
	.w6(32'hbb169fd8),
	.w7(32'h3c016195),
	.w8(32'h3b7f71ec),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91a9da),
	.w1(32'hbc43536a),
	.w2(32'hbce17e17),
	.w3(32'hbc8bd703),
	.w4(32'hbca8fdc3),
	.w5(32'hbad2248e),
	.w6(32'h39e3f29b),
	.w7(32'h3afa22a6),
	.w8(32'h3c2bf4df),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc741ea0),
	.w1(32'h3b7a1a3a),
	.w2(32'hbc7bc80c),
	.w3(32'hbc877436),
	.w4(32'hbc6a584d),
	.w5(32'hbcc5bb65),
	.w6(32'h3cd1f44a),
	.w7(32'h3b2182a6),
	.w8(32'hbc6ce458),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89108a),
	.w1(32'h3b0f8ed8),
	.w2(32'hbbe73aab),
	.w3(32'hbceef0d7),
	.w4(32'hbc37f13e),
	.w5(32'hbaa0afe2),
	.w6(32'hbcf5a902),
	.w7(32'hbca8c53f),
	.w8(32'h3bf0047d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe10583),
	.w1(32'hbc376d71),
	.w2(32'hbb891ecf),
	.w3(32'hbc009990),
	.w4(32'hbb6d7f1d),
	.w5(32'hbb992063),
	.w6(32'hbb3cb220),
	.w7(32'hbbc6e5a1),
	.w8(32'hbabf8c1f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5887e),
	.w1(32'hb99d9c2f),
	.w2(32'h3b8aa167),
	.w3(32'hbbc3b28a),
	.w4(32'hbc1cee7c),
	.w5(32'h3c8c2099),
	.w6(32'h3aad6975),
	.w7(32'h3a62f3b9),
	.w8(32'hbac255d2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5af818),
	.w1(32'h3c134cc0),
	.w2(32'h3abc9bb3),
	.w3(32'h3c3fe05b),
	.w4(32'h3c7cbd66),
	.w5(32'hb9f0e9de),
	.w6(32'h3991bc65),
	.w7(32'h3c7ae96c),
	.w8(32'hbae8fc41),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41f528),
	.w1(32'h39274818),
	.w2(32'hba470c5d),
	.w3(32'hbb8876f9),
	.w4(32'h3813e988),
	.w5(32'h3b691b0b),
	.w6(32'hbba15f6b),
	.w7(32'hba7f43b9),
	.w8(32'hba0e3bf3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904bfa),
	.w1(32'hbb141e58),
	.w2(32'hbab1e264),
	.w3(32'h3ae68845),
	.w4(32'h3adfcb26),
	.w5(32'h3b25aeff),
	.w6(32'hbba2d52c),
	.w7(32'h3b9a6d1a),
	.w8(32'hbb48187a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5787a4),
	.w1(32'h3bdbaaf9),
	.w2(32'hbb0eec27),
	.w3(32'h3c267610),
	.w4(32'hb9d7bfb9),
	.w5(32'hbb0dac60),
	.w6(32'h3bed36cf),
	.w7(32'h3bf6a2d1),
	.w8(32'hbb501318),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb522a8c),
	.w1(32'hbc0485c7),
	.w2(32'hbb2d49a1),
	.w3(32'hb8d1f284),
	.w4(32'h3bdc76d2),
	.w5(32'hbbef8ada),
	.w6(32'hbb2f54f8),
	.w7(32'hb8f57a32),
	.w8(32'hbb75a970),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14b4f1),
	.w1(32'hbb8adeb7),
	.w2(32'h3c102ecd),
	.w3(32'hbc202430),
	.w4(32'hbc1d0075),
	.w5(32'h3c4754cf),
	.w6(32'hbbf1d96a),
	.w7(32'hbbda7284),
	.w8(32'hba8daaec),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160e4b),
	.w1(32'h3be86c2c),
	.w2(32'h3b9370a4),
	.w3(32'hbac563ef),
	.w4(32'hbb864ee5),
	.w5(32'hbc964a92),
	.w6(32'h3bde9616),
	.w7(32'h3ba14f61),
	.w8(32'hbbf22819),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31bff1),
	.w1(32'h3c31b91a),
	.w2(32'h3bd66e09),
	.w3(32'hbc2e6658),
	.w4(32'h3bbce88f),
	.w5(32'h3c36a895),
	.w6(32'hbc87aa01),
	.w7(32'hbc25c62b),
	.w8(32'h3b907bb3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa659af),
	.w1(32'hbc15860b),
	.w2(32'hbbd02945),
	.w3(32'h3a161aa2),
	.w4(32'hbba47bb7),
	.w5(32'hbc59bd4a),
	.w6(32'h3ad1322e),
	.w7(32'hba962abf),
	.w8(32'hbc44ab05),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2da8bc),
	.w1(32'hba99b9e2),
	.w2(32'h383be44c),
	.w3(32'hbb3265fa),
	.w4(32'hbbafe4ff),
	.w5(32'h3ac6a358),
	.w6(32'hbc56167c),
	.w7(32'hbaad1a35),
	.w8(32'hbb31e21c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ddeb8),
	.w1(32'hba86c87d),
	.w2(32'h3ba6c43f),
	.w3(32'hba380e32),
	.w4(32'h3b602dec),
	.w5(32'h3b8c08e6),
	.w6(32'hbb87c697),
	.w7(32'h3a748f4e),
	.w8(32'h3b5caa27),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab694ea),
	.w1(32'hbaf942ac),
	.w2(32'h3bddc013),
	.w3(32'h3befacda),
	.w4(32'h3bdbbabe),
	.w5(32'h3c0ba51b),
	.w6(32'hbbe29539),
	.w7(32'h3b53c85f),
	.w8(32'h3b75120b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d7654),
	.w1(32'h3c41f927),
	.w2(32'h3c230baf),
	.w3(32'h3c9dbf1f),
	.w4(32'h3c804c9f),
	.w5(32'h3b08a1a9),
	.w6(32'h3c5f8e6b),
	.w7(32'h3bb3a16d),
	.w8(32'h3b089017),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5efc0f),
	.w1(32'h3c45fc33),
	.w2(32'h3b8268d6),
	.w3(32'h3babf013),
	.w4(32'h3c24deb9),
	.w5(32'h39a48731),
	.w6(32'h3ab542c3),
	.w7(32'h3c0a2370),
	.w8(32'h3c8af080),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0d31c),
	.w1(32'h3d11f581),
	.w2(32'hbadea6e4),
	.w3(32'h3ceac027),
	.w4(32'h3d2705e5),
	.w5(32'hbc197919),
	.w6(32'h3c82105f),
	.w7(32'h3c86b09f),
	.w8(32'hbaa957ae),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1816f),
	.w1(32'h3ad22141),
	.w2(32'hbb004662),
	.w3(32'hbc3ce1d6),
	.w4(32'hbb33d2b4),
	.w5(32'h3c38b06a),
	.w6(32'hbb7e5555),
	.w7(32'h399913c6),
	.w8(32'h3bcea628),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0d9c),
	.w1(32'hb8c7df3c),
	.w2(32'hbb84302e),
	.w3(32'hb7337a38),
	.w4(32'hbb69c000),
	.w5(32'hbb657453),
	.w6(32'h3b56a1cc),
	.w7(32'hb8f34ec7),
	.w8(32'h3a7726b9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfab939),
	.w1(32'hbbbeba95),
	.w2(32'h3be6bb04),
	.w3(32'hba616341),
	.w4(32'hbb628a62),
	.w5(32'hbbcdc0cd),
	.w6(32'h3bdd1aea),
	.w7(32'h3befa8af),
	.w8(32'hbb617af3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e7e8),
	.w1(32'hbb2814a9),
	.w2(32'hbca5d070),
	.w3(32'hbbb3cb08),
	.w4(32'hbb5ba015),
	.w5(32'hbc2b2260),
	.w6(32'h3a7ef567),
	.w7(32'h39ec6c9c),
	.w8(32'hbb4cea9b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc954f5f),
	.w1(32'h3bb68ec0),
	.w2(32'hbb5f0a45),
	.w3(32'hbd153f47),
	.w4(32'hbcd879f0),
	.w5(32'hbc0a6b70),
	.w6(32'hbccf483d),
	.w7(32'hbcee3888),
	.w8(32'hbb9d6c88),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc390ae8),
	.w1(32'hbcabbb39),
	.w2(32'h3b8afe39),
	.w3(32'hbc89eb87),
	.w4(32'h3a9451aa),
	.w5(32'hbb2750bd),
	.w6(32'hbc9a045e),
	.w7(32'hbc379a27),
	.w8(32'h3b81d06f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2852c6),
	.w1(32'hbc4b1611),
	.w2(32'h3be73350),
	.w3(32'hbc4eb05b),
	.w4(32'hbc8a3472),
	.w5(32'hbb1a3d1c),
	.w6(32'hbb77ae19),
	.w7(32'hbbfc0a5a),
	.w8(32'hbbc73e85),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828205),
	.w1(32'hbb358070),
	.w2(32'hbab71673),
	.w3(32'hbbda97fc),
	.w4(32'hbbf760a5),
	.w5(32'hba124e45),
	.w6(32'hbc074eef),
	.w7(32'hbc0c42a0),
	.w8(32'h39fc8598),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d2e05),
	.w1(32'hbbad194a),
	.w2(32'h3b9c1697),
	.w3(32'hbacea62e),
	.w4(32'hbb955edd),
	.w5(32'h3b8fc26e),
	.w6(32'h3a07a4aa),
	.w7(32'hbb30ac3b),
	.w8(32'h3c10a6aa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff3a30),
	.w1(32'hba8c615e),
	.w2(32'hbb9ed4cf),
	.w3(32'h3b9136ed),
	.w4(32'h3bb7fbb6),
	.w5(32'hbcb7dccb),
	.w6(32'h3c2e9d25),
	.w7(32'h3b6b4f2d),
	.w8(32'h3b051ec6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc669df),
	.w1(32'hb8932151),
	.w2(32'hbc44f556),
	.w3(32'hbcf11e0c),
	.w4(32'hbcc61b13),
	.w5(32'hbc54de8f),
	.w6(32'hbcc89cb5),
	.w7(32'hbcb67f2e),
	.w8(32'hbc03a335),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc68d44),
	.w1(32'hbd0103de),
	.w2(32'h3a0c0b1e),
	.w3(32'hbc5e2e6c),
	.w4(32'hbbbcffa8),
	.w5(32'h3c8ebe23),
	.w6(32'hbcc276ce),
	.w7(32'hbb3daaba),
	.w8(32'h3bdc24b4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873d43),
	.w1(32'hbc3074a2),
	.w2(32'hbc373abc),
	.w3(32'hbbb27ef3),
	.w4(32'hbc5d093c),
	.w5(32'hbb439b9e),
	.w6(32'hbb0f9ae9),
	.w7(32'h3ba1fa8a),
	.w8(32'h3ad273b6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826b09),
	.w1(32'hbb424e93),
	.w2(32'hba9a4403),
	.w3(32'hba1e87cc),
	.w4(32'hba57773a),
	.w5(32'hb886ce9a),
	.w6(32'hbb08737a),
	.w7(32'hbbb1c7f8),
	.w8(32'h3b3c0be2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100846),
	.w1(32'h3ba5f5d2),
	.w2(32'hbad988f4),
	.w3(32'hb94f54ed),
	.w4(32'h3a2fc9d7),
	.w5(32'hbb289bd1),
	.w6(32'h3b9f6fed),
	.w7(32'h3b0be795),
	.w8(32'h3939438d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2db5e),
	.w1(32'h3ac9c614),
	.w2(32'h3b545630),
	.w3(32'h3ace1860),
	.w4(32'hba9ef0ed),
	.w5(32'hbbef8fae),
	.w6(32'hbb1b222e),
	.w7(32'hba21795d),
	.w8(32'hbb00ff56),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2b79),
	.w1(32'hbc69216d),
	.w2(32'hbb2fd246),
	.w3(32'hbc4b1238),
	.w4(32'hbc8176f3),
	.w5(32'h3c02e650),
	.w6(32'hbbac05c0),
	.w7(32'hbbde35d3),
	.w8(32'h3b08f9f5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a190003),
	.w1(32'hbb2f647c),
	.w2(32'h3c2a7162),
	.w3(32'h3c289627),
	.w4(32'h3a522c02),
	.w5(32'h3b3a7031),
	.w6(32'hbc422c3f),
	.w7(32'hba933d56),
	.w8(32'h3c655797),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d1e3b),
	.w1(32'h3af5b7d8),
	.w2(32'h3b3cde0c),
	.w3(32'h3c9b6fbe),
	.w4(32'h3ce632a2),
	.w5(32'hbbbd947a),
	.w6(32'h394425e6),
	.w7(32'h3b9b2236),
	.w8(32'hbafdac0a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4587d1),
	.w1(32'hbbdbebd3),
	.w2(32'hbc13e332),
	.w3(32'hbc30c207),
	.w4(32'hbad188c0),
	.w5(32'h3ba345f7),
	.w6(32'hbc6b4af0),
	.w7(32'h3b2943c6),
	.w8(32'h3b029cb8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e38b1),
	.w1(32'hbc192a59),
	.w2(32'h3b579e94),
	.w3(32'hbbebf93b),
	.w4(32'hbc2f4229),
	.w5(32'hbbeb4788),
	.w6(32'hbae9eff8),
	.w7(32'hbb07fff4),
	.w8(32'h3b2c9e13),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e767c),
	.w1(32'h3aca0944),
	.w2(32'hbbc781b1),
	.w3(32'hbc09d4f9),
	.w4(32'h3aa8ecb4),
	.w5(32'hbbde7881),
	.w6(32'hbb9ee641),
	.w7(32'hbc6942c6),
	.w8(32'hbc0eb59f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2edee),
	.w1(32'h3c062e4a),
	.w2(32'hbbba60a4),
	.w3(32'hbc24a9f3),
	.w4(32'hbadfcb22),
	.w5(32'h3a75fcb5),
	.w6(32'hbb9a77c6),
	.w7(32'hbc150813),
	.w8(32'h3bf9d252),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc675bf3),
	.w1(32'hbc9f8a67),
	.w2(32'hbc6f1251),
	.w3(32'hbcbf397e),
	.w4(32'hbcaa73ca),
	.w5(32'hbc49f0a6),
	.w6(32'hbc0ebee5),
	.w7(32'hbb821678),
	.w8(32'h3b49e2e0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb958949),
	.w1(32'hbbcc2c6d),
	.w2(32'h3c017bc4),
	.w3(32'hbc02a13d),
	.w4(32'hbaf5ff94),
	.w5(32'h3b65da0f),
	.w6(32'hbb628b7b),
	.w7(32'hba5de50d),
	.w8(32'hbb1ca002),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b442c32),
	.w1(32'hbc2bf8b2),
	.w2(32'h3ad3de4e),
	.w3(32'h3c2d470d),
	.w4(32'h3a1249d8),
	.w5(32'hbbf384b9),
	.w6(32'h3c07f809),
	.w7(32'h3c25b34e),
	.w8(32'h3a90cb94),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d15d),
	.w1(32'hbb830d54),
	.w2(32'h3baa7e43),
	.w3(32'hbba8127d),
	.w4(32'hbb84a833),
	.w5(32'h3aecdad0),
	.w6(32'hbc18b5ff),
	.w7(32'hbc2ed2e7),
	.w8(32'h3b364c15),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f4dd8),
	.w1(32'h3b164b3b),
	.w2(32'hbbeddbc1),
	.w3(32'h3afcb5de),
	.w4(32'h3bb1e38e),
	.w5(32'hb97f9ab6),
	.w6(32'hbb488255),
	.w7(32'hbb4d7cf7),
	.w8(32'h3c093c4e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb336dd),
	.w1(32'hbc45c5d2),
	.w2(32'hbbc6a258),
	.w3(32'hbc369ba2),
	.w4(32'hbc513423),
	.w5(32'hbb2361aa),
	.w6(32'h3babec4d),
	.w7(32'hbb5e7c72),
	.w8(32'hbbd7c2aa),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c970),
	.w1(32'hbb6a5699),
	.w2(32'hbb0ae2b4),
	.w3(32'hbbc05976),
	.w4(32'hbc2a5bf2),
	.w5(32'hbc887ab6),
	.w6(32'hbc1648c8),
	.w7(32'hbaf53abe),
	.w8(32'hbb4de7ac),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38dd76),
	.w1(32'h3b1058c7),
	.w2(32'h3baa77e6),
	.w3(32'hbc915986),
	.w4(32'h3bcf2130),
	.w5(32'hbc2f6a4b),
	.w6(32'hbd03faff),
	.w7(32'hbca2aee0),
	.w8(32'h3c33449f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aacc7),
	.w1(32'h3a1f09e8),
	.w2(32'h3b1d4576),
	.w3(32'h3b44ace5),
	.w4(32'h3c84dd7c),
	.w5(32'h372057e6),
	.w6(32'hbb8fb1a6),
	.w7(32'hbb59a217),
	.w8(32'h3b4cd9c3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947a483),
	.w1(32'hbb94e425),
	.w2(32'h3b835354),
	.w3(32'hbaea6cc1),
	.w4(32'hbc026722),
	.w5(32'h3bdefdb7),
	.w6(32'h3a01e7ea),
	.w7(32'h3b21f2f3),
	.w8(32'h3bb6e622),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16bfe),
	.w1(32'h3b788368),
	.w2(32'h3bc8d52d),
	.w3(32'hbbd086f6),
	.w4(32'hbc14d8ad),
	.w5(32'hbc4c133e),
	.w6(32'hbbb810b2),
	.w7(32'hbb55136c),
	.w8(32'hbc52fc4b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41b2e2),
	.w1(32'h3bdc8c46),
	.w2(32'h3c23d9c2),
	.w3(32'hbbd6e467),
	.w4(32'h3c9e4707),
	.w5(32'h3bbac4db),
	.w6(32'hbca37158),
	.w7(32'hbc8e0a3c),
	.w8(32'hbbaf4e94),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8917bc),
	.w1(32'hbb234f2d),
	.w2(32'hbc42bfad),
	.w3(32'hbba32d96),
	.w4(32'hbb018e23),
	.w5(32'hbbb0c2ac),
	.w6(32'h3beb9d54),
	.w7(32'h3bb88fed),
	.w8(32'h3c253fd1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9109fc),
	.w1(32'hbc48124c),
	.w2(32'hbb0135cf),
	.w3(32'hbc85c809),
	.w4(32'hbca73181),
	.w5(32'hbbefb553),
	.w6(32'h3bc141a8),
	.w7(32'hbaf41443),
	.w8(32'h3b2c88f9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9b42),
	.w1(32'hb9afa88d),
	.w2(32'hbc58ab9b),
	.w3(32'hbc523279),
	.w4(32'h3afd41a7),
	.w5(32'h39878d7e),
	.w6(32'hbc6e6c48),
	.w7(32'hbc86b7a5),
	.w8(32'h3c2f2420),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc594dc7),
	.w1(32'hbb901ac9),
	.w2(32'h3bac2310),
	.w3(32'hbc1f3098),
	.w4(32'hbc52f75b),
	.w5(32'hbbca5742),
	.w6(32'h3c44483f),
	.w7(32'h3c0a8c96),
	.w8(32'h3b53bd1e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1949c5),
	.w1(32'hbb76fdae),
	.w2(32'hbaa095be),
	.w3(32'hbc186b81),
	.w4(32'h3b29530c),
	.w5(32'hbc06d0d4),
	.w6(32'hbc418b8e),
	.w7(32'hbbc0378a),
	.w8(32'hbb3d91de),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dfba3),
	.w1(32'hbb3b12e0),
	.w2(32'hbb8549b3),
	.w3(32'hbba65a9e),
	.w4(32'h3c536615),
	.w5(32'hbb836a53),
	.w6(32'hbb91526e),
	.w7(32'hbb0159df),
	.w8(32'h3c152130),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43b380),
	.w1(32'hbb86154f),
	.w2(32'hbba94772),
	.w3(32'hbbda49dd),
	.w4(32'hbafa42e1),
	.w5(32'h3a5faf76),
	.w6(32'hbbbfd7cf),
	.w7(32'hbbe64461),
	.w8(32'hbb2088af),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dbd7a),
	.w1(32'hbbaa4c0b),
	.w2(32'hb90c0674),
	.w3(32'h3b2c67a5),
	.w4(32'hba74f784),
	.w5(32'hba4de44c),
	.w6(32'h3b21da40),
	.w7(32'h3b4163c1),
	.w8(32'h3ac5e88a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ccc3a),
	.w1(32'h3999b446),
	.w2(32'h3c3221e7),
	.w3(32'hb9e0b5a5),
	.w4(32'h39f12b8b),
	.w5(32'hbc9a1471),
	.w6(32'hbb05c794),
	.w7(32'hba566281),
	.w8(32'h3ac8c5e2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89e221),
	.w1(32'h3a6252eb),
	.w2(32'hbb122d34),
	.w3(32'hbad2939f),
	.w4(32'h3c7bdea7),
	.w5(32'hb908045f),
	.w6(32'hbbd1456a),
	.w7(32'hbc20e200),
	.w8(32'h3a75bc80),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc3acd),
	.w1(32'h3a8fc2dc),
	.w2(32'h3b11405b),
	.w3(32'hbb978bde),
	.w4(32'hbb80b649),
	.w5(32'h3bf99453),
	.w6(32'hbb8049f7),
	.w7(32'h3a124e67),
	.w8(32'h3c8e63e9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be298),
	.w1(32'h39a12925),
	.w2(32'h3c1692dd),
	.w3(32'hbc883cd8),
	.w4(32'hba0556a9),
	.w5(32'h3c010df6),
	.w6(32'h3986607c),
	.w7(32'hbc0f6d67),
	.w8(32'h3c2fad66),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e55d),
	.w1(32'hbb41e6dc),
	.w2(32'h3c7d78ee),
	.w3(32'h3a4d433e),
	.w4(32'hba1ace41),
	.w5(32'h3bb3a5b7),
	.w6(32'h391f518e),
	.w7(32'hbb265e41),
	.w8(32'hbb5d53f4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2362c),
	.w1(32'hbb9f746b),
	.w2(32'h3b9e6de9),
	.w3(32'h3c05f8d0),
	.w4(32'h3b996396),
	.w5(32'hbc2044b3),
	.w6(32'h3ad8c619),
	.w7(32'h3c5dc753),
	.w8(32'hbcef8daa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule