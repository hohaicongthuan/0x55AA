module layer_8_featuremap_9(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a88d4),
	.w1(32'h3bdc58ec),
	.w2(32'hbbdcdcf5),
	.w3(32'h3c05151d),
	.w4(32'h3c11f65f),
	.w5(32'hba4eb4a5),
	.w6(32'h3ce17613),
	.w7(32'h3c31b796),
	.w8(32'h3bf3370f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a205269),
	.w1(32'hba6d7bd6),
	.w2(32'h3bba1648),
	.w3(32'h3bb39285),
	.w4(32'hb993b0d1),
	.w5(32'h3bb44311),
	.w6(32'h3c2091da),
	.w7(32'h3b222134),
	.w8(32'h3b603735),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f468),
	.w1(32'hbb91f18e),
	.w2(32'h3bbeee48),
	.w3(32'h3b8709c1),
	.w4(32'hbb612743),
	.w5(32'h3ba65d67),
	.w6(32'h3b09ae04),
	.w7(32'hbb61e34f),
	.w8(32'h3b879842),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92d697),
	.w1(32'hbc3b8a28),
	.w2(32'hba001119),
	.w3(32'h3b915397),
	.w4(32'hbbbda264),
	.w5(32'h3a2d25b3),
	.w6(32'h3bfc635c),
	.w7(32'hbba36004),
	.w8(32'h39e69de2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6913b),
	.w1(32'hbbc5cf85),
	.w2(32'hbc31c3d7),
	.w3(32'h3b6ccc40),
	.w4(32'hbc351590),
	.w5(32'hbc6e4609),
	.w6(32'h3c066326),
	.w7(32'hba1da928),
	.w8(32'hbb778f24),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ede5),
	.w1(32'h3bb5e966),
	.w2(32'hbbc5ef4f),
	.w3(32'hbc2df377),
	.w4(32'hbc42c579),
	.w5(32'hbc4a486c),
	.w6(32'hbb9de9c1),
	.w7(32'h3a994283),
	.w8(32'hbca0d687),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bea90),
	.w1(32'hbc24f071),
	.w2(32'h3baa7662),
	.w3(32'hbbcf3131),
	.w4(32'hbbe1f840),
	.w5(32'h3c09bce9),
	.w6(32'hbb66045e),
	.w7(32'hbc0be75b),
	.w8(32'h3bd79157),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57ce69),
	.w1(32'h3b4bd3fc),
	.w2(32'h3a12d6f9),
	.w3(32'h3a903891),
	.w4(32'hbbf65164),
	.w5(32'h3ac7efa0),
	.w6(32'h3bc9a45d),
	.w7(32'hbc226b2b),
	.w8(32'hbc750ba1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5f134),
	.w1(32'hbbc3249e),
	.w2(32'hbb84d2aa),
	.w3(32'hbbf3aa25),
	.w4(32'hbbb24909),
	.w5(32'hbc0c8f12),
	.w6(32'hbb5c011b),
	.w7(32'hbb5154a3),
	.w8(32'hbc01c7ed),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68486f),
	.w1(32'h3b77be4a),
	.w2(32'h3aab2e48),
	.w3(32'hba41bc7c),
	.w4(32'hbc1794d8),
	.w5(32'h3c59393c),
	.w6(32'h3a618e3b),
	.w7(32'h3bf81b53),
	.w8(32'hbb50c9af),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982729),
	.w1(32'hbceb25a8),
	.w2(32'hbb8978bf),
	.w3(32'h3ba9c742),
	.w4(32'hbc8f4ff5),
	.w5(32'hbbe9f496),
	.w6(32'h3c7f6bce),
	.w7(32'hbc8a01a6),
	.w8(32'hbbff10fc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06dd65),
	.w1(32'hbc597152),
	.w2(32'h3b1a4454),
	.w3(32'hbc4ade9a),
	.w4(32'hbbed7e8c),
	.w5(32'h3bdb8330),
	.w6(32'hbb56c550),
	.w7(32'h3c2bc2bc),
	.w8(32'h3c32257c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8952dd),
	.w1(32'hbcd37b7c),
	.w2(32'h3c692469),
	.w3(32'h3b749802),
	.w4(32'hbc6ad4a2),
	.w5(32'h3cb133d6),
	.w6(32'h3b7b311c),
	.w7(32'hbc051b1a),
	.w8(32'hbbb59b81),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb65fb2),
	.w1(32'hbbaa216b),
	.w2(32'h3b28ff68),
	.w3(32'hbbb03689),
	.w4(32'hbbabc2ad),
	.w5(32'h3b1131c1),
	.w6(32'h3c686f93),
	.w7(32'hbbdc9a12),
	.w8(32'h3b1a3cb1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc436e3),
	.w1(32'hbbf10a8c),
	.w2(32'h3b46a2b8),
	.w3(32'h3bbd2ccf),
	.w4(32'hb9169191),
	.w5(32'h3c0fd37f),
	.w6(32'h3c1ba128),
	.w7(32'hbbbf58dd),
	.w8(32'h3bd7bab0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c87b),
	.w1(32'hba3ced5e),
	.w2(32'hbba420be),
	.w3(32'h3b10a76e),
	.w4(32'hbb030708),
	.w5(32'hbb7a2770),
	.w6(32'hbad1b586),
	.w7(32'hbb68f596),
	.w8(32'hbc060a94),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f5fef),
	.w1(32'hbc943fee),
	.w2(32'h3c10d6be),
	.w3(32'hbba76b38),
	.w4(32'h3bd18afd),
	.w5(32'h3ae86bb5),
	.w6(32'hbbb2f541),
	.w7(32'h3aa58b3d),
	.w8(32'hbc1d5142),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69419),
	.w1(32'h3b14a976),
	.w2(32'h3ade568c),
	.w3(32'hbc11f60e),
	.w4(32'h399bdb29),
	.w5(32'hba7faacd),
	.w6(32'hba8284d2),
	.w7(32'h3afb2fed),
	.w8(32'hba816905),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68e65a),
	.w1(32'hbd28f564),
	.w2(32'hbc64b66e),
	.w3(32'hbb8ec900),
	.w4(32'hbd2ca8a5),
	.w5(32'h3c961e38),
	.w6(32'h3cca1f57),
	.w7(32'h3c87cc1c),
	.w8(32'hbb361d8a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba36d0f),
	.w1(32'hbccf9c89),
	.w2(32'hbc863e64),
	.w3(32'h3c363e2a),
	.w4(32'hbc856237),
	.w5(32'hbb829cd7),
	.w6(32'h3cd15eeb),
	.w7(32'hba12438c),
	.w8(32'h3b07908e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1af80c),
	.w1(32'hbcd711f1),
	.w2(32'h3af81610),
	.w3(32'h3c1b7cd2),
	.w4(32'hbc6f44e3),
	.w5(32'h3be27be4),
	.w6(32'h3c21892b),
	.w7(32'hbc9caac5),
	.w8(32'h3c189a2d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e1347c),
	.w1(32'h3c29c3bd),
	.w2(32'hbbb5efd9),
	.w3(32'h3abd3c64),
	.w4(32'hbc80c1c7),
	.w5(32'h3caa65c1),
	.w6(32'h3bc5a703),
	.w7(32'h3c01c946),
	.w8(32'hbb55dcf4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c814d94),
	.w1(32'hbcd2a282),
	.w2(32'hbc153472),
	.w3(32'h3c53e2f6),
	.w4(32'hbd01ca6b),
	.w5(32'h3cc0adfa),
	.w6(32'h3cd16f8f),
	.w7(32'h3cd7a076),
	.w8(32'hbb04833c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3a9df),
	.w1(32'hbcb0cb99),
	.w2(32'h3a908beb),
	.w3(32'hbb476ed7),
	.w4(32'hbc6dcb88),
	.w5(32'h3bc8f98a),
	.w6(32'h3ccbf824),
	.w7(32'hbc8babf8),
	.w8(32'h3b1e429e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4238ea),
	.w1(32'hbc54a577),
	.w2(32'h3b8cb2c2),
	.w3(32'h3b81d366),
	.w4(32'hb9b8ccb2),
	.w5(32'hbcab15ee),
	.w6(32'h3b881989),
	.w7(32'hbc531cfc),
	.w8(32'hbbaca348),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb548e),
	.w1(32'hbb25d145),
	.w2(32'h3ab450e9),
	.w3(32'hbbdae879),
	.w4(32'h3b8e35fa),
	.w5(32'hbbfe8680),
	.w6(32'h3c28f554),
	.w7(32'h3c835a32),
	.w8(32'h3bc23216),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5abcfb),
	.w1(32'hbc2e77ac),
	.w2(32'h3bf7b419),
	.w3(32'hbb18d51f),
	.w4(32'hbbd3f050),
	.w5(32'h3c47b490),
	.w6(32'hbac0d886),
	.w7(32'hbc195d2b),
	.w8(32'h3c23bd43),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82eea6),
	.w1(32'hbd604388),
	.w2(32'hbdb82188),
	.w3(32'hbd1f6b41),
	.w4(32'hbce1ba87),
	.w5(32'hbd68e559),
	.w6(32'hbc6dfd1e),
	.w7(32'h3d1d1d81),
	.w8(32'hbaa25559),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268a11),
	.w1(32'hbae0b8cf),
	.w2(32'hbc1c6ba6),
	.w3(32'h3c5f53a5),
	.w4(32'hbb1098c8),
	.w5(32'hbb94d8b1),
	.w6(32'h3b3fdb8a),
	.w7(32'h3afb61c5),
	.w8(32'hbc049b6d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075fdf),
	.w1(32'hba3198fe),
	.w2(32'h399af146),
	.w3(32'hbb8f3b7f),
	.w4(32'h3a50c0f0),
	.w5(32'hb91ec4bb),
	.w6(32'hbbdd93c9),
	.w7(32'hba9a8a9f),
	.w8(32'hbba92c00),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c280f),
	.w1(32'hbc3b5f49),
	.w2(32'hbc5ce659),
	.w3(32'h39a79ba9),
	.w4(32'hbc68838f),
	.w5(32'hbbd84ea1),
	.w6(32'hbac23946),
	.w7(32'hbbe4ca1e),
	.w8(32'hbb98c3e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba882e9),
	.w1(32'hbc099616),
	.w2(32'h3b8c83e4),
	.w3(32'hbc649b0e),
	.w4(32'hbb80c433),
	.w5(32'h3c22b0ee),
	.w6(32'hbc5a9c3f),
	.w7(32'hbb93ee10),
	.w8(32'h3bdb8c9d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb026c7),
	.w1(32'hbb430723),
	.w2(32'h3aa2f154),
	.w3(32'hba6ff42d),
	.w4(32'hbb2ceb0c),
	.w5(32'hba65d299),
	.w6(32'hbb3dbb4b),
	.w7(32'hbb1871f4),
	.w8(32'h3a02c9cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fcedf),
	.w1(32'hbb0e1ad0),
	.w2(32'h3c0eb38c),
	.w3(32'hba0d5fa6),
	.w4(32'hbac526a1),
	.w5(32'h3c8c167d),
	.w6(32'h395d18c8),
	.w7(32'hbb3e3bb7),
	.w8(32'hb9466ed0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c837a2a),
	.w1(32'h3babaa6c),
	.w2(32'h3a9efb48),
	.w3(32'h3c47c7a4),
	.w4(32'h3c136697),
	.w5(32'h3af73583),
	.w6(32'h3bdafd83),
	.w7(32'h3b9f9b6a),
	.w8(32'hbb07f4c2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac3532),
	.w1(32'hbac51796),
	.w2(32'hbc0aae66),
	.w3(32'hbb84b5ad),
	.w4(32'h3b876398),
	.w5(32'hbb454c21),
	.w6(32'h3b82918b),
	.w7(32'h3c914981),
	.w8(32'h3a042a32),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25e6b4),
	.w1(32'hbcaaf812),
	.w2(32'hb8e87d19),
	.w3(32'h3bb96882),
	.w4(32'hbc0b49f9),
	.w5(32'h3c7ced5a),
	.w6(32'h3c002ce0),
	.w7(32'h3a54cdd0),
	.w8(32'h3bfa763c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb980980),
	.w1(32'hbc278f04),
	.w2(32'hb9ba2a6c),
	.w3(32'hbb82891f),
	.w4(32'h3bd07bf4),
	.w5(32'h3b11fb12),
	.w6(32'h3acd5c5d),
	.w7(32'h3c116d65),
	.w8(32'hbbdcd14e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dec4f),
	.w1(32'h3aa78e3c),
	.w2(32'hbc73608d),
	.w3(32'hbc16c406),
	.w4(32'hbc195148),
	.w5(32'hbc3554f9),
	.w6(32'hbba8a986),
	.w7(32'hbb6d0a73),
	.w8(32'hbc55b290),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b94c8a),
	.w1(32'h3c8a61e8),
	.w2(32'h3bd65991),
	.w3(32'h3b4ade7a),
	.w4(32'h3c84e6bc),
	.w5(32'h3c044a41),
	.w6(32'hb8d0de5a),
	.w7(32'h3cb7cc50),
	.w8(32'h3c4b549e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b791),
	.w1(32'hbc57489a),
	.w2(32'h3c09ed38),
	.w3(32'h3c0e7018),
	.w4(32'h3c1f2ba5),
	.w5(32'h3b636619),
	.w6(32'h3bed6cdf),
	.w7(32'hbc0904d7),
	.w8(32'hbb67487d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc197fe4),
	.w1(32'hbc5831f1),
	.w2(32'hb8e8e244),
	.w3(32'hbbb46551),
	.w4(32'hbc4018f0),
	.w5(32'h3aa678d1),
	.w6(32'h3c901a9b),
	.w7(32'hbc04eb7c),
	.w8(32'h3b728c2e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e32cd),
	.w1(32'h3c00e287),
	.w2(32'hba278eda),
	.w3(32'h3b702bde),
	.w4(32'h3b995de9),
	.w5(32'hbb80f91d),
	.w6(32'h3bb9e1d7),
	.w7(32'h3b969a96),
	.w8(32'hbaea1219),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a00c0e),
	.w1(32'hbbd3b06e),
	.w2(32'hbc347fb6),
	.w3(32'hbb1e60a3),
	.w4(32'h3bb74f1f),
	.w5(32'h3ad93f6d),
	.w6(32'h391dd8f6),
	.w7(32'hbc85e945),
	.w8(32'h3bcbd171),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c738dc1),
	.w1(32'hbc22e627),
	.w2(32'hbc0fb97a),
	.w3(32'hbbdca2d0),
	.w4(32'hbd09ade5),
	.w5(32'h3c6f29b9),
	.w6(32'h3cfd2c47),
	.w7(32'h3c8fd0ac),
	.w8(32'hba0e1326),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68a41d),
	.w1(32'hbbca38a6),
	.w2(32'h3a2893c7),
	.w3(32'hbc770cfa),
	.w4(32'hbbeeb177),
	.w5(32'h3b56bddb),
	.w6(32'h3c5f53d3),
	.w7(32'hbc145802),
	.w8(32'h3bf8c979),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93b2b0),
	.w1(32'hbc122a88),
	.w2(32'hbc8578e3),
	.w3(32'h3af1b398),
	.w4(32'hbc85522b),
	.w5(32'h3bbaf133),
	.w6(32'h3b696f7f),
	.w7(32'hbc40c78b),
	.w8(32'hbbe24420),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c431c7c),
	.w1(32'h3b24d74c),
	.w2(32'h3d07b4f7),
	.w3(32'hbbfdf9d4),
	.w4(32'h3baa0094),
	.w5(32'h3d307aae),
	.w6(32'h3c7228d7),
	.w7(32'h3d155f1c),
	.w8(32'h3d17d72e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc7634),
	.w1(32'h39fbc91b),
	.w2(32'hbbde77f0),
	.w3(32'h3d32df88),
	.w4(32'hbb651bf9),
	.w5(32'hbbc75256),
	.w6(32'hbac38118),
	.w7(32'h3a95b61c),
	.w8(32'hbb2a730f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8d281),
	.w1(32'hbd91748a),
	.w2(32'h3e1947bd),
	.w3(32'hba68a47e),
	.w4(32'h3e1c3eb4),
	.w5(32'hbe5ea547),
	.w6(32'h3b805414),
	.w7(32'hbda9fffb),
	.w8(32'h3d668fdf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbd0391),
	.w1(32'h3a07e3fe),
	.w2(32'h3a9e55d6),
	.w3(32'h3d787b31),
	.w4(32'hbb30cf82),
	.w5(32'h3c39a4c4),
	.w6(32'h3d06c298),
	.w7(32'h3ac75ced),
	.w8(32'h3b9873cc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce4494),
	.w1(32'hbc3a0c94),
	.w2(32'hbc7393ce),
	.w3(32'hbc95c505),
	.w4(32'hbcd549e2),
	.w5(32'hbcb8bbc8),
	.w6(32'h3b33b7f2),
	.w7(32'hba6b1455),
	.w8(32'hbc2f1512),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b283ada),
	.w1(32'hba8fc1b6),
	.w2(32'hbc48d44c),
	.w3(32'hbb86d69a),
	.w4(32'hbd133202),
	.w5(32'hbafad9c1),
	.w6(32'h3be03be0),
	.w7(32'hbc1f32fb),
	.w8(32'hbc99ffd4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302114),
	.w1(32'hbc406f65),
	.w2(32'hbbaedb2f),
	.w3(32'hbc330132),
	.w4(32'hbc1233b6),
	.w5(32'h3bdad4ef),
	.w6(32'hbc810867),
	.w7(32'hbaf21496),
	.w8(32'h3cb0e98b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b9aa),
	.w1(32'hb709b5f5),
	.w2(32'hbbd3461b),
	.w3(32'h3c15db4d),
	.w4(32'hbc2da9ab),
	.w5(32'hbc52d825),
	.w6(32'h3b143f5b),
	.w7(32'hbc4bbc3d),
	.w8(32'h3c5f2eba),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec35ba),
	.w1(32'hbbda6d1d),
	.w2(32'hbc803c35),
	.w3(32'h3cae61da),
	.w4(32'h3a9ee1da),
	.w5(32'hbb051c1d),
	.w6(32'h3af68fbf),
	.w7(32'h3c20b167),
	.w8(32'h3b19ca04),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba640dc3),
	.w1(32'hba35658e),
	.w2(32'h3b640d77),
	.w3(32'hbaf3c643),
	.w4(32'h3b635f46),
	.w5(32'h3c149eee),
	.w6(32'hbb2200a0),
	.w7(32'h3a8ed515),
	.w8(32'h3bbcb08c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73387),
	.w1(32'h3aa61275),
	.w2(32'h3a8f4fd0),
	.w3(32'h3b5d83d0),
	.w4(32'hbc0b5ee8),
	.w5(32'hbc42dc7d),
	.w6(32'h3c21785f),
	.w7(32'hba575434),
	.w8(32'hbbfac5c9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba266651),
	.w1(32'hbacf4820),
	.w2(32'hbc076a86),
	.w3(32'hbc1f7ad8),
	.w4(32'hbaee9f5e),
	.w5(32'hbbf20b60),
	.w6(32'h3b85b4a4),
	.w7(32'h38f2570e),
	.w8(32'hbbbf8537),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b9f0c),
	.w1(32'hbd39e067),
	.w2(32'hbc29c1a2),
	.w3(32'hbb3c92ea),
	.w4(32'hbc98bdcf),
	.w5(32'hbd0dbf13),
	.w6(32'hbbf2825d),
	.w7(32'hbd03ad8a),
	.w8(32'hbd1b5f6f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca24696),
	.w1(32'hba71dcfd),
	.w2(32'hb970da17),
	.w3(32'hbd497fde),
	.w4(32'h3b9996d7),
	.w5(32'h3bdc4792),
	.w6(32'hbb9eb0f5),
	.w7(32'h3b8e81b4),
	.w8(32'h3c0fb072),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9866),
	.w1(32'hb9a88e6f),
	.w2(32'h3bff7562),
	.w3(32'h3bc4208c),
	.w4(32'hbb653b3c),
	.w5(32'h3bbdd7e5),
	.w6(32'hbb432267),
	.w7(32'hba737725),
	.w8(32'hbb6e97dd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4115),
	.w1(32'hbc0993d9),
	.w2(32'hbc697f28),
	.w3(32'hbbe32334),
	.w4(32'hbbccc72d),
	.w5(32'hbc53b89f),
	.w6(32'h3c05adb4),
	.w7(32'h3bcc6c14),
	.w8(32'hbb14ad33),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa00155),
	.w1(32'hbc37d210),
	.w2(32'hbb8f86e0),
	.w3(32'hbb18c35b),
	.w4(32'hbcfe4e4d),
	.w5(32'hbc26b00d),
	.w6(32'h3a90bb1c),
	.w7(32'hbcb218dd),
	.w8(32'h3c58d09d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4314da),
	.w1(32'h3b156112),
	.w2(32'h3c5f5fe7),
	.w3(32'h3c80da31),
	.w4(32'hbaca0470),
	.w5(32'h3c4bc07a),
	.w6(32'hba92b435),
	.w7(32'hba6f8fda),
	.w8(32'h3c3d8259),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ffc9),
	.w1(32'hba83062e),
	.w2(32'h3a13333c),
	.w3(32'hbba21e40),
	.w4(32'hba7e217e),
	.w5(32'h3973a105),
	.w6(32'hbaaeed45),
	.w7(32'h3b5f4659),
	.w8(32'h395ca54e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca99d2),
	.w1(32'h3adabc5a),
	.w2(32'hbbb0728b),
	.w3(32'h39655069),
	.w4(32'h3ab5de8b),
	.w5(32'hbbbfaca4),
	.w6(32'h3ab3f03d),
	.w7(32'h3b5c3dbf),
	.w8(32'hbbe4e792),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1efee6),
	.w1(32'hbc328a1b),
	.w2(32'hbc259d27),
	.w3(32'hba32d32b),
	.w4(32'hbc144731),
	.w5(32'h3b37a614),
	.w6(32'h3b8d15ce),
	.w7(32'hb7c092dc),
	.w8(32'h3c1b6b5b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2925c),
	.w1(32'hb86398ed),
	.w2(32'h3c033a37),
	.w3(32'h3c304b89),
	.w4(32'hba9f665b),
	.w5(32'h3c0cc67f),
	.w6(32'h3c248df9),
	.w7(32'hbb1a0097),
	.w8(32'h3c17403e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13a0a2),
	.w1(32'hbbf0054c),
	.w2(32'hbc256140),
	.w3(32'hbb8ef1bb),
	.w4(32'hbc37bd6f),
	.w5(32'hbb5a0a65),
	.w6(32'h3bfcb4b0),
	.w7(32'h3b093571),
	.w8(32'hbc0b119c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0d62),
	.w1(32'h3b7938a5),
	.w2(32'hb9e4e436),
	.w3(32'h3c240608),
	.w4(32'h3adc11a6),
	.w5(32'h3a04f036),
	.w6(32'hbb63d2eb),
	.w7(32'h3b0b6baf),
	.w8(32'hbb11b640),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a447d),
	.w1(32'hbb4e7d32),
	.w2(32'hbbd2f7ec),
	.w3(32'hbbf9212d),
	.w4(32'hbcf9c981),
	.w5(32'hbce2c3a8),
	.w6(32'h3b28c231),
	.w7(32'hbc88d3eb),
	.w8(32'hbd61c1b4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c356),
	.w1(32'hbb0408f6),
	.w2(32'hb8be3fe1),
	.w3(32'h3b2bdc73),
	.w4(32'hbb151cb9),
	.w5(32'hbb290dad),
	.w6(32'hbcb08486),
	.w7(32'h3a6b5195),
	.w8(32'h39aba712),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50523a),
	.w1(32'h3c11fc29),
	.w2(32'hbc721e65),
	.w3(32'h3b48b708),
	.w4(32'h3ad1f4ab),
	.w5(32'h3a0cbacb),
	.w6(32'h3bb6e99a),
	.w7(32'hba89b5d4),
	.w8(32'h3c5a7ecc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b7219),
	.w1(32'hbbd73eed),
	.w2(32'hbb612e67),
	.w3(32'hbb713500),
	.w4(32'hbb4cb747),
	.w5(32'hbc3c234c),
	.w6(32'hbc43f608),
	.w7(32'h3b19ba4c),
	.w8(32'hba87dd37),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4df9c0),
	.w1(32'h3b32b1a1),
	.w2(32'h3c53fe27),
	.w3(32'h3addf460),
	.w4(32'hbb9b0b00),
	.w5(32'h3b95945c),
	.w6(32'hbb220621),
	.w7(32'h3b8f59d8),
	.w8(32'hbc84521b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31a300),
	.w1(32'hbc883d43),
	.w2(32'hbd345dbc),
	.w3(32'h3ccd438d),
	.w4(32'h3d3ceb29),
	.w5(32'h3cf1ebd3),
	.w6(32'h3c092b93),
	.w7(32'hbc1afc88),
	.w8(32'h3d685f4f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce05c0e),
	.w1(32'hbc398b0e),
	.w2(32'hbca02715),
	.w3(32'hbd05e65a),
	.w4(32'h3a6db20a),
	.w5(32'hbc3ad42e),
	.w6(32'h3d228c7e),
	.w7(32'h3c4578ee),
	.w8(32'h3c0b6832),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba40920),
	.w1(32'h3b95a3cb),
	.w2(32'h3ba0c221),
	.w3(32'hbc1cd37d),
	.w4(32'hbafef602),
	.w5(32'h3b0c1d1f),
	.w6(32'h3a612722),
	.w7(32'hbb0ec4c1),
	.w8(32'hbc0a3031),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16c692),
	.w1(32'hbb7197be),
	.w2(32'hbba26667),
	.w3(32'h3c034cca),
	.w4(32'h3c5526a3),
	.w5(32'h3c60abf1),
	.w6(32'hbabc1e8f),
	.w7(32'hb9aafd45),
	.w8(32'hba9b5ce4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4796ff),
	.w1(32'hbc28cb05),
	.w2(32'h3c1745c7),
	.w3(32'h3c65331a),
	.w4(32'hbc5cf02b),
	.w5(32'hbd06b8f2),
	.w6(32'hbad217f9),
	.w7(32'h3be41f33),
	.w8(32'hbd34b82c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c997580),
	.w1(32'hb9eae9b6),
	.w2(32'hb8ae3686),
	.w3(32'h3c970c3f),
	.w4(32'h3b5267a3),
	.w5(32'h3a483fcd),
	.w6(32'hbb26d74f),
	.w7(32'h3b11fd92),
	.w8(32'h3b167c4b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195d7c),
	.w1(32'h3b5a5d2b),
	.w2(32'h3caac5d4),
	.w3(32'h3ab15a04),
	.w4(32'hbce7aaf6),
	.w5(32'h3cea4cde),
	.w6(32'h3c44b9cb),
	.w7(32'hbc3c3f23),
	.w8(32'hbd238dfd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87e81b),
	.w1(32'hbb187823),
	.w2(32'hbb0fd4f0),
	.w3(32'h3d00602e),
	.w4(32'hbb8be30f),
	.w5(32'hbb9094d4),
	.w6(32'hbb76966f),
	.w7(32'hbbb22b39),
	.w8(32'hbc7ca63e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f5026),
	.w1(32'hbbf8f41e),
	.w2(32'hbbfccfea),
	.w3(32'h3b99223c),
	.w4(32'h3bb5fa05),
	.w5(32'hbbc550fe),
	.w6(32'h3c89e447),
	.w7(32'h3cbf5d0d),
	.w8(32'h3c708a45),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8028),
	.w1(32'hbb751ff4),
	.w2(32'h3d18e95d),
	.w3(32'h3bc9e857),
	.w4(32'hbcc4f4b9),
	.w5(32'hbca57234),
	.w6(32'h3c3e522c),
	.w7(32'h3c42ee37),
	.w8(32'hbc3bc434),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1787cc),
	.w1(32'h3c9a487b),
	.w2(32'h3c0e3e5a),
	.w3(32'h3c99fef5),
	.w4(32'hbc9252a1),
	.w5(32'h3c18299d),
	.w6(32'hbc357732),
	.w7(32'hbd2ad03f),
	.w8(32'hbd1d6136),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb614af6),
	.w1(32'h3b59d463),
	.w2(32'h3b7eb03d),
	.w3(32'h3cd37125),
	.w4(32'hbabdc608),
	.w5(32'hbb8a8f33),
	.w6(32'h3b8629e9),
	.w7(32'h39cef18d),
	.w8(32'hbbcafb0f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f2508),
	.w1(32'h3bb062b5),
	.w2(32'h3c923bcc),
	.w3(32'hbb7d4de4),
	.w4(32'h3c14f928),
	.w5(32'h3a86b9c8),
	.w6(32'hbbdc376a),
	.w7(32'h3caa3bfb),
	.w8(32'h38050fbc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca68cc2),
	.w1(32'hbbc0b07d),
	.w2(32'hbc2a2525),
	.w3(32'h3ca1fc42),
	.w4(32'hbbe36dad),
	.w5(32'hbc58b74b),
	.w6(32'h3c2f0a9c),
	.w7(32'hbbd25631),
	.w8(32'hbc8a4992),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5254d8),
	.w1(32'hbb94436c),
	.w2(32'hbbbbded6),
	.w3(32'hbb9966c7),
	.w4(32'hba5801ca),
	.w5(32'hbc28a323),
	.w6(32'hbbf6d308),
	.w7(32'h3ad19a31),
	.w8(32'hbc0cbd88),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53965),
	.w1(32'h3bc36fb8),
	.w2(32'h3b7dc0a4),
	.w3(32'h3a4ce8f5),
	.w4(32'h3b7a92d6),
	.w5(32'h3c6654c9),
	.w6(32'hbb55761e),
	.w7(32'hbc9b5250),
	.w8(32'hbd0c1833),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb06fc8),
	.w1(32'hbc0887fc),
	.w2(32'hbc376228),
	.w3(32'h3cde66d9),
	.w4(32'hbb039f06),
	.w5(32'hbbb1ad14),
	.w6(32'hbaf5bf99),
	.w7(32'hbb8d9169),
	.w8(32'hbaf97ffd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd483),
	.w1(32'h3a89a63b),
	.w2(32'hbb3a7b0b),
	.w3(32'hbc0594c0),
	.w4(32'h3b94a3b4),
	.w5(32'h3b33faf1),
	.w6(32'hba45de9b),
	.w7(32'h3b88bd51),
	.w8(32'h39e1d9f5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27f7c9),
	.w1(32'hbbbfc754),
	.w2(32'h3c1ace60),
	.w3(32'h3b9b8457),
	.w4(32'hbc487858),
	.w5(32'hbb51eb8e),
	.w6(32'h3b95ed51),
	.w7(32'h3b8abe87),
	.w8(32'hbb4ca20c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2844dc),
	.w1(32'h3a2f01e7),
	.w2(32'h3b9186b0),
	.w3(32'h3bd283fe),
	.w4(32'hbb91e1d3),
	.w5(32'hbc0a6743),
	.w6(32'h3c46e978),
	.w7(32'hbb26fb86),
	.w8(32'hbbf8acba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a55e2),
	.w1(32'hbb1fc3d6),
	.w2(32'hba7845c4),
	.w3(32'h3a3d21d4),
	.w4(32'h3ae7954a),
	.w5(32'hbabb8bdc),
	.w6(32'h3c26846b),
	.w7(32'h3c8ae083),
	.w8(32'h3b383033),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b9aed),
	.w1(32'h3aa02caa),
	.w2(32'hbbea3099),
	.w3(32'hbbaf10b3),
	.w4(32'h3acb1e69),
	.w5(32'hbb86c718),
	.w6(32'hba1b7e2e),
	.w7(32'h3c086844),
	.w8(32'hbc6c4493),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafa190),
	.w1(32'h3b1a1e07),
	.w2(32'hba905ddc),
	.w3(32'hbc311972),
	.w4(32'h3abcfd30),
	.w5(32'h3b1f21ca),
	.w6(32'hbb5602e3),
	.w7(32'h3a65648d),
	.w8(32'h3aaf8db7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d5b4a),
	.w1(32'hbbfddce5),
	.w2(32'h3b69bfc2),
	.w3(32'h39d8d4a9),
	.w4(32'hbc61f202),
	.w5(32'hbad37db1),
	.w6(32'h3a570c01),
	.w7(32'hbca45c5f),
	.w8(32'hbc1cf17f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f43fd),
	.w1(32'h3c855908),
	.w2(32'h3bd92ccb),
	.w3(32'hbbfcfc62),
	.w4(32'hbb0a05a2),
	.w5(32'h3c844794),
	.w6(32'hbc02c784),
	.w7(32'hbc9c71f6),
	.w8(32'hbc1dcbbf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad4de6),
	.w1(32'h3b63990e),
	.w2(32'hbc955520),
	.w3(32'h3c3dd1ca),
	.w4(32'h3c905149),
	.w5(32'h3c279a7f),
	.w6(32'h3c9787b3),
	.w7(32'h3c1492bf),
	.w8(32'h3d1f5f0f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a564a5e),
	.w1(32'h3bbebcb4),
	.w2(32'hbc2e2b6d),
	.w3(32'hbd00e2b3),
	.w4(32'h3b4a5748),
	.w5(32'h3d0baeba),
	.w6(32'h3bb91b3c),
	.w7(32'hbd0b0ea1),
	.w8(32'hbcc9cda2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19f5f3),
	.w1(32'hb9d655af),
	.w2(32'h3c37e88f),
	.w3(32'h3c2dce6f),
	.w4(32'hbc28587d),
	.w5(32'h3c9ddf64),
	.w6(32'hbb7442d0),
	.w7(32'hbbce0fa1),
	.w8(32'hbbd7e1dc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14be42),
	.w1(32'h3b8d0f8c),
	.w2(32'h3b6ed090),
	.w3(32'hbb44aaad),
	.w4(32'h3b8e08ca),
	.w5(32'hbb356a0a),
	.w6(32'h3c2a3688),
	.w7(32'hbb82e149),
	.w8(32'h3bbf09bd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28726c),
	.w1(32'hbb425f28),
	.w2(32'hbba09064),
	.w3(32'hbb3b9e30),
	.w4(32'hb93862ac),
	.w5(32'hbb8134a3),
	.w6(32'h3c5a3815),
	.w7(32'h3bf08a9b),
	.w8(32'h3b97b489),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37b883),
	.w1(32'h3b26a911),
	.w2(32'h3b02a7b2),
	.w3(32'h3c09ace5),
	.w4(32'h3b3abbce),
	.w5(32'h3ae7fde3),
	.w6(32'h3c291bee),
	.w7(32'h3bb8d4d1),
	.w8(32'h3ab67e6c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fa8d7),
	.w1(32'h3bfb973c),
	.w2(32'hbc6ab324),
	.w3(32'h3ba7c99d),
	.w4(32'h3a843237),
	.w5(32'h3cb8bfd9),
	.w6(32'h3bb85689),
	.w7(32'hbc14863c),
	.w8(32'hb96bd574),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee89ab),
	.w1(32'h3b9f57c2),
	.w2(32'hba86b89a),
	.w3(32'h3b16648f),
	.w4(32'h3c8a0c5f),
	.w5(32'h3d301b46),
	.w6(32'h3ca3e339),
	.w7(32'hbca6ff2f),
	.w8(32'h3bf09e44),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbaf145),
	.w1(32'hbc037e75),
	.w2(32'h3cd304b5),
	.w3(32'h3c8dc7d0),
	.w4(32'hbd1fec62),
	.w5(32'hbc9a2ac9),
	.w6(32'h3ce4f945),
	.w7(32'hbc4b6171),
	.w8(32'hbce61d57),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cacd643),
	.w1(32'hba618859),
	.w2(32'hbc8069f1),
	.w3(32'h3cce4036),
	.w4(32'h3c11dcce),
	.w5(32'hbc00e3ea),
	.w6(32'hbc62f32a),
	.w7(32'h389fc36c),
	.w8(32'hbc907503),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca77fd1),
	.w1(32'h3a6a3fcc),
	.w2(32'h3c16aa9e),
	.w3(32'hbca09c3f),
	.w4(32'hbcc9168e),
	.w5(32'h3ca2e96d),
	.w6(32'h3af24d26),
	.w7(32'hbc8f1c56),
	.w8(32'hbcd6c03e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc494942),
	.w1(32'h3c6057ec),
	.w2(32'h3c3bd3fd),
	.w3(32'h3d195df4),
	.w4(32'h36ca25c8),
	.w5(32'h3bb60d67),
	.w6(32'h3cd2865b),
	.w7(32'hbc1072af),
	.w8(32'hbc18c581),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298099),
	.w1(32'hbac3a490),
	.w2(32'h3aaabece),
	.w3(32'hbae4cec9),
	.w4(32'hbb0f9c79),
	.w5(32'hbc43fb45),
	.w6(32'hbb60fc03),
	.w7(32'h3c0febcb),
	.w8(32'h387ae446),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f22ed),
	.w1(32'h3a989e54),
	.w2(32'hba2d4a6c),
	.w3(32'hbb976a13),
	.w4(32'hbad24449),
	.w5(32'h3bbe0414),
	.w6(32'hbb99fa50),
	.w7(32'hbbf5a190),
	.w8(32'hbc5bd11f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52e15),
	.w1(32'h3ada2361),
	.w2(32'hb7b89522),
	.w3(32'h3be3b7f6),
	.w4(32'h3b7e224d),
	.w5(32'h3b70de28),
	.w6(32'h3bdec6f0),
	.w7(32'h3b631ad4),
	.w8(32'h3a0d1829),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936ac99),
	.w1(32'h3b563914),
	.w2(32'h3b69acdd),
	.w3(32'h3b264244),
	.w4(32'h3bd28f98),
	.w5(32'h3aad13ca),
	.w6(32'h3a0454b7),
	.w7(32'hbb5e174d),
	.w8(32'hbc87fd6b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05069),
	.w1(32'hbb9bea0b),
	.w2(32'h38c5f80c),
	.w3(32'h3cb504f9),
	.w4(32'hbb193e9a),
	.w5(32'hbc53c2c2),
	.w6(32'hbb2a3fbd),
	.w7(32'hb9ac4ac6),
	.w8(32'hba772ec4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf47ab),
	.w1(32'h3bf8a14d),
	.w2(32'h3bf5b915),
	.w3(32'h37b576cf),
	.w4(32'hbc03fb52),
	.w5(32'hbc043a76),
	.w6(32'h3ab85c3a),
	.w7(32'hbce1a4f9),
	.w8(32'h3c6dfdd7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d32f8),
	.w1(32'hb7c0f1ff),
	.w2(32'hba942706),
	.w3(32'hbcb68ddf),
	.w4(32'h3a822c11),
	.w5(32'h3a0ddef4),
	.w6(32'h3be3809e),
	.w7(32'h3a4e0ba4),
	.w8(32'h3a1ccaa0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1948e9),
	.w1(32'h3b4a7aac),
	.w2(32'h3c05bec8),
	.w3(32'h3b6c21a1),
	.w4(32'hbc1ea335),
	.w5(32'h3b257520),
	.w6(32'hbb477a8c),
	.w7(32'hbc6e020c),
	.w8(32'hbca4a248),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31edf1),
	.w1(32'hbc3974d6),
	.w2(32'hbc46fd0d),
	.w3(32'h3c21975b),
	.w4(32'h3b1ebc2a),
	.w5(32'h3b540749),
	.w6(32'hb9b55c2a),
	.w7(32'h385bc692),
	.w8(32'hbc2b901a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a023),
	.w1(32'hbbe601c7),
	.w2(32'hbbbcecff),
	.w3(32'h3bc1f985),
	.w4(32'hbbc1a0cd),
	.w5(32'hbb3d4e70),
	.w6(32'hbbc6b882),
	.w7(32'hbbdda6df),
	.w8(32'hbbb8feef),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39660b),
	.w1(32'h3c05d0a6),
	.w2(32'h3c4f39c5),
	.w3(32'hb9d8e5e3),
	.w4(32'hbc122c72),
	.w5(32'h3bfa881b),
	.w6(32'hbbb1c5a4),
	.w7(32'hbcc2c3d7),
	.w8(32'hbca5d783),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c388f9),
	.w1(32'hbb583554),
	.w2(32'hbbfaff2a),
	.w3(32'h3c39b7dc),
	.w4(32'h3b2205ab),
	.w5(32'hbb8e39da),
	.w6(32'h3c076273),
	.w7(32'h3ac517c4),
	.w8(32'hbb8447a1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d236),
	.w1(32'h3c07677e),
	.w2(32'h3b8e76f1),
	.w3(32'hbbc036fb),
	.w4(32'hbbd247e0),
	.w5(32'h3be4a89c),
	.w6(32'hbbc01f0d),
	.w7(32'hbbb1d475),
	.w8(32'hbce327c5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba608fc0),
	.w1(32'hbaf6815e),
	.w2(32'h3ac2da59),
	.w3(32'h3c540181),
	.w4(32'hba80c4d6),
	.w5(32'hba1f611b),
	.w6(32'h3cc75eb9),
	.w7(32'hbb110ace),
	.w8(32'hbb93b17f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b426),
	.w1(32'h3b97e5e6),
	.w2(32'hbba3c760),
	.w3(32'h3ad116ee),
	.w4(32'h3abbb236),
	.w5(32'h3c5c95b4),
	.w6(32'hbb7d0b5d),
	.w7(32'hbc84e19f),
	.w8(32'hbcd5c8e5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule