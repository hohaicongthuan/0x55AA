module layer_10_featuremap_42(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc81a48),
	.w1(32'h3c5074cf),
	.w2(32'hbb53f416),
	.w3(32'h3c48379f),
	.w4(32'h3ca3a55a),
	.w5(32'h3c3c6d0a),
	.w6(32'h3c6f3523),
	.w7(32'h3c7ef596),
	.w8(32'h3abf01ac),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c8aaf),
	.w1(32'hbc392a4f),
	.w2(32'hbb4bfa15),
	.w3(32'hbb497144),
	.w4(32'hbc58471c),
	.w5(32'hbc2d1c75),
	.w6(32'hbbe59e82),
	.w7(32'hbc2fcc9a),
	.w8(32'hbbfa162f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab357),
	.w1(32'hba0e4609),
	.w2(32'hba70a8ff),
	.w3(32'hbc243c98),
	.w4(32'hbc1c93f2),
	.w5(32'hbb9500ab),
	.w6(32'hbae05913),
	.w7(32'h3b8afd26),
	.w8(32'hbbef6a1f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf87a),
	.w1(32'hbb84d6f9),
	.w2(32'hbc0ef99f),
	.w3(32'hbb3cc82f),
	.w4(32'h3b042046),
	.w5(32'hbc2e9f80),
	.w6(32'h3b93b9b5),
	.w7(32'h3c1c9e51),
	.w8(32'hbc14766b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f0abd),
	.w1(32'hbbf1aef8),
	.w2(32'hbc09ab3b),
	.w3(32'hbbaa0fcb),
	.w4(32'hbc64497c),
	.w5(32'hbbc31ff0),
	.w6(32'hbaae0077),
	.w7(32'hbafdc182),
	.w8(32'hb9242e67),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c0c43),
	.w1(32'hbc6927df),
	.w2(32'hbafcd4ed),
	.w3(32'hbc98848b),
	.w4(32'hbc8aa311),
	.w5(32'hbb0d2425),
	.w6(32'hbc0b50e0),
	.w7(32'hbc29972a),
	.w8(32'h3a8be57e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbcb98),
	.w1(32'hbb5243ca),
	.w2(32'h3c4a01f6),
	.w3(32'hbb9916f0),
	.w4(32'hbbf63612),
	.w5(32'h3c8b1ca5),
	.w6(32'hb8cd5b8a),
	.w7(32'hbae732e3),
	.w8(32'h3adafe0c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8831dc),
	.w1(32'h3be4c6e8),
	.w2(32'hbb9d2e89),
	.w3(32'h3b6792c2),
	.w4(32'hbae70a27),
	.w5(32'hbcc59ee1),
	.w6(32'hbadede81),
	.w7(32'hbbc9487f),
	.w8(32'hbcfe0a51),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d5542),
	.w1(32'h3bbee105),
	.w2(32'h3b0a78aa),
	.w3(32'h3bf446e2),
	.w4(32'h3c238c81),
	.w5(32'hba92f38d),
	.w6(32'hba91a9ea),
	.w7(32'h3c2fdd74),
	.w8(32'h3b233b3f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe6e10),
	.w1(32'h3ba4b1c5),
	.w2(32'h3ada2235),
	.w3(32'hbc092719),
	.w4(32'h3bb27748),
	.w5(32'h3b7aa4d2),
	.w6(32'hbbc6bfc6),
	.w7(32'h3a95718f),
	.w8(32'h3bccefa1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb69c),
	.w1(32'hb90744e1),
	.w2(32'hb9bbd480),
	.w3(32'hbc1738d7),
	.w4(32'hbb9b4bb8),
	.w5(32'hbb912f29),
	.w6(32'hbbb190f9),
	.w7(32'hbb68bc67),
	.w8(32'hbad341ce),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63ec6),
	.w1(32'h3a5aa770),
	.w2(32'hba847c28),
	.w3(32'hbb7b9ef7),
	.w4(32'hbc0b6a25),
	.w5(32'hbb1312ea),
	.w6(32'hbc2190da),
	.w7(32'h3afe64be),
	.w8(32'h3af03958),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7ec05),
	.w1(32'h383728a4),
	.w2(32'hbab0c565),
	.w3(32'hbc2baddd),
	.w4(32'hbb967483),
	.w5(32'hbacb24b6),
	.w6(32'hbbf4a4a6),
	.w7(32'hbb5e41ee),
	.w8(32'hbbdca468),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab038de),
	.w1(32'h3a39c036),
	.w2(32'hbbc82bfa),
	.w3(32'h3af967be),
	.w4(32'h3a64f92d),
	.w5(32'hbc6c9430),
	.w6(32'h3b29823f),
	.w7(32'h3859df7e),
	.w8(32'hbbda27b7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b9a2),
	.w1(32'hbb01f4b8),
	.w2(32'h3bfd4fd3),
	.w3(32'h3b4a17f9),
	.w4(32'h3a5771f8),
	.w5(32'h3c8f2754),
	.w6(32'hbbb51d29),
	.w7(32'hbae37284),
	.w8(32'h3c87e95c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0681a7),
	.w1(32'hbcd77113),
	.w2(32'h3b19167d),
	.w3(32'hbbe25a00),
	.w4(32'hbd263ba1),
	.w5(32'h3b890500),
	.w6(32'h3be2737b),
	.w7(32'hbcd885ab),
	.w8(32'h3bc7c97e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d9bfb),
	.w1(32'h3aee3b2d),
	.w2(32'hbb452b6e),
	.w3(32'hbbd86b18),
	.w4(32'hba8851f5),
	.w5(32'h39907acf),
	.w6(32'hbb831d83),
	.w7(32'hbac33832),
	.w8(32'h3c6f4813),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20b3fe),
	.w1(32'hbc962c3a),
	.w2(32'hbb4f373a),
	.w3(32'hbbe2b895),
	.w4(32'hbc9b216c),
	.w5(32'hbba9ba52),
	.w6(32'h3c98c85d),
	.w7(32'h3a9ec613),
	.w8(32'hb9ab3d06),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac22a3e),
	.w1(32'h3b259fff),
	.w2(32'hbc57ee48),
	.w3(32'hbaf61954),
	.w4(32'h3afecbbc),
	.w5(32'hbc787e41),
	.w6(32'hbba1a853),
	.w7(32'h39d33fb6),
	.w8(32'hbc426dd3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21bbea),
	.w1(32'hbc00e628),
	.w2(32'h3c2bf96d),
	.w3(32'h3b233005),
	.w4(32'h3a27857a),
	.w5(32'h3c38dea4),
	.w6(32'hbc8046fc),
	.w7(32'h3b268498),
	.w8(32'h3c5d6b30),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45c2fb),
	.w1(32'hbc4260e2),
	.w2(32'h3b26e0fc),
	.w3(32'h3b5131ff),
	.w4(32'hbc7b7ed9),
	.w5(32'hbb274db3),
	.w6(32'h3c0f9c6f),
	.w7(32'hbc3e048b),
	.w8(32'hbb37e2b7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06ee7),
	.w1(32'hba293116),
	.w2(32'h3acefc79),
	.w3(32'hbbf6aebb),
	.w4(32'hbc386f76),
	.w5(32'h3adc964b),
	.w6(32'hbc18efb2),
	.w7(32'hbbc4e573),
	.w8(32'h3a698aa8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91326b),
	.w1(32'hbc0bfe32),
	.w2(32'h3a7151a1),
	.w3(32'hb8e7bacf),
	.w4(32'hbc260df3),
	.w5(32'h3b219067),
	.w6(32'h3b810844),
	.w7(32'hb8780b94),
	.w8(32'h3bcbfe52),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974f45),
	.w1(32'hbb765f74),
	.w2(32'hbbf43877),
	.w3(32'hbbd52c9b),
	.w4(32'hbbc440d1),
	.w5(32'hbbe8b3d4),
	.w6(32'hbabe0f40),
	.w7(32'hb9e842c7),
	.w8(32'hbb719977),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe93776),
	.w1(32'hba9661c1),
	.w2(32'hbaa62953),
	.w3(32'h3b5102c0),
	.w4(32'h39893a3d),
	.w5(32'hbc5fc39e),
	.w6(32'hbb598d2e),
	.w7(32'h3b7106bc),
	.w8(32'hbc50d066),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862b20),
	.w1(32'hbc9d809a),
	.w2(32'hb9b645eb),
	.w3(32'h3c05bd02),
	.w4(32'hbc0cde71),
	.w5(32'hbb1b3c41),
	.w6(32'hbba36442),
	.w7(32'hbb753dbf),
	.w8(32'hbb0b576c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6ccf),
	.w1(32'h3b5fb9bb),
	.w2(32'h3a8acc4c),
	.w3(32'hbb9077af),
	.w4(32'hb9391147),
	.w5(32'h3a53fd4a),
	.w6(32'hbb3ad6f7),
	.w7(32'hbb136928),
	.w8(32'h3ab83487),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2926),
	.w1(32'h3a960749),
	.w2(32'hbd065207),
	.w3(32'hba726abe),
	.w4(32'hb4d8f7a8),
	.w5(32'hbd326cab),
	.w6(32'hbab8e0d7),
	.w7(32'h3a741b42),
	.w8(32'hbcf62815),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689baf),
	.w1(32'h3bb88d31),
	.w2(32'h3c2615a1),
	.w3(32'hbb9c3025),
	.w4(32'h3c7c8ec7),
	.w5(32'h3b05dccb),
	.w6(32'h3c00b30a),
	.w7(32'h3c2471fe),
	.w8(32'hbbd5e559),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8962),
	.w1(32'h3ac875ef),
	.w2(32'hbb03d1bd),
	.w3(32'h3a874672),
	.w4(32'hba162aa3),
	.w5(32'hb9a6bbd8),
	.w6(32'h3bfc17ba),
	.w7(32'hbb232307),
	.w8(32'hbadd2ccb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8895ac),
	.w1(32'hbc11e245),
	.w2(32'h3b9225ac),
	.w3(32'hbb24a0cf),
	.w4(32'hbbe60e80),
	.w5(32'h3b2ee7a2),
	.w6(32'hbbabdfa5),
	.w7(32'hbbe300bd),
	.w8(32'hbba39888),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d5c86),
	.w1(32'h3bc06797),
	.w2(32'hbbcbecef),
	.w3(32'hbbcc1702),
	.w4(32'hbbb09faf),
	.w5(32'hbb40a050),
	.w6(32'hbc289c06),
	.w7(32'h392ff2b3),
	.w8(32'h39af4be8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9177d6),
	.w1(32'h3b6d33e7),
	.w2(32'hb7b1257d),
	.w3(32'h3c0ee69f),
	.w4(32'h3bd78b4a),
	.w5(32'h3b2610c0),
	.w6(32'hbb5a74dd),
	.w7(32'hbbd356e4),
	.w8(32'h3b276472),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39921c6f),
	.w1(32'hbbf04805),
	.w2(32'hbc1bdc2a),
	.w3(32'h3aadc287),
	.w4(32'hbbb77b6d),
	.w5(32'hbc22b610),
	.w6(32'h3b1cead6),
	.w7(32'hbb604489),
	.w8(32'hbbca821a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8962e9),
	.w1(32'hbc8304d6),
	.w2(32'hbae67b22),
	.w3(32'hbd0be2fd),
	.w4(32'hbc4eca62),
	.w5(32'hba0fb9da),
	.w6(32'hbd002547),
	.w7(32'h3aadc823),
	.w8(32'hbab2cfe7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a326e),
	.w1(32'hbadd0f55),
	.w2(32'h3aeecb47),
	.w3(32'h3aa48d78),
	.w4(32'hba4bbc8b),
	.w5(32'hbc655ae5),
	.w6(32'h3ab6fca0),
	.w7(32'hba42ccb6),
	.w8(32'hbc0004e4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c621ffd),
	.w1(32'h3be27e87),
	.w2(32'hbbc53d70),
	.w3(32'h3bf593f7),
	.w4(32'h3ae5463a),
	.w5(32'hbb80cd51),
	.w6(32'h3bc1696c),
	.w7(32'hbb2552f3),
	.w8(32'hbaed729c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9628a),
	.w1(32'hbbd0447b),
	.w2(32'h3be32b00),
	.w3(32'h3c069c19),
	.w4(32'hbbf3f7cb),
	.w5(32'h3bccb585),
	.w6(32'h3bbe6d0e),
	.w7(32'hbbc9f125),
	.w8(32'hbaf201c9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d833),
	.w1(32'hbb9d6090),
	.w2(32'h3a3f2919),
	.w3(32'h3c30e087),
	.w4(32'h3c7f6ebb),
	.w5(32'h3c17cc33),
	.w6(32'h3c7ba51b),
	.w7(32'h3b68281a),
	.w8(32'h3bd533f8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee02e),
	.w1(32'h3bc73fcc),
	.w2(32'h39f0cf43),
	.w3(32'hbb366f06),
	.w4(32'h3bfd5bea),
	.w5(32'h3a5f754a),
	.w6(32'h3bbb5912),
	.w7(32'h3ad1cfd2),
	.w8(32'hbb78ecdb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6870fe),
	.w1(32'h3a65a232),
	.w2(32'h3be4a763),
	.w3(32'hbbc85019),
	.w4(32'h3ad007f3),
	.w5(32'h391e185b),
	.w6(32'hbbe5fd4c),
	.w7(32'hbbab8023),
	.w8(32'hbb07398d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f616b),
	.w1(32'h389cb951),
	.w2(32'hbb613045),
	.w3(32'h3b4150cd),
	.w4(32'h3bd1326d),
	.w5(32'h3bf8af3b),
	.w6(32'hbb89ba2b),
	.w7(32'hbaa6938c),
	.w8(32'h3c0b5f53),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880d6d),
	.w1(32'hb981ff7a),
	.w2(32'hbb948603),
	.w3(32'hbb93f658),
	.w4(32'hbbd6ae15),
	.w5(32'hbbed81b8),
	.w6(32'h3b052b43),
	.w7(32'h39b43e57),
	.w8(32'hbba54dfd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84163b),
	.w1(32'hbbeebcbf),
	.w2(32'hb9c90083),
	.w3(32'hbb9d8134),
	.w4(32'hbc1111bd),
	.w5(32'h3b1eaace),
	.w6(32'hbb05a6c5),
	.w7(32'hbbdfca93),
	.w8(32'h3b9f3484),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28821),
	.w1(32'hbaeb9451),
	.w2(32'hbbed4dae),
	.w3(32'h3b808c7d),
	.w4(32'hbc4f0202),
	.w5(32'hbc189580),
	.w6(32'hba011c99),
	.w7(32'hbc3cccbb),
	.w8(32'hbb5583f1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb751eff),
	.w1(32'h39e4fa16),
	.w2(32'h3b48493b),
	.w3(32'hbc4a805e),
	.w4(32'hbb7e2a00),
	.w5(32'h3afe8d16),
	.w6(32'h3bce8bc6),
	.w7(32'hbb0c8838),
	.w8(32'hbc1014fd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35b21b),
	.w1(32'hbc226262),
	.w2(32'h3c93476f),
	.w3(32'hbc53194d),
	.w4(32'hbc78bb8f),
	.w5(32'h3cef6797),
	.w6(32'hbc4b06fe),
	.w7(32'hbbcd4ceb),
	.w8(32'h3c9bc2e0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea603e),
	.w1(32'hbcada622),
	.w2(32'hbb7fe3f6),
	.w3(32'h3bba55a7),
	.w4(32'hbcbe2568),
	.w5(32'hbc18c294),
	.w6(32'h3c038b16),
	.w7(32'hbc71192d),
	.w8(32'hbbf0e25a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f01a3),
	.w1(32'h39311cd4),
	.w2(32'hbbc1ba5e),
	.w3(32'hbb15a790),
	.w4(32'hbb588941),
	.w5(32'hbb491a17),
	.w6(32'hbb16f1a2),
	.w7(32'hbacc8db0),
	.w8(32'hbacb3682),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b8505),
	.w1(32'h39881f6e),
	.w2(32'hba973a76),
	.w3(32'hbca70d55),
	.w4(32'h3bc4def8),
	.w5(32'h3b851f6a),
	.w6(32'hbb933497),
	.w7(32'h3bfe81b6),
	.w8(32'h3a87742b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b5f44),
	.w1(32'hbb89ab61),
	.w2(32'h3c63febd),
	.w3(32'hbbcfa61b),
	.w4(32'hbc10d9fe),
	.w5(32'h3c99b12f),
	.w6(32'hbc53d0e1),
	.w7(32'h3b3b9a80),
	.w8(32'h3b545d81),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9274b),
	.w1(32'hbb8ec04d),
	.w2(32'h3c421e5e),
	.w3(32'hbb9faf0a),
	.w4(32'h3c0b39e0),
	.w5(32'h3bdb154a),
	.w6(32'h3a43148b),
	.w7(32'h3b9bf84a),
	.w8(32'h3a2507e1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaedfe),
	.w1(32'h3af95788),
	.w2(32'hbb158f6d),
	.w3(32'hbba72b79),
	.w4(32'h3bb0e852),
	.w5(32'h3b4c431b),
	.w6(32'hbbb75b02),
	.w7(32'h3afc0151),
	.w8(32'h3c0f8afe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1ce8d),
	.w1(32'hbbf476f5),
	.w2(32'h3b01d953),
	.w3(32'hbc09b673),
	.w4(32'hbb5196ec),
	.w5(32'hba8064dd),
	.w6(32'hbbb84b15),
	.w7(32'h3b338dd9),
	.w8(32'hbbf0a2b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42d3b1),
	.w1(32'h3a8e8091),
	.w2(32'h3b42fa3e),
	.w3(32'hbb4018d5),
	.w4(32'h3c1d7f5e),
	.w5(32'hba9f4997),
	.w6(32'hb9a3ba6f),
	.w7(32'hbbab4d6d),
	.w8(32'h3c2d285a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27553),
	.w1(32'h3bc76795),
	.w2(32'hbca58ea2),
	.w3(32'h3a834e17),
	.w4(32'h3aadeae5),
	.w5(32'hbd33c02a),
	.w6(32'h3bf15beb),
	.w7(32'h3c012e06),
	.w8(32'hbcfd96a9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc547bbb),
	.w1(32'h3b0a1b28),
	.w2(32'h3c102eaf),
	.w3(32'hbc9b0228),
	.w4(32'h3a0d21cb),
	.w5(32'h3bdfc920),
	.w6(32'hbc9a9a8f),
	.w7(32'h3b000ab8),
	.w8(32'h3c646802),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadef8eb),
	.w1(32'h3b74a137),
	.w2(32'h3ad7c7b4),
	.w3(32'h3b6e9f66),
	.w4(32'h3c2205d7),
	.w5(32'h3b112b3d),
	.w6(32'h3b34d9b3),
	.w7(32'h3b567020),
	.w8(32'hba036c4c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12f18b),
	.w1(32'hb9bf7d54),
	.w2(32'h3c28b793),
	.w3(32'h3b8525f6),
	.w4(32'hb968f1d4),
	.w5(32'hbac717fd),
	.w6(32'h3b0d4eba),
	.w7(32'hbb65a899),
	.w8(32'hbbeeaf3f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a66d7),
	.w1(32'h3bba2c85),
	.w2(32'hbb3ecb2c),
	.w3(32'hbbc59fad),
	.w4(32'h3c0fc0a1),
	.w5(32'hb99c5dd2),
	.w6(32'hbb89404d),
	.w7(32'hbc023800),
	.w8(32'h3b04f556),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a071e),
	.w1(32'h3b3d7bc8),
	.w2(32'h3c55d51c),
	.w3(32'h3c3d0031),
	.w4(32'h3c4fe7c0),
	.w5(32'h3cc85ba6),
	.w6(32'h3c65c198),
	.w7(32'h3c373f31),
	.w8(32'h3c598d71),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86a01a),
	.w1(32'hbad52283),
	.w2(32'hbb8c110f),
	.w3(32'h3b07caf7),
	.w4(32'hbc28215d),
	.w5(32'h3abaf458),
	.w6(32'hbb0e3e06),
	.w7(32'hbbc7d7cb),
	.w8(32'hbc0e80b9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c28af),
	.w1(32'h3a2cd63b),
	.w2(32'hb96e0590),
	.w3(32'hbc4c7d92),
	.w4(32'hb97c6975),
	.w5(32'hbbb4b43c),
	.w6(32'hbc09ef18),
	.w7(32'hbbae574b),
	.w8(32'hbb2b9be6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a89bd),
	.w1(32'hbbbabe8b),
	.w2(32'hba4ae66c),
	.w3(32'hbb88dcdf),
	.w4(32'hb972a9e0),
	.w5(32'h3a3fd96b),
	.w6(32'hbbe57744),
	.w7(32'hbb3a48de),
	.w8(32'h3b4f36f8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a682a3c),
	.w1(32'h393e0232),
	.w2(32'hbc04f771),
	.w3(32'hba4eeab6),
	.w4(32'h3b35b4d4),
	.w5(32'hbc2ea0a2),
	.w6(32'h3b0cea5b),
	.w7(32'hba17289a),
	.w8(32'hbbaf3f0d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39724b4d),
	.w1(32'h3b414d66),
	.w2(32'hbb896fbf),
	.w3(32'hbb335073),
	.w4(32'h3a8de0e8),
	.w5(32'hbb9c6788),
	.w6(32'hbbc41a4f),
	.w7(32'hbbc82d7d),
	.w8(32'hbba48525),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e77a7),
	.w1(32'hbbc13e15),
	.w2(32'h3a65876b),
	.w3(32'h3a7bf5f4),
	.w4(32'hbbd467c0),
	.w5(32'hba823cf4),
	.w6(32'hba9b5775),
	.w7(32'hbbd14930),
	.w8(32'h3adac0a7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f83de),
	.w1(32'hbbc90e8a),
	.w2(32'hba5a7296),
	.w3(32'hbbd8b08a),
	.w4(32'hbbc73e10),
	.w5(32'hbb8901ad),
	.w6(32'hbc58feb3),
	.w7(32'hbb2a9a4f),
	.w8(32'hbc0eb82f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b9dde),
	.w1(32'hbb6aacb4),
	.w2(32'h3a33de4e),
	.w3(32'hbae0e024),
	.w4(32'h3ae4c1c2),
	.w5(32'hbaff98f7),
	.w6(32'hbb8e254c),
	.w7(32'hbba136f1),
	.w8(32'hba977a31),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc005df),
	.w1(32'h39f958f6),
	.w2(32'hb9d1a1c3),
	.w3(32'hbc1b15db),
	.w4(32'hbb063bb4),
	.w5(32'h3b96d3a0),
	.w6(32'hbbedd83f),
	.w7(32'hba95384b),
	.w8(32'hbb71069e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed012e),
	.w1(32'h3bd3ba8b),
	.w2(32'hbbec4f9d),
	.w3(32'hbc8487dd),
	.w4(32'h3ba33bac),
	.w5(32'hbc5fafd1),
	.w6(32'hbbd8d148),
	.w7(32'h3b4b5369),
	.w8(32'hbbf451bc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be100cd),
	.w1(32'h3c520a89),
	.w2(32'hbadf28b0),
	.w3(32'h3b3af1ef),
	.w4(32'h3c64dc28),
	.w5(32'h3c0d6e30),
	.w6(32'h3b6da960),
	.w7(32'h3c05e4ab),
	.w8(32'h3c09ad50),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90799),
	.w1(32'hbb2e8d05),
	.w2(32'hbc5b3c7b),
	.w3(32'hbbbb2bd8),
	.w4(32'hba73d0f2),
	.w5(32'hbc307480),
	.w6(32'hbba34a72),
	.w7(32'hbba141a7),
	.w8(32'h3a77653e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0e70),
	.w1(32'h3b2ee779),
	.w2(32'h3ac1e70b),
	.w3(32'h39a3d238),
	.w4(32'h3af41a49),
	.w5(32'hba2aa6a3),
	.w6(32'h39a045fa),
	.w7(32'hbb64bd3d),
	.w8(32'hba69d80d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5121),
	.w1(32'hbbf99f94),
	.w2(32'h3c1f0254),
	.w3(32'hbb9b3ed8),
	.w4(32'hbc24a140),
	.w5(32'h3c1ef3a3),
	.w6(32'hbb92e522),
	.w7(32'hbc03b10c),
	.w8(32'h3c3aac69),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926102),
	.w1(32'hbbbbc6f7),
	.w2(32'h3c7329c1),
	.w3(32'hbbf62a69),
	.w4(32'hbbea550f),
	.w5(32'h3c2d315c),
	.w6(32'h3ad08f24),
	.w7(32'hb9efdc35),
	.w8(32'h3b5f9803),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c3de4),
	.w1(32'h3bb688c2),
	.w2(32'h3be445ce),
	.w3(32'h3c0d8ee9),
	.w4(32'h3b50aab0),
	.w5(32'h3a2e5ed3),
	.w6(32'h3b9db629),
	.w7(32'h3a9aafa9),
	.w8(32'hbc16ec83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39886d54),
	.w1(32'hbb1a2971),
	.w2(32'hbca8a755),
	.w3(32'hbbc93d7d),
	.w4(32'h3ae1ad73),
	.w5(32'hbce3e513),
	.w6(32'hbb60c1d0),
	.w7(32'h3bb5e789),
	.w8(32'hbc8d2b47),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce5568),
	.w1(32'hbaddb02c),
	.w2(32'h3a77f67d),
	.w3(32'hbd3cdd13),
	.w4(32'hbb6f981c),
	.w5(32'h3b946a6e),
	.w6(32'hbd1c5075),
	.w7(32'hbc6946e7),
	.w8(32'h385ebb79),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969c3f8),
	.w1(32'h3afc37b0),
	.w2(32'h3b392b82),
	.w3(32'hba914e6f),
	.w4(32'h3acf011d),
	.w5(32'h3b7abfaa),
	.w6(32'hba1a1bf3),
	.w7(32'h3b2277e2),
	.w8(32'hba914966),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96caad),
	.w1(32'hbb7c8096),
	.w2(32'hbb384b51),
	.w3(32'hbc033c24),
	.w4(32'hbc1505ae),
	.w5(32'h3a53eed1),
	.w6(32'hbb699a45),
	.w7(32'hb9abfcd0),
	.w8(32'hb9dbc4f1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cf43c),
	.w1(32'hbb8cf298),
	.w2(32'h3b6abcec),
	.w3(32'h3abb9f93),
	.w4(32'hb9928b84),
	.w5(32'h3a9c0829),
	.w6(32'hbae7974d),
	.w7(32'hba6443d0),
	.w8(32'h3b782a05),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb576f),
	.w1(32'hbc257d06),
	.w2(32'h3cf2e066),
	.w3(32'hbc26add8),
	.w4(32'hbb0df2b1),
	.w5(32'h3d28decf),
	.w6(32'hbb8c9f17),
	.w7(32'hbb8e93d8),
	.w8(32'h3cc58ffe),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25faac),
	.w1(32'hbc69ef4f),
	.w2(32'h3b70a0e7),
	.w3(32'h3d01f168),
	.w4(32'hbc5dbbc0),
	.w5(32'h3b3bbf75),
	.w6(32'h3d06125c),
	.w7(32'hbb87099e),
	.w8(32'h3aef5749),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc242f1f),
	.w1(32'hbb639fec),
	.w2(32'hbcb11696),
	.w3(32'hbc22b8eb),
	.w4(32'hbb7435dd),
	.w5(32'hbd2ea02c),
	.w6(32'hbab39a93),
	.w7(32'hba96af8d),
	.w8(32'hbd1367b4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca32171),
	.w1(32'hba436349),
	.w2(32'hbc7e71e2),
	.w3(32'hbc1c5c63),
	.w4(32'h3c39534f),
	.w5(32'hbca45106),
	.w6(32'h3acccab6),
	.w7(32'hbb4033a7),
	.w8(32'hbc9963ea),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa73730),
	.w1(32'hba0d4d98),
	.w2(32'h39d0ea9d),
	.w3(32'hbae06c7b),
	.w4(32'h3b988ba7),
	.w5(32'h3b6199ff),
	.w6(32'hbb19a1c6),
	.w7(32'hbaa19048),
	.w8(32'h3af7c8cf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a3dca),
	.w1(32'hb9aafa28),
	.w2(32'hbabe4513),
	.w3(32'hbac918d6),
	.w4(32'h3a7dc06c),
	.w5(32'h3c804b17),
	.w6(32'hba4561a7),
	.w7(32'h3ac57eda),
	.w8(32'h39dcc719),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b0d7),
	.w1(32'hbb815bd2),
	.w2(32'h3bc00fdd),
	.w3(32'h3afded68),
	.w4(32'hbb9f0463),
	.w5(32'h3b5641b3),
	.w6(32'hbbebd628),
	.w7(32'hbb2bd744),
	.w8(32'h36992617),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187a31),
	.w1(32'hbc847c8e),
	.w2(32'h3bdcaac5),
	.w3(32'hbb5b9dc7),
	.w4(32'hba218db3),
	.w5(32'h3992d11f),
	.w6(32'h3c60f8f5),
	.w7(32'h3c1ebfa8),
	.w8(32'h3bde8e43),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73f4c0),
	.w1(32'h3c0e0278),
	.w2(32'hb91fd808),
	.w3(32'hbae5cc80),
	.w4(32'hbbc55fb7),
	.w5(32'hba485267),
	.w6(32'hbc3346b4),
	.w7(32'hbc06c914),
	.w8(32'h3b81c126),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27a347),
	.w1(32'h3c90a3cb),
	.w2(32'h3ba6317a),
	.w3(32'h3bfdfcc6),
	.w4(32'h3ca69484),
	.w5(32'h3bba6ed7),
	.w6(32'h3c0aa0d3),
	.w7(32'h3c8b970d),
	.w8(32'h3bfe1961),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4d671),
	.w1(32'h3bbe04b5),
	.w2(32'hbb9d494e),
	.w3(32'h3b9ff4e4),
	.w4(32'h3bf0d5fa),
	.w5(32'hbb6a5a3a),
	.w6(32'h3bc78a00),
	.w7(32'h3bde1616),
	.w8(32'hbb008926),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0d5ce),
	.w1(32'hbb384e14),
	.w2(32'h3a909e6a),
	.w3(32'hbbd5e4a9),
	.w4(32'hb9a45037),
	.w5(32'h3bf0649d),
	.w6(32'hbb8e070b),
	.w7(32'hbaea4d7c),
	.w8(32'h3a72538f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188c8b),
	.w1(32'h3b837083),
	.w2(32'hbc60b337),
	.w3(32'hbb392937),
	.w4(32'h3aa7601d),
	.w5(32'hb85fc68c),
	.w6(32'hbb1f627c),
	.w7(32'h39ede5c9),
	.w8(32'h3c2f1cb5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd58e43),
	.w1(32'hbad3e166),
	.w2(32'h3bf8c823),
	.w3(32'h3af1c34a),
	.w4(32'hbab4665f),
	.w5(32'hb92d65dd),
	.w6(32'hbb2747e0),
	.w7(32'hbbd0a699),
	.w8(32'h3aee979c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a305a),
	.w1(32'h3bcb2279),
	.w2(32'h3c134f25),
	.w3(32'hbc36c528),
	.w4(32'h3a163176),
	.w5(32'h3c407fce),
	.w6(32'hbaf9f54f),
	.w7(32'h3bca1eae),
	.w8(32'h3ba2f15c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0080c6),
	.w1(32'h3b8f83d5),
	.w2(32'h3b4f86bd),
	.w3(32'hbc0e6fe6),
	.w4(32'hbb9ebdb7),
	.w5(32'hbb4e9520),
	.w6(32'hba765463),
	.w7(32'hbbcb43c2),
	.w8(32'hb6f536a6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc056f84),
	.w1(32'hbc662a5f),
	.w2(32'hb9c039e3),
	.w3(32'hbc948e53),
	.w4(32'hbc7dad49),
	.w5(32'h3c0aabd0),
	.w6(32'hbc836380),
	.w7(32'hbaa7d0e7),
	.w8(32'h3bb8889f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7e0c3),
	.w1(32'hbbf1a390),
	.w2(32'h39c2f1ee),
	.w3(32'h3b8e4138),
	.w4(32'hbc3a15de),
	.w5(32'h3c2afa2c),
	.w6(32'h3c26907d),
	.w7(32'hbb4891bd),
	.w8(32'hb9f7802b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb45f5),
	.w1(32'hbb0977a0),
	.w2(32'h3835f1f5),
	.w3(32'h3a921f86),
	.w4(32'hbae8ff13),
	.w5(32'h3a40f644),
	.w6(32'h3bebdc14),
	.w7(32'h3c0ab6b9),
	.w8(32'h3c178821),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324f55),
	.w1(32'hbaba5c6c),
	.w2(32'hbc456364),
	.w3(32'h39f0cdab),
	.w4(32'hbba36332),
	.w5(32'hbc898499),
	.w6(32'h3b4e1af5),
	.w7(32'hba58effb),
	.w8(32'hbc62d5f5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239527),
	.w1(32'hbbbe7457),
	.w2(32'h3b1928e5),
	.w3(32'h3aa2f97a),
	.w4(32'h3c101182),
	.w5(32'h3bd09566),
	.w6(32'h3be6de4d),
	.w7(32'h3c157c8e),
	.w8(32'h3b0d4595),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df540),
	.w1(32'hbb4b07cb),
	.w2(32'hbc8ef780),
	.w3(32'hbb687424),
	.w4(32'h3729b2cd),
	.w5(32'hbcce91fa),
	.w6(32'h3acd768b),
	.w7(32'h3b63c9a9),
	.w8(32'hbc82aed4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5914),
	.w1(32'hb988e69e),
	.w2(32'hbba66080),
	.w3(32'hbbc7a558),
	.w4(32'h3aa295d4),
	.w5(32'hbcabb4b1),
	.w6(32'hbb8cfd75),
	.w7(32'hba84cf89),
	.w8(32'hbc28a51a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc86fbc),
	.w1(32'h3bb8b11e),
	.w2(32'hbc32f0c1),
	.w3(32'hbbeaca80),
	.w4(32'h3c84ba2e),
	.w5(32'hbc969c78),
	.w6(32'h3b3afc99),
	.w7(32'h3c6bca3a),
	.w8(32'hbc725b34),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb5c84),
	.w1(32'h3b8f1fb7),
	.w2(32'hbb45c19e),
	.w3(32'hbc36fb65),
	.w4(32'h3bc674ac),
	.w5(32'h3bc94c46),
	.w6(32'hbbd87ac8),
	.w7(32'h3b123f64),
	.w8(32'h3b086ef9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc019ce9),
	.w1(32'hbb12cf46),
	.w2(32'hbae801fe),
	.w3(32'hbc2b6b0d),
	.w4(32'hbbdd4e59),
	.w5(32'h3bb5b108),
	.w6(32'h3b967a21),
	.w7(32'h3aeb6149),
	.w8(32'h3b5104f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf249ee),
	.w1(32'hbb28e128),
	.w2(32'h3a306634),
	.w3(32'hbb6df16e),
	.w4(32'hbbbd90c7),
	.w5(32'hba0a2cd1),
	.w6(32'hbb9a4370),
	.w7(32'hbb7a8257),
	.w8(32'h3a95b280),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff8dc4),
	.w1(32'hbabd41fe),
	.w2(32'h3bb7d335),
	.w3(32'hbc243e24),
	.w4(32'hbbf1fcde),
	.w5(32'h3c5d8296),
	.w6(32'hbb3c580c),
	.w7(32'h3be6caef),
	.w8(32'h3bbf48c8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7da3),
	.w1(32'hb9361649),
	.w2(32'h38f5196a),
	.w3(32'h3b4acf28),
	.w4(32'hb8d5b896),
	.w5(32'hbbe30ee4),
	.w6(32'h3c006e16),
	.w7(32'hba6735d4),
	.w8(32'hba1f96cd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91bff0),
	.w1(32'hbbb142fc),
	.w2(32'h3c4fce1a),
	.w3(32'hbcc191ec),
	.w4(32'hba59045b),
	.w5(32'h3d00db14),
	.w6(32'hbc908bcb),
	.w7(32'hbb25d928),
	.w8(32'h3d11df15),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03a065),
	.w1(32'h3b83de18),
	.w2(32'hba56cfad),
	.w3(32'h3d3099bf),
	.w4(32'hbc445afc),
	.w5(32'h3ac98182),
	.w6(32'h3c8608ea),
	.w7(32'hbc878519),
	.w8(32'h3aef04a0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3969b8),
	.w1(32'hbb486e65),
	.w2(32'h3ba340a5),
	.w3(32'hbcb44f0c),
	.w4(32'hbc80cc9f),
	.w5(32'h3b31a79a),
	.w6(32'hbc4cbb6d),
	.w7(32'hbbe05984),
	.w8(32'h3ac3bf7c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3a6e),
	.w1(32'hbbabb992),
	.w2(32'h3bc34c9b),
	.w3(32'h3896ec24),
	.w4(32'hbbac2070),
	.w5(32'h3bc1859a),
	.w6(32'hbb2af861),
	.w7(32'h3bf2f2ce),
	.w8(32'h3b11cd26),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39957e6a),
	.w1(32'h3a982120),
	.w2(32'hbba68b10),
	.w3(32'h3b9e2d2e),
	.w4(32'h3bb58033),
	.w5(32'h3a969beb),
	.w6(32'h3be41069),
	.w7(32'h3ba095e2),
	.w8(32'h3b8a42c5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2463),
	.w1(32'hbbbf10dc),
	.w2(32'hb956c9bb),
	.w3(32'hbc4c9dd4),
	.w4(32'hbb719c0b),
	.w5(32'hbafab4f8),
	.w6(32'hbbcb5857),
	.w7(32'h3b8243ab),
	.w8(32'hbb0a4940),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb111786),
	.w1(32'hbb45601f),
	.w2(32'hba9241da),
	.w3(32'h3b0cad84),
	.w4(32'h3bad919d),
	.w5(32'h3c47aaf2),
	.w6(32'h3b7465de),
	.w7(32'hbb278d91),
	.w8(32'h3bba7ccd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8065de),
	.w1(32'h39aedcb8),
	.w2(32'h3b965a8e),
	.w3(32'hbc07f959),
	.w4(32'hbc01cc4e),
	.w5(32'h3c120714),
	.w6(32'h39cc0ee6),
	.w7(32'h3b375962),
	.w8(32'h3a17a2cb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2649e4),
	.w1(32'hbb178a06),
	.w2(32'hba2069f2),
	.w3(32'h3b834495),
	.w4(32'hbb0d90f5),
	.w5(32'h3bb64469),
	.w6(32'h3bd85de4),
	.w7(32'hba0f1d89),
	.w8(32'hbb77b3c5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39835fab),
	.w1(32'hbadb5a22),
	.w2(32'hba815e1d),
	.w3(32'h3b08a9f1),
	.w4(32'hbb91b406),
	.w5(32'hbaa591e3),
	.w6(32'h3b0f1483),
	.w7(32'hbbf42e48),
	.w8(32'h3a12e332),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcf4aa),
	.w1(32'hbb141f03),
	.w2(32'h3c01c1e0),
	.w3(32'hbaa05bc9),
	.w4(32'hbb2e76a7),
	.w5(32'h3c351ec7),
	.w6(32'hba594d03),
	.w7(32'hbb3d8b3d),
	.w8(32'h3be5ebdb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29fa18),
	.w1(32'hbb643d53),
	.w2(32'h3c553c65),
	.w3(32'hbb091e46),
	.w4(32'hbbade053),
	.w5(32'h3c32fd35),
	.w6(32'hbb4d14c5),
	.w7(32'hbb5e5de8),
	.w8(32'h3cfcbfdd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55ceac),
	.w1(32'hbb6d21ee),
	.w2(32'hbc0a4aa2),
	.w3(32'h3c3a3154),
	.w4(32'hbc68e3fb),
	.w5(32'hbc808670),
	.w6(32'h3b374590),
	.w7(32'hbc8266ba),
	.w8(32'hbc519d70),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7402),
	.w1(32'hb936e1b0),
	.w2(32'h3cb99dbf),
	.w3(32'hbb7a5285),
	.w4(32'h3b9f74b4),
	.w5(32'h3d234b13),
	.w6(32'hb9836276),
	.w7(32'h3b39aacd),
	.w8(32'h3cc7dd7a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5744eb),
	.w1(32'hbc2d4dde),
	.w2(32'h3bccbc10),
	.w3(32'hbbb157be),
	.w4(32'hbc7007dc),
	.w5(32'h3cd89fda),
	.w6(32'hbc81fae7),
	.w7(32'hbc20928b),
	.w8(32'h3c8baf4d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e1aa),
	.w1(32'hb9eda70d),
	.w2(32'hbbc811f2),
	.w3(32'h3c1f352c),
	.w4(32'hbc0f8afc),
	.w5(32'h3c281581),
	.w6(32'hbb62965b),
	.w7(32'h3ad7a1a1),
	.w8(32'hbad8f67b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba138072),
	.w1(32'hbb9493bf),
	.w2(32'hbc7e6de4),
	.w3(32'hbc7ae382),
	.w4(32'hba6620b8),
	.w5(32'hbc9b2b9b),
	.w6(32'hbc2b067e),
	.w7(32'hba0d0c4a),
	.w8(32'hbb820835),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68859),
	.w1(32'h3a7f058b),
	.w2(32'h3b81ca03),
	.w3(32'h3ba3057d),
	.w4(32'h3b83ce55),
	.w5(32'hbbb6e3d3),
	.w6(32'h3bd65fd4),
	.w7(32'h3be9c0b3),
	.w8(32'hbb8d197f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd97377),
	.w1(32'hbb662416),
	.w2(32'hbc7ab250),
	.w3(32'hbc44ed47),
	.w4(32'h3ad39102),
	.w5(32'hbcbc889a),
	.w6(32'hbbbdf560),
	.w7(32'hbb3afa47),
	.w8(32'h39574202),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874907),
	.w1(32'hbaa63f95),
	.w2(32'hbae0220e),
	.w3(32'h3cde73c0),
	.w4(32'hbb13b7bb),
	.w5(32'h3c1ce5c6),
	.w6(32'h3ca0745b),
	.w7(32'hbc2aba46),
	.w8(32'h3b88c125),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4353e4),
	.w1(32'hba8f2cbe),
	.w2(32'hbbcbcb62),
	.w3(32'hbb247092),
	.w4(32'h3a12d309),
	.w5(32'hbc829d8e),
	.w6(32'hbb104648),
	.w7(32'h396190a0),
	.w8(32'hbc586c2c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8eb7e9),
	.w1(32'hbb534f6b),
	.w2(32'h3bbdff2f),
	.w3(32'hbb91bc56),
	.w4(32'h3b9e042c),
	.w5(32'h3c7ea161),
	.w6(32'h3c19c2d4),
	.w7(32'h39c4a6bd),
	.w8(32'h3bede95a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac85bb6),
	.w1(32'hbc1afaa4),
	.w2(32'h3b98a078),
	.w3(32'hbc2b444a),
	.w4(32'hbc5ca74a),
	.w5(32'h3bbb722f),
	.w6(32'h3bdbbf2d),
	.w7(32'hbc7629b6),
	.w8(32'h3bb4c3fa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab743a2),
	.w1(32'h3a5f6faa),
	.w2(32'hbba8700e),
	.w3(32'h3b08a149),
	.w4(32'hbaae2319),
	.w5(32'hbb6dea9f),
	.w6(32'h3b602f29),
	.w7(32'h392bcd60),
	.w8(32'hbc15585d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44bd90),
	.w1(32'hbbd1c578),
	.w2(32'hbc353d87),
	.w3(32'hbc237569),
	.w4(32'h3adbda33),
	.w5(32'hbc840fee),
	.w6(32'h3b5b22be),
	.w7(32'h399ebafa),
	.w8(32'hbc39d85b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89587d),
	.w1(32'h3c51b0a1),
	.w2(32'hbbe2f3e4),
	.w3(32'hbbc62076),
	.w4(32'h3c178ec5),
	.w5(32'hbbe8a6b7),
	.w6(32'hbbf8109c),
	.w7(32'h39fdfcb8),
	.w8(32'hbbb30aee),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c3ba9),
	.w1(32'h398ecf72),
	.w2(32'h3a0016d0),
	.w3(32'hbb783b8a),
	.w4(32'h3bb591e2),
	.w5(32'h3b6ff5c8),
	.w6(32'hbac15e2a),
	.w7(32'h3b3ea747),
	.w8(32'h3a90152e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6466),
	.w1(32'hbb5f3e26),
	.w2(32'hb6c4f306),
	.w3(32'hba1fa246),
	.w4(32'hba9c1951),
	.w5(32'h3acbc07f),
	.w6(32'hbac999cb),
	.w7(32'hbb2e4d9f),
	.w8(32'h3a97b71e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0086d5),
	.w1(32'hbba0aab4),
	.w2(32'hbb5996cf),
	.w3(32'h3bc38a5f),
	.w4(32'hbb8a00f3),
	.w5(32'hbae5ac99),
	.w6(32'h394473ab),
	.w7(32'h3b2effb9),
	.w8(32'h3984b8c7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8449e7),
	.w1(32'hbb0e4f3e),
	.w2(32'hbaa71efe),
	.w3(32'hbbc8b5a8),
	.w4(32'hbb9b8791),
	.w5(32'hbaa29ea1),
	.w6(32'hbb7f40e5),
	.w7(32'hbb77ba50),
	.w8(32'hbb51a844),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76edb2),
	.w1(32'h3b2c98ec),
	.w2(32'h3b138013),
	.w3(32'h3b94a605),
	.w4(32'h3b63eecd),
	.w5(32'h3c3033c9),
	.w6(32'h3b85dbd2),
	.w7(32'h3bc4d831),
	.w8(32'h3bb4b2e2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c6f6),
	.w1(32'hbb8c74eb),
	.w2(32'h3b8a6460),
	.w3(32'hbba936d3),
	.w4(32'hbc006e78),
	.w5(32'h3aa898f8),
	.w6(32'hbc021b49),
	.w7(32'hbbd45f3f),
	.w8(32'h3b66ea0e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ffab4),
	.w1(32'h3ac18b79),
	.w2(32'h3a6f5ea4),
	.w3(32'h3b10e406),
	.w4(32'h3b681bf6),
	.w5(32'h3b545ef9),
	.w6(32'h3c083280),
	.w7(32'h3b593539),
	.w8(32'h3ae77177),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f7e7d),
	.w1(32'h3ac4085f),
	.w2(32'h3c1c61df),
	.w3(32'h39f09ae5),
	.w4(32'h3b8802ec),
	.w5(32'h3bdb380e),
	.w6(32'h3a0c8c06),
	.w7(32'h3b7de06e),
	.w8(32'h3ba21bad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba905a3d),
	.w1(32'hbb47f397),
	.w2(32'h3b27aeb0),
	.w3(32'hbb962ac8),
	.w4(32'hbb4d5368),
	.w5(32'h3ac5b7af),
	.w6(32'hbb808c12),
	.w7(32'hba95e1aa),
	.w8(32'h3b0f381e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d5d2f),
	.w1(32'h397f8f1a),
	.w2(32'hbc235691),
	.w3(32'h3b4a3fbc),
	.w4(32'hb9b5dc01),
	.w5(32'hbad1a08d),
	.w6(32'h3baee41d),
	.w7(32'h3b5aa2f1),
	.w8(32'h3a880214),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b580698),
	.w1(32'h3be13ec6),
	.w2(32'h3c6cd6a5),
	.w3(32'hbbc80998),
	.w4(32'h3ba5d05c),
	.w5(32'h3c4569e1),
	.w6(32'hbc212bbe),
	.w7(32'hbc3bdd11),
	.w8(32'h3b92d48c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed1b56),
	.w1(32'h3b443c6a),
	.w2(32'hbb9eacf3),
	.w3(32'hba2742aa),
	.w4(32'hbb81eee8),
	.w5(32'h3ad98bae),
	.w6(32'hbb957111),
	.w7(32'hbb87397c),
	.w8(32'hb9a6d4ba),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8926ac),
	.w1(32'h3bc26c13),
	.w2(32'h3c3cf028),
	.w3(32'hbc237a31),
	.w4(32'h3ae5c6a9),
	.w5(32'h3bb15e41),
	.w6(32'h3980d07d),
	.w7(32'hbae5db6d),
	.w8(32'h3b8df3be),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9168e0),
	.w1(32'hbb0fa4c9),
	.w2(32'h3a8e1bac),
	.w3(32'h3b777b96),
	.w4(32'h3b3f91cf),
	.w5(32'h3b0fb90b),
	.w6(32'h3c58f3a3),
	.w7(32'h3b8c9aeb),
	.w8(32'h3b01c1ed),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f05d2),
	.w1(32'hbb157c1a),
	.w2(32'h3ae8c343),
	.w3(32'hbaf5e0be),
	.w4(32'hba892011),
	.w5(32'hba8844c8),
	.w6(32'hba7a327e),
	.w7(32'hbb28d075),
	.w8(32'hb9a26ea9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a726446),
	.w1(32'h3ba6c317),
	.w2(32'h3b93eed4),
	.w3(32'hbbda603d),
	.w4(32'hbaf32d3a),
	.w5(32'hbc1fdcc4),
	.w6(32'h3b3aef63),
	.w7(32'h3c266903),
	.w8(32'h3b17d335),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecd5eb),
	.w1(32'h396ac1f2),
	.w2(32'h3c13a3f5),
	.w3(32'hbb152b19),
	.w4(32'hbb13ecc2),
	.w5(32'h3c780fd3),
	.w6(32'h3b859e76),
	.w7(32'hba9e5c83),
	.w8(32'h3bf51189),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0da0c8),
	.w1(32'h3bd0ebec),
	.w2(32'h3a72ad08),
	.w3(32'h3c451dfc),
	.w4(32'h3a90cd68),
	.w5(32'hb9a1ad32),
	.w6(32'h3b3771f6),
	.w7(32'h3b1d13fb),
	.w8(32'hba84a409),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b146c),
	.w1(32'h3acc0035),
	.w2(32'h3bdef935),
	.w3(32'hbbb8ca91),
	.w4(32'h3a34d9f4),
	.w5(32'h3bfb53cc),
	.w6(32'hbbf4ddb8),
	.w7(32'hb9a4c448),
	.w8(32'h3c4d82ad),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e0fc),
	.w1(32'h3c0a458e),
	.w2(32'hbb1b11ed),
	.w3(32'hbba3d01d),
	.w4(32'h39c4a202),
	.w5(32'hbb41dc61),
	.w6(32'h3bc08be9),
	.w7(32'h3b3e31a4),
	.w8(32'h3ba74de3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b987),
	.w1(32'hbabc540b),
	.w2(32'h3a09f8b5),
	.w3(32'hbb0262e0),
	.w4(32'hbb0db1a6),
	.w5(32'h3ac4c326),
	.w6(32'hbc22bc87),
	.w7(32'hbb4575fc),
	.w8(32'h3b5b5687),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9509b),
	.w1(32'hba308587),
	.w2(32'hbc5b5358),
	.w3(32'hbbbc93c8),
	.w4(32'h3ace8587),
	.w5(32'hbb42dfcd),
	.w6(32'hbbdbf5c2),
	.w7(32'h3aac307d),
	.w8(32'hbb961cd6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40faeb),
	.w1(32'hbc322dea),
	.w2(32'hbb9f6c53),
	.w3(32'hbc232b1a),
	.w4(32'hbc1d0a31),
	.w5(32'hbc7b85bc),
	.w6(32'hbc24f4a2),
	.w7(32'hbb47cb78),
	.w8(32'hbc268430),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb227),
	.w1(32'h3ba07d99),
	.w2(32'h3c2efb68),
	.w3(32'hbc88f0a5),
	.w4(32'hbc38afb3),
	.w5(32'h3bc4f1d9),
	.w6(32'hbc9496a9),
	.w7(32'hbc00729e),
	.w8(32'hbbffa25d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80c474),
	.w1(32'h3cb21678),
	.w2(32'hbb5445f5),
	.w3(32'h3bd29950),
	.w4(32'h3c74bd3b),
	.w5(32'h3c1e11ff),
	.w6(32'hbc849708),
	.w7(32'hbb106ae9),
	.w8(32'h3c11a38b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dd665),
	.w1(32'h3c726c28),
	.w2(32'hbabd34a0),
	.w3(32'h3c816256),
	.w4(32'h3bf11e70),
	.w5(32'hbb40a5d5),
	.w6(32'h3b8fc7a2),
	.w7(32'hb96d2e37),
	.w8(32'hbc13d597),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd34e1a),
	.w1(32'h3aeda41f),
	.w2(32'h3b459b5e),
	.w3(32'h3b7dd82e),
	.w4(32'hbaf37892),
	.w5(32'h3af7fcf9),
	.w6(32'hbba7333f),
	.w7(32'hbbd2416f),
	.w8(32'h3b6485fb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a593d2c),
	.w1(32'hbbcc7e4a),
	.w2(32'h3bc2b012),
	.w3(32'h3b66f340),
	.w4(32'h3917b93e),
	.w5(32'h3ab8d6ce),
	.w6(32'h3b81412f),
	.w7(32'h3c0c117a),
	.w8(32'hbca5b819),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8661ef),
	.w1(32'h3c98a233),
	.w2(32'hbc230c5f),
	.w3(32'h3ac1af0c),
	.w4(32'h3c73f8ac),
	.w5(32'h3bb1d6e3),
	.w6(32'hbd003701),
	.w7(32'hbc4b229a),
	.w8(32'h3c23098d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d0770),
	.w1(32'hbc642131),
	.w2(32'h3c1daab9),
	.w3(32'h3a0dd1a7),
	.w4(32'h3a15c602),
	.w5(32'h3c6383b0),
	.w6(32'h3bef1b19),
	.w7(32'h3bc43833),
	.w8(32'h3ac80a60),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8222dd),
	.w1(32'hbc6d377d),
	.w2(32'h393b584c),
	.w3(32'h3c791d57),
	.w4(32'h3bbd0c18),
	.w5(32'hbabd96e2),
	.w6(32'h3bb93ebf),
	.w7(32'h3b671b0c),
	.w8(32'hba3d1b88),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a85ab),
	.w1(32'hbc19997b),
	.w2(32'hbb6f63ba),
	.w3(32'hbbba8d4b),
	.w4(32'hbbe02a4f),
	.w5(32'hbb9fa3eb),
	.w6(32'h3b51ebce),
	.w7(32'h3b1a110e),
	.w8(32'hbc3b92b1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdb3f3),
	.w1(32'h3c197a1c),
	.w2(32'hbab7a193),
	.w3(32'hbb9afbd8),
	.w4(32'hbbd0337c),
	.w5(32'h3b9db6c2),
	.w6(32'hbc4fbe2c),
	.w7(32'hbc3cc558),
	.w8(32'h3ad2de37),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c250),
	.w1(32'hbc1192e9),
	.w2(32'h3b83b80d),
	.w3(32'hba2478d7),
	.w4(32'h3aa7ccce),
	.w5(32'h3b8647aa),
	.w6(32'hbac09a6b),
	.w7(32'hbaa13df8),
	.w8(32'hbc127705),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71751c),
	.w1(32'h3c188fab),
	.w2(32'h3aa0b723),
	.w3(32'h3c21fa67),
	.w4(32'h3bfdb287),
	.w5(32'h3aab2a09),
	.w6(32'hbb8475c8),
	.w7(32'hbb899a51),
	.w8(32'h3b6f0ba2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f95cb),
	.w1(32'hb9cd21d2),
	.w2(32'hbab78486),
	.w3(32'h3bb5184e),
	.w4(32'h3c2eaf9a),
	.w5(32'hbbafdda0),
	.w6(32'h3b9fd2a4),
	.w7(32'hb99f9a7c),
	.w8(32'hbbf6b151),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f294),
	.w1(32'hbb791e30),
	.w2(32'hbb192bd8),
	.w3(32'hbbfb0194),
	.w4(32'hbba87e2e),
	.w5(32'h3c23a5fc),
	.w6(32'hbb1faa3e),
	.w7(32'h3a91d25f),
	.w8(32'h3c572123),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5b56e),
	.w1(32'hbb4823bc),
	.w2(32'hbb132ad3),
	.w3(32'h3b516147),
	.w4(32'hbb31e16f),
	.w5(32'h3b9a9598),
	.w6(32'h399acdd4),
	.w7(32'hbb55469b),
	.w8(32'h3c159fc8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33a9cc),
	.w1(32'h3b572c5e),
	.w2(32'h3bea2f33),
	.w3(32'h3b6ec367),
	.w4(32'h3bac59b7),
	.w5(32'h3b75c384),
	.w6(32'hbb47af4d),
	.w7(32'hbc1fc1ac),
	.w8(32'hbb72f9d6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4647ee),
	.w1(32'h3c0b15a7),
	.w2(32'hbc10f4af),
	.w3(32'h3c02bd32),
	.w4(32'h3b8adc2c),
	.w5(32'hba9c28d3),
	.w6(32'hbb4a9754),
	.w7(32'hbc023b3e),
	.w8(32'h3ba30fa8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3e873),
	.w1(32'h3ab2efb9),
	.w2(32'hba851d32),
	.w3(32'h3b8de415),
	.w4(32'h3ba1977b),
	.w5(32'h3c04a0c5),
	.w6(32'h3c19803b),
	.w7(32'h3b46e79b),
	.w8(32'hbb38d132),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73e8c3),
	.w1(32'h3b251712),
	.w2(32'h3bf67f19),
	.w3(32'h3a120955),
	.w4(32'h3bc407e4),
	.w5(32'h39f47aeb),
	.w6(32'hbb228150),
	.w7(32'h3b36624a),
	.w8(32'hbc0a5944),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0014a7),
	.w1(32'hbba5ef2e),
	.w2(32'hbbd87178),
	.w3(32'hbc0e3e3a),
	.w4(32'h3a922e71),
	.w5(32'h3ad206bd),
	.w6(32'hbbc56dec),
	.w7(32'hbaad5b1c),
	.w8(32'h3a1eef63),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2064),
	.w1(32'hbbc98dd2),
	.w2(32'hbc9783a3),
	.w3(32'h3bfa9b58),
	.w4(32'hbb5a8584),
	.w5(32'hbd14f37c),
	.w6(32'h3ab3593f),
	.w7(32'hbb1239a1),
	.w8(32'hbce643ea),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c5b41),
	.w1(32'hbd1c32e0),
	.w2(32'hbb138fae),
	.w3(32'hbd552d67),
	.w4(32'hbd2957fa),
	.w5(32'hbba39b1a),
	.w6(32'hbcd5d2da),
	.w7(32'hbcaf4647),
	.w8(32'hba958cf4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bdb21),
	.w1(32'hbaf821d1),
	.w2(32'h3c21f0fa),
	.w3(32'hbc68172e),
	.w4(32'hbb1bac98),
	.w5(32'h3b3cb75e),
	.w6(32'hbb4eee86),
	.w7(32'hbbbd40fe),
	.w8(32'h3a86e32d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2fd8),
	.w1(32'hbc057d94),
	.w2(32'hbc81a5f6),
	.w3(32'hbbcfa16d),
	.w4(32'h3ac2d0b7),
	.w5(32'hbc41b869),
	.w6(32'h38540dee),
	.w7(32'h3b924199),
	.w8(32'h3ad7bd65),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d814d),
	.w1(32'hbbc79a57),
	.w2(32'hbcdead5c),
	.w3(32'hbb3a1896),
	.w4(32'h3ae1a045),
	.w5(32'h39b53a50),
	.w6(32'hbb82f94c),
	.w7(32'hba43e591),
	.w8(32'h3c418248),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9490aa),
	.w1(32'h3c1a8711),
	.w2(32'h3af95aa3),
	.w3(32'hbb2c24d6),
	.w4(32'h3bc79ec0),
	.w5(32'h3b88ae7b),
	.w6(32'h3c3aa1c1),
	.w7(32'hbafc0139),
	.w8(32'h3c1ae912),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e550a),
	.w1(32'h3bcc3e2e),
	.w2(32'h3c6f1a19),
	.w3(32'hba4463ac),
	.w4(32'h3c58cc93),
	.w5(32'h3cb5a6f3),
	.w6(32'h3b39c3ac),
	.w7(32'h3c897798),
	.w8(32'h3c5b2b71),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce96b44),
	.w1(32'h3c2fdd5b),
	.w2(32'hbb7cafbe),
	.w3(32'h3d270f48),
	.w4(32'h3ca61b25),
	.w5(32'h3bec1124),
	.w6(32'h3d082f19),
	.w7(32'h3caa582d),
	.w8(32'hbafa14f6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0711a6),
	.w1(32'hbc3b0c7d),
	.w2(32'h3ad123d9),
	.w3(32'h3c2f3cfb),
	.w4(32'h3a202e6a),
	.w5(32'h3c4000f7),
	.w6(32'h3b325f86),
	.w7(32'hbc09ab73),
	.w8(32'h3aec04e6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165fa0),
	.w1(32'hbb1c4724),
	.w2(32'hbb6e8077),
	.w3(32'h3bfbc7d6),
	.w4(32'hb908d3ab),
	.w5(32'h3b911034),
	.w6(32'hb9aecfd3),
	.w7(32'h3a969732),
	.w8(32'hba23337e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcf9d2),
	.w1(32'hbc096509),
	.w2(32'h3be6a6e8),
	.w3(32'hba89f61f),
	.w4(32'h3b90ae5f),
	.w5(32'h3c9d5b1a),
	.w6(32'hba0ff8f5),
	.w7(32'hbb80c1ee),
	.w8(32'hbb9a12fd),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f022b),
	.w1(32'hbc040d1b),
	.w2(32'h3b17a78c),
	.w3(32'h3cb737af),
	.w4(32'h3cd7deac),
	.w5(32'hbb0c3c63),
	.w6(32'hbabe70af),
	.w7(32'h3b8f73d2),
	.w8(32'h3b1abb6a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5eeb5),
	.w1(32'hbb0b2087),
	.w2(32'hbcedef22),
	.w3(32'h3b03e9ae),
	.w4(32'h3b74875c),
	.w5(32'hbcc9c702),
	.w6(32'h3bc2fe87),
	.w7(32'h3b3769eb),
	.w8(32'hbcab205b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd104780),
	.w1(32'hbcec5bca),
	.w2(32'hbb051adf),
	.w3(32'hbd059acb),
	.w4(32'hbccb22c3),
	.w5(32'h3bd31d00),
	.w6(32'hbcd82cf2),
	.w7(32'hbcb7a406),
	.w8(32'hbb533349),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f1b15),
	.w1(32'h3b81a06c),
	.w2(32'h3b662e3b),
	.w3(32'h3c3103e2),
	.w4(32'h3c3790a4),
	.w5(32'h3bc81627),
	.w6(32'hbb7fba8a),
	.w7(32'h3a91771e),
	.w8(32'h3ae05db7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25d356),
	.w1(32'hbb882447),
	.w2(32'hbb4377df),
	.w3(32'h3c3b62aa),
	.w4(32'h3b08e4a3),
	.w5(32'hba9077b4),
	.w6(32'hb910873c),
	.w7(32'h3b6a6a67),
	.w8(32'hbc2bcf05),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4308cc),
	.w1(32'h3b4b58ba),
	.w2(32'h3ae9060f),
	.w3(32'hbb35e13f),
	.w4(32'hb968a5d7),
	.w5(32'hb9237dc5),
	.w6(32'hbc067a8b),
	.w7(32'hbb44cf8c),
	.w8(32'h3ae4c126),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bddbf1),
	.w1(32'h3ad3e7bb),
	.w2(32'h3ccbd3d6),
	.w3(32'hb986f058),
	.w4(32'hbb168da8),
	.w5(32'h3cea2e3e),
	.w6(32'h3bcfd6d7),
	.w7(32'h3b026e93),
	.w8(32'h3c09fe71),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6397c),
	.w1(32'hbce79db1),
	.w2(32'hbc5e06c8),
	.w3(32'h3ccb9be9),
	.w4(32'h3c1ea9c5),
	.w5(32'hbc840239),
	.w6(32'h3cb44861),
	.w7(32'h3c7dc6b5),
	.w8(32'hbc2b9eb3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd379f8),
	.w1(32'hbc9f715e),
	.w2(32'h3b748839),
	.w3(32'hbd0d5359),
	.w4(32'hbc9c12aa),
	.w5(32'h3c21aeb2),
	.w6(32'hbcaa49e7),
	.w7(32'hbc1006bb),
	.w8(32'h3c1b0e68),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4886b2),
	.w1(32'h3a1c7ccc),
	.w2(32'h3a5a0fa1),
	.w3(32'h3b854441),
	.w4(32'h3b59d19b),
	.w5(32'h3a550ef9),
	.w6(32'h3bca324e),
	.w7(32'h3be60853),
	.w8(32'hbadc4014),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add22b4),
	.w1(32'h3ab808a5),
	.w2(32'h3c074bde),
	.w3(32'h3bdb1e28),
	.w4(32'h3c13c49c),
	.w5(32'h3ba68c8a),
	.w6(32'hba51db31),
	.w7(32'h3beedb2a),
	.w8(32'h3b16b94b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8a28),
	.w1(32'h3b8b5f05),
	.w2(32'hbba41153),
	.w3(32'hbb4700d7),
	.w4(32'h3b9856fd),
	.w5(32'hbbbea985),
	.w6(32'hbb9c0bd3),
	.w7(32'h3b1bfae2),
	.w8(32'hbc24cc21),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c512f),
	.w1(32'h3b67ad9e),
	.w2(32'hba815af8),
	.w3(32'hbbb7a937),
	.w4(32'h3ac82537),
	.w5(32'h3b631d94),
	.w6(32'hbc927336),
	.w7(32'hbc1bd839),
	.w8(32'hba803c6c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0548ba),
	.w1(32'h3c27ab35),
	.w2(32'h3bb05f81),
	.w3(32'h3ba88203),
	.w4(32'h3bd2e397),
	.w5(32'h3b4faa3a),
	.w6(32'h3bbeb9cf),
	.w7(32'h38f16d5b),
	.w8(32'h3b70afda),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c159339),
	.w1(32'hb9db1662),
	.w2(32'hba15fb84),
	.w3(32'h3b986582),
	.w4(32'h3bd1dab4),
	.w5(32'hbaeca164),
	.w6(32'h3b4430f3),
	.w7(32'h3b41f876),
	.w8(32'h3b19dc1f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7638e),
	.w1(32'h3c80744c),
	.w2(32'h3b790b09),
	.w3(32'hbb23d2de),
	.w4(32'h3b398f35),
	.w5(32'hbc0b3ee0),
	.w6(32'hbba66c36),
	.w7(32'hbad7b684),
	.w8(32'hbaf458a2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae9ed2),
	.w1(32'h3bc71a4c),
	.w2(32'h3bf25036),
	.w3(32'hbc49a804),
	.w4(32'hbc42ce01),
	.w5(32'h3bf6f689),
	.w6(32'h3a2ea7ae),
	.w7(32'h3a938af2),
	.w8(32'hbb944d1a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99eade5),
	.w1(32'hbc2fdc77),
	.w2(32'h3b656592),
	.w3(32'hbb6e49fd),
	.w4(32'hba44e04b),
	.w5(32'h3b26cf9c),
	.w6(32'hbc2dcbfb),
	.w7(32'hba00dc15),
	.w8(32'hbc0a3b00),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eea8d),
	.w1(32'h3c067c9b),
	.w2(32'h3c037a06),
	.w3(32'h3a8d97a2),
	.w4(32'h3c188d80),
	.w5(32'h3c10f193),
	.w6(32'hbc6b2afa),
	.w7(32'hbac5a2c9),
	.w8(32'h3c141e47),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19f82f),
	.w1(32'h3ad9a194),
	.w2(32'hbaeb5977),
	.w3(32'h3bdf8d3c),
	.w4(32'h3ba491bb),
	.w5(32'h3c121468),
	.w6(32'h3c2c6e22),
	.w7(32'h3b8be82e),
	.w8(32'h3baf2eef),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafd377),
	.w1(32'hbc286a4c),
	.w2(32'h3aab9d30),
	.w3(32'h3c0deed8),
	.w4(32'h3be0f617),
	.w5(32'h3a8aeb81),
	.w6(32'h3baf2056),
	.w7(32'h3bd7de70),
	.w8(32'h3b31560a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde546),
	.w1(32'h3b62fad1),
	.w2(32'h3b4d30dd),
	.w3(32'h3b2f53d6),
	.w4(32'h3bbfef59),
	.w5(32'hba9f9f1a),
	.w6(32'h3c4ff2d3),
	.w7(32'h3bfb97f8),
	.w8(32'hb99bf459),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9605cb),
	.w1(32'hbafd953d),
	.w2(32'hbc633dc3),
	.w3(32'h3bd6dc21),
	.w4(32'h366302c9),
	.w5(32'hbc0da0d7),
	.w6(32'h3bc8aaf7),
	.w7(32'hbbc1625a),
	.w8(32'hbc2d5206),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64d654),
	.w1(32'hbc1eee40),
	.w2(32'hbb97f67b),
	.w3(32'hbcdcd85f),
	.w4(32'hbc265d51),
	.w5(32'hbbd9c668),
	.w6(32'hbcf38427),
	.w7(32'hbc451d01),
	.w8(32'hbbb54370),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32d68),
	.w1(32'hbbf0f5f0),
	.w2(32'hb9fb29ba),
	.w3(32'hbba0bfbf),
	.w4(32'hbbc601c1),
	.w5(32'h3ba17747),
	.w6(32'hbb7e5f72),
	.w7(32'hbbc24fd2),
	.w8(32'h3abf069c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63d1c4),
	.w1(32'hbbf88566),
	.w2(32'hbbd4f0c3),
	.w3(32'hbb325f91),
	.w4(32'h3816b998),
	.w5(32'h3bd538b5),
	.w6(32'h3bdfd748),
	.w7(32'h3b5d0227),
	.w8(32'hbb0e3c80),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847d5b),
	.w1(32'hbb0fbe63),
	.w2(32'hbd30e9cf),
	.w3(32'hbae5d40c),
	.w4(32'h3c406134),
	.w5(32'hbc9a48bd),
	.w6(32'hbb0c4343),
	.w7(32'h3bb79dbc),
	.w8(32'hbc9db8ea),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5d3f8e),
	.w1(32'hbd2fb4e0),
	.w2(32'hbc823330),
	.w3(32'hbd1b56a2),
	.w4(32'hbc9423d8),
	.w5(32'h3cb4dbfd),
	.w6(32'hbd186bb0),
	.w7(32'hbcde8c50),
	.w8(32'h3cfbfb6e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc5673),
	.w1(32'hbcdc8f4d),
	.w2(32'hbbe73124),
	.w3(32'h3cd859ff),
	.w4(32'h3c01928c),
	.w5(32'hbc8d7030),
	.w6(32'h3d127292),
	.w7(32'h3c9f0d55),
	.w8(32'hbca0a5bb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05d10),
	.w1(32'hbbbeb0c0),
	.w2(32'hbbda1cc9),
	.w3(32'hbc8042b8),
	.w4(32'hbc809fd2),
	.w5(32'hba31c657),
	.w6(32'hbca5430d),
	.w7(32'hbca224e7),
	.w8(32'h3b84377d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc175978),
	.w1(32'hbc08df0f),
	.w2(32'hbaade85c),
	.w3(32'hb9abc7df),
	.w4(32'hbb6616ce),
	.w5(32'hbb270729),
	.w6(32'h3c264fca),
	.w7(32'h3ba441a8),
	.w8(32'hbb2f2d2b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8fb5b),
	.w1(32'hbb7d7cbc),
	.w2(32'h3bfc44bc),
	.w3(32'hbb477b2b),
	.w4(32'h3a5ec343),
	.w5(32'hbb7b101c),
	.w6(32'h39b4cd7b),
	.w7(32'hbb4f86fe),
	.w8(32'h3a6f377e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645830),
	.w1(32'hbb9edcac),
	.w2(32'h3bd21713),
	.w3(32'hbc198fbc),
	.w4(32'hbbc3c809),
	.w5(32'h3aee0ebc),
	.w6(32'h3b2aaf2e),
	.w7(32'h3b2c7f7f),
	.w8(32'hbbd1f3de),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae66b61),
	.w1(32'h3c1ce098),
	.w2(32'hbb94c1be),
	.w3(32'hbbfe9d4a),
	.w4(32'h3b41b38c),
	.w5(32'hbbc71385),
	.w6(32'hbc2142ce),
	.w7(32'h3a67cf03),
	.w8(32'hbbb3dab5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdbfe2),
	.w1(32'hbbd0000c),
	.w2(32'hba560007),
	.w3(32'h3ac7a505),
	.w4(32'hba8035d6),
	.w5(32'h3bcf12bb),
	.w6(32'h3b22ba82),
	.w7(32'h3b4c7e08),
	.w8(32'hbb3ea15c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae33716),
	.w1(32'h3a48fe2e),
	.w2(32'hba95b9b3),
	.w3(32'h3b378919),
	.w4(32'hbb004c20),
	.w5(32'hbb69a1bb),
	.w6(32'hbc2fe21f),
	.w7(32'hbc0c46a8),
	.w8(32'hbc831d6f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d393d),
	.w1(32'hbb4adfdc),
	.w2(32'hbbaea30b),
	.w3(32'h3c14ad56),
	.w4(32'h3c2982ab),
	.w5(32'hbaff953f),
	.w6(32'hb9cc3fac),
	.w7(32'h3c466d8b),
	.w8(32'h3be68b72),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff4f26),
	.w1(32'hb9038d10),
	.w2(32'h3acbe527),
	.w3(32'hbbdb7df2),
	.w4(32'h3a57f865),
	.w5(32'h38295e74),
	.w6(32'hbba0c04e),
	.w7(32'h3a8658bf),
	.w8(32'h3b0613c1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72bdf2),
	.w1(32'hbbc41c7b),
	.w2(32'h3c37f227),
	.w3(32'hbbda4ab0),
	.w4(32'hbc0464f8),
	.w5(32'h3b9e905e),
	.w6(32'hba13e499),
	.w7(32'h3968e407),
	.w8(32'h3c0beaed),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88b46c),
	.w1(32'h3c3ab235),
	.w2(32'hbc29804f),
	.w3(32'hbbbd4c08),
	.w4(32'h3ba26f2f),
	.w5(32'hbcd65bd5),
	.w6(32'hbb9bdbb4),
	.w7(32'h3bfd45b0),
	.w8(32'hbcc42426),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd042fd6),
	.w1(32'hbd0c88bf),
	.w2(32'hbb31070f),
	.w3(32'hbd3b6537),
	.w4(32'hbcce4816),
	.w5(32'hb9bad6cd),
	.w6(32'hbcf9d099),
	.w7(32'hbc276b6f),
	.w8(32'hba05615a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39a358),
	.w1(32'h3ba96add),
	.w2(32'hbb811e0e),
	.w3(32'h3c00a9ca),
	.w4(32'h3b5a3212),
	.w5(32'hbb6880c2),
	.w6(32'hbb0fd722),
	.w7(32'hbb10faae),
	.w8(32'hba9d3eb0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f13c),
	.w1(32'h39cb92ad),
	.w2(32'hbbd783d1),
	.w3(32'hbc98512a),
	.w4(32'h3b4ce23a),
	.w5(32'hbc26d400),
	.w6(32'hbc54434e),
	.w7(32'hb9a3556b),
	.w8(32'hbc4726c0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dcc10),
	.w1(32'hbb420267),
	.w2(32'h3b2890f7),
	.w3(32'hbcc6dfd6),
	.w4(32'hbab93c60),
	.w5(32'h3aad5dd9),
	.w6(32'hbc907faf),
	.w7(32'hbbb4ae35),
	.w8(32'hbbf3f25c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6eff3),
	.w1(32'h3c6f8138),
	.w2(32'hbc1a5bb9),
	.w3(32'h3c81e827),
	.w4(32'h3c229c82),
	.w5(32'h3ae1a793),
	.w6(32'h3b733a70),
	.w7(32'h3be74b2c),
	.w8(32'h3b36d290),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad86239),
	.w1(32'h3b945b71),
	.w2(32'hbc130184),
	.w3(32'h3b4fd695),
	.w4(32'h3bceea4a),
	.w5(32'h3b6b1078),
	.w6(32'hbb063731),
	.w7(32'h3b8529c7),
	.w8(32'hbb9f1821),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb307d59),
	.w1(32'hbad80822),
	.w2(32'hbc01dd91),
	.w3(32'hbb8c152c),
	.w4(32'hbab4fdd7),
	.w5(32'h3bb14a12),
	.w6(32'hbbc4c155),
	.w7(32'hbc407248),
	.w8(32'hba151968),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee003b),
	.w1(32'h3bb7f40a),
	.w2(32'hbc11af54),
	.w3(32'h3b452b93),
	.w4(32'h3beec5c2),
	.w5(32'h3a762488),
	.w6(32'h3aee746c),
	.w7(32'h3b9e15c0),
	.w8(32'h3b161ca7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03cbbb),
	.w1(32'hbb9692b8),
	.w2(32'hbae92b96),
	.w3(32'h3a62ca44),
	.w4(32'h3b38cc45),
	.w5(32'h39e6baf7),
	.w6(32'hb865cf75),
	.w7(32'hbb432fec),
	.w8(32'hb96f2736),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa40cb7),
	.w1(32'hbbadb74a),
	.w2(32'h3b2b8899),
	.w3(32'hba895e86),
	.w4(32'hbbdac7d1),
	.w5(32'hbab5648e),
	.w6(32'h3bb6f095),
	.w7(32'h3bce14d0),
	.w8(32'hbc291b2f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc9cd),
	.w1(32'h38a63f08),
	.w2(32'h3b8a3fbc),
	.w3(32'hbab89fc0),
	.w4(32'hbac9e439),
	.w5(32'hbadf3223),
	.w6(32'hbc22a01e),
	.w7(32'hbbbffbcb),
	.w8(32'hbc307143),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65da25),
	.w1(32'h3cc0ee47),
	.w2(32'h3cb77e1d),
	.w3(32'h3b04769b),
	.w4(32'h3c115360),
	.w5(32'h3cb431d6),
	.w6(32'hbc05d097),
	.w7(32'hba93a20e),
	.w8(32'h3c89b957),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0eed2a),
	.w1(32'h3cbc65e4),
	.w2(32'hbd7bd90f),
	.w3(32'h3d068f2f),
	.w4(32'h3cbf2123),
	.w5(32'hbd685200),
	.w6(32'h3cf951b1),
	.w7(32'h3ce7f6d4),
	.w8(32'hbd250dfb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb3cb8d),
	.w1(32'hbd934534),
	.w2(32'h3cc6af9f),
	.w3(32'hbdab551c),
	.w4(32'hbd8a419e),
	.w5(32'h3cee71a8),
	.w6(32'hbd7bd94d),
	.w7(32'hbd756eb4),
	.w8(32'h3c88cd58),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1a8c6d),
	.w1(32'h3cec9d09),
	.w2(32'hbbf8d7c0),
	.w3(32'h3d362ed4),
	.w4(32'h3d1f9991),
	.w5(32'h3c0429a7),
	.w6(32'h3d066670),
	.w7(32'h3cf77ef2),
	.w8(32'hbaee9f9f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d722c),
	.w1(32'hbb247cf1),
	.w2(32'hbb81a952),
	.w3(32'hbb24468f),
	.w4(32'h3940689a),
	.w5(32'hbb8db052),
	.w6(32'hbaebf913),
	.w7(32'hb92af04a),
	.w8(32'h399858ed),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022f87),
	.w1(32'hb9e824c7),
	.w2(32'hba6cd870),
	.w3(32'hbb741ecf),
	.w4(32'hbb9e5998),
	.w5(32'h3bc2a041),
	.w6(32'hbaf88f1e),
	.w7(32'hbb1385f3),
	.w8(32'hba0b472b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558044),
	.w1(32'h3c0283bb),
	.w2(32'h39627862),
	.w3(32'h3ba87b89),
	.w4(32'hba17be01),
	.w5(32'h3a77819a),
	.w6(32'h3ab2846d),
	.w7(32'h3b01092f),
	.w8(32'h3b943434),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3c19),
	.w1(32'hbb8fb35b),
	.w2(32'hbb7e16d0),
	.w3(32'h3a296b62),
	.w4(32'h3a1b84af),
	.w5(32'h3b045c24),
	.w6(32'h3a9fdf32),
	.w7(32'h3abfef5b),
	.w8(32'h3bd3f458),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321f63),
	.w1(32'hbbd1b20f),
	.w2(32'h3bb06f6b),
	.w3(32'hbb946228),
	.w4(32'hbb08f3ca),
	.w5(32'h3c08c68f),
	.w6(32'h3a20f857),
	.w7(32'h3a9fe4a0),
	.w8(32'hbb441e8e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb120c0d),
	.w1(32'hbb9e37d4),
	.w2(32'h3bc32497),
	.w3(32'hbc253537),
	.w4(32'hbbcf6c37),
	.w5(32'h3b17f363),
	.w6(32'hbcab6e7d),
	.w7(32'hbb9df396),
	.w8(32'h3c08688f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3373e8),
	.w1(32'h3c6e6af8),
	.w2(32'h3c2ac456),
	.w3(32'h3b6c7bd9),
	.w4(32'h3bc3e99e),
	.w5(32'h3b35839f),
	.w6(32'h3c40c757),
	.w7(32'h3be6d5e4),
	.w8(32'h3bea00a5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06c103),
	.w1(32'hbb2492fd),
	.w2(32'h3b0ac106),
	.w3(32'h3b9d6a0e),
	.w4(32'h3b824d0a),
	.w5(32'h3c22d0f1),
	.w6(32'h3c664c86),
	.w7(32'h3c8cbeaa),
	.w8(32'h3c306f40),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1264b8),
	.w1(32'hbb880be9),
	.w2(32'hbb52a577),
	.w3(32'h3c0987ce),
	.w4(32'h3b3305ae),
	.w5(32'h3bcedf78),
	.w6(32'h3c140d20),
	.w7(32'h3c3ec704),
	.w8(32'h3b8e07b8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a825e44),
	.w1(32'h3bcabf95),
	.w2(32'hb945b73f),
	.w3(32'h3c0abeb3),
	.w4(32'h3bc05c85),
	.w5(32'h3b8e42af),
	.w6(32'h39a7f759),
	.w7(32'h3a81d75a),
	.w8(32'hbc18e763),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule