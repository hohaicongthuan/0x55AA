module layer_10_featuremap_143(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e9b5b2),
	.w1(32'h36f371c0),
	.w2(32'h3706e022),
	.w3(32'h37a81673),
	.w4(32'h379aaa80),
	.w5(32'h3798dc5e),
	.w6(32'h37c79fe9),
	.w7(32'h37c1b064),
	.w8(32'h37051af5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974afe4),
	.w1(32'h395ce137),
	.w2(32'hba093100),
	.w3(32'h3a758d36),
	.w4(32'h3a99a4a0),
	.w5(32'hb8d44331),
	.w6(32'h3a67b503),
	.w7(32'h3a4c8783),
	.w8(32'h37fd2fd0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ba2bcf),
	.w1(32'h36d1cc1c),
	.w2(32'h36c5a96a),
	.w3(32'h36634aa8),
	.w4(32'h36431d71),
	.w5(32'h366cdabf),
	.w6(32'h370b78d2),
	.w7(32'h36bb99c9),
	.w8(32'h3700ddcf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38312f0f),
	.w1(32'h37e7a250),
	.w2(32'h383c2089),
	.w3(32'h380602b8),
	.w4(32'hb80b6b23),
	.w5(32'h38c58647),
	.w6(32'hb818c84d),
	.w7(32'hb84de4d4),
	.w8(32'hb892c30a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fb60c),
	.w1(32'h3974b7fb),
	.w2(32'h381174fe),
	.w3(32'h39b344da),
	.w4(32'h39af9a3b),
	.w5(32'h38993aa6),
	.w6(32'h39b4f37c),
	.w7(32'h39bec8c1),
	.w8(32'h390e2f79),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb688e156),
	.w1(32'hb74601df),
	.w2(32'h36a22f81),
	.w3(32'hb501306b),
	.w4(32'hb723d91b),
	.w5(32'h3600e218),
	.w6(32'h370c12f0),
	.w7(32'h371883ca),
	.w8(32'h37a01634),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae54b94),
	.w1(32'h3a8a83d5),
	.w2(32'h3aa0dd41),
	.w3(32'h3b32dcca),
	.w4(32'h3a2ae271),
	.w5(32'h385d523e),
	.w6(32'h38d48e59),
	.w7(32'hba9338f0),
	.w8(32'hbaf31d5a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ef78),
	.w1(32'hbb599872),
	.w2(32'hbb533273),
	.w3(32'hbbfaee87),
	.w4(32'hbba64c6e),
	.w5(32'hbb1fbd5a),
	.w6(32'hbac46fa1),
	.w7(32'hbb70710b),
	.w8(32'hba86e375),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afb57c),
	.w1(32'hb8564b25),
	.w2(32'hb9d5eab5),
	.w3(32'h3a03bf52),
	.w4(32'h3a1b79df),
	.w5(32'h37b4828e),
	.w6(32'h38dc05b0),
	.w7(32'hb7c08ccf),
	.w8(32'hba0ccf44),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76aa7c),
	.w1(32'hbab893d3),
	.w2(32'h3ab86dca),
	.w3(32'hbb6dd9ac),
	.w4(32'hba907d48),
	.w5(32'hba4f2f82),
	.w6(32'hbb514027),
	.w7(32'hba2a93a2),
	.w8(32'hbac34da3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947a7ab),
	.w1(32'hb715c313),
	.w2(32'hb8f5ebd3),
	.w3(32'hba143e99),
	.w4(32'hb909a346),
	.w5(32'hb9f9c17e),
	.w6(32'hb9cf59e0),
	.w7(32'hb869878d),
	.w8(32'hb983f582),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b210212),
	.w1(32'h3b08c5e2),
	.w2(32'h3b188205),
	.w3(32'h3b7f8670),
	.w4(32'h3b0b9048),
	.w5(32'h3b440e13),
	.w6(32'h3b587929),
	.w7(32'h3a7e7454),
	.w8(32'h3aa7f2e8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2459cd),
	.w1(32'h3a38ace8),
	.w2(32'h3aedd9cb),
	.w3(32'hbb421257),
	.w4(32'hb9dbc0be),
	.w5(32'hbaa32987),
	.w6(32'hba389044),
	.w7(32'h3a5bcba1),
	.w8(32'hba51c64b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b3bc2),
	.w1(32'h3ab466d4),
	.w2(32'h3a498421),
	.w3(32'h3910e08e),
	.w4(32'h3a519a38),
	.w5(32'h384b072d),
	.w6(32'h3a2b2d35),
	.w7(32'h3a832590),
	.w8(32'h381e0b86),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f05d25),
	.w1(32'hba17ee1b),
	.w2(32'hbab4e751),
	.w3(32'h3a2e2e01),
	.w4(32'h3a4e4b47),
	.w5(32'h393a09c4),
	.w6(32'hba07fde3),
	.w7(32'hb9222d2a),
	.w8(32'h39fccfc3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2883aa),
	.w1(32'h3abfc8af),
	.w2(32'h3ad11670),
	.w3(32'hbb8d32a6),
	.w4(32'hba3a1564),
	.w5(32'hb6d59032),
	.w6(32'hbb7a0c95),
	.w7(32'hba312963),
	.w8(32'hbad2b6f5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9af4d),
	.w1(32'h388aa11d),
	.w2(32'h364ab248),
	.w3(32'h397daa39),
	.w4(32'h38226416),
	.w5(32'h391d48c0),
	.w6(32'h3972e3e7),
	.w7(32'h380d6fc8),
	.w8(32'h3933d576),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bcac3),
	.w1(32'hbad26357),
	.w2(32'hbab17f1a),
	.w3(32'hbbe8ca02),
	.w4(32'hbba72dd5),
	.w5(32'hbb1a76c9),
	.w6(32'hbb790ae9),
	.w7(32'hbbb07a62),
	.w8(32'hbbaa4d34),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaed546),
	.w1(32'h398ccd3b),
	.w2(32'h3a823190),
	.w3(32'hbb59d32a),
	.w4(32'hbaf3ca5d),
	.w5(32'hb9d80894),
	.w6(32'hbacdca76),
	.w7(32'hbaeb68a5),
	.w8(32'hbadbe40e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35937f4a),
	.w1(32'hb7822d85),
	.w2(32'h384fd095),
	.w3(32'h37e3a405),
	.w4(32'h37b7f159),
	.w5(32'h38937302),
	.w6(32'hb6c7bd69),
	.w7(32'h3859a292),
	.w8(32'h37bfc42e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5f2a2),
	.w1(32'hb8f0889e),
	.w2(32'h36ae2433),
	.w3(32'h37860747),
	.w4(32'hb8f4cb9b),
	.w5(32'hb7348b1e),
	.w6(32'hb6e4e76b),
	.w7(32'hb7b38b9e),
	.w8(32'h388620a7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab61d73),
	.w1(32'h3a53cdcf),
	.w2(32'h3956df88),
	.w3(32'h3ac541b6),
	.w4(32'h3a96888e),
	.w5(32'h3a2018bc),
	.w6(32'h3a9b4c61),
	.w7(32'h3a60c3b7),
	.w8(32'h3a5ae0a7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ceab),
	.w1(32'hbb02e6bd),
	.w2(32'h39aa26bc),
	.w3(32'hbb5f2f79),
	.w4(32'hba5ad81a),
	.w5(32'hbaa240c9),
	.w6(32'hbbe516f6),
	.w7(32'hbb5d7047),
	.w8(32'hbbbc2cfc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafad1ff),
	.w1(32'hba3a08e3),
	.w2(32'h39ba5f42),
	.w3(32'hba994fc8),
	.w4(32'hba1e3822),
	.w5(32'hba53e355),
	.w6(32'hbab54d58),
	.w7(32'hb9e06495),
	.w8(32'hba8ed9bc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b9d86),
	.w1(32'hba80d406),
	.w2(32'hbb00195d),
	.w3(32'hb8d371d9),
	.w4(32'h3a964097),
	.w5(32'hba47ab55),
	.w6(32'hba52786b),
	.w7(32'h3a15d200),
	.w8(32'h3a5d5b1d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964ba6e),
	.w1(32'h3a3c65a2),
	.w2(32'h3a0b072d),
	.w3(32'hb9426f91),
	.w4(32'h3a016caf),
	.w5(32'h39686d29),
	.w6(32'hb9fef161),
	.w7(32'h39da82b5),
	.w8(32'h399fcfff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a403c1),
	.w1(32'h37cc340c),
	.w2(32'h38933693),
	.w3(32'h38801146),
	.w4(32'h37210b32),
	.w5(32'h3876d8e3),
	.w6(32'h38e52d82),
	.w7(32'h3865af1b),
	.w8(32'h390df098),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0c699),
	.w1(32'h3b1a1be0),
	.w2(32'hba4e1836),
	.w3(32'h3990af44),
	.w4(32'h3b398bad),
	.w5(32'hb98695d9),
	.w6(32'h3a7506e0),
	.w7(32'h3a93b0c7),
	.w8(32'hba174736),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ec1b4),
	.w1(32'h3a13a7e4),
	.w2(32'h3a8f56e3),
	.w3(32'h3a9b71d6),
	.w4(32'h3a6ebf8a),
	.w5(32'h3aa6b2de),
	.w6(32'h3a74ac5a),
	.w7(32'h39e3e1a1),
	.w8(32'h3abb0ed4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88bb85),
	.w1(32'h3b261edb),
	.w2(32'hb90fe22d),
	.w3(32'hb981ef7c),
	.w4(32'h3b75113d),
	.w5(32'hb9b79d1a),
	.w6(32'h3aa0523a),
	.w7(32'h3b80efaa),
	.w8(32'hba25cfca),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384f04cd),
	.w1(32'h3804bb88),
	.w2(32'h3839c31a),
	.w3(32'h38249d5e),
	.w4(32'h37e5ec78),
	.w5(32'h3811dc32),
	.w6(32'h38622be8),
	.w7(32'h38428acb),
	.w8(32'h386ba74f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0822a),
	.w1(32'hb92feca7),
	.w2(32'hb7dc2f84),
	.w3(32'hb8b68a8d),
	.w4(32'hb92b127d),
	.w5(32'h391bec39),
	.w6(32'hb86a4d90),
	.w7(32'h379c796c),
	.w8(32'h39aaaf1a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9841c53),
	.w1(32'hb9868aef),
	.w2(32'hb8c3271f),
	.w3(32'hb9ed54a8),
	.w4(32'hb9971574),
	.w5(32'hb9e8510c),
	.w6(32'hb9c47f56),
	.w7(32'hb8c5e098),
	.w8(32'hba0393dc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ffaef),
	.w1(32'hb9d0fedd),
	.w2(32'hba4d7a71),
	.w3(32'hb950a02a),
	.w4(32'h39aaaa45),
	.w5(32'hb9bd6d80),
	.w6(32'hb9b2f53a),
	.w7(32'h3982b5fd),
	.w8(32'hb999ba33),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c61da),
	.w1(32'hb810480c),
	.w2(32'h39a92216),
	.w3(32'h38bc394e),
	.w4(32'h393623e4),
	.w5(32'h39bf51ca),
	.w6(32'h38faa38d),
	.w7(32'hb9211349),
	.w8(32'h38946ee3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadcb45),
	.w1(32'h39a6eb9a),
	.w2(32'h3a9903e4),
	.w3(32'h399a0d6a),
	.w4(32'hba98a88a),
	.w5(32'h37a9ff2f),
	.w6(32'h3a337dc8),
	.w7(32'h3916b671),
	.w8(32'hb9af9bb7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da0c17),
	.w1(32'hbb93f4c4),
	.w2(32'h3afe0095),
	.w3(32'h3b2946c8),
	.w4(32'hbb99639d),
	.w5(32'h3b80cc37),
	.w6(32'h39b9c8cb),
	.w7(32'hbb14d8bc),
	.w8(32'hb9842043),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f88872),
	.w1(32'h3a72bd39),
	.w2(32'hbb174331),
	.w3(32'h3b4f7e8c),
	.w4(32'h3b9acde3),
	.w5(32'h3adc8712),
	.w6(32'h39becb0c),
	.w7(32'h3b2f9a58),
	.w8(32'h3b45391d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be181a1),
	.w1(32'h3bf01b75),
	.w2(32'h3ad46df6),
	.w3(32'h3c04d66a),
	.w4(32'h3c048ab1),
	.w5(32'h3b25b1c0),
	.w6(32'h3bcc38fb),
	.w7(32'h3b5fb7d5),
	.w8(32'h3a4ab505),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dced9),
	.w1(32'hba0382aa),
	.w2(32'hba8a8c84),
	.w3(32'hb8da65cc),
	.w4(32'hb9501462),
	.w5(32'hb9a71dc7),
	.w6(32'hb998d5f9),
	.w7(32'hb96b2b4f),
	.w8(32'hb98d3248),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d810e1),
	.w1(32'hb99b18a1),
	.w2(32'hb841ed20),
	.w3(32'hb9d9d555),
	.w4(32'hb9289454),
	.w5(32'hb8dcf28d),
	.w6(32'hb97c9e00),
	.w7(32'hb8a82b0f),
	.w8(32'h37f26ebd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f9531a),
	.w1(32'hb76ce770),
	.w2(32'hb8c49795),
	.w3(32'h392e8581),
	.w4(32'h370874c5),
	.w5(32'hb90c1d66),
	.w6(32'h398c9656),
	.w7(32'hb7f580aa),
	.w8(32'hb9830316),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896f7e4),
	.w1(32'h3ac0c8e5),
	.w2(32'h3ae3b7ac),
	.w3(32'h3866abd9),
	.w4(32'h3ab3f95b),
	.w5(32'h3a917545),
	.w6(32'hba2cf491),
	.w7(32'h3a598822),
	.w8(32'h3a3de02d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fcee8),
	.w1(32'h39f31f6b),
	.w2(32'h3abf0cab),
	.w3(32'hbbb79184),
	.w4(32'hb9aa140a),
	.w5(32'hbb46b249),
	.w6(32'hbb6876b3),
	.w7(32'hba2c0a08),
	.w8(32'hbb4b33f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6614cd),
	.w1(32'hba5e871e),
	.w2(32'hba4c7de9),
	.w3(32'hbb132227),
	.w4(32'h3a49430c),
	.w5(32'hb8cfdf95),
	.w6(32'hbaa58800),
	.w7(32'h3a952ace),
	.w8(32'h39a35385),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f613),
	.w1(32'hbafc8c99),
	.w2(32'h3a294343),
	.w3(32'hbb0bedfb),
	.w4(32'hba47e855),
	.w5(32'h384adc81),
	.w6(32'hbaaa4a9b),
	.w7(32'h3aa21578),
	.w8(32'h39c2a831),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185aea),
	.w1(32'h389cacc1),
	.w2(32'h397be52b),
	.w3(32'hba2b450b),
	.w4(32'h3a8a10f4),
	.w5(32'h3a7926e8),
	.w6(32'hbab5ac7c),
	.w7(32'h39025600),
	.w8(32'hba8c7501),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86d8f1e),
	.w1(32'h38720803),
	.w2(32'h39f16631),
	.w3(32'hbbb07239),
	.w4(32'hbb8508f6),
	.w5(32'hba457343),
	.w6(32'hbb82e1aa),
	.w7(32'hbb7f876b),
	.w8(32'hbb3711d3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b9665),
	.w1(32'hba094ce7),
	.w2(32'hb91a2800),
	.w3(32'hba05a915),
	.w4(32'hb909694a),
	.w5(32'hb90117b2),
	.w6(32'hb9b70d1e),
	.w7(32'h376f0688),
	.w8(32'hb9b0f91b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa17eef),
	.w1(32'hb9e483d9),
	.w2(32'hb9977d1e),
	.w3(32'hba21e050),
	.w4(32'hb9449267),
	.w5(32'hba744f34),
	.w6(32'hb9f9f530),
	.w7(32'hba18fb9b),
	.w8(32'hbac729b0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afa2c0),
	.w1(32'hb9b31e04),
	.w2(32'hb971c180),
	.w3(32'h39a7b5b0),
	.w4(32'h39a4ec24),
	.w5(32'hb901b45b),
	.w6(32'h39965acf),
	.w7(32'h399128a2),
	.w8(32'hb6b266af),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f41cc),
	.w1(32'hb9b04463),
	.w2(32'hba24e3f1),
	.w3(32'hbb0d9dec),
	.w4(32'hb880562b),
	.w5(32'hba9f2f89),
	.w6(32'hba9b5e53),
	.w7(32'h3a1a6953),
	.w8(32'hba8140e8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78c516),
	.w1(32'hba48530b),
	.w2(32'hba1f102f),
	.w3(32'hba211e86),
	.w4(32'hba303e00),
	.w5(32'hb9a488a0),
	.w6(32'h38a138db),
	.w7(32'hb998b5eb),
	.w8(32'hba1c9385),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3618),
	.w1(32'hbb1e78a1),
	.w2(32'hb8f37d1b),
	.w3(32'hbbcad193),
	.w4(32'hbb781c0c),
	.w5(32'hb81d0744),
	.w6(32'hbb70fe68),
	.w7(32'hbb53a903),
	.w8(32'hbafca55d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e8d19),
	.w1(32'hb92e7d76),
	.w2(32'hb9574dfe),
	.w3(32'hb951cc23),
	.w4(32'hb91b8833),
	.w5(32'hb8b5e8ef),
	.w6(32'h3a0efe64),
	.w7(32'hb92d7c03),
	.w8(32'hb90cddea),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2ee66),
	.w1(32'h390e525f),
	.w2(32'hb7b4df67),
	.w3(32'h384149fb),
	.w4(32'h3921fbb6),
	.w5(32'hb7b1ffce),
	.w6(32'h37a42e2b),
	.w7(32'h392e608f),
	.w8(32'h372f70b9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e8f165),
	.w1(32'hb81b0b9a),
	.w2(32'hb8338d1e),
	.w3(32'h37c89824),
	.w4(32'hb7c4e6c9),
	.w5(32'hb7d5d60f),
	.w6(32'h382210b5),
	.w7(32'h374d4338),
	.w8(32'h369cf7b7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965832b),
	.w1(32'h38d90e5b),
	.w2(32'hb8ffd4eb),
	.w3(32'h3998757e),
	.w4(32'h3917878d),
	.w5(32'hb9362aad),
	.w6(32'h3999f7b9),
	.w7(32'hb78d4a69),
	.w8(32'hb83a0d7d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a705984),
	.w1(32'h3a68d655),
	.w2(32'h3a182043),
	.w3(32'h3a4fa107),
	.w4(32'h3a5d01c4),
	.w5(32'h3a091275),
	.w6(32'h3a1c7590),
	.w7(32'h3a1f2f30),
	.w8(32'h39f6d4bb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a38f6d),
	.w1(32'h39b06f8f),
	.w2(32'h3989cd9d),
	.w3(32'hb9b14b3d),
	.w4(32'h38733644),
	.w5(32'hb8dbf55f),
	.w6(32'hb90538b2),
	.w7(32'h384e5848),
	.w8(32'hb96e8b09),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca611),
	.w1(32'hb8480d00),
	.w2(32'h39f0b453),
	.w3(32'hbaec1cd2),
	.w4(32'hba34d736),
	.w5(32'hb9adb70f),
	.w6(32'h3658018d),
	.w7(32'hb7d5f476),
	.w8(32'hbaaaf9a5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdf2a),
	.w1(32'h348633b4),
	.w2(32'hb8c66af1),
	.w3(32'hbb98f06e),
	.w4(32'hba087b83),
	.w5(32'hba7833f0),
	.w6(32'hbb3b7af7),
	.w7(32'hb9f64182),
	.w8(32'hba08d877),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90738f9),
	.w1(32'hb8a94cbe),
	.w2(32'hb675070e),
	.w3(32'hb88c3a1e),
	.w4(32'hb675b6b2),
	.w5(32'h37ea4d4a),
	.w6(32'hb63cda42),
	.w7(32'h382a9a67),
	.w8(32'h3874207c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cf29b),
	.w1(32'hb6ce3117),
	.w2(32'h36704ef3),
	.w3(32'hb7ae6253),
	.w4(32'hb75d8610),
	.w5(32'h36beec5b),
	.w6(32'hb6ca36c8),
	.w7(32'h3626ab38),
	.w8(32'h37b6436d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cbccfc),
	.w1(32'hb801f862),
	.w2(32'h381fb8cc),
	.w3(32'hb7493422),
	.w4(32'hb8bd3b6d),
	.w5(32'hb8996ac5),
	.w6(32'h389cc8f6),
	.w7(32'hb6690dea),
	.w8(32'h37021b12),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37555d81),
	.w1(32'hb8004e83),
	.w2(32'h3813dba8),
	.w3(32'h3777fc05),
	.w4(32'hb6ec013a),
	.w5(32'h38599fa1),
	.w6(32'h387d6ec8),
	.w7(32'h384a2206),
	.w8(32'h38e477e0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5cae),
	.w1(32'h39c43c53),
	.w2(32'h3a6f914f),
	.w3(32'hbb06fee3),
	.w4(32'hba02f518),
	.w5(32'h3ab51c85),
	.w6(32'hbb5f165d),
	.w7(32'hbb2008ab),
	.w8(32'hba37f9c6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2962c8),
	.w1(32'hbb26b92d),
	.w2(32'hba8b3694),
	.w3(32'hba4b65b2),
	.w4(32'hbb678611),
	.w5(32'hbb23f983),
	.w6(32'hb8f9131d),
	.w7(32'hba07f3aa),
	.w8(32'hbadc08fd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ce31),
	.w1(32'hbb0059e2),
	.w2(32'hbadf9826),
	.w3(32'hbae1c4e0),
	.w4(32'hba9c9e13),
	.w5(32'hba9ed3bc),
	.w6(32'hbae3f8ad),
	.w7(32'hbadb1995),
	.w8(32'hbb0a57f8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf577f1),
	.w1(32'hba428851),
	.w2(32'hbb3454f7),
	.w3(32'h3a30a4f7),
	.w4(32'h3b307499),
	.w5(32'hb9acd66b),
	.w6(32'hb97082b1),
	.w7(32'h3b09013c),
	.w8(32'h3a912738),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a4545a),
	.w1(32'hb72812e2),
	.w2(32'h37c062eb),
	.w3(32'h3683a19b),
	.w4(32'hb6a12622),
	.w5(32'h37baab20),
	.w6(32'h380b529d),
	.w7(32'h37d9e7c0),
	.w8(32'h38588785),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3771d540),
	.w1(32'hb6d19ba8),
	.w2(32'h380b6f49),
	.w3(32'hb6cb5da0),
	.w4(32'hb7813ca6),
	.w5(32'h37dfa9d3),
	.w6(32'h38283eb3),
	.w7(32'h38173851),
	.w8(32'h38a50f54),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378a7245),
	.w1(32'h37d05e7a),
	.w2(32'h386501ed),
	.w3(32'hb7e90324),
	.w4(32'h363c6d04),
	.w5(32'h3814e4f5),
	.w6(32'h382abeb2),
	.w7(32'h382086da),
	.w8(32'h3881053b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847af1f),
	.w1(32'hb800b858),
	.w2(32'hb903ceb2),
	.w3(32'hb9f35df8),
	.w4(32'hb9b3b188),
	.w5(32'h382f5f4e),
	.w6(32'hb9188c70),
	.w7(32'hba580404),
	.w8(32'hba28728b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c2cbf),
	.w1(32'hb8877d5f),
	.w2(32'hb87bc108),
	.w3(32'h3917ebef),
	.w4(32'h38c5bcf7),
	.w5(32'hb8b179f3),
	.w6(32'h396d5c75),
	.w7(32'h38720ca7),
	.w8(32'hb91ca156),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad36d7b),
	.w1(32'hbb3441cf),
	.w2(32'hba18e405),
	.w3(32'hbabaf18a),
	.w4(32'hbb0d0b2b),
	.w5(32'h39a915c1),
	.w6(32'hba93a150),
	.w7(32'hbb0fb369),
	.w8(32'hba4afdbb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d69f5),
	.w1(32'hbb274812),
	.w2(32'hba148f0a),
	.w3(32'hbb4b94a1),
	.w4(32'hbbafd05e),
	.w5(32'hb714e77c),
	.w6(32'hbac6ec9f),
	.w7(32'hbb4c2ced),
	.w8(32'hbaa5f7d3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030445),
	.w1(32'h3971e302),
	.w2(32'hb8ac75a0),
	.w3(32'hbb05a9cc),
	.w4(32'h3a068b72),
	.w5(32'hba0d6791),
	.w6(32'hb9f3ef8a),
	.w7(32'h3aca4dcb),
	.w8(32'h3a456b24),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0b629),
	.w1(32'hba658403),
	.w2(32'hba30321c),
	.w3(32'hbae6b967),
	.w4(32'hba8e2b0a),
	.w5(32'hba4d2961),
	.w6(32'hbac00e42),
	.w7(32'hbaab1e46),
	.w8(32'hbaa357ab),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb095fb6),
	.w1(32'hbadd1fe9),
	.w2(32'h3a2a5089),
	.w3(32'hba4b1d29),
	.w4(32'hba2982c2),
	.w5(32'h3a83fd09),
	.w6(32'hba0d8c9b),
	.w7(32'hba03a0b4),
	.w8(32'hb951d4c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad13cfd),
	.w1(32'hb96c1028),
	.w2(32'hba290be9),
	.w3(32'hba4cf778),
	.w4(32'h3a101b57),
	.w5(32'hb999ce83),
	.w6(32'hba646f73),
	.w7(32'h3807b16d),
	.w8(32'hb9987ca8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c81ccd),
	.w1(32'hb92c999d),
	.w2(32'h39668981),
	.w3(32'hbaacbb3d),
	.w4(32'hba589336),
	.w5(32'hb98981a7),
	.w6(32'hba86e27b),
	.w7(32'hbac021f3),
	.w8(32'hbabb649a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f02ddb),
	.w1(32'hb704149a),
	.w2(32'h36c2975f),
	.w3(32'hb6afc4e5),
	.w4(32'hb6873150),
	.w5(32'h3696c917),
	.w6(32'h37378079),
	.w7(32'h374b733a),
	.w8(32'h37a4631d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75133d6),
	.w1(32'hb713c3b2),
	.w2(32'h3710f66c),
	.w3(32'h36f6bfca),
	.w4(32'h34ec2130),
	.w5(32'hb7346e22),
	.w6(32'hb5f4c1c7),
	.w7(32'hb76d014a),
	.w8(32'hb7315398),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b42e7),
	.w1(32'h389e2594),
	.w2(32'h38d344cf),
	.w3(32'h38c59c3d),
	.w4(32'h38325d57),
	.w5(32'h384a787f),
	.w6(32'h39067dbe),
	.w7(32'h388ef0e4),
	.w8(32'h3895e57d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39228714),
	.w1(32'h368e639e),
	.w2(32'hb8b7b902),
	.w3(32'h3962d274),
	.w4(32'h38ec23d7),
	.w5(32'h3860959a),
	.w6(32'h397fa907),
	.w7(32'h384b76ae),
	.w8(32'h38c01370),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ed8c8),
	.w1(32'hbaa48d02),
	.w2(32'hbad41a2c),
	.w3(32'h3a57d25e),
	.w4(32'h3a773d38),
	.w5(32'h3a07d106),
	.w6(32'hb9f87dbc),
	.w7(32'hb7bcc5e0),
	.w8(32'h3a1f0f91),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997eb51),
	.w1(32'h390cc35b),
	.w2(32'h39c699a7),
	.w3(32'h38c02f36),
	.w4(32'h39783e57),
	.w5(32'h39751d4c),
	.w6(32'hb88788d0),
	.w7(32'hb807a970),
	.w8(32'h399558cf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb286ecf),
	.w1(32'hbb0e81bd),
	.w2(32'hba935e4c),
	.w3(32'hbafaed07),
	.w4(32'hba84c85f),
	.w5(32'hb9ea66e1),
	.w6(32'hb9d0b6dd),
	.w7(32'h3a56d9c3),
	.w8(32'hb901096a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc19b),
	.w1(32'hbb65f3b0),
	.w2(32'hba8dae4c),
	.w3(32'hbbc2974d),
	.w4(32'hbbb29100),
	.w5(32'hbac99557),
	.w6(32'hbbadc164),
	.w7(32'hbbd2c3c8),
	.w8(32'hbb55f6ba),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab97086),
	.w1(32'h3aaf86bf),
	.w2(32'h38eb3cbd),
	.w3(32'h3b23bfec),
	.w4(32'h3b248704),
	.w5(32'h3ada68f5),
	.w6(32'h3a682666),
	.w7(32'h3a5f396d),
	.w8(32'h3aa8dd76),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f47da),
	.w1(32'hb9a1d49b),
	.w2(32'h3add7972),
	.w3(32'hb93cc5be),
	.w4(32'h38d259ea),
	.w5(32'h3b50edc5),
	.w6(32'hbadb22f0),
	.w7(32'h3a9cfbd7),
	.w8(32'hbaa8cf10),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507c5c),
	.w1(32'h3a7690df),
	.w2(32'h391297a6),
	.w3(32'h3b19dc66),
	.w4(32'h3ade73af),
	.w5(32'hb9b68a7d),
	.w6(32'h3afa3c2a),
	.w7(32'h3a484ec0),
	.w8(32'hb9eafdce),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2e9f),
	.w1(32'hbb528044),
	.w2(32'hbb321148),
	.w3(32'hbb928ae9),
	.w4(32'hbb195637),
	.w5(32'h37308952),
	.w6(32'hbb79029c),
	.w7(32'hbb3dd6f4),
	.w8(32'hbae7af74),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c66c4),
	.w1(32'hb9d6e2ae),
	.w2(32'h3908cb2c),
	.w3(32'hb95a3799),
	.w4(32'h3a13122e),
	.w5(32'h3a83b3f3),
	.w6(32'h3991af02),
	.w7(32'h3a155277),
	.w8(32'hb96a1bf4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104e7a),
	.w1(32'hba6c0e18),
	.w2(32'hbb41f64a),
	.w3(32'h3981fc80),
	.w4(32'h3b111405),
	.w5(32'h38ef2d66),
	.w6(32'hb948e70f),
	.w7(32'h3a8a2011),
	.w8(32'h399dd0c7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c1971),
	.w1(32'h38b7da78),
	.w2(32'hba13949b),
	.w3(32'hb9d83ff0),
	.w4(32'hb8b923ae),
	.w5(32'hba5ace4b),
	.w6(32'hb9e49617),
	.w7(32'hb9e88123),
	.w8(32'hba804088),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8d92),
	.w1(32'h3a1447a7),
	.w2(32'h380f70f0),
	.w3(32'hbb58c470),
	.w4(32'hba0b3c62),
	.w5(32'hba9a4342),
	.w6(32'hbb1c269f),
	.w7(32'hbae29090),
	.w8(32'hbb3911ae),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb269a9f),
	.w1(32'hbafb988c),
	.w2(32'h3aa4b11d),
	.w3(32'h3ac1f034),
	.w4(32'h3a92fb56),
	.w5(32'h3b250945),
	.w6(32'h3aaffa7d),
	.w7(32'hb9e71820),
	.w8(32'hba616390),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fc4fb),
	.w1(32'hbb852b5b),
	.w2(32'hbab73128),
	.w3(32'h397c772f),
	.w4(32'hbbd69deb),
	.w5(32'hba3bc2f5),
	.w6(32'h399f088b),
	.w7(32'hbafe0319),
	.w8(32'hbabb81e2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319b6a),
	.w1(32'hbad64c43),
	.w2(32'hbb8c961d),
	.w3(32'h3b41da0b),
	.w4(32'h3bd53509),
	.w5(32'h3b104be7),
	.w6(32'hbad92079),
	.w7(32'h3ae871d1),
	.w8(32'hb960ccc1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6da5),
	.w1(32'h3980984b),
	.w2(32'h389bacbc),
	.w3(32'hbb0e33a4),
	.w4(32'h39b4fb8f),
	.w5(32'hbac1b7b3),
	.w6(32'hba9e3fc8),
	.w7(32'h3aa86738),
	.w8(32'hba3a6b31),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcb350),
	.w1(32'hba8cb611),
	.w2(32'h3b06377d),
	.w3(32'h3b1100be),
	.w4(32'h3aad3de9),
	.w5(32'h3b358334),
	.w6(32'hb8882317),
	.w7(32'h3ad3a0d5),
	.w8(32'hbaf87e0e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf176c),
	.w1(32'hb9ade801),
	.w2(32'hba007630),
	.w3(32'hb8bf1ebe),
	.w4(32'h3a5d975d),
	.w5(32'h38ebef2a),
	.w6(32'h3a132b02),
	.w7(32'h3a8ad8e4),
	.w8(32'hb881d54c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e677),
	.w1(32'hbc145354),
	.w2(32'hbbc89375),
	.w3(32'hbb7487a0),
	.w4(32'hbbc0a68b),
	.w5(32'hbada6fec),
	.w6(32'hbb15a501),
	.w7(32'hbb3844ae),
	.w8(32'h395939aa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e10a98),
	.w1(32'hbabadc7c),
	.w2(32'hba222365),
	.w3(32'h3b170bfb),
	.w4(32'hba4415bf),
	.w5(32'hba13b07b),
	.w6(32'h3ac7ac25),
	.w7(32'h39d8c3c1),
	.w8(32'h3a4056b9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397884c7),
	.w1(32'h38b3dbe4),
	.w2(32'hb88da08e),
	.w3(32'h3975adc6),
	.w4(32'h3940c4f6),
	.w5(32'hb7c9b58f),
	.w6(32'h3991609a),
	.w7(32'h39034f0c),
	.w8(32'h363dc5db),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f1889),
	.w1(32'hb98ea667),
	.w2(32'hba2a2aff),
	.w3(32'hba543663),
	.w4(32'h3a0f1635),
	.w5(32'h3859d1d6),
	.w6(32'hbaeb3585),
	.w7(32'hb936e6b1),
	.w8(32'hb8a80ede),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba215425),
	.w1(32'h3ac38b23),
	.w2(32'h3b096bf6),
	.w3(32'hbacfc669),
	.w4(32'h3786059f),
	.w5(32'hba5403ef),
	.w6(32'hba933727),
	.w7(32'hb993c05c),
	.w8(32'hbabe04f0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c211a),
	.w1(32'h3955bae5),
	.w2(32'h39370a6c),
	.w3(32'hbad50cc4),
	.w4(32'h3a9e0f7d),
	.w5(32'hba4ad53a),
	.w6(32'hba833f1f),
	.w7(32'h3a8f439a),
	.w8(32'h39bfd009),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9f56e),
	.w1(32'h3aa0edca),
	.w2(32'hbb1062a3),
	.w3(32'h398d12fe),
	.w4(32'h3ac9e08e),
	.w5(32'hba668e84),
	.w6(32'hb8e26f1b),
	.w7(32'hb94172c6),
	.w8(32'hb9463d92),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ec7b),
	.w1(32'hbaaf1b64),
	.w2(32'hba929e2b),
	.w3(32'hba907e15),
	.w4(32'h3a344946),
	.w5(32'h387c54e9),
	.w6(32'hba23b721),
	.w7(32'hb92f0d2e),
	.w8(32'hba9eeecb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba674dce),
	.w1(32'hba5aff57),
	.w2(32'h3b0da7de),
	.w3(32'hbb2b06df),
	.w4(32'hbadf1ce3),
	.w5(32'h3ab38eb4),
	.w6(32'hb8dbe60b),
	.w7(32'h3b050bb8),
	.w8(32'h3b33b752),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e3664),
	.w1(32'h37e05590),
	.w2(32'hb8db4724),
	.w3(32'hbb727635),
	.w4(32'hba5b379c),
	.w5(32'h39850e3e),
	.w6(32'hbb56ab65),
	.w7(32'hba55b5dd),
	.w8(32'hbaa80989),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6348),
	.w1(32'h384266d0),
	.w2(32'h39bc23ea),
	.w3(32'hba9030c5),
	.w4(32'hb8005a85),
	.w5(32'hb9b1c85c),
	.w6(32'hb91fab46),
	.w7(32'h3a2b19ad),
	.w8(32'h38e18f8c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d36196),
	.w1(32'hb80e773e),
	.w2(32'hb7e5946a),
	.w3(32'hb8000445),
	.w4(32'hb73c55b4),
	.w5(32'hb5fad823),
	.w6(32'hb85c7a88),
	.w7(32'hb7da65c3),
	.w8(32'h37a8a0c8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95caa65),
	.w1(32'h378324de),
	.w2(32'hb8bdfc70),
	.w3(32'hb8f62e9f),
	.w4(32'h37d70d6a),
	.w5(32'h39314452),
	.w6(32'h3885bcf0),
	.w7(32'h3946af64),
	.w8(32'h380dd374),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f487a6),
	.w1(32'hb8499cb0),
	.w2(32'hb70951a6),
	.w3(32'h379ba2c7),
	.w4(32'hb8019172),
	.w5(32'hb81b81be),
	.w6(32'h3806363a),
	.w7(32'h3727ce4f),
	.w8(32'h37df4073),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1aa54),
	.w1(32'h3a3a4d45),
	.w2(32'h3a2e0da7),
	.w3(32'h39b6afaf),
	.w4(32'h3a1900cb),
	.w5(32'h3a300162),
	.w6(32'h393ac4e0),
	.w7(32'h39d4b9db),
	.w8(32'h38fc21ef),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb3b01),
	.w1(32'h39cae23c),
	.w2(32'h39e88cff),
	.w3(32'hba3d21f4),
	.w4(32'h3a295229),
	.w5(32'h393a75e5),
	.w6(32'hb905a7c7),
	.w7(32'h3a830549),
	.w8(32'hb759f81f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3855eb75),
	.w1(32'hb94ac4cc),
	.w2(32'hb8e4f69c),
	.w3(32'h380b4a26),
	.w4(32'h391b914b),
	.w5(32'h39582844),
	.w6(32'h38c42ccf),
	.w7(32'h39a6c43f),
	.w8(32'h38dc0137),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac241ef),
	.w1(32'hb98c1bb8),
	.w2(32'h3a5caafa),
	.w3(32'hbabc2637),
	.w4(32'hba93b173),
	.w5(32'h3a51131a),
	.w6(32'hba8050ac),
	.w7(32'hba8e09a4),
	.w8(32'hba16ab73),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2ee78),
	.w1(32'h3a1271c0),
	.w2(32'hbaeb16da),
	.w3(32'hb6dae3e3),
	.w4(32'h3b07f1b5),
	.w5(32'hba111162),
	.w6(32'hba45ebff),
	.w7(32'h397dd3c2),
	.w8(32'hbaca91ce),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca31e4),
	.w1(32'h388cb4c8),
	.w2(32'hb55c3815),
	.w3(32'h38198b9c),
	.w4(32'hb60bc24a),
	.w5(32'hb891d4db),
	.w6(32'h388f9057),
	.w7(32'hb769aeea),
	.w8(32'h371116c6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39891cc5),
	.w1(32'h398108be),
	.w2(32'h38ce1ae4),
	.w3(32'h39824b75),
	.w4(32'h393c8750),
	.w5(32'hb724742a),
	.w6(32'h3977fbf4),
	.w7(32'h38d6d947),
	.w8(32'hb8cd64d7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3816f114),
	.w1(32'h37bae2e3),
	.w2(32'h3803181b),
	.w3(32'h387a8f45),
	.w4(32'h382b0bc6),
	.w5(32'h38474b6f),
	.w6(32'h38be7c83),
	.w7(32'h387fe32e),
	.w8(32'h388556a7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a4c25),
	.w1(32'h39c2d396),
	.w2(32'h396f871a),
	.w3(32'h3989b981),
	.w4(32'h39b6773f),
	.w5(32'h38f4b245),
	.w6(32'h396b15d9),
	.w7(32'h3983a7a3),
	.w8(32'h382a1d8b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84c96f),
	.w1(32'h3a2b7937),
	.w2(32'h3ab53d57),
	.w3(32'hba835419),
	.w4(32'hbb786bc4),
	.w5(32'hbae28282),
	.w6(32'hbaaec797),
	.w7(32'h3a146ef5),
	.w8(32'hba4bcaaa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf193e9),
	.w1(32'hb9ce5b80),
	.w2(32'h3923541a),
	.w3(32'hbb55af09),
	.w4(32'hbad15c9e),
	.w5(32'hb9f7e357),
	.w6(32'hbacf0cc3),
	.w7(32'hbaa6fb1c),
	.w8(32'hbaa33198),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910bbe9),
	.w1(32'hb98b1df4),
	.w2(32'hb8fe4583),
	.w3(32'hb942850a),
	.w4(32'hb974f2a1),
	.w5(32'h38efbb14),
	.w6(32'hb9d78803),
	.w7(32'hb9c24edd),
	.w8(32'hb9956cd8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084827),
	.w1(32'hbaabcd85),
	.w2(32'hb9f6bda9),
	.w3(32'hbaa11e99),
	.w4(32'hba9f6f9f),
	.w5(32'h39d700e2),
	.w6(32'hb9c1efb0),
	.w7(32'hb8a45e59),
	.w8(32'h3a018bc1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba151b62),
	.w1(32'hb94bf4c6),
	.w2(32'hb99b582f),
	.w3(32'hb971e045),
	.w4(32'hb8e7ba39),
	.w5(32'hb892b718),
	.w6(32'h3821c116),
	.w7(32'hb8b12e26),
	.w8(32'h38876864),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf9d89),
	.w1(32'hb98d55d0),
	.w2(32'h392aa1fe),
	.w3(32'hbaedf60f),
	.w4(32'hba680292),
	.w5(32'hb8d55fb4),
	.w6(32'hba7c6618),
	.w7(32'hba1df973),
	.w8(32'h390ff63b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032841),
	.w1(32'hb99a0ced),
	.w2(32'hba8d6f7a),
	.w3(32'hba6c06b4),
	.w4(32'h3a4db485),
	.w5(32'h39a0035b),
	.w6(32'hb76f3eda),
	.w7(32'h393c8216),
	.w8(32'hb983d844),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8258),
	.w1(32'hbaa6448e),
	.w2(32'hb973e408),
	.w3(32'hbb51245f),
	.w4(32'hbad2cf49),
	.w5(32'hb8b28093),
	.w6(32'hbb8dd533),
	.w7(32'hbb7d56ad),
	.w8(32'hbb39eefc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8f011),
	.w1(32'hba0a8e38),
	.w2(32'hba51e5e3),
	.w3(32'hb9be0f24),
	.w4(32'h3a2a3339),
	.w5(32'hba0fbcd4),
	.w6(32'hba12fbb9),
	.w7(32'h3a2925f1),
	.w8(32'hb916b696),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5caad0),
	.w1(32'hba9899b5),
	.w2(32'hba8439d7),
	.w3(32'hbb07dc25),
	.w4(32'hb8e3a55d),
	.w5(32'h39c55cc7),
	.w6(32'hbb0537c6),
	.w7(32'hb9b3a756),
	.w8(32'hbaa36f5a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f5eb),
	.w1(32'hbad07a4c),
	.w2(32'h39b3d2a3),
	.w3(32'hbb5395e2),
	.w4(32'hbaee33a1),
	.w5(32'h391d1a35),
	.w6(32'hbb2b8c79),
	.w7(32'hbaf17409),
	.w8(32'hbaba1218),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffd22b),
	.w1(32'hba96aa30),
	.w2(32'hb9537355),
	.w3(32'hba9c7bcb),
	.w4(32'hba0c9100),
	.w5(32'hb8499844),
	.w6(32'hba3db890),
	.w7(32'h3a797127),
	.w8(32'h3a86d9cc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044940),
	.w1(32'hb99cf0c8),
	.w2(32'h3a169e5e),
	.w3(32'hbacfed95),
	.w4(32'hb98b4d50),
	.w5(32'hb83cbb1b),
	.w6(32'hbaa4a7a7),
	.w7(32'hb8e6481b),
	.w8(32'hbab4718d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afa5a3),
	.w1(32'h388d50b9),
	.w2(32'h38f54b28),
	.w3(32'hb9a01155),
	.w4(32'h390530be),
	.w5(32'hb8cd4136),
	.w6(32'hb82ed34a),
	.w7(32'h39dc3699),
	.w8(32'h3842bace),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20bac7),
	.w1(32'hbafe3261),
	.w2(32'hbb3cf7ff),
	.w3(32'h39f93f28),
	.w4(32'h3b0c2c8d),
	.w5(32'hbb12a8da),
	.w6(32'h3a9afb84),
	.w7(32'h3ac514a2),
	.w8(32'hbafcfd40),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f671a),
	.w1(32'hba972361),
	.w2(32'hba778c35),
	.w3(32'hba9de9fe),
	.w4(32'hba0bee33),
	.w5(32'hba446d4a),
	.w6(32'hbab5f978),
	.w7(32'hba553184),
	.w8(32'hba3bda10),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb803cad4),
	.w1(32'hb8240d77),
	.w2(32'h375e3494),
	.w3(32'h37039870),
	.w4(32'hb7153940),
	.w5(32'h3811858f),
	.w6(32'h37ba0677),
	.w7(32'h3884a1d2),
	.w8(32'h384970c6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7140e85),
	.w1(32'hb84c1f6c),
	.w2(32'h371c7876),
	.w3(32'h382e4e78),
	.w4(32'h36d6ecec),
	.w5(32'h34ed363f),
	.w6(32'h3717bdc0),
	.w7(32'h368d4036),
	.w8(32'hb78dfd5c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e8391),
	.w1(32'hba06296f),
	.w2(32'hb9d57e5a),
	.w3(32'hb92025ef),
	.w4(32'hba35ab7a),
	.w5(32'hb9a4992c),
	.w6(32'h39b65999),
	.w7(32'h38c3ddcd),
	.w8(32'h39a41ef9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d8a7a),
	.w1(32'hbae3a0b8),
	.w2(32'hbb470fca),
	.w3(32'hba0519e9),
	.w4(32'hb9128570),
	.w5(32'hba89afe5),
	.w6(32'hbb1d4c0b),
	.w7(32'hbb096acf),
	.w8(32'hbb044737),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3651),
	.w1(32'h3a0535ee),
	.w2(32'h3ae763b9),
	.w3(32'hbacbeeb6),
	.w4(32'hba70407e),
	.w5(32'hb5f86558),
	.w6(32'h3a8ae8b8),
	.w7(32'h3a32d5b4),
	.w8(32'h37a1d5ec),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85de359),
	.w1(32'hb77b0eff),
	.w2(32'hb7ce8e91),
	.w3(32'hb83e72c0),
	.w4(32'hb7c08c1d),
	.w5(32'hb80fd7f8),
	.w6(32'hb6ffc57b),
	.w7(32'hb7f060b7),
	.w8(32'hb7fdf40b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf77a12),
	.w1(32'hb9f0a1ee),
	.w2(32'h3a42d890),
	.w3(32'hba92e151),
	.w4(32'hba217cce),
	.w5(32'hba1fed9c),
	.w6(32'hba964a49),
	.w7(32'hba55c552),
	.w8(32'hbaba0854),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d20bbb),
	.w1(32'h3946b443),
	.w2(32'h39844ed2),
	.w3(32'hb9314bb4),
	.w4(32'hb9f10efb),
	.w5(32'hbad54ceb),
	.w6(32'hbab40eee),
	.w7(32'hba44944b),
	.w8(32'hbb06d78e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144a61),
	.w1(32'h3992c70f),
	.w2(32'h3a41dec2),
	.w3(32'hba9c4e48),
	.w4(32'hba0f1a82),
	.w5(32'h3a494708),
	.w6(32'hbb3bef3d),
	.w7(32'hbb22424d),
	.w8(32'hbb13d81f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d813),
	.w1(32'h3a50d623),
	.w2(32'hbafa7209),
	.w3(32'h3ab779bc),
	.w4(32'h3b60b175),
	.w5(32'hba7279a3),
	.w6(32'h3a190a0e),
	.w7(32'h3a5398bf),
	.w8(32'hba01e12f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05220a),
	.w1(32'h393756b7),
	.w2(32'hba1f75cb),
	.w3(32'h3987f4d9),
	.w4(32'h3981d23e),
	.w5(32'hba2d2d3c),
	.w6(32'hb8ac2598),
	.w7(32'hb9f14e8c),
	.w8(32'hb9c850d6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63bdad),
	.w1(32'hba9a1cca),
	.w2(32'hb9aed82e),
	.w3(32'hb9c76eb9),
	.w4(32'h388a19f2),
	.w5(32'h3a578bbb),
	.w6(32'h3922e4b7),
	.w7(32'h39cba53a),
	.w8(32'h3a09d836),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad236a3),
	.w1(32'h39bf6d43),
	.w2(32'h3a55d096),
	.w3(32'hba6b1a89),
	.w4(32'h3a83eb1a),
	.w5(32'h39da4e73),
	.w6(32'hb9cc007b),
	.w7(32'h3aaea029),
	.w8(32'h39d0a3d8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef6182),
	.w1(32'hb993924a),
	.w2(32'hb9346a0c),
	.w3(32'h3aa0a964),
	.w4(32'h3a38e927),
	.w5(32'h3a4fcb4e),
	.w6(32'h3a078eb4),
	.w7(32'hbab51f27),
	.w8(32'hba37b475),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0cf07),
	.w1(32'h3aa4c6e6),
	.w2(32'h39d0bd3a),
	.w3(32'h3af66e27),
	.w4(32'h3ad7f739),
	.w5(32'h3a938fdf),
	.w6(32'h3a91057b),
	.w7(32'h3a511cec),
	.w8(32'h3a8ead61),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f12cd),
	.w1(32'hba211c81),
	.w2(32'h38b60f53),
	.w3(32'hb9cec43e),
	.w4(32'hb9be207a),
	.w5(32'h392298f9),
	.w6(32'hba2b2ea9),
	.w7(32'hba29eafc),
	.w8(32'hba188c0b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38979d2b),
	.w1(32'h3907acd3),
	.w2(32'h38686c4f),
	.w3(32'hb7271a6e),
	.w4(32'h3941af90),
	.w5(32'h38a0249b),
	.w6(32'hb90c2bfb),
	.w7(32'h3717dcf1),
	.w8(32'hb88af082),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8587),
	.w1(32'hba7be4d5),
	.w2(32'h37c49ffa),
	.w3(32'hbabe4ddc),
	.w4(32'hba87dedd),
	.w5(32'h39ea5055),
	.w6(32'hbafff4d0),
	.w7(32'hbad3a46a),
	.w8(32'hba0dc6eb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397db703),
	.w1(32'hb88ffddb),
	.w2(32'h36d367e2),
	.w3(32'h39a7b60e),
	.w4(32'h39110d7a),
	.w5(32'h39901f76),
	.w6(32'h38c7fd98),
	.w7(32'h39026948),
	.w8(32'h393a2a6f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30d27a),
	.w1(32'hb962d1ee),
	.w2(32'hba0dc79f),
	.w3(32'hbb17aaaa),
	.w4(32'h39061ed9),
	.w5(32'hba76bac8),
	.w6(32'hbade9e10),
	.w7(32'h3a99cea7),
	.w8(32'h39414065),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934d0fb),
	.w1(32'hb7ad346f),
	.w2(32'h38002e06),
	.w3(32'hb89f04a8),
	.w4(32'h381ad21b),
	.w5(32'h38ec7ff6),
	.w6(32'hb90ff3fa),
	.w7(32'h38ef02e0),
	.w8(32'h3930d98f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1f032),
	.w1(32'h3b05e324),
	.w2(32'h3ad6f341),
	.w3(32'h3b9ef323),
	.w4(32'h3a77c3d2),
	.w5(32'h3a5ea468),
	.w6(32'h3b85f550),
	.w7(32'h39452daa),
	.w8(32'hb9f8e8e9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c7e72),
	.w1(32'hb913a922),
	.w2(32'hb92cd66f),
	.w3(32'hb955e231),
	.w4(32'hb94977fc),
	.w5(32'hb9669b82),
	.w6(32'hb91ad7df),
	.w7(32'hb8c45f29),
	.w8(32'hb92e2832),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f506ed),
	.w1(32'hb99e810a),
	.w2(32'hb98b6d23),
	.w3(32'h39746f70),
	.w4(32'hb90aca27),
	.w5(32'hb9155f80),
	.w6(32'h3980a529),
	.w7(32'hb9057001),
	.w8(32'hb91efee2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacecdb0),
	.w1(32'hba8dcef6),
	.w2(32'hbaa09a5f),
	.w3(32'hb9a92141),
	.w4(32'h3ac0baaf),
	.w5(32'h39a11f97),
	.w6(32'hbadb4a54),
	.w7(32'h3a1bd72c),
	.w8(32'h39c6b197),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec288e),
	.w1(32'hb9d7e255),
	.w2(32'h3aa3265a),
	.w3(32'hbb0fa5fa),
	.w4(32'hbb034ef3),
	.w5(32'h39105f05),
	.w6(32'hbb583dce),
	.w7(32'hbb0612fb),
	.w8(32'hbb253fd7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8fe50),
	.w1(32'h3a75b593),
	.w2(32'h3a8a2fdb),
	.w3(32'h3aaed9a8),
	.w4(32'h3a117acf),
	.w5(32'h3a3c5da0),
	.w6(32'h3a9044a6),
	.w7(32'h3a08c52c),
	.w8(32'h3a735871),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73b16),
	.w1(32'h39f87378),
	.w2(32'hba61724d),
	.w3(32'hbabd9581),
	.w4(32'h3a1c71f0),
	.w5(32'hba64e276),
	.w6(32'h39c1c594),
	.w7(32'h3b0dea0c),
	.w8(32'hb985d296),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb806f),
	.w1(32'h3aa068c5),
	.w2(32'h399042e6),
	.w3(32'h36f9055f),
	.w4(32'h3a15ec2a),
	.w5(32'h39528bac),
	.w6(32'h395ac2cd),
	.w7(32'hb93de4a0),
	.w8(32'h39a1232f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805a8f),
	.w1(32'hb9886dc1),
	.w2(32'h3a994edd),
	.w3(32'hbb14c5b6),
	.w4(32'h3757700f),
	.w5(32'hb808ce8d),
	.w6(32'hba206895),
	.w7(32'h37f810df),
	.w8(32'hba2812f9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae13e5c),
	.w1(32'hbad68b3c),
	.w2(32'hbacc92fe),
	.w3(32'hba0dd6c0),
	.w4(32'hba90f135),
	.w5(32'hb9856946),
	.w6(32'hba917a97),
	.w7(32'hba9599ad),
	.w8(32'hba0489a7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67580f),
	.w1(32'hba1fdd27),
	.w2(32'h39e25f90),
	.w3(32'hbb6e6399),
	.w4(32'hba60820d),
	.w5(32'hb9e948b4),
	.w6(32'hbb2d4593),
	.w7(32'hba95aea4),
	.w8(32'hbb2f125c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e0c5c),
	.w1(32'hb91308b0),
	.w2(32'h38e871d3),
	.w3(32'hb91a110c),
	.w4(32'hb83f7474),
	.w5(32'h398a7f64),
	.w6(32'hb98c7bfe),
	.w7(32'h398cf471),
	.w8(32'h3a18db5d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058b94),
	.w1(32'hb9714233),
	.w2(32'hb9cbcbce),
	.w3(32'hbb0b211c),
	.w4(32'hba0a1933),
	.w5(32'h38721427),
	.w6(32'hbaf53a6b),
	.w7(32'hba621bf5),
	.w8(32'hba565826),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37854270),
	.w1(32'h37ce2dbf),
	.w2(32'h381d2ce4),
	.w3(32'h37ab12e3),
	.w4(32'h37312f3f),
	.w5(32'h37879ba3),
	.w6(32'h388c13c4),
	.w7(32'h382e2cf0),
	.w8(32'h380aacaf),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804ae02),
	.w1(32'h38433c9b),
	.w2(32'h398bc84b),
	.w3(32'h39029c56),
	.w4(32'h396cf51d),
	.w5(32'h39a14aa2),
	.w6(32'h39ab7aec),
	.w7(32'h397f7492),
	.w8(32'h39555caa),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ca74b),
	.w1(32'hb97a56a8),
	.w2(32'hb98a9c59),
	.w3(32'hb7861a67),
	.w4(32'h38803e77),
	.w5(32'hb934e65f),
	.w6(32'hb8f724a9),
	.w7(32'hb93065a3),
	.w8(32'hb98f392c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21e397),
	.w1(32'hb962f896),
	.w2(32'hb9f67794),
	.w3(32'hbb2b0f58),
	.w4(32'hbac8b30f),
	.w5(32'hb9f5b70e),
	.w6(32'hbb097974),
	.w7(32'hbac13c13),
	.w8(32'hba997093),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7344688),
	.w1(32'hb70b233a),
	.w2(32'h36b1b42a),
	.w3(32'hb73bb107),
	.w4(32'hb6d95fd9),
	.w5(32'h35e1414d),
	.w6(32'h349eb9eb),
	.w7(32'hb4e632ed),
	.w8(32'h36037e21),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984d166),
	.w1(32'hb94f34bb),
	.w2(32'hb837fb9f),
	.w3(32'hb953971c),
	.w4(32'hb7ffecb5),
	.w5(32'h376efe4d),
	.w6(32'hb93a01d1),
	.w7(32'hb87447af),
	.w8(32'hb82c4221),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a24b2),
	.w1(32'h39a136f7),
	.w2(32'h38fafd69),
	.w3(32'hba6b6561),
	.w4(32'h3938fe5f),
	.w5(32'h399006b2),
	.w6(32'hba688de6),
	.w7(32'h37c01c76),
	.w8(32'h399ae154),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6de34),
	.w1(32'hb98432dc),
	.w2(32'h3a38eafe),
	.w3(32'h3b274373),
	.w4(32'hb8eb9984),
	.w5(32'h3aa9beac),
	.w6(32'h3abbc755),
	.w7(32'hb986dbe7),
	.w8(32'hba2489a4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ace680),
	.w1(32'hba9e9615),
	.w2(32'h3911c976),
	.w3(32'h395f565b),
	.w4(32'h394e717e),
	.w5(32'h3ab93a1b),
	.w6(32'hba4dfe73),
	.w7(32'hb9f275a3),
	.w8(32'h38f27751),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c439e8),
	.w1(32'hba2efa68),
	.w2(32'hba010576),
	.w3(32'hb932d999),
	.w4(32'hb904a9f8),
	.w5(32'hb9e2821d),
	.w6(32'h3890c441),
	.w7(32'hb9b508c9),
	.w8(32'hb95dbfde),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9132e0),
	.w1(32'hbab37e10),
	.w2(32'h3ae92734),
	.w3(32'hbb9511cf),
	.w4(32'hbb89d7a3),
	.w5(32'hbb44f4fa),
	.w6(32'h3aa42d77),
	.w7(32'h3b01748b),
	.w8(32'hbb40424f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d149),
	.w1(32'h3a80fae0),
	.w2(32'hba29a8b7),
	.w3(32'hba3798b7),
	.w4(32'h3ba03446),
	.w5(32'h3ae022d2),
	.w6(32'hba82487d),
	.w7(32'h3996afff),
	.w8(32'hb8fce53e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac7089),
	.w1(32'hb9bf3dfd),
	.w2(32'h3a3c2da5),
	.w3(32'h391439c6),
	.w4(32'hb9d66ca8),
	.w5(32'h3a2f64a4),
	.w6(32'h389b676d),
	.w7(32'hb903d18b),
	.w8(32'h37c36237),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a44718),
	.w1(32'hb8700009),
	.w2(32'hb72802a8),
	.w3(32'hb84f45b2),
	.w4(32'hb83af23c),
	.w5(32'hb5a77d3e),
	.w6(32'h3782f148),
	.w7(32'hb745719d),
	.w8(32'hb725437c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e45893),
	.w1(32'hb9499e81),
	.w2(32'hb8313739),
	.w3(32'hb9276b95),
	.w4(32'h39bd911d),
	.w5(32'h38f533d9),
	.w6(32'h39806d22),
	.w7(32'h3a1f91a3),
	.w8(32'h395cbf03),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3816a0fb),
	.w1(32'h37b4b09c),
	.w2(32'h37da2daf),
	.w3(32'h37ff05e0),
	.w4(32'h36f150c1),
	.w5(32'h3710fdde),
	.w6(32'h3855fc23),
	.w7(32'h3788a4b1),
	.w8(32'h379b46ac),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e3160),
	.w1(32'h3a810780),
	.w2(32'h3a9e5102),
	.w3(32'h3a8c22ef),
	.w4(32'h3994abb8),
	.w5(32'h39d04ad0),
	.w6(32'h39868d6a),
	.w7(32'hb9814002),
	.w8(32'hba236411),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ccf36),
	.w1(32'hbae8d08d),
	.w2(32'hbac5bf9d),
	.w3(32'hba23afc1),
	.w4(32'hba3015f2),
	.w5(32'hb8a92d85),
	.w6(32'hba3e2916),
	.w7(32'hbae5a4db),
	.w8(32'hbab50639),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3b1ab),
	.w1(32'hba859ccb),
	.w2(32'hb9e81b3f),
	.w3(32'hb9854f69),
	.w4(32'h39199021),
	.w5(32'hb9d2659b),
	.w6(32'h3a29e6bf),
	.w7(32'h3acee5d3),
	.w8(32'h3a8e02e0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eff2a),
	.w1(32'hb9f9e8aa),
	.w2(32'h3735bda6),
	.w3(32'hb9b50cd1),
	.w4(32'hb920b96d),
	.w5(32'h39007fcc),
	.w6(32'hb9a2d95e),
	.w7(32'h39744f02),
	.w8(32'h393488c2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae68f1d),
	.w1(32'h3a28e825),
	.w2(32'h3a6a5b5f),
	.w3(32'hbaf91194),
	.w4(32'h37a26bd5),
	.w5(32'hba6b7fc3),
	.w6(32'hbabbf210),
	.w7(32'h399a8b30),
	.w8(32'hba1f58c4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981d9cc),
	.w1(32'hba12b1dc),
	.w2(32'hb8c36396),
	.w3(32'h390272dd),
	.w4(32'hb9d27d2a),
	.w5(32'h34d92058),
	.w6(32'h3a018c67),
	.w7(32'h3a232786),
	.w8(32'h392ba3a1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79eba5a),
	.w1(32'hb7902bfb),
	.w2(32'h37bbf516),
	.w3(32'hb79a0b25),
	.w4(32'hb730c683),
	.w5(32'h37f598aa),
	.w6(32'hb632334d),
	.w7(32'h36f1365e),
	.w8(32'h3837c634),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e4654),
	.w1(32'hbaa4282c),
	.w2(32'hb9eee0f6),
	.w3(32'hba863628),
	.w4(32'hba8bf54d),
	.w5(32'hb9e0af45),
	.w6(32'h398b5376),
	.w7(32'h39eecc86),
	.w8(32'hb8451403),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b6251),
	.w1(32'hb7a98c02),
	.w2(32'h3805a249),
	.w3(32'h3797d07c),
	.w4(32'hb7c9e884),
	.w5(32'h37fd74f4),
	.w6(32'h38a3c9ed),
	.w7(32'h37e5b6cc),
	.w8(32'h38b06dad),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918452c),
	.w1(32'h3aab9007),
	.w2(32'h39fc9d74),
	.w3(32'hba682662),
	.w4(32'h3a8658c3),
	.w5(32'hb987f4fc),
	.w6(32'hb889cdaa),
	.w7(32'h39f847fc),
	.w8(32'hba89f897),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a3870),
	.w1(32'hba3a556b),
	.w2(32'hbb088d13),
	.w3(32'h3a8dcd6c),
	.w4(32'h3ab451bd),
	.w5(32'h3a20f857),
	.w6(32'hb7d4e279),
	.w7(32'hb9e90b18),
	.w8(32'h3a278e14),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a09c0),
	.w1(32'hb8ee829d),
	.w2(32'hba1b27ba),
	.w3(32'hb9395afd),
	.w4(32'h39dde1f8),
	.w5(32'hb9a5d215),
	.w6(32'hb9c02424),
	.w7(32'h392ffa43),
	.w8(32'hb97462fe),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a0ce6),
	.w1(32'h3a1e533e),
	.w2(32'h398f03ce),
	.w3(32'h3a3d7283),
	.w4(32'h3a05f255),
	.w5(32'h396194b2),
	.w6(32'h38e24f09),
	.w7(32'h37e3aa21),
	.w8(32'h3916aeac),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84639b),
	.w1(32'h39605b94),
	.w2(32'hba379684),
	.w3(32'hb9d252c8),
	.w4(32'h3a8e263b),
	.w5(32'hb9e8c0b8),
	.w6(32'h394da581),
	.w7(32'h3a86ccc1),
	.w8(32'h3930483a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f573),
	.w1(32'hb9bc4c44),
	.w2(32'h3a1900a2),
	.w3(32'hbb1886a4),
	.w4(32'hba7b5af9),
	.w5(32'hb9932be9),
	.w6(32'hbaf7f00a),
	.w7(32'hb9ba2efa),
	.w8(32'hb9ccd6c9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa68e2a),
	.w1(32'hb94da700),
	.w2(32'h3aa5da28),
	.w3(32'hbb12ceea),
	.w4(32'hbab3678e),
	.w5(32'hb9931c78),
	.w6(32'hb97b64c3),
	.w7(32'h38f2173c),
	.w8(32'hb9c8a4be),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e05c65),
	.w1(32'h3797052e),
	.w2(32'h37fdc3ca),
	.w3(32'h3814144b),
	.w4(32'h388547ab),
	.w5(32'h38df3ca8),
	.w6(32'h38c9bdb8),
	.w7(32'h390355da),
	.w8(32'h3924f9e5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e4631b),
	.w1(32'h37dfa7a2),
	.w2(32'h37c99c19),
	.w3(32'hb917a3a6),
	.w4(32'hb8db6352),
	.w5(32'h37ecd526),
	.w6(32'h390edd28),
	.w7(32'hb6bb29eb),
	.w8(32'h37972bc9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15bf6a),
	.w1(32'hbabef478),
	.w2(32'h39cbaa46),
	.w3(32'h3a63b2be),
	.w4(32'hbacce903),
	.w5(32'h3a063195),
	.w6(32'h3a330943),
	.w7(32'h3a0f47d1),
	.w8(32'h3a9745a0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e75f3),
	.w1(32'hbaf5d9f8),
	.w2(32'hba5afc15),
	.w3(32'hbb191784),
	.w4(32'hbb03394d),
	.w5(32'hbad45562),
	.w6(32'hbb63a5e9),
	.w7(32'hbb04d0f9),
	.w8(32'hbb712fff),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28073),
	.w1(32'hba423b4e),
	.w2(32'h398d760e),
	.w3(32'hbaa8e5a8),
	.w4(32'hba66a528),
	.w5(32'hb960a4ab),
	.w6(32'hba776284),
	.w7(32'hb9c66cd2),
	.w8(32'hb8b4793c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e548),
	.w1(32'hba817757),
	.w2(32'h3aaf7e47),
	.w3(32'hba5526bd),
	.w4(32'h38639adc),
	.w5(32'h3b19d164),
	.w6(32'h39a65886),
	.w7(32'h3996330c),
	.w8(32'hb947e00b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908246d),
	.w1(32'hb889bd3d),
	.w2(32'hb6ae8dc9),
	.w3(32'hb92c15b1),
	.w4(32'hb8fbd57c),
	.w5(32'hb991d3eb),
	.w6(32'hb901c0df),
	.w7(32'hb7d9a6a4),
	.w8(32'hb937e9de),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fc9e5),
	.w1(32'hba4b1f74),
	.w2(32'hb928d0d4),
	.w3(32'hba4f574a),
	.w4(32'hba467388),
	.w5(32'hb984939a),
	.w6(32'hba1ca7f6),
	.w7(32'hb94f32ad),
	.w8(32'hb90abc86),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850ef0),
	.w1(32'h3a35f350),
	.w2(32'h3ac265be),
	.w3(32'h3b6be31c),
	.w4(32'hba902462),
	.w5(32'h3a35035b),
	.w6(32'h3a967523),
	.w7(32'h3a4dc735),
	.w8(32'hb8ae5dc9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836742),
	.w1(32'hbadf72fd),
	.w2(32'h37654d00),
	.w3(32'hbbcf5fd6),
	.w4(32'hbb994d57),
	.w5(32'hbaa1641d),
	.w6(32'hbb2d1935),
	.w7(32'hbb5eab0d),
	.w8(32'hbb06c235),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eef98),
	.w1(32'h398cd978),
	.w2(32'h3aacc719),
	.w3(32'h38a75a2a),
	.w4(32'hbb07e266),
	.w5(32'h3a892352),
	.w6(32'hba8f0b6a),
	.w7(32'hbaa28309),
	.w8(32'hbb04cc1d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecb8fe),
	.w1(32'h37235136),
	.w2(32'hbaa04d5b),
	.w3(32'h39b26535),
	.w4(32'h3a50eff8),
	.w5(32'hb9e220d8),
	.w6(32'h37b50c1c),
	.w7(32'h39964127),
	.w8(32'h3935ce1c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa8d6),
	.w1(32'hba02e2ef),
	.w2(32'hbaf1143e),
	.w3(32'hba847a61),
	.w4(32'h3abc8850),
	.w5(32'hb82a2873),
	.w6(32'hbaf0d687),
	.w7(32'hb80bbcd4),
	.w8(32'hb8c1562a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac97e8),
	.w1(32'h370e6865),
	.w2(32'h37c05c8c),
	.w3(32'h3774ce9c),
	.w4(32'h366476de),
	.w5(32'h37a3533e),
	.w6(32'h37d97bf6),
	.w7(32'h377153a6),
	.w8(32'h3803927a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375d1929),
	.w1(32'h373d8e0e),
	.w2(32'h37b1c57d),
	.w3(32'h377ea550),
	.w4(32'h37466c48),
	.w5(32'h37b5073b),
	.w6(32'h37d6ac6c),
	.w7(32'h37ad10c8),
	.w8(32'h380cade4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981033c),
	.w1(32'h3995b6d7),
	.w2(32'h3a26f8cb),
	.w3(32'hb95cc51a),
	.w4(32'h39d66579),
	.w5(32'hb8884942),
	.w6(32'hb9d429bc),
	.w7(32'hb9790ab4),
	.w8(32'hb9582b7f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb752b73d),
	.w1(32'hb7472fbe),
	.w2(32'h3781a1a6),
	.w3(32'hb7d99540),
	.w4(32'hb78d77ae),
	.w5(32'h3639d894),
	.w6(32'hb705db6f),
	.w7(32'h377dd648),
	.w8(32'h37bf0283),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0024f),
	.w1(32'h3a2d3f3d),
	.w2(32'h3993c3ce),
	.w3(32'h3a87bc54),
	.w4(32'h39c11bcd),
	.w5(32'h3a092e85),
	.w6(32'h39b3d200),
	.w7(32'h38ec2136),
	.w8(32'h3a0b77df),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5b9f),
	.w1(32'hbb434da2),
	.w2(32'hbaafb214),
	.w3(32'hbab40771),
	.w4(32'hbb19be2c),
	.w5(32'hbaf62139),
	.w6(32'hbb106ce6),
	.w7(32'hba8fbfdb),
	.w8(32'hbb426191),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba300623),
	.w1(32'hb7caf259),
	.w2(32'hb91cdabd),
	.w3(32'hba03c989),
	.w4(32'hb6be9d07),
	.w5(32'h383d6584),
	.w6(32'hba51313b),
	.w7(32'hb9015265),
	.w8(32'hb99fca93),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb2a09),
	.w1(32'h37ee440a),
	.w2(32'h384c951e),
	.w3(32'h3719a4a3),
	.w4(32'h37e80def),
	.w5(32'h382a6a91),
	.w6(32'h37b30110),
	.w7(32'h382db9c6),
	.w8(32'h38776bdf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6da71a),
	.w1(32'hb95ae5a5),
	.w2(32'h3af1171e),
	.w3(32'hbb014af6),
	.w4(32'hbb439e7a),
	.w5(32'h3b106981),
	.w6(32'hbaf434b8),
	.w7(32'hbb1d565c),
	.w8(32'hbb07b516),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba879e16),
	.w1(32'h388e1974),
	.w2(32'h3a6d82ff),
	.w3(32'hba919a48),
	.w4(32'hb92be276),
	.w5(32'h394bdad0),
	.w6(32'hba0addb8),
	.w7(32'hba1c148f),
	.w8(32'hba52caef),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cd229),
	.w1(32'h37b41007),
	.w2(32'h36abcb63),
	.w3(32'hb9166ca2),
	.w4(32'hb7e1d33f),
	.w5(32'hb81ea587),
	.w6(32'hb8bbbc10),
	.w7(32'hb801667b),
	.w8(32'hb89e5053),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaced8bd),
	.w1(32'hba483512),
	.w2(32'h39ad2dfb),
	.w3(32'hbb099243),
	.w4(32'hba88137c),
	.w5(32'h370b080c),
	.w6(32'hbadff370),
	.w7(32'hba75adb5),
	.w8(32'hba5bd9b0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39877fa7),
	.w1(32'h39948166),
	.w2(32'h39107e17),
	.w3(32'h398649be),
	.w4(32'h3983d953),
	.w5(32'h382e69aa),
	.w6(32'h395b332b),
	.w7(32'h39384aaa),
	.w8(32'hb6c3db22),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388215cc),
	.w1(32'h3908a64b),
	.w2(32'hb8daf6a8),
	.w3(32'h374d28e4),
	.w4(32'hb799477d),
	.w5(32'hb8cdf0b5),
	.w6(32'h37dc5697),
	.w7(32'h3833c5f8),
	.w8(32'hb96d7d0c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb625b21c),
	.w1(32'hb7097d46),
	.w2(32'hb6b2ef51),
	.w3(32'h3679c223),
	.w4(32'h37d2c1ae),
	.w5(32'h378e96ef),
	.w6(32'h37e8a6ad),
	.w7(32'h38235e78),
	.w8(32'h378f4119),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cabe3c),
	.w1(32'h37dc0d7a),
	.w2(32'h381a44f9),
	.w3(32'h389feafc),
	.w4(32'h3810379d),
	.w5(32'h374925e4),
	.w6(32'h381a1555),
	.w7(32'h38661582),
	.w8(32'h380bc13e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1ab14),
	.w1(32'h3a3b8901),
	.w2(32'h3a3e4183),
	.w3(32'h393d8b2f),
	.w4(32'h3a056baf),
	.w5(32'h3a19ea2c),
	.w6(32'hb913bd1f),
	.w7(32'h39550d57),
	.w8(32'h3a535719),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389ab2),
	.w1(32'h3a6c7303),
	.w2(32'h3abdd47e),
	.w3(32'hbae835fc),
	.w4(32'h3a398a20),
	.w5(32'h392f513e),
	.w6(32'hbb5af64b),
	.w7(32'hbad60a3f),
	.w8(32'hba7b8560),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530238),
	.w1(32'hbab0993c),
	.w2(32'hb96d5496),
	.w3(32'hbb5187eb),
	.w4(32'hbaafe108),
	.w5(32'h38a13d1a),
	.w6(32'hbafd989a),
	.w7(32'hba4a1c43),
	.w8(32'hba3ad396),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9b3f5),
	.w1(32'h398f7889),
	.w2(32'h3ae11cb2),
	.w3(32'hbb0c6d40),
	.w4(32'hb8dc3e88),
	.w5(32'h3a662fca),
	.w6(32'hbb1079b4),
	.w7(32'hbaa03240),
	.w8(32'hba053234),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f8d16),
	.w1(32'h39b1da7a),
	.w2(32'h399b9ec0),
	.w3(32'h398e439c),
	.w4(32'h39b89bad),
	.w5(32'h398ff763),
	.w6(32'h3985ae90),
	.w7(32'h39a27da3),
	.w8(32'h3997dce6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c62b2f),
	.w1(32'h384bbbb2),
	.w2(32'hb89a16f7),
	.w3(32'hb8467271),
	.w4(32'h37c890fe),
	.w5(32'hb7ae261e),
	.w6(32'h39112f80),
	.w7(32'h38999eac),
	.w8(32'h36c2c3b5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e0fb83),
	.w1(32'hb886eae5),
	.w2(32'hb7ffa5b9),
	.w3(32'hb83ef5ca),
	.w4(32'hb884effe),
	.w5(32'hb697be3c),
	.w6(32'hb7b0ecb9),
	.w7(32'hb8b06c49),
	.w8(32'hb77082b5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ec25c),
	.w1(32'hb776524e),
	.w2(32'hb7fcd407),
	.w3(32'h38627326),
	.w4(32'h37faff81),
	.w5(32'h37d8f05a),
	.w6(32'h38961367),
	.w7(32'h38683458),
	.w8(32'h387ddfd3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53eddd),
	.w1(32'hbadbb761),
	.w2(32'hbb2be8be),
	.w3(32'hbb88b39e),
	.w4(32'hbb245cc5),
	.w5(32'hbb0f011f),
	.w6(32'hbb1c7adf),
	.w7(32'hbb1595c9),
	.w8(32'hbb30248d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2e465),
	.w1(32'hb91ce6db),
	.w2(32'h3890a7d9),
	.w3(32'hb979f2fc),
	.w4(32'h38c7764e),
	.w5(32'h38a3ec09),
	.w6(32'hb88bf4c7),
	.w7(32'h388535ec),
	.w8(32'hb594c803),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dcbab),
	.w1(32'h39f452da),
	.w2(32'h3a300f5c),
	.w3(32'h3a92bf9c),
	.w4(32'h3a2ac42d),
	.w5(32'h3a440743),
	.w6(32'h39c15eb6),
	.w7(32'h39a91cb6),
	.w8(32'h3a0f72c8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39831d1b),
	.w1(32'hb8801a52),
	.w2(32'hb9cf29eb),
	.w3(32'h394b66ad),
	.w4(32'hb8f9abc4),
	.w5(32'h39acb4d8),
	.w6(32'h39aa65e0),
	.w7(32'h39786096),
	.w8(32'h39b226b6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0b68b),
	.w1(32'h388db9df),
	.w2(32'h37f0ca93),
	.w3(32'h3836ece8),
	.w4(32'h3904d025),
	.w5(32'h3400855b),
	.w6(32'h390df141),
	.w7(32'h38ba45f0),
	.w8(32'hb8260f39),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972fa5f),
	.w1(32'h398fe24d),
	.w2(32'h3988afcd),
	.w3(32'hb91b74cf),
	.w4(32'hb90ba2ad),
	.w5(32'hb932a80e),
	.w6(32'h392d0aa9),
	.w7(32'hb8d55b02),
	.w8(32'hba087469),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb834a12e),
	.w1(32'h3851edc6),
	.w2(32'hb8a42210),
	.w3(32'h390fcb65),
	.w4(32'hb76edd2f),
	.w5(32'hb83ad823),
	.w6(32'h399d612f),
	.w7(32'h390acfec),
	.w8(32'hb8f11cd3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb714fef),
	.w1(32'h3a45eafa),
	.w2(32'hbae4a426),
	.w3(32'hbb872af7),
	.w4(32'hb9a017f4),
	.w5(32'hb8e5b1b5),
	.w6(32'hbbb8a80d),
	.w7(32'hbb66d87c),
	.w8(32'hba17d033),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df03a8),
	.w1(32'hb91beabd),
	.w2(32'h39aa74b4),
	.w3(32'h389c5ce9),
	.w4(32'hb9973af0),
	.w5(32'h3a1fb557),
	.w6(32'hbac0a3b4),
	.w7(32'hb9ef7401),
	.w8(32'hbab2c379),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a6536),
	.w1(32'hbaa324b8),
	.w2(32'h3b39e4c8),
	.w3(32'hb9e42f21),
	.w4(32'hbb5190e2),
	.w5(32'h3a916127),
	.w6(32'hbae5a25b),
	.w7(32'h3b0c19dd),
	.w8(32'h394357cb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule