module layer_10_featuremap_186(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5079903),
	.w1(32'h357d3109),
	.w2(32'h3645965d),
	.w3(32'hb1b71d4a),
	.w4(32'h32cf4050),
	.w5(32'h33faa0e6),
	.w6(32'hb641d0c4),
	.w7(32'h360d4f22),
	.w8(32'h36a6f7b4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369f2d17),
	.w1(32'hb747e0d8),
	.w2(32'hb72d7755),
	.w3(32'h36fccdd5),
	.w4(32'h3700324c),
	.w5(32'h36844ef7),
	.w6(32'h383fd964),
	.w7(32'h3852a6d2),
	.w8(32'h38220a51),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34d10457),
	.w1(32'hb5997941),
	.w2(32'h34d29263),
	.w3(32'h3532a8b1),
	.w4(32'hb54e3c2c),
	.w5(32'h34aee31a),
	.w6(32'hb5c53391),
	.w7(32'hb42b8ed7),
	.w8(32'hb4295e10),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34daa6b8),
	.w1(32'hb60670c6),
	.w2(32'hb535f619),
	.w3(32'hb55165e2),
	.w4(32'h361ac954),
	.w5(32'hb568d78e),
	.w6(32'h36a9123f),
	.w7(32'h3561b4a4),
	.w8(32'hb629d34a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb49827f1),
	.w1(32'h3583656b),
	.w2(32'hb51ecd25),
	.w3(32'hb5873653),
	.w4(32'h351d5e07),
	.w5(32'hb61c3d2a),
	.w6(32'h36018159),
	.w7(32'hb19487b3),
	.w8(32'h34ae8b32),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5aedf03),
	.w1(32'h33fd249a),
	.w2(32'hb52a1a8b),
	.w3(32'hb647f206),
	.w4(32'h34bf4e64),
	.w5(32'hb492eb81),
	.w6(32'hb560f216),
	.w7(32'hb51a1bc2),
	.w8(32'hb4af1755),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da1bc8),
	.w1(32'h37cb3ccf),
	.w2(32'h37a28d65),
	.w3(32'h360ac3c2),
	.w4(32'hb6f0f2eb),
	.w5(32'h377a61b9),
	.w6(32'h36b3d100),
	.w7(32'hb657cc3d),
	.w8(32'h3745199b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e0e0b3),
	.w1(32'hb88825a1),
	.w2(32'hb8c5bb4d),
	.w3(32'hb803bf4e),
	.w4(32'hb810ac35),
	.w5(32'hb59f5062),
	.w6(32'hb8a2dc78),
	.w7(32'hb8be26ca),
	.w8(32'hb84f2e50),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3790107b),
	.w1(32'h37725618),
	.w2(32'h36b0a0bb),
	.w3(32'h3809443b),
	.w4(32'hb5d46869),
	.w5(32'hb79b581b),
	.w6(32'h3834509e),
	.w7(32'h383eba15),
	.w8(32'h37803bd7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38721f17),
	.w1(32'h3760c66f),
	.w2(32'hb5295fb2),
	.w3(32'h3685463b),
	.w4(32'hb8149754),
	.w5(32'hb876fbe2),
	.w6(32'hb804a479),
	.w7(32'hb74faafd),
	.w8(32'hb6cfac71),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bc5684),
	.w1(32'hb5975847),
	.w2(32'hb750b74d),
	.w3(32'h369b5f1f),
	.w4(32'h35a13467),
	.w5(32'hb6b63694),
	.w6(32'h36d15283),
	.w7(32'h36d951b8),
	.w8(32'h3701d9eb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372704ed),
	.w1(32'h373a6e4f),
	.w2(32'hb5bc2af4),
	.w3(32'hb72db933),
	.w4(32'hb763305e),
	.w5(32'hb808e7ce),
	.w6(32'h38193d05),
	.w7(32'h3723f219),
	.w8(32'hb6b8575e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c5dfc),
	.w1(32'h37f12d22),
	.w2(32'hb7bd70f4),
	.w3(32'hb73a7a73),
	.w4(32'hb7b1a644),
	.w5(32'hb85e5b0c),
	.w6(32'hb91027aa),
	.w7(32'hb915312b),
	.w8(32'hb8f387a0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b42467),
	.w1(32'h36689dfb),
	.w2(32'hb49ab3f7),
	.w3(32'h37086eb4),
	.w4(32'hb4f6ecd5),
	.w5(32'hb73ec47f),
	.w6(32'h37828432),
	.w7(32'h37318519),
	.w8(32'hb68a6788),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36aa84f1),
	.w1(32'h36c4f6e5),
	.w2(32'h375f02cc),
	.w3(32'h36ce75fc),
	.w4(32'h36f53379),
	.w5(32'hb68db263),
	.w6(32'h3840d8f9),
	.w7(32'h38055fae),
	.w8(32'h3804d4b5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f59362),
	.w1(32'hb8154a26),
	.w2(32'h369b2ab1),
	.w3(32'hb7c73863),
	.w4(32'hb7faa193),
	.w5(32'hb7e855a8),
	.w6(32'hb72b5d79),
	.w7(32'h36614b87),
	.w8(32'hb63093ee),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dd707c),
	.w1(32'h36506add),
	.w2(32'hb6215d2e),
	.w3(32'hb716867e),
	.w4(32'hb7d0c0f1),
	.w5(32'hb7e85e51),
	.w6(32'h36c63dad),
	.w7(32'h361c558d),
	.w8(32'h361cb2df),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383fe82f),
	.w1(32'h38337f41),
	.w2(32'h37b524fa),
	.w3(32'h380f4bc9),
	.w4(32'hb760b018),
	.w5(32'hb7de0730),
	.w6(32'hb8ad3b5d),
	.w7(32'hb85ff5dd),
	.w8(32'hb6bea97f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb601aa19),
	.w1(32'hb8147da9),
	.w2(32'hb74c25b2),
	.w3(32'h353a2fa7),
	.w4(32'hb8232805),
	.w5(32'hb83519fc),
	.w6(32'hb886d436),
	.w7(32'hb8834d2f),
	.w8(32'hb8675608),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb551b9aa),
	.w1(32'hb5645a33),
	.w2(32'hb464d9d5),
	.w3(32'hb5c0db7d),
	.w4(32'hb5084abd),
	.w5(32'h33ef9cb0),
	.w6(32'hb4f96b82),
	.w7(32'h3484c5f8),
	.w8(32'hb5409c52),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4870742),
	.w1(32'hb58df38c),
	.w2(32'hb5870a69),
	.w3(32'h34d935a7),
	.w4(32'h3552ec4e),
	.w5(32'h35b900ce),
	.w6(32'hb5ce9ac4),
	.w7(32'hb5b255ec),
	.w8(32'hb577386d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5685007),
	.w1(32'hb59d6158),
	.w2(32'hb63b7b91),
	.w3(32'hb4f58886),
	.w4(32'hb69e6959),
	.w5(32'hb70bdc46),
	.w6(32'hb65302cc),
	.w7(32'hb63a62a9),
	.w8(32'hb53ae228),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393610fe),
	.w1(32'h3846dfc7),
	.w2(32'h38fba36b),
	.w3(32'h391ce3db),
	.w4(32'hb812240e),
	.w5(32'h37e12232),
	.w6(32'h392aff52),
	.w7(32'h3931ffeb),
	.w8(32'h3927a22d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f78b6),
	.w1(32'h3717cbb9),
	.w2(32'hb577afd9),
	.w3(32'h37d4f34b),
	.w4(32'hb734802c),
	.w5(32'hb7925286),
	.w6(32'h38895526),
	.w7(32'h38851f49),
	.w8(32'h388f4d03),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c1b4e),
	.w1(32'h376caf72),
	.w2(32'h3778a9a6),
	.w3(32'h380a8175),
	.w4(32'h33119d12),
	.w5(32'hb749a5dc),
	.w6(32'h38474ea9),
	.w7(32'h3817be99),
	.w8(32'h3883dddb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6204213),
	.w1(32'hb5e3c2db),
	.w2(32'hb6986e1d),
	.w3(32'hb6e314f6),
	.w4(32'hb6697b81),
	.w5(32'hb5a1e9fd),
	.w6(32'hb5c5fd81),
	.w7(32'h34722955),
	.w8(32'hb6af74a4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb606f52c),
	.w1(32'hb5574cc9),
	.w2(32'hb51f0111),
	.w3(32'h36c74ef4),
	.w4(32'h35a0f799),
	.w5(32'h358b85f4),
	.w6(32'hb609657a),
	.w7(32'hb562178b),
	.w8(32'hb5c7ba72),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dc580c),
	.w1(32'hb6d5a681),
	.w2(32'hb709c13d),
	.w3(32'hb6fbe605),
	.w4(32'hb7119e1d),
	.w5(32'hb778a6ca),
	.w6(32'h36d81682),
	.w7(32'hb634c9d0),
	.w8(32'hb649759c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60f040c),
	.w1(32'h3679ad5d),
	.w2(32'h370336ec),
	.w3(32'h36de7e04),
	.w4(32'hb65434b3),
	.w5(32'hb6a3a741),
	.w6(32'h37741e0a),
	.w7(32'h3763bb7c),
	.w8(32'h3743db25),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37273380),
	.w1(32'hb74da5c1),
	.w2(32'hb7beef89),
	.w3(32'hb6dbcd7a),
	.w4(32'hb7fe99e2),
	.w5(32'hb827c097),
	.w6(32'h383d8b84),
	.w7(32'h381d9732),
	.w8(32'h37cbfaf3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3602b1d9),
	.w1(32'hb59f128a),
	.w2(32'hb5f35de8),
	.w3(32'h358c0b7e),
	.w4(32'hb5667f43),
	.w5(32'hb621daf0),
	.w6(32'hb519dde6),
	.w7(32'hb464ee2a),
	.w8(32'hb44e9206),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350d7c03),
	.w1(32'hb61512eb),
	.w2(32'hb587a9a2),
	.w3(32'hb5d754ec),
	.w4(32'hb70b131d),
	.w5(32'hb6fd69b1),
	.w6(32'h35992ef7),
	.w7(32'h3490c97b),
	.w8(32'h35e1c4ad),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d09276),
	.w1(32'h37305cea),
	.w2(32'h37472d25),
	.w3(32'h37c6bffc),
	.w4(32'h370d9e28),
	.w5(32'hb621538b),
	.w6(32'h37ad5e18),
	.w7(32'h37cfab5c),
	.w8(32'h37df8837),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36855cfc),
	.w1(32'h35bbe3bd),
	.w2(32'h370bb93d),
	.w3(32'h369c46c0),
	.w4(32'h3601b9d4),
	.w5(32'h36dee6cb),
	.w6(32'h37b5541b),
	.w7(32'h37f0b2ff),
	.w8(32'h37c474f6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360c8a94),
	.w1(32'hb4a834ea),
	.w2(32'hb3df5fc6),
	.w3(32'hb5e08200),
	.w4(32'hb6947937),
	.w5(32'hb66d2e47),
	.w6(32'hb642e555),
	.w7(32'hb352491e),
	.w8(32'hb58e6f38),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ba6c6),
	.w1(32'h362ac01f),
	.w2(32'h370bc228),
	.w3(32'h37503508),
	.w4(32'hb5b7ced7),
	.w5(32'h36132b73),
	.w6(32'hb80fec42),
	.w7(32'hb813b391),
	.w8(32'hb75c2bbc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827fb7b),
	.w1(32'h34284642),
	.w2(32'h3806bf70),
	.w3(32'h37eb4276),
	.w4(32'hb6c711f9),
	.w5(32'h381bc95f),
	.w6(32'h3753e179),
	.w7(32'h380cf303),
	.w8(32'h380c7b53),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e1cca5),
	.w1(32'hb787607d),
	.w2(32'hb806480e),
	.w3(32'h364d42e3),
	.w4(32'hb7d5f194),
	.w5(32'hb7fa9c6f),
	.w6(32'h3941fdee),
	.w7(32'h3940229e),
	.w8(32'h390d62ae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fe7fbd),
	.w1(32'h361910ec),
	.w2(32'h37a421fb),
	.w3(32'h37c223f1),
	.w4(32'h3788ca5a),
	.w5(32'h37bde123),
	.w6(32'h394061d1),
	.w7(32'h39316648),
	.w8(32'h3913b2e7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69b8bcb),
	.w1(32'hb743a81b),
	.w2(32'hb7f674c9),
	.w3(32'hb7a28f42),
	.w4(32'hb7ca0a49),
	.w5(32'hb82f6374),
	.w6(32'hb6cce21c),
	.w7(32'hb724a506),
	.w8(32'hb6d728ca),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4592ab9),
	.w1(32'hb62f9aa8),
	.w2(32'h363db1ee),
	.w3(32'hb6a014ad),
	.w4(32'hb6d379a5),
	.w5(32'hb6a62fc6),
	.w6(32'hb672f300),
	.w7(32'h356fec85),
	.w8(32'hb646e36b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h340e5485),
	.w1(32'hb4df9748),
	.w2(32'h354ef88f),
	.w3(32'h35ea1430),
	.w4(32'hb4db42af),
	.w5(32'h33234f6f),
	.w6(32'hb6391e2d),
	.w7(32'hb22a78c6),
	.w8(32'hb44f9a41),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57ed2a4),
	.w1(32'h35de63ef),
	.w2(32'hb76909ce),
	.w3(32'hb72326a3),
	.w4(32'hb7180a34),
	.w5(32'hb8003c6e),
	.w6(32'hb6884ccc),
	.w7(32'hb6867f5b),
	.w8(32'hb7661a88),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384fe9a7),
	.w1(32'hb5e84635),
	.w2(32'h38056ded),
	.w3(32'h37581406),
	.w4(32'hb852365c),
	.w5(32'hb883db5b),
	.w6(32'h379a842b),
	.w7(32'hb6b9bb6f),
	.w8(32'h3635a66e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c809ed),
	.w1(32'hb66a5188),
	.w2(32'hb6925b2a),
	.w3(32'h37929809),
	.w4(32'hb6dfc38d),
	.w5(32'hb77f86bc),
	.w6(32'h38b7b74d),
	.w7(32'h38995c11),
	.w8(32'h38947556),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c05d8),
	.w1(32'h37a99b47),
	.w2(32'h3610440a),
	.w3(32'h37e4fb8c),
	.w4(32'hb7ae9c54),
	.w5(32'hb7c894a4),
	.w6(32'h384e1cd9),
	.w7(32'h386b84a0),
	.w8(32'h3896e6d5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fc29d6),
	.w1(32'hb74d33fd),
	.w2(32'hb78fb2ff),
	.w3(32'h375c5ef3),
	.w4(32'hb3ee1db1),
	.w5(32'hb75a9dc5),
	.w6(32'h38cddd49),
	.w7(32'h3854859e),
	.w8(32'h38498b3a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38737e4c),
	.w1(32'hb75d733e),
	.w2(32'hb6f428f1),
	.w3(32'h36aa35a8),
	.w4(32'hb878f4cf),
	.w5(32'hb8982aed),
	.w6(32'hb903d802),
	.w7(32'hb8f2f382),
	.w8(32'hb8b64c75),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373e6c44),
	.w1(32'h360efebe),
	.w2(32'hb598574d),
	.w3(32'h36e37d6b),
	.w4(32'h35f48ad8),
	.w5(32'h3626428a),
	.w6(32'h36d3ecff),
	.w7(32'h369d1905),
	.w8(32'h35d0d9a2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb18e54c6),
	.w1(32'h330647a0),
	.w2(32'h36815ec3),
	.w3(32'h35c3a0e0),
	.w4(32'h357ec2ae),
	.w5(32'h3729e4f6),
	.w6(32'h37478b1e),
	.w7(32'h3756d5ff),
	.w8(32'h37765d93),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a68f7d),
	.w1(32'hb70714a7),
	.w2(32'hb6819a2a),
	.w3(32'hb4e91b8e),
	.w4(32'hb6e4b550),
	.w5(32'h363e92b0),
	.w6(32'h36a4203f),
	.w7(32'h369959fa),
	.w8(32'h36ca00b7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375bf17b),
	.w1(32'hb7052267),
	.w2(32'hb6928afa),
	.w3(32'h35c8684a),
	.w4(32'h37a96c23),
	.w5(32'hb7b1538e),
	.w6(32'hb683a1a3),
	.w7(32'hb78cf4d5),
	.w8(32'h37a1e297),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d6ed18),
	.w1(32'h3690c454),
	.w2(32'h360fe71a),
	.w3(32'h35d44673),
	.w4(32'hb62876c5),
	.w5(32'hb6ae8449),
	.w6(32'h373bf272),
	.w7(32'h3742e0c5),
	.w8(32'h375511dc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384ccd71),
	.w1(32'h381017c8),
	.w2(32'h387c34ac),
	.w3(32'h36ff0821),
	.w4(32'hb5f01f34),
	.w5(32'hb83af5e9),
	.w6(32'hb8148340),
	.w7(32'hb7fe9a57),
	.w8(32'h37b76500),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59dea37),
	.w1(32'hb66bf4bb),
	.w2(32'h3614309a),
	.w3(32'h368288c4),
	.w4(32'h34060577),
	.w5(32'h36136a86),
	.w6(32'h37a19785),
	.w7(32'h372c22eb),
	.w8(32'h374bee07),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b8b72a),
	.w1(32'hb65f66de),
	.w2(32'hb58d62a3),
	.w3(32'hb5abcc7c),
	.w4(32'hb66596f4),
	.w5(32'hb5945473),
	.w6(32'hb601fd1f),
	.w7(32'h34ae7726),
	.w8(32'hb65c101a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb611f3fe),
	.w1(32'h35c6f92c),
	.w2(32'h35e9c254),
	.w3(32'hb625703f),
	.w4(32'h347cfac5),
	.w5(32'h35e606ed),
	.w6(32'hb414f936),
	.w7(32'h35c5fbe3),
	.w8(32'h356ba32c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3392dfc0),
	.w1(32'hb52f0244),
	.w2(32'hb53d06cf),
	.w3(32'hb510a954),
	.w4(32'hb504d872),
	.w5(32'hb6ad3a90),
	.w6(32'hb4eb60cf),
	.w7(32'h34d2cb78),
	.w8(32'h351db33f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63124dd),
	.w1(32'hb6b96df9),
	.w2(32'hb7081bfb),
	.w3(32'hb6e82bf2),
	.w4(32'hb70b85bf),
	.w5(32'hb7259ca1),
	.w6(32'h378b426b),
	.w7(32'h3735d349),
	.w8(32'h372d7b3d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a0843b),
	.w1(32'hb64bfceb),
	.w2(32'hb6f0bb9a),
	.w3(32'hb70d93ca),
	.w4(32'hb6d5978c),
	.w5(32'hb74396b1),
	.w6(32'h362d3091),
	.w7(32'h361dc5d2),
	.w8(32'h352ec7bd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6936c38),
	.w1(32'hb5379c58),
	.w2(32'hb7e8794a),
	.w3(32'hb7957b7f),
	.w4(32'hb7c71a95),
	.w5(32'hb8256569),
	.w6(32'hb8787aca),
	.w7(32'hb897280a),
	.w8(32'hb8279ceb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3778cee6),
	.w1(32'h36300654),
	.w2(32'h37053154),
	.w3(32'h37496305),
	.w4(32'h369a6369),
	.w5(32'hb62e9a38),
	.w6(32'h377043fe),
	.w7(32'h37a6ab58),
	.w8(32'h37a216e9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3577656d),
	.w1(32'hb65418a6),
	.w2(32'hb3e73102),
	.w3(32'h34930ff5),
	.w4(32'hb62fc09f),
	.w5(32'hb5cbbaac),
	.w6(32'hb655be09),
	.w7(32'h358d0333),
	.w8(32'hb53eaa98),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d6ddf6),
	.w1(32'hb4736220),
	.w2(32'h34daaa6d),
	.w3(32'hb61dcb6c),
	.w4(32'hb51c3497),
	.w5(32'h35128a91),
	.w6(32'hb36d33e9),
	.w7(32'hb412bf17),
	.w8(32'hb514d7e6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350f7439),
	.w1(32'h355db480),
	.w2(32'hb2ec4762),
	.w3(32'h35be67ad),
	.w4(32'hb4d00adc),
	.w5(32'hb55785ad),
	.w6(32'h35e27d5d),
	.w7(32'h365e0f75),
	.w8(32'h36177cb5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359401b9),
	.w1(32'hb4fa8659),
	.w2(32'hb5d60a11),
	.w3(32'h3415a080),
	.w4(32'hb5821440),
	.w5(32'hb60b8ceb),
	.w6(32'hb5f08774),
	.w7(32'h345d0091),
	.w8(32'h340d6b67),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ae8c14),
	.w1(32'hb7b9de31),
	.w2(32'hb706d3ea),
	.w3(32'hb8059040),
	.w4(32'hb8577bf8),
	.w5(32'hb82e7435),
	.w6(32'hb7ab6b72),
	.w7(32'hb73d049e),
	.w8(32'hb69a405c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37022176),
	.w1(32'hb6f2d800),
	.w2(32'h381ae1db),
	.w3(32'h3777c02a),
	.w4(32'hb782c847),
	.w5(32'h37941d68),
	.w6(32'h38e8c569),
	.w7(32'h39094259),
	.w8(32'h390cd88a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3824ea1f),
	.w1(32'h37ba6ddc),
	.w2(32'h37f86f6d),
	.w3(32'h3842738e),
	.w4(32'h380f4f99),
	.w5(32'h380d8bc4),
	.w6(32'h38d14cd1),
	.w7(32'h38c172a1),
	.w8(32'h38d6f704),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f89fc),
	.w1(32'hb899ba0f),
	.w2(32'hb860f803),
	.w3(32'h365ccf3f),
	.w4(32'hb80ccefd),
	.w5(32'hb6757c58),
	.w6(32'h390ac6c8),
	.w7(32'h389c1a8a),
	.w8(32'h3888a517),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb28651da),
	.w1(32'hb3ff98bc),
	.w2(32'h34fe07a8),
	.w3(32'hb5ce466f),
	.w4(32'hb49108aa),
	.w5(32'h344bb3e2),
	.w6(32'hb5ed42b7),
	.w7(32'hb5396a04),
	.w8(32'hb5fc7d84),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4c45755),
	.w1(32'hb49a0a99),
	.w2(32'hb40b320e),
	.w3(32'hb523610d),
	.w4(32'h3509b1ef),
	.w5(32'h351baea1),
	.w6(32'hb673b6af),
	.w7(32'hb60b9ef7),
	.w8(32'hb5ea9257),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5487454),
	.w1(32'hb420508d),
	.w2(32'hb5646555),
	.w3(32'hb46d8d7d),
	.w4(32'hb48c49e0),
	.w5(32'hb525c84f),
	.w6(32'hb6930b62),
	.w7(32'hb631ccf7),
	.w8(32'hb66f540b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68e63b9),
	.w1(32'h3732cded),
	.w2(32'hb7132be4),
	.w3(32'hb71094f2),
	.w4(32'hb7366922),
	.w5(32'hb7c728a6),
	.w6(32'hb7bdd949),
	.w7(32'hb7a091e2),
	.w8(32'hb7b35bdc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b97bd2),
	.w1(32'hb60061fe),
	.w2(32'hb49e625b),
	.w3(32'hb445418d),
	.w4(32'hb5f9322f),
	.w5(32'h3601a368),
	.w6(32'hb655e304),
	.w7(32'hb5e00351),
	.w8(32'h34e117b9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dd38c7),
	.w1(32'h381c78ae),
	.w2(32'h381d2232),
	.w3(32'h371968e1),
	.w4(32'h363f57fd),
	.w5(32'hb7943b90),
	.w6(32'hb7d772bc),
	.w7(32'hb7c5ecc8),
	.w8(32'hb714766f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f9bbe),
	.w1(32'hb64f146f),
	.w2(32'hb75029a2),
	.w3(32'hb898514a),
	.w4(32'hb8819ebe),
	.w5(32'hb7bd4ae5),
	.w6(32'hb86064ec),
	.w7(32'hb8a778eb),
	.w8(32'hb8b59908),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810aebe),
	.w1(32'h375325b3),
	.w2(32'hb70605dd),
	.w3(32'hb72a887c),
	.w4(32'hb799548c),
	.w5(32'hb7e1f3d4),
	.w6(32'hb893f07f),
	.w7(32'hb8ab09aa),
	.w8(32'hb8a2d7b3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377931a0),
	.w1(32'h3719fe7f),
	.w2(32'h3768bc88),
	.w3(32'h3735d49a),
	.w4(32'h36c79560),
	.w5(32'h3671dbfb),
	.w6(32'h37d82e20),
	.w7(32'h37dad964),
	.w8(32'h37f79f6a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373eca06),
	.w1(32'h362731da),
	.w2(32'hb495f77f),
	.w3(32'h3632ff71),
	.w4(32'hb752d634),
	.w5(32'hb7538f75),
	.w6(32'hb4857ad6),
	.w7(32'h3710952b),
	.w8(32'h37324c3c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37382cf2),
	.w1(32'h363861e0),
	.w2(32'h3724c418),
	.w3(32'h3747ff0b),
	.w4(32'h35cbdc49),
	.w5(32'h364ae55b),
	.w6(32'h3808d18c),
	.w7(32'h38159e39),
	.w8(32'h37efa5ce),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807297c),
	.w1(32'h37990788),
	.w2(32'h37f54b17),
	.w3(32'h37887f78),
	.w4(32'h36d9e31e),
	.w5(32'hb70fd881),
	.w6(32'hb7c8b08d),
	.w7(32'hb7a71b62),
	.w8(32'hb7b3d45b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b5ff1f),
	.w1(32'hb5136350),
	.w2(32'hb531bfb9),
	.w3(32'hb62cb543),
	.w4(32'hb45f9e8f),
	.w5(32'hb581cf6a),
	.w6(32'hb54ebec4),
	.w7(32'h3334db4e),
	.w8(32'hb59f243d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fef5d2),
	.w1(32'h34c33347),
	.w2(32'h3498cf4e),
	.w3(32'hb60e0e3a),
	.w4(32'hb5b13ac0),
	.w5(32'hb48122e1),
	.w6(32'h3487c120),
	.w7(32'h35b0b48d),
	.w8(32'h35a6d851),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34afb6b5),
	.w1(32'hb6b72ca0),
	.w2(32'h353fd815),
	.w3(32'h344b063d),
	.w4(32'hb6f666c9),
	.w5(32'hb6005815),
	.w6(32'hb6d5518f),
	.w7(32'hb5b1db07),
	.w8(32'hb506aacd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c83b92),
	.w1(32'h3580c469),
	.w2(32'h35ad9e00),
	.w3(32'hb3df29a5),
	.w4(32'h350416b9),
	.w5(32'h359ca00a),
	.w6(32'h35391aa5),
	.w7(32'h3597ced6),
	.w8(32'hb48c992c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cea1d),
	.w1(32'hb6cdcb07),
	.w2(32'hb6f5886e),
	.w3(32'h366a48b8),
	.w4(32'h3727c4f5),
	.w5(32'h365422c1),
	.w6(32'h38ae434e),
	.w7(32'h38886778),
	.w8(32'h38263cd5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb633d11c),
	.w1(32'hb4ec3b1b),
	.w2(32'h358b6bba),
	.w3(32'hb656450d),
	.w4(32'hb682cbd7),
	.w5(32'hb605f831),
	.w6(32'h36f9a1ed),
	.w7(32'h365e0e12),
	.w8(32'h36593d0f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37176df1),
	.w1(32'hb668ac90),
	.w2(32'hb6ae8379),
	.w3(32'h37427b5e),
	.w4(32'h360f4890),
	.w5(32'hb618cb7a),
	.w6(32'h38387374),
	.w7(32'h38075ddb),
	.w8(32'h37ac8c6b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b8c3f4),
	.w1(32'h384a3f08),
	.w2(32'h384604fa),
	.w3(32'hb72dce4f),
	.w4(32'hb8077d44),
	.w5(32'h35b6e84b),
	.w6(32'hb7fade86),
	.w7(32'hb82c6715),
	.w8(32'h379def58),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366105f7),
	.w1(32'h36aaa150),
	.w2(32'h36a32886),
	.w3(32'h36b0ebe4),
	.w4(32'h35dab69c),
	.w5(32'h36852f30),
	.w6(32'h38803e03),
	.w7(32'h38427b3f),
	.w8(32'h3828e772),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5560a),
	.w1(32'h37507f08),
	.w2(32'h376d1537),
	.w3(32'h37b4fe8e),
	.w4(32'h35812482),
	.w5(32'h34f3628b),
	.w6(32'h382b486b),
	.w7(32'h37eadc7f),
	.w8(32'h3756bbc0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c29d4d),
	.w1(32'h361bbb7e),
	.w2(32'h35d3caac),
	.w3(32'h36f2fd55),
	.w4(32'h369a9bcc),
	.w5(32'h36e411f2),
	.w6(32'h3846390b),
	.w7(32'h3830c60d),
	.w8(32'h384c161f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bd1e52),
	.w1(32'hb5a9c496),
	.w2(32'hb817acf6),
	.w3(32'hb5927221),
	.w4(32'hb7205f89),
	.w5(32'hb8618cf3),
	.w6(32'h38b630bb),
	.w7(32'h3893ddf5),
	.w8(32'h3818ecff),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5e622),
	.w1(32'h3787f60a),
	.w2(32'h3751d5de),
	.w3(32'h37c91ffc),
	.w4(32'h36f687da),
	.w5(32'h37a91dbf),
	.w6(32'h387f6385),
	.w7(32'h386b92a0),
	.w8(32'h383f9cc1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68db45f),
	.w1(32'h37a63a61),
	.w2(32'h37057b50),
	.w3(32'h378ad6bc),
	.w4(32'hb6ab4b52),
	.w5(32'hb8155624),
	.w6(32'h3834bb46),
	.w7(32'h38543645),
	.w8(32'h388dc200),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36006386),
	.w1(32'hb5e4d6d9),
	.w2(32'h368f8595),
	.w3(32'h371f56b7),
	.w4(32'h36e659ab),
	.w5(32'h37639dc0),
	.w6(32'h364616a2),
	.w7(32'h377552da),
	.w8(32'h36f5f062),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380cd372),
	.w1(32'h37255f2d),
	.w2(32'hb6f516a9),
	.w3(32'h37e07e62),
	.w4(32'h3792881d),
	.w5(32'h367784f9),
	.w6(32'h37c5a31f),
	.w7(32'h380eb2b0),
	.w8(32'h3855ddee),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a8cc9),
	.w1(32'h3715e8c9),
	.w2(32'h37f4cdd8),
	.w3(32'h3800be6a),
	.w4(32'h378682d7),
	.w5(32'h37ae905b),
	.w6(32'h384ff865),
	.w7(32'h38808695),
	.w8(32'h3895e912),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38503907),
	.w1(32'h383c732f),
	.w2(32'h38a8af0b),
	.w3(32'h38267c10),
	.w4(32'h379797e6),
	.w5(32'h36c43a5f),
	.w6(32'hb7c1be38),
	.w7(32'hb7415160),
	.w8(32'h37f7fd24),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3702279c),
	.w1(32'h35d33da6),
	.w2(32'hb81084f9),
	.w3(32'h366aae90),
	.w4(32'h377d32fd),
	.w5(32'h37294741),
	.w6(32'h398289d5),
	.w7(32'h3971c501),
	.w8(32'h3930049c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c9c3e),
	.w1(32'h37932c5f),
	.w2(32'hb7910d38),
	.w3(32'h3753131c),
	.w4(32'hb70b7a48),
	.w5(32'hb81b857c),
	.w6(32'h38021504),
	.w7(32'h37ce6036),
	.w8(32'h37c71c4b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3721a8ce),
	.w1(32'hb665797b),
	.w2(32'hb5e3c3ab),
	.w3(32'h37940a69),
	.w4(32'h3555e476),
	.w5(32'hb6f38d42),
	.w6(32'h3869ede8),
	.w7(32'h3845cf2b),
	.w8(32'h3809ff81),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71a6e00),
	.w1(32'hb764d7a3),
	.w2(32'hb7470978),
	.w3(32'hb784035e),
	.w4(32'hb7c6d4ab),
	.w5(32'hb75471ec),
	.w6(32'h37266164),
	.w7(32'h3708b64c),
	.w8(32'h372aa8c8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383ac213),
	.w1(32'h37370f7e),
	.w2(32'h384ba6f3),
	.w3(32'h37abbd35),
	.w4(32'h371cc384),
	.w5(32'hb7117d61),
	.w6(32'hb73ff8ba),
	.w7(32'hb86991fa),
	.w8(32'hb847c8b2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370988d9),
	.w1(32'hb79bc919),
	.w2(32'h35d26eb6),
	.w3(32'hb7c902e0),
	.w4(32'hb79e337d),
	.w5(32'hb5ace0cb),
	.w6(32'hb71ce863),
	.w7(32'hb7fac343),
	.w8(32'hb7ff7b01),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b3f37d),
	.w1(32'hb5caf651),
	.w2(32'h34b0957c),
	.w3(32'h35f9b749),
	.w4(32'hb5e92b7a),
	.w5(32'hb5b51b99),
	.w6(32'h369fcc92),
	.w7(32'h369d0dbd),
	.w8(32'h3691b27a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35edc925),
	.w1(32'hb5c1a7e6),
	.w2(32'hb71a38f1),
	.w3(32'hb724db10),
	.w4(32'hb70939d6),
	.w5(32'hb746f2d9),
	.w6(32'h367197b0),
	.w7(32'h361505c0),
	.w8(32'h35e252c8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35df0031),
	.w1(32'hb71f0a21),
	.w2(32'hb766835e),
	.w3(32'hb6f3ee23),
	.w4(32'hb790935d),
	.w5(32'hb7fbb0db),
	.w6(32'hb81183b6),
	.w7(32'hb808915a),
	.w8(32'hb8301494),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f099fd),
	.w1(32'h37a90791),
	.w2(32'h3816e866),
	.w3(32'h381b9f23),
	.w4(32'h37d5a367),
	.w5(32'h3714bcb4),
	.w6(32'hb6b86762),
	.w7(32'h379fca5b),
	.w8(32'h3802da41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb834419a),
	.w1(32'hb80ddcd1),
	.w2(32'hb55ee60c),
	.w3(32'h369d1158),
	.w4(32'hb74829e0),
	.w5(32'hb6ca3d82),
	.w6(32'h3814b403),
	.w7(32'h383092c4),
	.w8(32'h38393abd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3753a817),
	.w1(32'hb794ec5d),
	.w2(32'h37e177c9),
	.w3(32'h37ac5776),
	.w4(32'h374683bb),
	.w5(32'h382a125d),
	.w6(32'h38a82141),
	.w7(32'h38a57de7),
	.w8(32'h38a4f9ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37054a83),
	.w1(32'h371aeaa7),
	.w2(32'h3722c138),
	.w3(32'h36c067ae),
	.w4(32'hb75ad11e),
	.w5(32'hb7139554),
	.w6(32'h37ae6f5f),
	.w7(32'h3642a1ed),
	.w8(32'h37151893),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f0e010),
	.w1(32'h372f16f6),
	.w2(32'h378c733d),
	.w3(32'h36e11128),
	.w4(32'hb6de0f9f),
	.w5(32'hb7caf4e9),
	.w6(32'h384528fa),
	.w7(32'h381285a8),
	.w8(32'h379bc1cb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a273c2),
	.w1(32'h35eba3c5),
	.w2(32'hb64c1959),
	.w3(32'h348dbe3c),
	.w4(32'hb447acd7),
	.w5(32'hb6c29aaa),
	.w6(32'h37f5a694),
	.w7(32'h37e17577),
	.w8(32'h37cd5faf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366f6f51),
	.w1(32'hb3b3dd40),
	.w2(32'hb4bc13b7),
	.w3(32'h365e16da),
	.w4(32'h350b874a),
	.w5(32'h3470504b),
	.w6(32'h3466f47e),
	.w7(32'h3574d1ca),
	.w8(32'hb4892d23),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb589269b),
	.w1(32'h3505e281),
	.w2(32'hb4856b7b),
	.w3(32'h33b8978c),
	.w4(32'h35746e20),
	.w5(32'h34a18ad7),
	.w6(32'h35ba21d3),
	.w7(32'h35d22e65),
	.w8(32'h359be215),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5914dda),
	.w1(32'h35926893),
	.w2(32'h36146f29),
	.w3(32'h34eb206b),
	.w4(32'h36059034),
	.w5(32'h359a4465),
	.w6(32'hb1af70ee),
	.w7(32'h34af5bad),
	.w8(32'h350f43ea),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b53b30),
	.w1(32'h344c0042),
	.w2(32'h365658f2),
	.w3(32'hb4ada93f),
	.w4(32'hb5933b20),
	.w5(32'h35681441),
	.w6(32'hb65b5094),
	.w7(32'hb5d05071),
	.w8(32'h3595cc46),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ddfd48),
	.w1(32'h351fe8b5),
	.w2(32'hb71e3b4e),
	.w3(32'h37a113a0),
	.w4(32'hb724a731),
	.w5(32'hb79f6e0d),
	.w6(32'h37d7e14a),
	.w7(32'h37974ff2),
	.w8(32'h37983502),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366399fe),
	.w1(32'h34e64811),
	.w2(32'h33fe39f5),
	.w3(32'h3669008a),
	.w4(32'h35923f34),
	.w5(32'hb2ad5010),
	.w6(32'h368d1c43),
	.w7(32'h3620b0ce),
	.w8(32'h3624ce3c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378224cd),
	.w1(32'h340f16c8),
	.w2(32'hb7c63e78),
	.w3(32'hb79cf1ce),
	.w4(32'hb76779ee),
	.w5(32'hb62b23f8),
	.w6(32'hb841228d),
	.w7(32'hb879d910),
	.w8(32'hb83d6030),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38312c74),
	.w1(32'h373ff86b),
	.w2(32'h380ef0c7),
	.w3(32'h3880009f),
	.w4(32'h383e3f5b),
	.w5(32'h37a547ee),
	.w6(32'h38669ab5),
	.w7(32'h3879bb83),
	.w8(32'h38b240a4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f88955),
	.w1(32'h36110f48),
	.w2(32'h36689c45),
	.w3(32'h33502bac),
	.w4(32'hb5fa7948),
	.w5(32'h3488a5a0),
	.w6(32'hb6a8cdc9),
	.w7(32'hb5433fb6),
	.w8(32'h360a87c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a2a589),
	.w1(32'hb62898ec),
	.w2(32'hb64288f1),
	.w3(32'h3576b4c4),
	.w4(32'hb58f3cdc),
	.w5(32'hb56800cb),
	.w6(32'hb57ecf6d),
	.w7(32'hb5e26326),
	.w8(32'hb563b266),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61791f4),
	.w1(32'hb5d1644e),
	.w2(32'hb62b8d87),
	.w3(32'hb65a12f8),
	.w4(32'hb6097a49),
	.w5(32'hb5b7bccc),
	.w6(32'hb5ebd434),
	.w7(32'hb5435d86),
	.w8(32'h34a87bb8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360f70dd),
	.w1(32'h3c02060d),
	.w2(32'h3c033032),
	.w3(32'hb576ffd7),
	.w4(32'h3c9f95d9),
	.w5(32'h3d014c22),
	.w6(32'hbc838437),
	.w7(32'hbc975ecd),
	.w8(32'hbc35ce9b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af06933),
	.w1(32'h3c111615),
	.w2(32'h3b8cb4a4),
	.w3(32'h3c4e0c3b),
	.w4(32'h3c285212),
	.w5(32'h3c971632),
	.w6(32'hbb55cf61),
	.w7(32'hbc572c3f),
	.w8(32'hbba0c594),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd7c44),
	.w1(32'hbb1307dc),
	.w2(32'h3c66569c),
	.w3(32'h3ba0f7f8),
	.w4(32'hbb16f531),
	.w5(32'hbb99a8cf),
	.w6(32'h3c56b17a),
	.w7(32'h3c008927),
	.w8(32'hbb17635c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90f44c),
	.w1(32'hbbc7862a),
	.w2(32'h3b5a3846),
	.w3(32'hbb151330),
	.w4(32'hbb684b9c),
	.w5(32'hbbf6accf),
	.w6(32'h395286e4),
	.w7(32'h3c2c64c3),
	.w8(32'hbb109f0d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf503a0),
	.w1(32'hbc150f25),
	.w2(32'hbb9cc193),
	.w3(32'hbb95f3b6),
	.w4(32'h379d494a),
	.w5(32'h3a03d010),
	.w6(32'hb9f57503),
	.w7(32'h3bf1609f),
	.w8(32'h3b544470),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904fc3),
	.w1(32'h3b43079a),
	.w2(32'hbb87b3c4),
	.w3(32'h3a380622),
	.w4(32'hbba23d18),
	.w5(32'hbb90841d),
	.w6(32'h3b18b5a5),
	.w7(32'h3b895f42),
	.w8(32'h3bd22d5a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad116e9),
	.w1(32'h3b4d64b0),
	.w2(32'hbbd45f18),
	.w3(32'hbb9d02c7),
	.w4(32'h3ba6d246),
	.w5(32'hba06df33),
	.w6(32'hb8489366),
	.w7(32'h3be70d15),
	.w8(32'h3c6bdb72),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3c3a),
	.w1(32'h3bc3d080),
	.w2(32'h3b140921),
	.w3(32'hbc097547),
	.w4(32'h3b321a93),
	.w5(32'h3c249059),
	.w6(32'hba88ba53),
	.w7(32'hbbcde01c),
	.w8(32'hba801e1f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b2b05),
	.w1(32'hbb2890f2),
	.w2(32'h3c02a351),
	.w3(32'hba8e8166),
	.w4(32'h3b731636),
	.w5(32'hb9bc5df3),
	.w6(32'h3b432040),
	.w7(32'h3c664dc2),
	.w8(32'h3aebe41e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b239bf7),
	.w1(32'h3c3a725f),
	.w2(32'h3a98c52a),
	.w3(32'hbb663196),
	.w4(32'h3ca89097),
	.w5(32'h3d007577),
	.w6(32'hbc7baca8),
	.w7(32'hbd014d3b),
	.w8(32'hbc9e8e3a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d4a11),
	.w1(32'h3bf063f6),
	.w2(32'h3b8c8529),
	.w3(32'h3c6a75f2),
	.w4(32'h3c12819f),
	.w5(32'h3c6816d4),
	.w6(32'hbb702af2),
	.w7(32'hbc216bf0),
	.w8(32'hbb12a4c3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6825),
	.w1(32'hbcabfaa2),
	.w2(32'hbaf175a4),
	.w3(32'h3b07b802),
	.w4(32'hbca0390e),
	.w5(32'hbcecf050),
	.w6(32'h3c1cc264),
	.w7(32'h3d22056e),
	.w8(32'h3c68974f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00737e),
	.w1(32'hbc832e84),
	.w2(32'hbca36a87),
	.w3(32'hbc6d7ada),
	.w4(32'h3a9e8341),
	.w5(32'h3b51372d),
	.w6(32'h390c5c69),
	.w7(32'hba6fcfae),
	.w8(32'h3b1701cc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82c89c),
	.w1(32'hbb01595f),
	.w2(32'hbbfc11b4),
	.w3(32'h3b58a6f6),
	.w4(32'h3b3e00d2),
	.w5(32'h3b167427),
	.w6(32'hbbfa2d94),
	.w7(32'hbc58b678),
	.w8(32'hbc2abcf8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41e1d5),
	.w1(32'h3b05f46f),
	.w2(32'hb9341436),
	.w3(32'hbbbebb84),
	.w4(32'h3c499953),
	.w5(32'h3c92898b),
	.w6(32'hbbf06846),
	.w7(32'hbc639738),
	.w8(32'hbc3ba38f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb9aff),
	.w1(32'h3c82802f),
	.w2(32'hba86cec8),
	.w3(32'h3bbe001a),
	.w4(32'h3d372c7e),
	.w5(32'h3d85a692),
	.w6(32'hbcfc5b48),
	.w7(32'hbd784925),
	.w8(32'hbd1d69a5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07bbd1),
	.w1(32'hbc3e736c),
	.w2(32'hbc9966d7),
	.w3(32'h3d229083),
	.w4(32'hbc50c811),
	.w5(32'hbc07d545),
	.w6(32'h3b05fc19),
	.w7(32'h3aab8df1),
	.w8(32'hbbd43622),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d7de),
	.w1(32'h3bfe4aa2),
	.w2(32'h3b5533f4),
	.w3(32'hbc37c0cd),
	.w4(32'h3b80843c),
	.w5(32'h3c0e184e),
	.w6(32'hba8b72bf),
	.w7(32'hbc111408),
	.w8(32'hbb65044f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e404),
	.w1(32'hbb79fef9),
	.w2(32'hbafd6955),
	.w3(32'hbb1dc30d),
	.w4(32'hbb8336d4),
	.w5(32'h3add5909),
	.w6(32'hbb685fcd),
	.w7(32'hbb9e2ac1),
	.w8(32'hbb2960c3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1d5fd),
	.w1(32'hbc95f975),
	.w2(32'hba94a481),
	.w3(32'hbbd43c62),
	.w4(32'hbc9981a1),
	.w5(32'hbccc8d45),
	.w6(32'h3ba09ad2),
	.w7(32'h3ccc445c),
	.w8(32'h3c098972),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ba05),
	.w1(32'hbb7328c8),
	.w2(32'hbaf612de),
	.w3(32'hbc7fa13d),
	.w4(32'hbb7365a1),
	.w5(32'hbbe1b7a5),
	.w6(32'h38a3353a),
	.w7(32'h3b8dfa06),
	.w8(32'hbb24e7e5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0a62),
	.w1(32'h3b570374),
	.w2(32'hb744c060),
	.w3(32'hbb9532f7),
	.w4(32'h3c00a875),
	.w5(32'h3c33f805),
	.w6(32'hbbd80bd1),
	.w7(32'hbc3f491d),
	.w8(32'hbbb13356),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907897),
	.w1(32'h3c324777),
	.w2(32'h3b18489e),
	.w3(32'hb75a616a),
	.w4(32'h3c6aae0d),
	.w5(32'h3cbf5375),
	.w6(32'hbc2de67f),
	.w7(32'hbcbc4140),
	.w8(32'hbc5e26ae),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e6a5),
	.w1(32'hbca10f9b),
	.w2(32'hbd06f0e0),
	.w3(32'h3c001013),
	.w4(32'h3ae99676),
	.w5(32'hbb6bc5ca),
	.w6(32'h3bd1a7c4),
	.w7(32'hbbcc1eac),
	.w8(32'hbb25dc7f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf64aee),
	.w1(32'h3b888498),
	.w2(32'h3bb4d875),
	.w3(32'hbbb2cf21),
	.w4(32'hb917d74f),
	.w5(32'h3b4fcd7f),
	.w6(32'h3aba80fe),
	.w7(32'h3b241087),
	.w8(32'hbaf62bea),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d7ae),
	.w1(32'h3c273c2a),
	.w2(32'h3b44db3e),
	.w3(32'hba291452),
	.w4(32'h3c9ec8fc),
	.w5(32'h3cfb72cb),
	.w6(32'hbc77949a),
	.w7(32'hbcfc6ba7),
	.w8(32'hbc996e26),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e53a),
	.w1(32'h3b7ecf13),
	.w2(32'h3bc166d5),
	.w3(32'h3c57148a),
	.w4(32'h3acbf141),
	.w5(32'hb61ce8c4),
	.w6(32'h3bc149b3),
	.w7(32'h3c0e1a92),
	.w8(32'h3b48abaf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867714),
	.w1(32'h3b8278e4),
	.w2(32'hbb501ece),
	.w3(32'hba61ce56),
	.w4(32'h39f8904b),
	.w5(32'h3a637d71),
	.w6(32'hbb97a08d),
	.w7(32'hbc507568),
	.w8(32'hbbd319f1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d047),
	.w1(32'h3b018ffd),
	.w2(32'h3982a3d8),
	.w3(32'hbaf4af9a),
	.w4(32'h3bc15bc7),
	.w5(32'h3c43ec81),
	.w6(32'hbc0e8d76),
	.w7(32'hbc8efc9f),
	.w8(32'hbc558c88),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc2ed5),
	.w1(32'hbb60ce33),
	.w2(32'h3b2a94e3),
	.w3(32'h3a002637),
	.w4(32'hbbac5582),
	.w5(32'hbbb72048),
	.w6(32'h3b1bef36),
	.w7(32'h3c388e43),
	.w8(32'h3b3dc4c4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb917fd),
	.w1(32'hbc123e70),
	.w2(32'h3b189acf),
	.w3(32'hbc0cc5aa),
	.w4(32'hbb90257b),
	.w5(32'h3c2f33f9),
	.w6(32'hbc3636e8),
	.w7(32'hbb074d0e),
	.w8(32'hbb6929bd),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6cd11),
	.w1(32'hbbd7aaa0),
	.w2(32'hbb577fcb),
	.w3(32'h3b0ee9c5),
	.w4(32'hbbcb6926),
	.w5(32'h3a69fb4f),
	.w6(32'hbbf1db76),
	.w7(32'hbb47da24),
	.w8(32'hbb4c0bf3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba858e),
	.w1(32'h3bb8b6b1),
	.w2(32'h3b5dc04f),
	.w3(32'h3b587800),
	.w4(32'h3c144d02),
	.w5(32'h3c74dc47),
	.w6(32'hbbedc36c),
	.w7(32'hbc644765),
	.w8(32'hbc348216),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb398949),
	.w1(32'h3b86afd2),
	.w2(32'h3b0fd024),
	.w3(32'h3b4de845),
	.w4(32'h3bf180c2),
	.w5(32'h3c5f8ce7),
	.w6(32'hbbc6c968),
	.w7(32'hbc79a6ac),
	.w8(32'hbc3bee20),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98172c),
	.w1(32'h3b8582f2),
	.w2(32'hbb488292),
	.w3(32'h3b73b752),
	.w4(32'h3c02a132),
	.w5(32'h3c457a67),
	.w6(32'hbb828c8f),
	.w7(32'hbc3f2614),
	.w8(32'hbc0e9e58),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b952),
	.w1(32'h3b402646),
	.w2(32'h3bcbcedd),
	.w3(32'h3c15ce57),
	.w4(32'h3bb334de),
	.w5(32'h3b8971b8),
	.w6(32'h3b7b494d),
	.w7(32'h3991bcad),
	.w8(32'hbbfb739f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da116),
	.w1(32'hbcaafb05),
	.w2(32'hbb34c7cd),
	.w3(32'h3a2876ef),
	.w4(32'hbce00ef9),
	.w5(32'hbd0e9f36),
	.w6(32'h3bba176b),
	.w7(32'h3cdda8ba),
	.w8(32'h3c09be43),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0e2ed),
	.w1(32'h3bd4c9d8),
	.w2(32'h3bcbc7eb),
	.w3(32'hbce011ae),
	.w4(32'h3ba1081e),
	.w5(32'h3c202025),
	.w6(32'hbb3c7c2e),
	.w7(32'hbc1b7fdf),
	.w8(32'hbc0da8e1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb11eb),
	.w1(32'hbc368bee),
	.w2(32'hbbcbf27d),
	.w3(32'h39befff1),
	.w4(32'hbc247f55),
	.w5(32'hbc9eb1c5),
	.w6(32'h3b0e2e0c),
	.w7(32'h3c30b043),
	.w8(32'hbac251a0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc165a51),
	.w1(32'hbbd28fc6),
	.w2(32'h3b707357),
	.w3(32'hbc9028bb),
	.w4(32'hbae6c0e8),
	.w5(32'hbb819a7f),
	.w6(32'hbac94d3f),
	.w7(32'h3c1ecd53),
	.w8(32'hbac7d5ab),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd4c52),
	.w1(32'h3c010f1b),
	.w2(32'h3b4268d1),
	.w3(32'hbb6e1317),
	.w4(32'h3c45859e),
	.w5(32'h3caf884d),
	.w6(32'hbc14920a),
	.w7(32'hbcaf9047),
	.w8(32'hbc4dec76),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bde2f),
	.w1(32'hbb6144ee),
	.w2(32'h3a023a81),
	.w3(32'h3bc0cd06),
	.w4(32'hb96086db),
	.w5(32'hbbadace0),
	.w6(32'hbb4ce7a4),
	.w7(32'h3b73aa3f),
	.w8(32'hbb9e79cf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12cbc1),
	.w1(32'hbb90dd9d),
	.w2(32'hbacfeac4),
	.w3(32'hbb9c106d),
	.w4(32'hbbad0fce),
	.w5(32'hb9ff9450),
	.w6(32'hbbef335f),
	.w7(32'hbb7f8da1),
	.w8(32'hba5a07dd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0a615),
	.w1(32'h39e7d194),
	.w2(32'h3b2e7695),
	.w3(32'h3b558b91),
	.w4(32'h3ae5c9fe),
	.w5(32'hbb452f32),
	.w6(32'h39638074),
	.w7(32'h3b169fcc),
	.w8(32'h3aaa236b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa11c),
	.w1(32'h3baf70ed),
	.w2(32'h3b68aeb6),
	.w3(32'hb763c3ac),
	.w4(32'h3c760066),
	.w5(32'h3cafb389),
	.w6(32'hbbdfea4a),
	.w7(32'hbc793278),
	.w8(32'hbc45f00b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f98d7),
	.w1(32'hbcd74597),
	.w2(32'h3a9e7f4b),
	.w3(32'h3c3df650),
	.w4(32'hbcbe7128),
	.w5(32'hbcd44d73),
	.w6(32'h3c900d23),
	.w7(32'h3d5b45d6),
	.w8(32'h3cae4f27),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c2524),
	.w1(32'h3a9eecf2),
	.w2(32'h3c36c9df),
	.w3(32'hbc0ea11b),
	.w4(32'h3c21f2d7),
	.w5(32'h3c3f7ade),
	.w6(32'h3ba0e3a7),
	.w7(32'h3bf9e909),
	.w8(32'hbb20e3d7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c36b),
	.w1(32'h3b75877d),
	.w2(32'h3bf4c335),
	.w3(32'h3c495fbe),
	.w4(32'h3bed48b0),
	.w5(32'h3be5109a),
	.w6(32'h3c154500),
	.w7(32'h3c398ed8),
	.w8(32'h3bb85e73),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a68c),
	.w1(32'hb8998ca1),
	.w2(32'hbc92422a),
	.w3(32'h3b886d78),
	.w4(32'h3bd0adc3),
	.w5(32'hbb9e0b23),
	.w6(32'h3b6466b2),
	.w7(32'hba9a6d5d),
	.w8(32'h3a0e75fc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd23d),
	.w1(32'hbb8ce2ad),
	.w2(32'h38c0f036),
	.w3(32'hbc41db55),
	.w4(32'hbb6d7da5),
	.w5(32'hb8ad1ed5),
	.w6(32'hbbad8c86),
	.w7(32'hbaedde26),
	.w8(32'hbabb858e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c7ac),
	.w1(32'h3b8480dd),
	.w2(32'h3aee8133),
	.w3(32'h3b21e205),
	.w4(32'h3c3de5b6),
	.w5(32'h3c7dd011),
	.w6(32'hbb9c050e),
	.w7(32'hbc545e51),
	.w8(32'hbc0dd028),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32cd83),
	.w1(32'h3c4824cd),
	.w2(32'h3aa481d2),
	.w3(32'h3bd80ff8),
	.w4(32'h3cbad8ab),
	.w5(32'h3d07f51a),
	.w6(32'hbc7d915d),
	.w7(32'hbd08a150),
	.w8(32'hbca73f4f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796265),
	.w1(32'h38d9733c),
	.w2(32'hbb0885fd),
	.w3(32'h3c85c1f8),
	.w4(32'h3c1ba088),
	.w5(32'h3b94a920),
	.w6(32'hba0a4f08),
	.w7(32'h3ad8ec8b),
	.w8(32'hbb31ee78),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a934a),
	.w1(32'h3b9e209c),
	.w2(32'h3bde974d),
	.w3(32'h3b1e1e20),
	.w4(32'h387205ab),
	.w5(32'hbb00a707),
	.w6(32'h3c0c8ee0),
	.w7(32'h3c45b2df),
	.w8(32'h39d5c70c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7be596),
	.w1(32'h3b93880f),
	.w2(32'h3b204d3f),
	.w3(32'hbbe7b2ea),
	.w4(32'h3b5370a2),
	.w5(32'h3bf8da1c),
	.w6(32'hbb7a9817),
	.w7(32'hbc6821ad),
	.w8(32'hbc4c79bf),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98d21),
	.w1(32'h3c201f0d),
	.w2(32'h3b92b1ef),
	.w3(32'hbb3521ae),
	.w4(32'h3b9fde7d),
	.w5(32'h39ead89d),
	.w6(32'h3c32d3a4),
	.w7(32'h3be4a88b),
	.w8(32'hbb5839ea),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b304451),
	.w1(32'hbb950744),
	.w2(32'hb952bbf8),
	.w3(32'hbb84ff55),
	.w4(32'hbbe939bb),
	.w5(32'hbc1b8890),
	.w6(32'h3b2b2247),
	.w7(32'h3c10e559),
	.w8(32'h3b27e3f6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b51b0),
	.w1(32'h3ac0799b),
	.w2(32'h3bc4830d),
	.w3(32'hbbb08613),
	.w4(32'hbb92fc13),
	.w5(32'h3b8764a1),
	.w6(32'hbae3f86b),
	.w7(32'h3ad893cd),
	.w8(32'h3aa1e6ca),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66af79),
	.w1(32'h3bb31d8a),
	.w2(32'h3bd0e71e),
	.w3(32'h3a45f3c4),
	.w4(32'h3c4ce6bd),
	.w5(32'h3c70849b),
	.w6(32'h3abc8d8e),
	.w7(32'hbb860d15),
	.w8(32'hbb2e2f50),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d1bd4),
	.w1(32'h3b69d3ac),
	.w2(32'hbc0fe4c5),
	.w3(32'h3c2b0326),
	.w4(32'h3ada62f6),
	.w5(32'h3bcf5f54),
	.w6(32'hbb98b730),
	.w7(32'hbc205184),
	.w8(32'hbc33540d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cc543),
	.w1(32'hbb931718),
	.w2(32'h3c04ef31),
	.w3(32'h3b73611a),
	.w4(32'h3a3a2f94),
	.w5(32'h39273347),
	.w6(32'h3b4854f4),
	.w7(32'h3c73e459),
	.w8(32'hbb02fdc6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81aa50),
	.w1(32'h3c0add9c),
	.w2(32'h3b5b9943),
	.w3(32'h3a05a0e5),
	.w4(32'h3c7723be),
	.w5(32'h3cc8ee25),
	.w6(32'hbc3a5562),
	.w7(32'hbccf59cd),
	.w8(32'hbc80dde0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb777a22),
	.w1(32'hbc26d1bf),
	.w2(32'hbb25ad1e),
	.w3(32'h3c0e97ba),
	.w4(32'hbb931156),
	.w5(32'hbc0a37c4),
	.w6(32'hbbd43782),
	.w7(32'h3b6320ac),
	.w8(32'hbb9bf15d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8272),
	.w1(32'h3b8dc956),
	.w2(32'hba404c02),
	.w3(32'hbb37ab4f),
	.w4(32'h3c76250b),
	.w5(32'h3ca1ed0c),
	.w6(32'hbc098a43),
	.w7(32'hbcaf3dd9),
	.w8(32'hbc4a837f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83c08),
	.w1(32'h3ae2bd7d),
	.w2(32'hbc1c88bb),
	.w3(32'h3be10085),
	.w4(32'h3c29fadf),
	.w5(32'h3b06630f),
	.w6(32'hbc0179ee),
	.w7(32'hbc0c0eaf),
	.w8(32'h3b05f850),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b825),
	.w1(32'hbc9ad8da),
	.w2(32'h3a4c3d70),
	.w3(32'h3aaf5a35),
	.w4(32'hbc95ac09),
	.w5(32'hbcb43fb6),
	.w6(32'h3c5aac60),
	.w7(32'h3d231c80),
	.w8(32'h3c8879f0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a296b),
	.w1(32'hbbaaece9),
	.w2(32'hbb4d8db5),
	.w3(32'hbc1a1bf6),
	.w4(32'hbb6ea059),
	.w5(32'hbbfa2a6a),
	.w6(32'h3b529a43),
	.w7(32'h3c077791),
	.w8(32'h3b982fdf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e737),
	.w1(32'h3c013c92),
	.w2(32'hbb6b2a9f),
	.w3(32'hbc195ba2),
	.w4(32'h3c1b0a53),
	.w5(32'h3c3f91b9),
	.w6(32'hbbb9f454),
	.w7(32'hbbde2d1b),
	.w8(32'hbbb72fa2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f2536),
	.w1(32'hbbe00c50),
	.w2(32'hbbe616e5),
	.w3(32'h3b94565b),
	.w4(32'hbc369bd4),
	.w5(32'hbc280469),
	.w6(32'hbbcbb8f5),
	.w7(32'hbb9aaf58),
	.w8(32'h3b171ae5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983b76e),
	.w1(32'h3a924da8),
	.w2(32'hb92e4f27),
	.w3(32'hba8e8b95),
	.w4(32'h3af7b49c),
	.w5(32'h3b75d8cb),
	.w6(32'hbac540b7),
	.w7(32'hba6b2b29),
	.w8(32'hbb4749da),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00737c),
	.w1(32'h3b8da10a),
	.w2(32'h3af2f09a),
	.w3(32'h3bafa7b4),
	.w4(32'hbaa98ab0),
	.w5(32'h3bed0875),
	.w6(32'hbb70b53a),
	.w7(32'hbc837fa5),
	.w8(32'hbc1e7c23),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae696),
	.w1(32'h3bcc0563),
	.w2(32'hbb506d23),
	.w3(32'hbb2e3d70),
	.w4(32'h3cb8a11c),
	.w5(32'h3c9dc0d7),
	.w6(32'hbbb389b7),
	.w7(32'hbbd0c0f0),
	.w8(32'hbb824451),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96ffae),
	.w1(32'hbc510f94),
	.w2(32'h3a2db38e),
	.w3(32'h3c4871db),
	.w4(32'hbc425443),
	.w5(32'hbc6fba3e),
	.w6(32'h3b1a21a0),
	.w7(32'h3c800c7f),
	.w8(32'h3b204af5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ec91),
	.w1(32'h3bb37bf0),
	.w2(32'h3aed15be),
	.w3(32'hbc23e3d2),
	.w4(32'h3c10c293),
	.w5(32'h3c9bd1f4),
	.w6(32'hbc32df85),
	.w7(32'hbcb533dd),
	.w8(32'hbc402c51),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512d91),
	.w1(32'h3bcd18b7),
	.w2(32'h3b33701e),
	.w3(32'h3b96fd9b),
	.w4(32'h3c30e58b),
	.w5(32'h3c9dd8a4),
	.w6(32'hbc12e8af),
	.w7(32'hbca5e6b6),
	.w8(32'hbc477958),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f99e0),
	.w1(32'h3b5d2ab5),
	.w2(32'h3b44f97c),
	.w3(32'h3bb0cdd2),
	.w4(32'h3b8c01ab),
	.w5(32'h3c59c0b1),
	.w6(32'hbbe4b28d),
	.w7(32'hbc92371e),
	.w8(32'hbc6d2bbe),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6e66),
	.w1(32'hbbc260db),
	.w2(32'hb96ce8e5),
	.w3(32'h3a8f8847),
	.w4(32'hbb7e07e8),
	.w5(32'hbbcf3aa9),
	.w6(32'hbaf9c527),
	.w7(32'h3ba84cc6),
	.w8(32'hbba49ff1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16cefb),
	.w1(32'h3b45e29e),
	.w2(32'hbaecb52d),
	.w3(32'hbbc62be8),
	.w4(32'h3c6028a0),
	.w5(32'h3c27e56c),
	.w6(32'hbc4c5c39),
	.w7(32'hbbdaf0ab),
	.w8(32'hbb6222e5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac769c7),
	.w1(32'h3c324d49),
	.w2(32'hba70e506),
	.w3(32'h3aae8595),
	.w4(32'h3cc81f62),
	.w5(32'h3d21f02d),
	.w6(32'hbc81c283),
	.w7(32'hbd07f4d4),
	.w8(32'hbc934410),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba76269),
	.w1(32'hba9e0118),
	.w2(32'h3a044e56),
	.w3(32'h3ca1cbce),
	.w4(32'hb9f22218),
	.w5(32'hbc17c9e9),
	.w6(32'h3a8624e2),
	.w7(32'h3bd9c560),
	.w8(32'hba92945d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adb95f),
	.w1(32'hb949d0d6),
	.w2(32'h3a45d073),
	.w3(32'hbb06575f),
	.w4(32'hbb6e739a),
	.w5(32'hbb3857d2),
	.w6(32'h3a3cdec0),
	.w7(32'h3ae2de82),
	.w8(32'h3a6676cb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b45d1),
	.w1(32'h3c138d22),
	.w2(32'h3bfa8de6),
	.w3(32'hbba2f903),
	.w4(32'h3c77ccbf),
	.w5(32'h3ce23e49),
	.w6(32'hbc6cfb8e),
	.w7(32'hbca84ba7),
	.w8(32'hbc47becb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7bd8a),
	.w1(32'h390dabad),
	.w2(32'h3b2f39c6),
	.w3(32'h3bf4fe1a),
	.w4(32'hbb2314c6),
	.w5(32'h3a9755ff),
	.w6(32'hbacb29db),
	.w7(32'h3a98be0e),
	.w8(32'hb9c401a8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b101ec9),
	.w1(32'h3b7894bf),
	.w2(32'h3c1e005a),
	.w3(32'h3b94b7d3),
	.w4(32'h3bbfa796),
	.w5(32'h374124d5),
	.w6(32'h3b684568),
	.w7(32'h3c025794),
	.w8(32'h3afdf1f9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd34bbd),
	.w1(32'h3b7f1a15),
	.w2(32'h3bac8734),
	.w3(32'h3aeed6c2),
	.w4(32'h3a27ee52),
	.w5(32'h3ad16d1e),
	.w6(32'h3adf6d11),
	.w7(32'h3b40e274),
	.w8(32'h39a9224e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c23d5),
	.w1(32'hbb222b29),
	.w2(32'h3bb27f41),
	.w3(32'h3b390f10),
	.w4(32'h3a933940),
	.w5(32'hbae07f76),
	.w6(32'hbb8f85d2),
	.w7(32'h3b339af5),
	.w8(32'hbc00f69e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f40d94),
	.w1(32'h382eafd3),
	.w2(32'hbba99304),
	.w3(32'hba0df9b9),
	.w4(32'hb914b161),
	.w5(32'hbb87c5e7),
	.w6(32'hba21cce5),
	.w7(32'hba864916),
	.w8(32'h3aaf9595),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83582d9),
	.w1(32'hbab0d235),
	.w2(32'h3ae735b9),
	.w3(32'hbb670afd),
	.w4(32'hba541286),
	.w5(32'h3a4e5adb),
	.w6(32'hbae28bb8),
	.w7(32'hbae44862),
	.w8(32'hbb48e2ae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acab9ba),
	.w1(32'h3ab24413),
	.w2(32'h3bfaab74),
	.w3(32'h3ba7e136),
	.w4(32'h3c4fe7b5),
	.w5(32'h3c74567a),
	.w6(32'hba36357e),
	.w7(32'hbb81e3a5),
	.w8(32'hbc11357f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b758dd),
	.w1(32'h3b98e6a9),
	.w2(32'h3b271724),
	.w3(32'h3c7a5d46),
	.w4(32'h3bab1bab),
	.w5(32'h3c3bdd4f),
	.w6(32'hbbcc87ab),
	.w7(32'hbc63dfe6),
	.w8(32'hbc22f4b2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb519c07),
	.w1(32'hba4e6b5a),
	.w2(32'h3bb768b6),
	.w3(32'h3ada1bb5),
	.w4(32'hbb32808d),
	.w5(32'hbafb1c2d),
	.w6(32'h3b58a5aa),
	.w7(32'h3c0a45d1),
	.w8(32'h3b221e4d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8159bf),
	.w1(32'h3c087fa3),
	.w2(32'h3b9c9259),
	.w3(32'hbaafa91c),
	.w4(32'h3c42c102),
	.w5(32'h3caeb843),
	.w6(32'hbc326154),
	.w7(32'hbcaee24f),
	.w8(32'hbc6899fa),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb531c60),
	.w1(32'h3b47adb0),
	.w2(32'hba07ba20),
	.w3(32'h3bdbdcec),
	.w4(32'h3c02168d),
	.w5(32'h3c4c7d65),
	.w6(32'hbbebd14d),
	.w7(32'hbc784934),
	.w8(32'hbc4e0111),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0fadb),
	.w1(32'hbc7109f3),
	.w2(32'hbb722ce1),
	.w3(32'h3b3a658f),
	.w4(32'hbc166cbd),
	.w5(32'hbc5f64d4),
	.w6(32'hbb155990),
	.w7(32'h3c48fb91),
	.w8(32'h3b6bf1ef),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9369cf),
	.w1(32'hbb8725a9),
	.w2(32'h3bca9731),
	.w3(32'hbbec7c5c),
	.w4(32'hbc29af9b),
	.w5(32'hbc489c5b),
	.w6(32'h3beca9bf),
	.w7(32'h3c67026c),
	.w8(32'h3bdfb44a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6e575),
	.w1(32'h3b903da1),
	.w2(32'h3c0c0579),
	.w3(32'hbc1425b5),
	.w4(32'h3a5aabde),
	.w5(32'h3c044027),
	.w6(32'h3b1b569b),
	.w7(32'h3bc8925d),
	.w8(32'hbb13dc3b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392382a7),
	.w1(32'hbc2d6cea),
	.w2(32'hbbd9bc30),
	.w3(32'h3b477f36),
	.w4(32'hbb9b55b1),
	.w5(32'hbbe816ba),
	.w6(32'hbbd355d5),
	.w7(32'hba05fa40),
	.w8(32'hbbb1afbb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1f0c9),
	.w1(32'h3bb2f5ae),
	.w2(32'h3ba01989),
	.w3(32'hbb8983dd),
	.w4(32'h3be5b4a6),
	.w5(32'h3bae304d),
	.w6(32'h3c5602f7),
	.w7(32'h3bab7e36),
	.w8(32'h3a7a12fd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75dd37),
	.w1(32'h3a95269a),
	.w2(32'h3b5b8cbd),
	.w3(32'h3aeb596a),
	.w4(32'hbb17c7dd),
	.w5(32'hbb7b5f21),
	.w6(32'hbb05052c),
	.w7(32'h3b149819),
	.w8(32'h3b14b5c8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d33ca),
	.w1(32'hb9b0b907),
	.w2(32'h3bc07af8),
	.w3(32'hbb53c7ab),
	.w4(32'h3a184624),
	.w5(32'h3b9bbc1d),
	.w6(32'h3b36f018),
	.w7(32'h3c0308b6),
	.w8(32'h3b69b957),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943a699),
	.w1(32'hbb15fb0d),
	.w2(32'h3b7fee19),
	.w3(32'h3bee5ff6),
	.w4(32'h3a5b24a0),
	.w5(32'hbbca79a6),
	.w6(32'hba774caa),
	.w7(32'h3b958cfd),
	.w8(32'hbbcc5400),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03bf7b),
	.w1(32'h3b1e3283),
	.w2(32'h3bf1f27a),
	.w3(32'hbbe68517),
	.w4(32'hbbd06933),
	.w5(32'hbb89c6bd),
	.w6(32'h3c0f8624),
	.w7(32'h3c50f57b),
	.w8(32'h3b85479c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ece39c),
	.w1(32'h391cd40a),
	.w2(32'hbab8e664),
	.w3(32'hbb977496),
	.w4(32'h3af7968a),
	.w5(32'h3c515c99),
	.w6(32'h3b31affd),
	.w7(32'h3abc5c71),
	.w8(32'hbbac211f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb19bf6),
	.w1(32'h3c6ec3a9),
	.w2(32'h3bf4705e),
	.w3(32'h3bc407ab),
	.w4(32'h3ba7bd4b),
	.w5(32'hb9a80bd0),
	.w6(32'h3b6abb3e),
	.w7(32'h3b911188),
	.w8(32'h3c760845),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2fcad),
	.w1(32'h3c8bad76),
	.w2(32'hba963a0a),
	.w3(32'hbbc3dfb4),
	.w4(32'h3d1a0a21),
	.w5(32'h3d783655),
	.w6(32'hbcc5c408),
	.w7(32'hbd4fce9d),
	.w8(32'hbce2f4f9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf41358),
	.w1(32'h3bb9c197),
	.w2(32'h3a9b871a),
	.w3(32'h3cfa84ab),
	.w4(32'h3baf2fd3),
	.w5(32'h3c911fb0),
	.w6(32'hbc3e9fbd),
	.w7(32'hbcbd04bb),
	.w8(32'hbc6d21b1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b0f9),
	.w1(32'h3beed9c2),
	.w2(32'hba50e76f),
	.w3(32'h3b452aaa),
	.w4(32'h3c8bcd5c),
	.w5(32'h3ce98d8a),
	.w6(32'hbc3f52b2),
	.w7(32'hbcc4a83a),
	.w8(32'hbc537881),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e8cd),
	.w1(32'h3bd8dbc8),
	.w2(32'h3b863fdf),
	.w3(32'h3c5f14c9),
	.w4(32'h3c3963d6),
	.w5(32'h3c872cff),
	.w6(32'hbbe7bcc4),
	.w7(32'hbc664422),
	.w8(32'hbc2cc40d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24aa7a),
	.w1(32'hbbf05018),
	.w2(32'hbbeeffe9),
	.w3(32'h3bb3e0fe),
	.w4(32'h3af64ace),
	.w5(32'hbb0c53a5),
	.w6(32'hbac06190),
	.w7(32'h3bb424ab),
	.w8(32'hbab7691c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb714ec),
	.w1(32'h3be4a3c7),
	.w2(32'h3a6644cc),
	.w3(32'hbb131d5d),
	.w4(32'h3c215f39),
	.w5(32'h3c82a92f),
	.w6(32'hbbe32b37),
	.w7(32'hbc9474ce),
	.w8(32'hbc6785da),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91cafa),
	.w1(32'h3c1b433c),
	.w2(32'hba1f49fd),
	.w3(32'h3baadd08),
	.w4(32'h3ca87084),
	.w5(32'h3d059848),
	.w6(32'hbc551bcd),
	.w7(32'hbce1a7fd),
	.w8(32'hbc73dace),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7117ea),
	.w1(32'h3ae73957),
	.w2(32'h3bfe58dc),
	.w3(32'h3c880ac8),
	.w4(32'h3ba55487),
	.w5(32'h3a1eaf8a),
	.w6(32'h3b88ebd1),
	.w7(32'h3c1ff85f),
	.w8(32'h3b1ddd70),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5001e8),
	.w1(32'h3bef1ec4),
	.w2(32'h3a98ae43),
	.w3(32'h3ba525a5),
	.w4(32'h3b9771b0),
	.w5(32'h3c02f269),
	.w6(32'hbb87ae44),
	.w7(32'hbc6538c0),
	.w8(32'hbc2756c2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c84c9),
	.w1(32'hbb8b4c61),
	.w2(32'hbba80a44),
	.w3(32'hbb120f49),
	.w4(32'h3b8eb64b),
	.w5(32'h3a177e7b),
	.w6(32'hbb7952a8),
	.w7(32'hbc087fcd),
	.w8(32'hbb4f75d4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac34ce3),
	.w1(32'h3becb443),
	.w2(32'h3b755d72),
	.w3(32'h3b35f10b),
	.w4(32'hbaa005ab),
	.w5(32'h3bccce1a),
	.w6(32'h3a30c274),
	.w7(32'hbbe82d76),
	.w8(32'hbbaf64a2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f4cd),
	.w1(32'hbbe15c4b),
	.w2(32'hbb5d0588),
	.w3(32'hbb9c9a5e),
	.w4(32'hba9cfb9f),
	.w5(32'hbbf01946),
	.w6(32'h3bb46b3c),
	.w7(32'h3c26aa6e),
	.w8(32'hba0c26ed),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdec17a),
	.w1(32'h3bc3e89e),
	.w2(32'h3affa2d2),
	.w3(32'hbbb73cc6),
	.w4(32'h3cd1292a),
	.w5(32'h3d133dac),
	.w6(32'hbc9f8de4),
	.w7(32'hbd0020b7),
	.w8(32'hbc93e693),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54c7ee),
	.w1(32'h3c4a3c97),
	.w2(32'hba858cd4),
	.w3(32'h3ca3d669),
	.w4(32'h3ce2a264),
	.w5(32'h3d375e05),
	.w6(32'hbc933ffe),
	.w7(32'hbd1a0e01),
	.w8(32'hbca6d251),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd81d),
	.w1(32'h3b8e0857),
	.w2(32'hbacb5371),
	.w3(32'h3cb73efe),
	.w4(32'h3c423e4e),
	.w5(32'h3caba7a8),
	.w6(32'hbc3d0ddf),
	.w7(32'hbcb94687),
	.w8(32'hbc4582d7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7bf8),
	.w1(32'h3b9f70a2),
	.w2(32'hba31e67b),
	.w3(32'h3bf58897),
	.w4(32'h3c246df5),
	.w5(32'h3ca264f2),
	.w6(32'hbc1b0835),
	.w7(32'hbc9c4616),
	.w8(32'hbc0e0c16),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789337),
	.w1(32'hbb71c613),
	.w2(32'hbba51535),
	.w3(32'h3bbbacec),
	.w4(32'h3c1a10b2),
	.w5(32'h3c1da44c),
	.w6(32'h3c0683a4),
	.w7(32'h3bb260e1),
	.w8(32'h3a2434b6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fce82),
	.w1(32'hbc31fb8d),
	.w2(32'hbbefeece),
	.w3(32'h3b20f368),
	.w4(32'hbc11e704),
	.w5(32'hbc43f6b7),
	.w6(32'hbb768178),
	.w7(32'h3aa8f9d6),
	.w8(32'hbbbead4b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c94e1),
	.w1(32'h3c045be0),
	.w2(32'h3bb33905),
	.w3(32'hbbffd1fe),
	.w4(32'h3bfa50f2),
	.w5(32'h3c7eaf09),
	.w6(32'hbb861be6),
	.w7(32'hbc4270c3),
	.w8(32'hbc8ce5ad),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8622a4),
	.w1(32'h3bd29652),
	.w2(32'h38a7dbf8),
	.w3(32'h3b8bbbe3),
	.w4(32'h3c3aa8f7),
	.w5(32'h3c2fb3b4),
	.w6(32'hbb748460),
	.w7(32'hbc295ab8),
	.w8(32'hbbbb4bf5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780c15),
	.w1(32'h3c2b7555),
	.w2(32'h3b81f2fe),
	.w3(32'h38dec164),
	.w4(32'h3c9b065a),
	.w5(32'h3cf6c15a),
	.w6(32'hbc5828fe),
	.w7(32'hbced9d48),
	.w8(32'hbc8e1e1f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6020a9),
	.w1(32'h3bb79aff),
	.w2(32'h3b833d1c),
	.w3(32'h3c4b200c),
	.w4(32'hba9bd977),
	.w5(32'hbb8484af),
	.w6(32'h3c07cafa),
	.w7(32'h3c094bfe),
	.w8(32'h3c024f54),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97d51),
	.w1(32'h3ae8e044),
	.w2(32'h3abe6f26),
	.w3(32'hbbd20dd9),
	.w4(32'hbb2b5d39),
	.w5(32'h3b8e9a2f),
	.w6(32'h3a895acd),
	.w7(32'hbb91670a),
	.w8(32'hbc059c25),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0faf83),
	.w1(32'h3be73b12),
	.w2(32'h3bb8ece1),
	.w3(32'hbc15d93e),
	.w4(32'h3c4100a4),
	.w5(32'h3cac7fc9),
	.w6(32'hbc2827c8),
	.w7(32'hbc8824b6),
	.w8(32'hbc51d6ed),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57f532),
	.w1(32'hb606ee53),
	.w2(32'hb626c551),
	.w3(32'h3bb10782),
	.w4(32'hb487befd),
	.w5(32'hb51e554a),
	.w6(32'hb4b51216),
	.w7(32'h3591f198),
	.w8(32'h35eeff6c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60e564c),
	.w1(32'hb7a53346),
	.w2(32'hb79c93d5),
	.w3(32'h3780dc72),
	.w4(32'h37a5d09f),
	.w5(32'h3794c89e),
	.w6(32'h38345e9d),
	.w7(32'h3804f05e),
	.w8(32'h380e9a58),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule