module layer_10_featuremap_217(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382edad3),
	.w1(32'hb6ff0997),
	.w2(32'h374f56aa),
	.w3(32'h384b21f2),
	.w4(32'hb6643eca),
	.w5(32'h372dc10b),
	.w6(32'h38447e76),
	.w7(32'h3566a76a),
	.w8(32'h37b7399a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4953cb),
	.w1(32'hb8304ad7),
	.w2(32'hba780f3a),
	.w3(32'hbb06ea99),
	.w4(32'h3a4a127c),
	.w5(32'hb8e6ec34),
	.w6(32'hbabfc915),
	.w7(32'h3a71963b),
	.w8(32'hba92a43c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37adb7d3),
	.w1(32'h37179e0b),
	.w2(32'h3789fd4a),
	.w3(32'h37710c69),
	.w4(32'hb68c757e),
	.w5(32'h36f7fe33),
	.w6(32'h373145fd),
	.w7(32'hb6b8e478),
	.w8(32'h36d5f8a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288a44),
	.w1(32'h3a1b2042),
	.w2(32'h3a3b9178),
	.w3(32'h37b063c4),
	.w4(32'hb94bc110),
	.w5(32'h38a8ec94),
	.w6(32'h39ae3695),
	.w7(32'h39585cd4),
	.w8(32'h3884abbd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391eb4b9),
	.w1(32'hb93e6146),
	.w2(32'hb9958c6f),
	.w3(32'h3976236f),
	.w4(32'hb8103440),
	.w5(32'hb933cbd4),
	.w6(32'h395ee294),
	.w7(32'h37a07f26),
	.w8(32'hb88491c3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d2b9b),
	.w1(32'h35ef85c8),
	.w2(32'h37fa15dc),
	.w3(32'h37fec3a5),
	.w4(32'hb6252a2e),
	.w5(32'h37df7355),
	.w6(32'h38228572),
	.w7(32'hb70e7d53),
	.w8(32'h3808186e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f56d39),
	.w1(32'hbaff6777),
	.w2(32'hbb8d12f7),
	.w3(32'hb8d6141f),
	.w4(32'hbb3e652e),
	.w5(32'hbbab1789),
	.w6(32'h39c055b2),
	.w7(32'hbb202b85),
	.w8(32'hbb9bab0b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfe1ed),
	.w1(32'hbb80d9c7),
	.w2(32'hbb5dc8d5),
	.w3(32'hbbfdf77e),
	.w4(32'hbba7a62c),
	.w5(32'hbb143913),
	.w6(32'hbbf89829),
	.w7(32'hbb960921),
	.w8(32'hbb67dc37),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7347da),
	.w1(32'h39065b30),
	.w2(32'hb9e9782c),
	.w3(32'hb9e37f1f),
	.w4(32'h39849736),
	.w5(32'hb9b5f7f6),
	.w6(32'hba0f1b7c),
	.w7(32'hb8a18992),
	.w8(32'hba17086a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc84c),
	.w1(32'hbb0db6e5),
	.w2(32'hbc2beda4),
	.w3(32'hbbcf6a27),
	.w4(32'hba6bbe83),
	.w5(32'hbbeccc79),
	.w6(32'hbb99274c),
	.w7(32'h3a9b2edf),
	.w8(32'hbbbd6b46),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911b21e),
	.w1(32'hba2404bd),
	.w2(32'hba0a62ed),
	.w3(32'h38c466a2),
	.w4(32'hb9d38c98),
	.w5(32'hb99fc088),
	.w6(32'hb5e9a761),
	.w7(32'hb9904b3a),
	.w8(32'hb97fcb57),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e5936),
	.w1(32'h3b526c8b),
	.w2(32'hb842bf98),
	.w3(32'hb907f5d3),
	.w4(32'h3af1d767),
	.w5(32'hba599808),
	.w6(32'h38985082),
	.w7(32'h3b1d0173),
	.w8(32'hbb4683dd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4621),
	.w1(32'hba8120d3),
	.w2(32'hbc1964d3),
	.w3(32'hbb486abe),
	.w4(32'hba429ae2),
	.w5(32'hbc0255c4),
	.w6(32'hbaa05728),
	.w7(32'h3a0f8f7d),
	.w8(32'hbbb9f590),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096c25),
	.w1(32'hba394dc1),
	.w2(32'hbaecc294),
	.w3(32'hbaf77a87),
	.w4(32'hb9e03cc4),
	.w5(32'hbab987b1),
	.w6(32'hbb1d43f1),
	.w7(32'hba30be8d),
	.w8(32'hbabe878a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386aaf),
	.w1(32'hb9d121bc),
	.w2(32'hbb3dc21f),
	.w3(32'hbafa9ef6),
	.w4(32'h3ad18695),
	.w5(32'hb9eeee43),
	.w6(32'hbb167267),
	.w7(32'h3b2d0027),
	.w8(32'hba29c073),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98884f),
	.w1(32'hbb28dc0f),
	.w2(32'hbc05fe85),
	.w3(32'hbb5a74a6),
	.w4(32'h39c960d0),
	.w5(32'hbb9c2f4c),
	.w6(32'hbb343815),
	.w7(32'hb9347f8d),
	.w8(32'hbb878f8b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c07023),
	.w1(32'h39c74bed),
	.w2(32'h3a0b5e1c),
	.w3(32'hb914d82b),
	.w4(32'h39800727),
	.w5(32'h3a25318a),
	.w6(32'hb9439657),
	.w7(32'h37b48567),
	.w8(32'h39ab39c8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d22f),
	.w1(32'hbaddc227),
	.w2(32'hbbf4fe62),
	.w3(32'hbbb3df4f),
	.w4(32'hbb22eefa),
	.w5(32'hbbdc8dfa),
	.w6(32'hbb878a8c),
	.w7(32'hbb5251a4),
	.w8(32'hbbd135be),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadefff3),
	.w1(32'hba40b7c2),
	.w2(32'hbba0eabc),
	.w3(32'hbb073209),
	.w4(32'hbad5e8a6),
	.w5(32'hbb9a7293),
	.w6(32'hba83d0c0),
	.w7(32'hbab4c1ba),
	.w8(32'hbb58f1d4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ed71ea),
	.w1(32'h38e69053),
	.w2(32'h385df29e),
	.w3(32'h381ca520),
	.w4(32'h390eada3),
	.w5(32'h386abd13),
	.w6(32'h387dd123),
	.w7(32'h39146379),
	.w8(32'h3732be4d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f42fa),
	.w1(32'hb623f3bb),
	.w2(32'h37b76358),
	.w3(32'h38804536),
	.w4(32'hb7d90276),
	.w5(32'h36b0ecc4),
	.w6(32'h38bd3a89),
	.w7(32'hb801983e),
	.w8(32'h3836dd12),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f9dd5),
	.w1(32'h3ab4d9c3),
	.w2(32'hb9ebad73),
	.w3(32'h3974707a),
	.w4(32'h3abe2a0a),
	.w5(32'hb9a8e64f),
	.w6(32'h369a6316),
	.w7(32'h3ae5e5ed),
	.w8(32'h37b6cc65),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03cd8b),
	.w1(32'hb795d7ed),
	.w2(32'hbb84c021),
	.w3(32'hbc114c9c),
	.w4(32'h3a553c76),
	.w5(32'hbbddd792),
	.w6(32'hbbc2f33f),
	.w7(32'h3a265759),
	.w8(32'hbc2d70f6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7ba81),
	.w1(32'hb99846f3),
	.w2(32'hbbf61442),
	.w3(32'hbb7e25da),
	.w4(32'h3b025614),
	.w5(32'hbb9fc3ea),
	.w6(32'hbb183d21),
	.w7(32'h3b938721),
	.w8(32'hbb241d46),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bb26),
	.w1(32'h3b31401f),
	.w2(32'hbb5fbf3c),
	.w3(32'hbbadc786),
	.w4(32'h3b3cc642),
	.w5(32'hbb1c4b1e),
	.w6(32'hbb927de0),
	.w7(32'h3baf1bf7),
	.w8(32'hb98bff77),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66654fa),
	.w1(32'hb8c528bb),
	.w2(32'hb9448526),
	.w3(32'h391facec),
	.w4(32'h38e4a2e1),
	.w5(32'hb8ea2903),
	.w6(32'hb76d681b),
	.w7(32'hb7802ea2),
	.w8(32'hb9823c4d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945830),
	.w1(32'h390abd7a),
	.w2(32'h3942debf),
	.w3(32'h39880afa),
	.w4(32'h38da325a),
	.w5(32'h391aa61b),
	.w6(32'h3964ec1f),
	.w7(32'h38bb8e31),
	.w8(32'h392ae679),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b887f),
	.w1(32'h3b3a121a),
	.w2(32'hbac38cc7),
	.w3(32'h36e8153e),
	.w4(32'h3b22272e),
	.w5(32'h3ac3a0e0),
	.w6(32'hb90fac89),
	.w7(32'h3b2234c6),
	.w8(32'h3b1c26a1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e43f54),
	.w1(32'h3ac4bab8),
	.w2(32'h399749da),
	.w3(32'hb7b00d8b),
	.w4(32'h3ab3850b),
	.w5(32'h3a3dc039),
	.w6(32'hba860a1b),
	.w7(32'h3aac5484),
	.w8(32'h3a294bf9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0280),
	.w1(32'h3b372efc),
	.w2(32'hbb59889e),
	.w3(32'hbaf4ef60),
	.w4(32'h3b31b0c5),
	.w5(32'hbb22d7e9),
	.w6(32'hbaefaae1),
	.w7(32'h3b699b2a),
	.w8(32'hba1f1501),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0cef7),
	.w1(32'h3897b615),
	.w2(32'h38970b2d),
	.w3(32'h388ce0f6),
	.w4(32'h38852f09),
	.w5(32'h38a79782),
	.w6(32'h37f5cc79),
	.w7(32'h3783d5c1),
	.w8(32'h38348474),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37847bf1),
	.w1(32'h385668e4),
	.w2(32'h38dd3e46),
	.w3(32'hb81b2bd8),
	.w4(32'hb7ccf3d9),
	.w5(32'h392b86f5),
	.w6(32'hb885147a),
	.w7(32'hb8099496),
	.w8(32'h38fffdb6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb220b23),
	.w1(32'hba4f84ac),
	.w2(32'hbb6e3fc6),
	.w3(32'hbae9a584),
	.w4(32'h39ce69fe),
	.w5(32'hbb18098f),
	.w6(32'hba4af466),
	.w7(32'h3aae3e93),
	.w8(32'hbaa7d90f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1da08),
	.w1(32'h3a51690e),
	.w2(32'hb97a50f7),
	.w3(32'hbab9db59),
	.w4(32'h3a934415),
	.w5(32'h398ebca6),
	.w6(32'hbad3a4cd),
	.w7(32'h3a8817d6),
	.w8(32'hb767be11),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a754b5),
	.w1(32'hb8fd46d4),
	.w2(32'hb9559d37),
	.w3(32'hba43f4b0),
	.w4(32'hba11ca16),
	.w5(32'hb94785ba),
	.w6(32'hba06208b),
	.w7(32'hba0d3f1b),
	.w8(32'hba214b8d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179c4f),
	.w1(32'hbaa5ea84),
	.w2(32'hbb32eac3),
	.w3(32'hb999aba2),
	.w4(32'hbaa1a438),
	.w5(32'hbb166848),
	.w6(32'h3a386c71),
	.w7(32'hba1bf8b7),
	.w8(32'hbb050424),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fe92),
	.w1(32'h3a4d7c0d),
	.w2(32'hbbb559e6),
	.w3(32'hbb80577d),
	.w4(32'h3b145c04),
	.w5(32'hbb2056c2),
	.w6(32'hb99517c2),
	.w7(32'h3bb8c58a),
	.w8(32'hbb9802b6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc054869),
	.w1(32'h3b964fea),
	.w2(32'h3b4bb212),
	.w3(32'hbbd50d9b),
	.w4(32'h3bc5ec28),
	.w5(32'h3b8c2d84),
	.w6(32'hbc223358),
	.w7(32'h3ba10211),
	.w8(32'h3a634731),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94ff14),
	.w1(32'h3c0ef2e2),
	.w2(32'h3b65caa4),
	.w3(32'hbb42969c),
	.w4(32'h3bc2e8bf),
	.w5(32'hba489eca),
	.w6(32'hbbdb701a),
	.w7(32'h3b2465a4),
	.w8(32'hbb2d6ae6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaf6c3),
	.w1(32'h3a8b3138),
	.w2(32'h3a880702),
	.w3(32'hbad07854),
	.w4(32'h3aabec13),
	.w5(32'h3aaf4b7f),
	.w6(32'hbb141934),
	.w7(32'h3a763b21),
	.w8(32'h39d5cfa9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815f047),
	.w1(32'hb895617e),
	.w2(32'h38a72b66),
	.w3(32'hb7e40a40),
	.w4(32'hb893c84f),
	.w5(32'h38a31f97),
	.w6(32'hb8f515b8),
	.w7(32'hb881184b),
	.w8(32'h388e76cc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e8f52),
	.w1(32'h3915b296),
	.w2(32'h392b7ed6),
	.w3(32'h39b72474),
	.w4(32'h3973a9f0),
	.w5(32'h3964cd90),
	.w6(32'h399bf48d),
	.w7(32'h39444e08),
	.w8(32'h39932ee2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92514),
	.w1(32'h3ae1802b),
	.w2(32'h38851804),
	.w3(32'hba3b9112),
	.w4(32'h3b00957c),
	.w5(32'hb931a63d),
	.w6(32'hba991589),
	.w7(32'h3a154ada),
	.w8(32'hbabc300b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd678f2),
	.w1(32'hb98b1e82),
	.w2(32'hbc1dcb4b),
	.w3(32'hbbc42ea7),
	.w4(32'h3781792d),
	.w5(32'hbc0164e6),
	.w6(32'hbb955f0a),
	.w7(32'hbb12c8f0),
	.w8(32'hbbf41a57),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb631f2),
	.w1(32'h39681411),
	.w2(32'hbbdb6097),
	.w3(32'hbb74d9ff),
	.w4(32'h3b2dd56a),
	.w5(32'hbb85f903),
	.w6(32'hbb405ddb),
	.w7(32'h3b974936),
	.w8(32'hbaf3bf87),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf048d9),
	.w1(32'h38dff46b),
	.w2(32'hbbfbffc0),
	.w3(32'hbba7ea8c),
	.w4(32'h3b004dd0),
	.w5(32'hbbb402ea),
	.w6(32'hbb538f11),
	.w7(32'h3ba7e288),
	.w8(32'hbb11571b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde220f),
	.w1(32'h3a0845a9),
	.w2(32'hbb4e8ca7),
	.w3(32'hbbb4f786),
	.w4(32'h3b253f60),
	.w5(32'hba5a3de0),
	.w6(32'hbb8228f4),
	.w7(32'h3b7b66a0),
	.w8(32'hba3d6143),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5986eb),
	.w1(32'hbb627857),
	.w2(32'hbc15723d),
	.w3(32'hbb74e24a),
	.w4(32'hbbae38b6),
	.w5(32'hbc0c66d2),
	.w6(32'hba9098ca),
	.w7(32'hbb9fee1b),
	.w8(32'hbc134649),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f35e0),
	.w1(32'h39f5f3d4),
	.w2(32'h3910be02),
	.w3(32'h39c4ae14),
	.w4(32'h39f742ca),
	.w5(32'h35e9b5bf),
	.w6(32'h39c0dc8b),
	.w7(32'h39eac9e2),
	.w8(32'h3967ae78),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a931),
	.w1(32'h3ae43819),
	.w2(32'h3a826baf),
	.w3(32'h3a9b9f56),
	.w4(32'h3a9fb74a),
	.w5(32'h3a7fd3d0),
	.w6(32'h3a9994d0),
	.w7(32'h3ab21eff),
	.w8(32'h3a705dfe),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eaf08),
	.w1(32'h3a8af266),
	.w2(32'h3891260e),
	.w3(32'h3a62d0b7),
	.w4(32'h3a80c7d7),
	.w5(32'h39a269d9),
	.w6(32'h3a89e977),
	.w7(32'h3a5c42a9),
	.w8(32'h3a1cf315),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e2b12),
	.w1(32'hb9c4ea42),
	.w2(32'hbb6dc368),
	.w3(32'hbac1fec3),
	.w4(32'h3a9a2d29),
	.w5(32'hbb06427c),
	.w6(32'hb963e9a4),
	.w7(32'h3b100b55),
	.w8(32'hb8d95869),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1275b7),
	.w1(32'h37f48ba2),
	.w2(32'hbacdd47d),
	.w3(32'hba2ddaab),
	.w4(32'hb7926857),
	.w5(32'hbac3ed93),
	.w6(32'hb9af4b92),
	.w7(32'h3983b39d),
	.w8(32'hbaa15dc9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb557a50),
	.w1(32'hbaa637d1),
	.w2(32'hbc09b389),
	.w3(32'hbb4f27f7),
	.w4(32'hbb09af57),
	.w5(32'hbbe2aaef),
	.w6(32'hbb56a325),
	.w7(32'hba3e33d4),
	.w8(32'hbba05b22),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddd29f),
	.w1(32'h39e5a398),
	.w2(32'hb9310a1e),
	.w3(32'hba1b9b9f),
	.w4(32'hb8e404d6),
	.w5(32'hb9bb1494),
	.w6(32'hb9f24765),
	.w7(32'hb8d6e4d0),
	.w8(32'hba16acc8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c42e0),
	.w1(32'h3787196f),
	.w2(32'hb842469e),
	.w3(32'h389e6daa),
	.w4(32'h38ff4089),
	.w5(32'h38aaca63),
	.w6(32'hb7ac4dca),
	.w7(32'h38af05bf),
	.w8(32'h38b7b687),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383fc319),
	.w1(32'h38185a48),
	.w2(32'h37f020e9),
	.w3(32'h38520825),
	.w4(32'h382480b8),
	.w5(32'h380aaf17),
	.w6(32'h38120fb0),
	.w7(32'h380dd47d),
	.w8(32'h3764028f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947aac0),
	.w1(32'h39bf3261),
	.w2(32'h38fd14a2),
	.w3(32'h38583ddf),
	.w4(32'h3906a48b),
	.w5(32'h37aeb1f4),
	.w6(32'hb87ff9d7),
	.w7(32'h3903b34b),
	.w8(32'h379d1c27),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900ccea),
	.w1(32'h3a722e74),
	.w2(32'h3a147b24),
	.w3(32'hb8d41627),
	.w4(32'h3a4d7d3c),
	.w5(32'h39b15ac0),
	.w6(32'hba57079a),
	.w7(32'h3916b38a),
	.w8(32'hb9bf1ed1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c6856),
	.w1(32'h38fd0d48),
	.w2(32'hb86dd565),
	.w3(32'h3713fec0),
	.w4(32'h39453004),
	.w5(32'hb888414d),
	.w6(32'h392344a5),
	.w7(32'hb8dd6f6d),
	.w8(32'hb9b29a7b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37ebd4),
	.w1(32'hba73e0a0),
	.w2(32'hbb6d1d5a),
	.w3(32'hbb2c2480),
	.w4(32'hba9a2c53),
	.w5(32'hbb4f43ca),
	.w6(32'hbaa4d7d1),
	.w7(32'hb9f1bd3a),
	.w8(32'hbafb8b82),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315e06),
	.w1(32'hba20d6bb),
	.w2(32'hbb1a130b),
	.w3(32'hbb048e23),
	.w4(32'hb9acfb27),
	.w5(32'hba84e1c5),
	.w6(32'hbad6fb3a),
	.w7(32'hbab3aa6a),
	.w8(32'hbaeb74fd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899e5c9),
	.w1(32'hb665a9c3),
	.w2(32'h3795dbe9),
	.w3(32'h38a01cca),
	.w4(32'h37428927),
	.w5(32'h38a9c1e5),
	.w6(32'h389921bc),
	.w7(32'h3725f84b),
	.w8(32'h38f5e610),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381626c0),
	.w1(32'hb6ce3191),
	.w2(32'h37c0be89),
	.w3(32'h3826ea22),
	.w4(32'hb6f4ed57),
	.w5(32'h377b7624),
	.w6(32'h384c2457),
	.w7(32'hb5e6b164),
	.w8(32'h37eedf14),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39217d82),
	.w1(32'h3904a430),
	.w2(32'h38dab284),
	.w3(32'h39438937),
	.w4(32'h38efe9db),
	.w5(32'h3898e7b6),
	.w6(32'h391808ea),
	.w7(32'h38f3f6a1),
	.w8(32'h3910dde6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e43cc1),
	.w1(32'h37d80df7),
	.w2(32'h38b1080f),
	.w3(32'h38ca7d0a),
	.w4(32'h377bffe5),
	.w5(32'h387fddba),
	.w6(32'h38a7bb7f),
	.w7(32'h360a929f),
	.w8(32'h3861df87),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb334fba),
	.w1(32'hbb42f255),
	.w2(32'hbbbf5b5d),
	.w3(32'hbba3527e),
	.w4(32'hbb8d3ef6),
	.w5(32'hbb58f654),
	.w6(32'hbb83bd2e),
	.w7(32'hbb83df6e),
	.w8(32'hbb8c8cc3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9589b6),
	.w1(32'hb9c3abec),
	.w2(32'hbbe0a649),
	.w3(32'hbb92ce6f),
	.w4(32'hbaa77986),
	.w5(32'hbc037dd0),
	.w6(32'hb8cba099),
	.w7(32'h3b328251),
	.w8(32'hbbb5bff4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c4749),
	.w1(32'h3b033bfe),
	.w2(32'hbb059496),
	.w3(32'hbb3fc6e0),
	.w4(32'h3b3cf312),
	.w5(32'hba688bd5),
	.w6(32'hbb3a2f8d),
	.w7(32'h3b0d933b),
	.w8(32'hbab14f8c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6f6b),
	.w1(32'h3b651fc0),
	.w2(32'hbc0af269),
	.w3(32'hbb7262b3),
	.w4(32'h3be62fc5),
	.w5(32'hbadc5630),
	.w6(32'hbb9739fa),
	.w7(32'h3c324f98),
	.w8(32'hba448e11),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9af73),
	.w1(32'hb7c0a4f2),
	.w2(32'h380d7f63),
	.w3(32'h38f5096c),
	.w4(32'hb80a97d6),
	.w5(32'h37cf578e),
	.w6(32'h38dbbb3c),
	.w7(32'hb7e69903),
	.w8(32'h380e53f9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39450084),
	.w1(32'h3758db44),
	.w2(32'h38f80803),
	.w3(32'h393e7de6),
	.w4(32'h335cdd37),
	.w5(32'h38debfd9),
	.w6(32'h3938cda7),
	.w7(32'h371617f7),
	.w8(32'h390c9b38),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902a44b),
	.w1(32'hb88b13b4),
	.w2(32'h380e5677),
	.w3(32'h38f50cba),
	.w4(32'hb8c03357),
	.w5(32'h33e7ab27),
	.w6(32'h39111e61),
	.w7(32'hb8cfd2f2),
	.w8(32'h380ebd9b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba568c87),
	.w1(32'h396e1261),
	.w2(32'hba4fc582),
	.w3(32'hba757b42),
	.w4(32'hba38c19b),
	.w5(32'hbab9c58a),
	.w6(32'hba85fe3f),
	.w7(32'hba884dfd),
	.w8(32'hba8db8de),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bcfd2),
	.w1(32'h37e970c1),
	.w2(32'h38d3cb0f),
	.w3(32'h392c7250),
	.w4(32'h38b37583),
	.w5(32'h3912d448),
	.w6(32'h39424600),
	.w7(32'h38c21f49),
	.w8(32'h39388025),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad51048),
	.w1(32'hba4dbfe7),
	.w2(32'hbafe4311),
	.w3(32'hbaea1a69),
	.w4(32'hbafc2520),
	.w5(32'hbb041843),
	.w6(32'hb97e2da5),
	.w7(32'hb9b996fd),
	.w8(32'hba8d68b1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef6b7),
	.w1(32'hbaedee77),
	.w2(32'hbba00136),
	.w3(32'hbb912e2c),
	.w4(32'hbab5b479),
	.w5(32'hbb17c267),
	.w6(32'hbb26385b),
	.w7(32'hba0cd549),
	.w8(32'hbb71840f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba039ce),
	.w1(32'hbb23f8cf),
	.w2(32'hbbda755c),
	.w3(32'hbb82e69b),
	.w4(32'hba4e3162),
	.w5(32'hbb7c0d89),
	.w6(32'hbb0d17ed),
	.w7(32'h3b00f7ed),
	.w8(32'hba939e3e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdc6a4),
	.w1(32'hb97542e9),
	.w2(32'hbb780616),
	.w3(32'hbaad9349),
	.w4(32'h3a1b9938),
	.w5(32'hbb148664),
	.w6(32'hbb00344a),
	.w7(32'h39318142),
	.w8(32'hbacf7d63),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954b8fc),
	.w1(32'h3976c937),
	.w2(32'hbb350379),
	.w3(32'hbb03c432),
	.w4(32'hbab6a922),
	.w5(32'hbb199e40),
	.w6(32'h39453d93),
	.w7(32'h3a8831c6),
	.w8(32'hbacc69d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29b90c),
	.w1(32'hba6815b4),
	.w2(32'hbb60f986),
	.w3(32'hbafc86f3),
	.w4(32'h395aa8c5),
	.w5(32'hbafb2893),
	.w6(32'hbad183d4),
	.w7(32'h3a4a6844),
	.w8(32'hba757b02),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63288f),
	.w1(32'h38d2fb75),
	.w2(32'hbb56675f),
	.w3(32'hbab068bf),
	.w4(32'hbad7128b),
	.w5(32'hbb87a657),
	.w6(32'hb9817ef3),
	.w7(32'hb99d53e1),
	.w8(32'hbb35fc26),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379760f6),
	.w1(32'hb693832b),
	.w2(32'h37482f6b),
	.w3(32'h3798e69d),
	.w4(32'hb6c8a645),
	.w5(32'h372170f4),
	.w6(32'h376bfe0a),
	.w7(32'hb6ee2756),
	.w8(32'h373ab1cb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a475b4),
	.w1(32'hb6cd9bb6),
	.w2(32'h36892aa1),
	.w3(32'h37a69938),
	.w4(32'h3719e241),
	.w5(32'h37974165),
	.w6(32'h376ac1ff),
	.w7(32'h370d8850),
	.w8(32'h37a2b1bf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb612fac7),
	.w1(32'h35b49c1f),
	.w2(32'h37531e8b),
	.w3(32'hb808e156),
	.w4(32'hb7f496ba),
	.w5(32'h35c4fea2),
	.w6(32'h371f5178),
	.w7(32'h3773763f),
	.w8(32'hb64551b3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b813b0),
	.w1(32'h39ebfcda),
	.w2(32'h39a4143f),
	.w3(32'h37e79465),
	.w4(32'h39a521ce),
	.w5(32'h39434cf1),
	.w6(32'h38be128b),
	.w7(32'h3a072910),
	.w8(32'h39c9c06a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0a894),
	.w1(32'hb9b1be40),
	.w2(32'h3a77c79a),
	.w3(32'hbba51063),
	.w4(32'h3a87f25b),
	.w5(32'h3b3af17b),
	.w6(32'hbb9b98c2),
	.w7(32'h3b161c4e),
	.w8(32'h3acb84d4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03a332),
	.w1(32'h3a62dcec),
	.w2(32'h39f4d608),
	.w3(32'h3a2d407c),
	.w4(32'h3aad3b3d),
	.w5(32'h39d0429a),
	.w6(32'hb987f862),
	.w7(32'h3a29e619),
	.w8(32'hb93079cc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6afa88),
	.w1(32'hb989a429),
	.w2(32'hbb7dfc7c),
	.w3(32'hbb1dcf20),
	.w4(32'h3a2ac68e),
	.w5(32'hbb4be6da),
	.w6(32'hbadb76bb),
	.w7(32'h3af4faa7),
	.w8(32'hbb08dadf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0aab),
	.w1(32'hb9ce4a78),
	.w2(32'hbb41688b),
	.w3(32'hbbdd0b4a),
	.w4(32'hbadd37b0),
	.w5(32'hbb27e7ea),
	.w6(32'hbbbb948e),
	.w7(32'hbb238a45),
	.w8(32'hbb31ee9e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91cee3f),
	.w1(32'h3b4b6217),
	.w2(32'h3a1bae67),
	.w3(32'hba5face5),
	.w4(32'h3b079fc1),
	.w5(32'h3965beb5),
	.w6(32'hbb051d11),
	.w7(32'h3b1b788b),
	.w8(32'hb95f4378),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32c387),
	.w1(32'hbb31b961),
	.w2(32'hbbdadb60),
	.w3(32'hbb824884),
	.w4(32'hbb1c5310),
	.w5(32'hbba7838f),
	.w6(32'hba9bc9cc),
	.w7(32'hbac31149),
	.w8(32'hbbe23b8c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08b603),
	.w1(32'h3b8a458e),
	.w2(32'h39a4d08d),
	.w3(32'h3a5bea5d),
	.w4(32'h3b4ae39a),
	.w5(32'hba536a23),
	.w6(32'h3ab99c3a),
	.w7(32'h3b933daf),
	.w8(32'h3ad93951),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd75b),
	.w1(32'hba8c4269),
	.w2(32'hbb8d6512),
	.w3(32'hbb91dc31),
	.w4(32'h392f3e2b),
	.w5(32'hbafa4986),
	.w6(32'hbba598dc),
	.w7(32'hb964ecb4),
	.w8(32'hbb12ff28),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c899),
	.w1(32'h3a14f857),
	.w2(32'hbb0ebe27),
	.w3(32'hbb2f8879),
	.w4(32'h3afe1f9a),
	.w5(32'h3a225806),
	.w6(32'hbae66df1),
	.w7(32'h3b0bd976),
	.w8(32'h3a0b5ec2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae8f6),
	.w1(32'h3b17171b),
	.w2(32'hba3b4322),
	.w3(32'hbb6cc571),
	.w4(32'h3b44adc5),
	.w5(32'hba889249),
	.w6(32'hbb642562),
	.w7(32'h3b9290fa),
	.w8(32'h3a54a1d4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855398),
	.w1(32'h3afa3d84),
	.w2(32'h3a0f11be),
	.w3(32'h3a9e01da),
	.w4(32'h3a964435),
	.w5(32'h39b7331f),
	.w6(32'h3a757aa9),
	.w7(32'h3a88c007),
	.w8(32'h3a70d7cd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4878b2),
	.w1(32'h3ae4f52e),
	.w2(32'hbbc358a0),
	.w3(32'hbb4040c4),
	.w4(32'h3b1c2383),
	.w5(32'hbb817a15),
	.w6(32'hbb0bb0ef),
	.w7(32'h3a255a68),
	.w8(32'hbb77f416),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e0a6),
	.w1(32'h3ab558c6),
	.w2(32'hbadd6b69),
	.w3(32'hbb2fa93e),
	.w4(32'h3adcca44),
	.w5(32'h397bb325),
	.w6(32'hb9f24dba),
	.w7(32'h3aede365),
	.w8(32'hbb17782a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a37a),
	.w1(32'hb9e0d264),
	.w2(32'hbbdcc4fd),
	.w3(32'hbb69faf8),
	.w4(32'h39f7648b),
	.w5(32'hbbc9c346),
	.w6(32'h3b1e90c9),
	.w7(32'h3b8a928e),
	.w8(32'hbbe7547a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc579000),
	.w1(32'h3b1c9b31),
	.w2(32'h3baaa447),
	.w3(32'hbc4bd2bf),
	.w4(32'h3b77d5c4),
	.w5(32'h3bcd0c52),
	.w6(32'hbc54f789),
	.w7(32'h3aaf43a6),
	.w8(32'hbb1a8d4f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d98b),
	.w1(32'h3a49ed27),
	.w2(32'hbc04f331),
	.w3(32'hbb2efe77),
	.w4(32'h3a9b0dee),
	.w5(32'hbbd645c9),
	.w6(32'hba987ab4),
	.w7(32'h3b86f655),
	.w8(32'hbb471730),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db5fb),
	.w1(32'hb8ec6663),
	.w2(32'hbb42a863),
	.w3(32'hbb6da3e0),
	.w4(32'h3a619e58),
	.w5(32'hbad2e71a),
	.w6(32'h3abd96ff),
	.w7(32'h3b28c5e8),
	.w8(32'hbb5cca46),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ac472),
	.w1(32'h3aa4ef46),
	.w2(32'h39b8b963),
	.w3(32'hba251bca),
	.w4(32'h39ce9747),
	.w5(32'hbabb855e),
	.w6(32'h3781dfd4),
	.w7(32'hb91532e5),
	.w8(32'hbaaca09b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bae65),
	.w1(32'hbbb6a47e),
	.w2(32'hbc00895b),
	.w3(32'hbbb61c10),
	.w4(32'hbb65ee5f),
	.w5(32'hbbd6fc6b),
	.w6(32'hba710602),
	.w7(32'h3b60475f),
	.w8(32'hbb17aee2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb9cb4),
	.w1(32'hba91a072),
	.w2(32'hbb5a1c11),
	.w3(32'hba94acbf),
	.w4(32'hba812f81),
	.w5(32'hbb504570),
	.w6(32'h3a7e8c72),
	.w7(32'h3a559be3),
	.w8(32'hbb337e70),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384dce01),
	.w1(32'h38e78474),
	.w2(32'hb87c1bd1),
	.w3(32'h37a6654e),
	.w4(32'h39070125),
	.w5(32'h3792c1ba),
	.w6(32'h38b75fb9),
	.w7(32'h3935e5e0),
	.w8(32'h37986c12),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946cd1),
	.w1(32'hba5600ad),
	.w2(32'hba81530c),
	.w3(32'hba0105f3),
	.w4(32'hb976347c),
	.w5(32'hba13eb4b),
	.w6(32'hba4769d3),
	.w7(32'hb9aeba79),
	.w8(32'hba2ef884),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588446),
	.w1(32'h391179d5),
	.w2(32'hbb9f2467),
	.w3(32'hbb2d7d4f),
	.w4(32'hba7855b8),
	.w5(32'hbba72bb3),
	.w6(32'hbae40ace),
	.w7(32'hbaebcbc3),
	.w8(32'hbba475d2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508279),
	.w1(32'h3b714385),
	.w2(32'hbb51228f),
	.w3(32'h3a45a1d5),
	.w4(32'h3b384aa9),
	.w5(32'hbb415db2),
	.w6(32'h3a8cec1c),
	.w7(32'h3b9419db),
	.w8(32'hb8afe5ab),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb425a85),
	.w1(32'h3984a639),
	.w2(32'hbad3f2bc),
	.w3(32'hbb3a9a46),
	.w4(32'h3a0d2d80),
	.w5(32'hbab4cc4c),
	.w6(32'hbb661c76),
	.w7(32'hba3c50a3),
	.w8(32'hbb29930b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2905fc),
	.w1(32'h3ae4fb8e),
	.w2(32'hba51ede0),
	.w3(32'hbb0a1aa7),
	.w4(32'h3b0fef18),
	.w5(32'hb8c82a07),
	.w6(32'hbaa5ca05),
	.w7(32'h3af4a995),
	.w8(32'hba131320),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8244c5),
	.w1(32'h3a9bcbbc),
	.w2(32'hb9fdc33c),
	.w3(32'hbafe8d5a),
	.w4(32'h39fa078e),
	.w5(32'hba852f78),
	.w6(32'hbab55dd5),
	.w7(32'h3a505064),
	.w8(32'hbae07d6f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6229e0),
	.w1(32'hbaa3c92a),
	.w2(32'hbb89186f),
	.w3(32'hbb4468c8),
	.w4(32'h3965e8fd),
	.w5(32'hbb2b551e),
	.w6(32'hbad2c047),
	.w7(32'h393bba5c),
	.w8(32'hbb1800f0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206b8b),
	.w1(32'h38d6bef5),
	.w2(32'hbb1ccdb4),
	.w3(32'hbb0782dd),
	.w4(32'h39fce539),
	.w5(32'hbb0a3167),
	.w6(32'hbacd8359),
	.w7(32'h3ab4723a),
	.w8(32'hbabd435a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9217571),
	.w1(32'hb896b9ab),
	.w2(32'hb81ddbe8),
	.w3(32'hb92ecf8e),
	.w4(32'hb8a9cdff),
	.w5(32'hb653127f),
	.w6(32'hb92a48a7),
	.w7(32'hb90a03ba),
	.w8(32'hb8c05573),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98228e8),
	.w1(32'hb8e6c8ca),
	.w2(32'hb8885553),
	.w3(32'hb8accb78),
	.w4(32'h386830b2),
	.w5(32'h38b37141),
	.w6(32'hb942957d),
	.w7(32'h384753a5),
	.w8(32'hb858e06b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38848e74),
	.w1(32'h391cc2c6),
	.w2(32'h3901ed78),
	.w3(32'hb8103fc6),
	.w4(32'h38b5870e),
	.w5(32'h388b5c9b),
	.w6(32'hb52deab3),
	.w7(32'h38339869),
	.w8(32'h3768af95),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954ea3a),
	.w1(32'h363af656),
	.w2(32'h38c1dc04),
	.w3(32'h39804521),
	.w4(32'h391c2ece),
	.w5(32'h3992c5e2),
	.w6(32'h398e2264),
	.w7(32'h390df5a1),
	.w8(32'h3a0988d6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cfb49),
	.w1(32'h376832a4),
	.w2(32'hbb8b9f6f),
	.w3(32'hbb05c7de),
	.w4(32'h3aa627e2),
	.w5(32'hbb417818),
	.w6(32'hbaba18bd),
	.w7(32'h3b38505c),
	.w8(32'hbaa9bf6a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba453d3b),
	.w1(32'hba8f5a20),
	.w2(32'hba9feeca),
	.w3(32'hb9cc4d84),
	.w4(32'hba3212be),
	.w5(32'hba85387a),
	.w6(32'hba165e2f),
	.w7(32'hba2c95f0),
	.w8(32'hba224847),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff76cc),
	.w1(32'hba668dde),
	.w2(32'hbb2a33eb),
	.w3(32'hba93d57d),
	.w4(32'hbaa30c3b),
	.w5(32'hbad36c1c),
	.w6(32'h390188ff),
	.w7(32'hb9a0f15e),
	.w8(32'hbabe716d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb138f4),
	.w1(32'h3a1665a8),
	.w2(32'hb9b65235),
	.w3(32'hbbb2041a),
	.w4(32'h396bce3a),
	.w5(32'hba47844e),
	.w6(32'hbba423ef),
	.w7(32'h3958a246),
	.w8(32'hbb216ca3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907a27b),
	.w1(32'hb5cdf404),
	.w2(32'hb8490078),
	.w3(32'h392ada25),
	.w4(32'h38a93ccd),
	.w5(32'h389b5f32),
	.w6(32'h39571f9c),
	.w7(32'h39252bd3),
	.w8(32'h38c14e91),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c49e73),
	.w1(32'h39820e05),
	.w2(32'h3917ea66),
	.w3(32'h393ac0b2),
	.w4(32'h39ce69c9),
	.w5(32'h3989e576),
	.w6(32'hb90cd61f),
	.w7(32'hb74b738e),
	.w8(32'hb89cf010),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843dff3),
	.w1(32'h37f0a243),
	.w2(32'h386c5f22),
	.w3(32'h380062a1),
	.w4(32'h37a85253),
	.w5(32'h388828b1),
	.w6(32'hb778be76),
	.w7(32'hb7a64e0e),
	.w8(32'h37bec1b0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba818c04),
	.w1(32'hba479c04),
	.w2(32'hba228408),
	.w3(32'hba988be4),
	.w4(32'hb9f9738b),
	.w5(32'hb97a739b),
	.w6(32'hbabc1836),
	.w7(32'hbaa0a3c0),
	.w8(32'hba8c1d81),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9737a),
	.w1(32'hbb34c76d),
	.w2(32'hbb74c1f9),
	.w3(32'hb9e269ae),
	.w4(32'hbb783091),
	.w5(32'hbbc7d31c),
	.w6(32'h3ab4eb19),
	.w7(32'hbb1ee11d),
	.w8(32'hbb85feb3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e6ef),
	.w1(32'hbb3f570a),
	.w2(32'hbbeed70d),
	.w3(32'hbb34bc71),
	.w4(32'hbb27c7a3),
	.w5(32'hbbcf3f4a),
	.w6(32'hbb2a0f81),
	.w7(32'hba4f14f6),
	.w8(32'hbba18102),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8bd75),
	.w1(32'h3879d285),
	.w2(32'hb90e3640),
	.w3(32'hba2085b8),
	.w4(32'h3977cea7),
	.w5(32'h3998f8af),
	.w6(32'h3a24c667),
	.w7(32'h39f2ca9d),
	.w8(32'hb92c139a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb01c3),
	.w1(32'hba36e447),
	.w2(32'hbaaa1447),
	.w3(32'hbadcce4f),
	.w4(32'hba43744b),
	.w5(32'hba8c60f6),
	.w6(32'hbb0fec09),
	.w7(32'hba9a48e4),
	.w8(32'hbaf0d911),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb9a84),
	.w1(32'h39be4187),
	.w2(32'hba615eab),
	.w3(32'hbb1270f2),
	.w4(32'h3a66e392),
	.w5(32'hba3fb41e),
	.w6(32'hba93f413),
	.w7(32'h39ff8272),
	.w8(32'hba853aca),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c1a51),
	.w1(32'hba94a906),
	.w2(32'hbb4eb4a0),
	.w3(32'hba5a0ae5),
	.w4(32'h39865315),
	.w5(32'hbb19306c),
	.w6(32'hbb2f9842),
	.w7(32'hbac329be),
	.w8(32'hbab9d836),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839e0d),
	.w1(32'hbb0415ed),
	.w2(32'hbb7fecb8),
	.w3(32'hbb4d6037),
	.w4(32'hb915cf83),
	.w5(32'hba9cfc39),
	.w6(32'hbb47524f),
	.w7(32'hb9b59609),
	.w8(32'hba322b35),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ce6d),
	.w1(32'hba8b159e),
	.w2(32'hbbaf8377),
	.w3(32'hbb892d3d),
	.w4(32'hbb081d13),
	.w5(32'hbbb8bc35),
	.w6(32'hba8f20ba),
	.w7(32'hba6882a3),
	.w8(32'hbbb45b61),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75671e),
	.w1(32'h398e3629),
	.w2(32'hbb10f602),
	.w3(32'hbb39abbe),
	.w4(32'h3a9d58a4),
	.w5(32'hbac1de64),
	.w6(32'hbb5865b5),
	.w7(32'h3a282458),
	.w8(32'hbb1bd36c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fd17),
	.w1(32'hbb1da38f),
	.w2(32'hbb5963ec),
	.w3(32'hbb6ad1b4),
	.w4(32'h391a9a0c),
	.w5(32'hba831166),
	.w6(32'hbaa698a7),
	.w7(32'h3addbdaa),
	.w8(32'hba92fd79),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a238),
	.w1(32'hb9ce5bb2),
	.w2(32'hbb798281),
	.w3(32'hbb757129),
	.w4(32'h3a29df8d),
	.w5(32'hbb3e5d87),
	.w6(32'hbaa95b38),
	.w7(32'h3a0c11fd),
	.w8(32'hbb25bf80),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0505e2),
	.w1(32'h395e98ca),
	.w2(32'h39e5de12),
	.w3(32'hba8eae25),
	.w4(32'h3a03cb5a),
	.w5(32'h3a15ba10),
	.w6(32'hbb2155d4),
	.w7(32'h3acc810d),
	.w8(32'hb91e2d23),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d87b),
	.w1(32'hb9a056f5),
	.w2(32'hbb80b479),
	.w3(32'hbb36294f),
	.w4(32'h3a15b8d4),
	.w5(32'hbb2def4e),
	.w6(32'hbac9460c),
	.w7(32'h39afd6cf),
	.w8(32'hbb5e71ff),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad8d44),
	.w1(32'hb9fde7b2),
	.w2(32'hbad67b66),
	.w3(32'hbace1b76),
	.w4(32'h381ef4a2),
	.w5(32'hbaa2baac),
	.w6(32'hba8a5275),
	.w7(32'h39447b07),
	.w8(32'hba647005),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95374f),
	.w1(32'h3b82b18a),
	.w2(32'h39ea3c01),
	.w3(32'hbbb7918d),
	.w4(32'h3b3a33fc),
	.w5(32'hba071511),
	.w6(32'hbb9278b1),
	.w7(32'h3b4c9bba),
	.w8(32'hba91516e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb610a85),
	.w1(32'h3a4192b9),
	.w2(32'h3b061a37),
	.w3(32'hbb32f4d9),
	.w4(32'h3ae70f4a),
	.w5(32'h3ab0556e),
	.w6(32'hbb547da7),
	.w7(32'h3a7e9dcc),
	.w8(32'h397fa8b0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2410c),
	.w1(32'hba8e90a3),
	.w2(32'hba60a022),
	.w3(32'hb9a1c845),
	.w4(32'hba52ebe9),
	.w5(32'hba3640d4),
	.w6(32'hba82607b),
	.w7(32'hba537a39),
	.w8(32'hb9f7f508),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2213bf),
	.w1(32'h39cf3ab9),
	.w2(32'h398d77e8),
	.w3(32'hb9db9db9),
	.w4(32'hb98aeab8),
	.w5(32'h3963db9a),
	.w6(32'hb833b29e),
	.w7(32'h398b7b22),
	.w8(32'h3a3f2fc2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2ce9a),
	.w1(32'hb9c59891),
	.w2(32'hba8caab0),
	.w3(32'hbab66235),
	.w4(32'h3a4416e0),
	.w5(32'h3a3a56da),
	.w6(32'hb9e6b296),
	.w7(32'h394f2cfe),
	.w8(32'hba509276),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcc2c),
	.w1(32'h394388d1),
	.w2(32'hba2bbfba),
	.w3(32'hbb5383a6),
	.w4(32'h3b1e0c3f),
	.w5(32'h3a4377ed),
	.w6(32'hbb1f12a6),
	.w7(32'h3b38bea5),
	.w8(32'hb92054b8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8771d1),
	.w1(32'hba9ea1ec),
	.w2(32'hbbf70961),
	.w3(32'hbb9ebb39),
	.w4(32'hba237afb),
	.w5(32'hbbd452e8),
	.w6(32'hbb32d570),
	.w7(32'hb9046e90),
	.w8(32'hbb85ecee),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9a3b2),
	.w1(32'hb85fb821),
	.w2(32'hb9360f67),
	.w3(32'h38f3cbaf),
	.w4(32'hb739c8fe),
	.w5(32'hb8f97445),
	.w6(32'h37470d5a),
	.w7(32'hb9b2a9a3),
	.w8(32'h386c212b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842637),
	.w1(32'hbb13bdf6),
	.w2(32'hbbe096d5),
	.w3(32'hbb727a2f),
	.w4(32'hba85c3bb),
	.w5(32'hbbb1ba68),
	.w6(32'hbb2f26ec),
	.w7(32'h3a689e07),
	.w8(32'hbb5a7065),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26e9c5),
	.w1(32'hb93da2aa),
	.w2(32'hbb74fdf0),
	.w3(32'hbb338a17),
	.w4(32'h39e5df50),
	.w5(32'hbb6574a4),
	.w6(32'hba2b6b06),
	.w7(32'h3a9e8c00),
	.w8(32'hbaaec594),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db2f9),
	.w1(32'hbb77c7cc),
	.w2(32'hbbdbf823),
	.w3(32'hbb4afc6c),
	.w4(32'hbb404abd),
	.w5(32'hbb98a447),
	.w6(32'hbaf272bd),
	.w7(32'hbaf69dfd),
	.w8(32'hbb8938f2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a007a),
	.w1(32'h3b5c5102),
	.w2(32'hbb89dccf),
	.w3(32'hbadca4bb),
	.w4(32'h3b7834bc),
	.w5(32'hbab034bb),
	.w6(32'hb9b0ede6),
	.w7(32'h3be0ad16),
	.w8(32'h3addcf1d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974ea3),
	.w1(32'h3adabaa3),
	.w2(32'h3aa2dbcb),
	.w3(32'hba4708e4),
	.w4(32'h3a8e709d),
	.w5(32'h3a09b9fe),
	.w6(32'hbb054241),
	.w7(32'h3a3ac6ec),
	.w8(32'hbab3e9e8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0c0b2),
	.w1(32'h3ad56b02),
	.w2(32'h39d1410e),
	.w3(32'h3ae35247),
	.w4(32'h3a901b8b),
	.w5(32'hb9178962),
	.w6(32'h3aae6949),
	.w7(32'h3a201b1d),
	.w8(32'h39d7ea77),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506799),
	.w1(32'h3a2c2d42),
	.w2(32'h39bee95e),
	.w3(32'hbac1ce8d),
	.w4(32'h3b31784e),
	.w5(32'h3ac98ab9),
	.w6(32'hbb85a158),
	.w7(32'h3b07d5e7),
	.w8(32'h3a97ca95),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb274fc),
	.w1(32'h3aa6fc9d),
	.w2(32'h39ac97e9),
	.w3(32'hbb63afc4),
	.w4(32'h3b200b6b),
	.w5(32'h3ac7ff21),
	.w6(32'hbb70c1bf),
	.w7(32'h3a8450ab),
	.w8(32'hbac72acf),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39875afc),
	.w1(32'h3b57e731),
	.w2(32'h3a8894b6),
	.w3(32'hb9d0889a),
	.w4(32'h3b363ddd),
	.w5(32'h3a81c04b),
	.w6(32'hba69644d),
	.w7(32'h3b4871d1),
	.w8(32'h385b22ce),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d614ed),
	.w1(32'hba0c9fc8),
	.w2(32'hba68368a),
	.w3(32'hba539e3c),
	.w4(32'hbaa400b4),
	.w5(32'hba8f3d8a),
	.w6(32'hb97f3d3e),
	.w7(32'hb9f21813),
	.w8(32'hba4f2e30),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a57f58),
	.w1(32'hba3a84bf),
	.w2(32'hba0fed79),
	.w3(32'hb9487adf),
	.w4(32'hb9c061a3),
	.w5(32'hb9ab996a),
	.w6(32'hba550ca8),
	.w7(32'hba692497),
	.w8(32'hba4df786),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68567c),
	.w1(32'hbaf63797),
	.w2(32'hbafc4b1f),
	.w3(32'hbb500ceb),
	.w4(32'hba9c1e8a),
	.w5(32'hbaab04d7),
	.w6(32'hbb0a6434),
	.w7(32'h3a7d3c12),
	.w8(32'hbb0d8d0b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20c1bf),
	.w1(32'hb905800b),
	.w2(32'hba54f738),
	.w3(32'h3a1f60f4),
	.w4(32'h399f23a1),
	.w5(32'hba777f2a),
	.w6(32'hb9a763be),
	.w7(32'hba7aafc0),
	.w8(32'hba6e9de1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101e64),
	.w1(32'h3aa2af1c),
	.w2(32'hba763456),
	.w3(32'hbac75988),
	.w4(32'h3aca3103),
	.w5(32'hba6551c6),
	.w6(32'hba69b0ab),
	.w7(32'h3aec3c9c),
	.w8(32'h39758cf8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a078389),
	.w1(32'h39f524b8),
	.w2(32'h39640f11),
	.w3(32'h39da1c54),
	.w4(32'h3a0444f2),
	.w5(32'h396bb191),
	.w6(32'hb7264235),
	.w7(32'h388f46cb),
	.w8(32'h39d7b597),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d83935),
	.w1(32'h3abdc60e),
	.w2(32'hbb06287a),
	.w3(32'hbb07d8cc),
	.w4(32'hba58c611),
	.w5(32'hbb62b2cb),
	.w6(32'h397d4235),
	.w7(32'h3a3fe0fb),
	.w8(32'hbb0394bb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fab13e),
	.w1(32'h3a21ecbc),
	.w2(32'h3a112005),
	.w3(32'h3a1fe4ec),
	.w4(32'h3a6c1b61),
	.w5(32'h3a4dac44),
	.w6(32'h3a6be199),
	.w7(32'h3a36969d),
	.w8(32'h39a1e9d5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39810ea0),
	.w1(32'hba7fe1a1),
	.w2(32'hba7de9f0),
	.w3(32'h397e0371),
	.w4(32'hba46e843),
	.w5(32'hba6eada9),
	.w6(32'hba7011bd),
	.w7(32'hba8a5e03),
	.w8(32'hba686994),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9973e7),
	.w1(32'hba65d2d4),
	.w2(32'hbaccb028),
	.w3(32'hbb5d99e3),
	.w4(32'h3aa2b837),
	.w5(32'h38ce6360),
	.w6(32'hbb82e726),
	.w7(32'hba029c19),
	.w8(32'hbaf3790c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5a3fe),
	.w1(32'hb9d3cce1),
	.w2(32'hbbc19e90),
	.w3(32'hbba26d88),
	.w4(32'hba7e8532),
	.w5(32'hbc10ae3f),
	.w6(32'hba89cf40),
	.w7(32'h3b5c0d30),
	.w8(32'hbbbf6417),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f37f2),
	.w1(32'h3b149fb6),
	.w2(32'h39e578fd),
	.w3(32'h395e686f),
	.w4(32'h3ae02000),
	.w5(32'h39c9869b),
	.w6(32'hb9f77def),
	.w7(32'h3abfa480),
	.w8(32'hb9681258),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33ef40),
	.w1(32'h38700756),
	.w2(32'hbb77dd5c),
	.w3(32'hbb12b62a),
	.w4(32'h3a9bed0f),
	.w5(32'hbb4e05c5),
	.w6(32'hbb05b3a7),
	.w7(32'h3b096bf4),
	.w8(32'hbb2ffbdb),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996a178),
	.w1(32'h3b22fa75),
	.w2(32'h3994dc8c),
	.w3(32'hba3db692),
	.w4(32'h3b178032),
	.w5(32'h3aaccd15),
	.w6(32'h3af44acc),
	.w7(32'h3b0a7196),
	.w8(32'h3ac476ed),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba94a8),
	.w1(32'hbac7041c),
	.w2(32'hbc128940),
	.w3(32'hbba47946),
	.w4(32'h3ad710dd),
	.w5(32'hbb940b31),
	.w6(32'hbb4b0a82),
	.w7(32'h39e853e1),
	.w8(32'hbbae7cbe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6778d8),
	.w1(32'hba8abcc1),
	.w2(32'hbb9cd114),
	.w3(32'hbb5754e9),
	.w4(32'hb8895bc2),
	.w5(32'hbb48035e),
	.w6(32'hbb4f005a),
	.w7(32'h3a636bba),
	.w8(32'hbb1fbad4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b73f9),
	.w1(32'h3966416b),
	.w2(32'hbbd92da0),
	.w3(32'hbb5f9562),
	.w4(32'h3a49f5dd),
	.w5(32'hbbda5726),
	.w6(32'hbaa6da18),
	.w7(32'h3ab9a40d),
	.w8(32'hbb6febbb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8ff15),
	.w1(32'h3a37e295),
	.w2(32'hb911fe81),
	.w3(32'hba19b6cf),
	.w4(32'h39dfb06d),
	.w5(32'h39b78bbe),
	.w6(32'h3939a699),
	.w7(32'hb99f6d76),
	.w8(32'h3a135428),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac521ec),
	.w1(32'hb9b90867),
	.w2(32'hbb1130a3),
	.w3(32'hba9c1719),
	.w4(32'h3a5e75d8),
	.w5(32'hba1e0403),
	.w6(32'hb9d57cbe),
	.w7(32'h3adfad37),
	.w8(32'hb92e8734),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e4068c),
	.w1(32'hba15eb74),
	.w2(32'hba1a5a2c),
	.w3(32'h39bee703),
	.w4(32'hb9ca73e0),
	.w5(32'hb9ded7d9),
	.w6(32'hb9eafa3a),
	.w7(32'hba248fb8),
	.w8(32'hb9fb2ecb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9a40e),
	.w1(32'h396c9471),
	.w2(32'hbb0856e1),
	.w3(32'h39027c6e),
	.w4(32'h39cb61a2),
	.w5(32'hba85be52),
	.w6(32'h3a859b9b),
	.w7(32'h39b433b0),
	.w8(32'hba57c633),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba234f91),
	.w1(32'h3aa028b1),
	.w2(32'h3a366f59),
	.w3(32'hba81c8a2),
	.w4(32'h39ab4ec9),
	.w5(32'h3a158f55),
	.w6(32'hb9b66f28),
	.w7(32'h3a983e21),
	.w8(32'h3937de88),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea0522),
	.w1(32'hba79f7f2),
	.w2(32'hbb6d6b97),
	.w3(32'hbabb895b),
	.w4(32'hb8cb4f8d),
	.w5(32'hbad13346),
	.w6(32'hbb2bed60),
	.w7(32'h399016a6),
	.w8(32'hbaabb756),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31496b),
	.w1(32'hba0c2792),
	.w2(32'hb9a7e93b),
	.w3(32'h3a49471e),
	.w4(32'hb95e0a16),
	.w5(32'hb9a108f1),
	.w6(32'hb9f82387),
	.w7(32'hba85aee5),
	.w8(32'hba148163),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c41bf7),
	.w1(32'h37db8b1f),
	.w2(32'h3923af9d),
	.w3(32'hb9a43e23),
	.w4(32'h38933e73),
	.w5(32'h392da429),
	.w6(32'hb9832527),
	.w7(32'h39047052),
	.w8(32'h38ea6df9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ea6b),
	.w1(32'h3a3d2a33),
	.w2(32'h39359a0b),
	.w3(32'hba326a42),
	.w4(32'h3a98df1b),
	.w5(32'h3a44ac45),
	.w6(32'hb8360eec),
	.w7(32'h3a42271f),
	.w8(32'h3a1d0653),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ba4ee),
	.w1(32'h39f61cd3),
	.w2(32'hba7fdf5b),
	.w3(32'hbafdf244),
	.w4(32'h39ea1e58),
	.w5(32'hb9570b48),
	.w6(32'hbb2509a7),
	.w7(32'hb9db0bd5),
	.w8(32'hbb020b76),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa563b1),
	.w1(32'hb6992601),
	.w2(32'hbb24ee1f),
	.w3(32'hbb0266ab),
	.w4(32'hb96767cb),
	.w5(32'hbb31a60a),
	.w6(32'hba45b918),
	.w7(32'hb9a758eb),
	.w8(32'hbb1ed068),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba628b15),
	.w1(32'h38a293f9),
	.w2(32'hba1db91f),
	.w3(32'hba76433c),
	.w4(32'hb8ecae6c),
	.w5(32'hb935f8be),
	.w6(32'hb9ed7d04),
	.w7(32'h390e6ae4),
	.w8(32'hba5ba63c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0fc53),
	.w1(32'hbb61c211),
	.w2(32'hbc8539d2),
	.w3(32'hbb93c842),
	.w4(32'hbb3292cd),
	.w5(32'hbc4231a6),
	.w6(32'hba8596fd),
	.w7(32'hbabecb80),
	.w8(32'hbbb94924),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185453),
	.w1(32'h3a377aba),
	.w2(32'hbb4f64d7),
	.w3(32'hbbf7d85a),
	.w4(32'h3b751609),
	.w5(32'h3a86688f),
	.w6(32'hbbad721b),
	.w7(32'h3badde30),
	.w8(32'hba889b24),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39213b6c),
	.w1(32'hba2a48d4),
	.w2(32'hba2e3e9e),
	.w3(32'h39bd0ab7),
	.w4(32'hba82a339),
	.w5(32'hba6bccbf),
	.w6(32'h399d60d4),
	.w7(32'hb9cd6074),
	.w8(32'hba98542c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9886c43),
	.w1(32'hb896a607),
	.w2(32'h3b12a598),
	.w3(32'hb940241d),
	.w4(32'hba049ea8),
	.w5(32'h3a2fadb5),
	.w6(32'h38ee7ed8),
	.w7(32'h3a40788b),
	.w8(32'h38c46d84),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb7dbf),
	.w1(32'h3ac21503),
	.w2(32'h3a7991e9),
	.w3(32'h39b4b498),
	.w4(32'h3aa41df5),
	.w5(32'h3a58b5f3),
	.w6(32'h3ab21a6b),
	.w7(32'h3a598f2f),
	.w8(32'h3a6c48ee),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60f1ff),
	.w1(32'hba1146c7),
	.w2(32'h37cd940e),
	.w3(32'h3a618e34),
	.w4(32'hba1cb973),
	.w5(32'hb8c57bb5),
	.w6(32'hb929409c),
	.w7(32'hb8f752fc),
	.w8(32'hb63308b1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f76c6),
	.w1(32'hba9228c4),
	.w2(32'hbb16303c),
	.w3(32'hb9346c0a),
	.w4(32'hbaa29e9b),
	.w5(32'hbb2f274f),
	.w6(32'hb9c4c8cb),
	.w7(32'hbb27d9aa),
	.w8(32'hbb73963f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e696a),
	.w1(32'h3a4b1382),
	.w2(32'hb9b21991),
	.w3(32'hbb7341dc),
	.w4(32'h3a8724a4),
	.w5(32'hba9beeb6),
	.w6(32'hbaef9501),
	.w7(32'h3a94d5f0),
	.w8(32'hbb534207),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06058),
	.w1(32'hba61a0cc),
	.w2(32'hbbc376c0),
	.w3(32'hbb6dd3ec),
	.w4(32'h3a57af0b),
	.w5(32'hbb8950a2),
	.w6(32'hbb3b9e53),
	.w7(32'h3b2024e0),
	.w8(32'hba49d4dc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983a77c),
	.w1(32'hb9867979),
	.w2(32'hb9fedf85),
	.w3(32'hba00cdf9),
	.w4(32'hb96d8317),
	.w5(32'hb997ae6d),
	.w6(32'hbac9ba3d),
	.w7(32'hb990396c),
	.w8(32'hba425e87),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83fd58),
	.w1(32'hbb21d27a),
	.w2(32'hbbfbde25),
	.w3(32'hbb800e54),
	.w4(32'hbabf5d92),
	.w5(32'hbbc069f0),
	.w6(32'hbb27b751),
	.w7(32'hbae9d3b1),
	.w8(32'hbb91a6c7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95de90),
	.w1(32'hba92a09b),
	.w2(32'hbb0f638c),
	.w3(32'hba14a830),
	.w4(32'hba0ddd8c),
	.w5(32'hbac186da),
	.w6(32'h39678525),
	.w7(32'hb9efef8c),
	.w8(32'hbab3dae3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0ee0a),
	.w1(32'hba37b876),
	.w2(32'hba22d78f),
	.w3(32'h38795839),
	.w4(32'hba070f12),
	.w5(32'hba262373),
	.w6(32'hba3b0995),
	.w7(32'hba637221),
	.w8(32'hba3073e9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad31c42),
	.w1(32'hbb0c8c8b),
	.w2(32'hbaae2535),
	.w3(32'hbac48408),
	.w4(32'hbaadfdf6),
	.w5(32'hb9d959ce),
	.w6(32'hbad723f7),
	.w7(32'hba8c3d98),
	.w8(32'hba7ef680),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43a642),
	.w1(32'hb9a5e957),
	.w2(32'hb8d5d030),
	.w3(32'hb9f83ee8),
	.w4(32'hb9149c7d),
	.w5(32'hb7052253),
	.w6(32'hb92c5128),
	.w7(32'hb9c8cae2),
	.w8(32'h3805f3b3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18ff03),
	.w1(32'h3a994e88),
	.w2(32'hb9d762b9),
	.w3(32'hbae5369d),
	.w4(32'h39fb2481),
	.w5(32'hb98eb623),
	.w6(32'hba6a7347),
	.w7(32'h3a5feeb8),
	.w8(32'hb9ab610d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db686),
	.w1(32'h3b727d6b),
	.w2(32'h3a261691),
	.w3(32'hbb04be39),
	.w4(32'h3b7f14cf),
	.w5(32'h3aaf5d1e),
	.w6(32'hbb3ecb52),
	.w7(32'h3b88f614),
	.w8(32'hbac55f2b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92aab4),
	.w1(32'hba96206a),
	.w2(32'hbb89cad3),
	.w3(32'hbb21afd2),
	.w4(32'h3a472e68),
	.w5(32'hbb280a91),
	.w6(32'hbb43bd7e),
	.w7(32'h3a6633ff),
	.w8(32'hbb282a32),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6572c0),
	.w1(32'h39e141d3),
	.w2(32'h3aad9aac),
	.w3(32'hba658167),
	.w4(32'h388dae45),
	.w5(32'h3a479875),
	.w6(32'hbaca5410),
	.w7(32'hba277762),
	.w8(32'hba552d5d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97436),
	.w1(32'hb9d06153),
	.w2(32'hbb2b45e0),
	.w3(32'hbb678b92),
	.w4(32'h3abfe9ac),
	.w5(32'hba4107ed),
	.w6(32'hbb8c536a),
	.w7(32'h3a8d25dd),
	.w8(32'hbb38fa7b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa10709),
	.w1(32'hb808233b),
	.w2(32'hbb419b71),
	.w3(32'hbaca4190),
	.w4(32'h3955f272),
	.w5(32'hbb112ada),
	.w6(32'hbb096c41),
	.w7(32'hb654faa9),
	.w8(32'hba98aacf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4f6ad),
	.w1(32'h39542575),
	.w2(32'hbbfd43c7),
	.w3(32'hbbb01893),
	.w4(32'h3a8ca04c),
	.w5(32'hbbc31fcc),
	.w6(32'hbad25dab),
	.w7(32'h3b34e629),
	.w8(32'hbb5f15c3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31ecd9),
	.w1(32'h38edc438),
	.w2(32'h396d6749),
	.w3(32'h39903f2c),
	.w4(32'h3881e9f0),
	.w5(32'h39bd146b),
	.w6(32'h39d6b47e),
	.w7(32'h3a0095e1),
	.w8(32'h39b7dba9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d63bf3),
	.w1(32'h3a024d08),
	.w2(32'h39b00019),
	.w3(32'h38f82965),
	.w4(32'h39eebf83),
	.w5(32'h39be87ac),
	.w6(32'h39c2bd55),
	.w7(32'h39a81bba),
	.w8(32'h39a5ee03),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e85e),
	.w1(32'h3a6a388d),
	.w2(32'hbb260103),
	.w3(32'hbb014d3f),
	.w4(32'h3a8bcf3c),
	.w5(32'hbb358d0b),
	.w6(32'hb9b20909),
	.w7(32'h3b341a9d),
	.w8(32'hbb3c941c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79e06b),
	.w1(32'h3ab8497e),
	.w2(32'hbbc22ffe),
	.w3(32'hbb5389f2),
	.w4(32'h3a872431),
	.w5(32'hbbf01320),
	.w6(32'hba336df2),
	.w7(32'h3b7fea55),
	.w8(32'hbb367d5d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969d2c),
	.w1(32'h391d24c0),
	.w2(32'hbb6e5d10),
	.w3(32'hbb75925d),
	.w4(32'h3add013f),
	.w5(32'hbaecc1ea),
	.w6(32'hbacd52c1),
	.w7(32'h3b6e5b74),
	.w8(32'hba3bc2b0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ef8ae),
	.w1(32'hbaa7ec16),
	.w2(32'hbac88472),
	.w3(32'hbb17a50a),
	.w4(32'hbb5bda64),
	.w5(32'hbaf81a33),
	.w6(32'h3a98ce14),
	.w7(32'hbaa9205e),
	.w8(32'hbb5fae7a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fbcdc),
	.w1(32'hb9f81d01),
	.w2(32'hb9c80f4f),
	.w3(32'hbaa1794c),
	.w4(32'hba0d0b75),
	.w5(32'hb9b6042c),
	.w6(32'hb9987e25),
	.w7(32'hba1f97c7),
	.w8(32'hb91c3ac1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e9114),
	.w1(32'hb9c47d89),
	.w2(32'hb744b8be),
	.w3(32'hba2adf20),
	.w4(32'hb985f66a),
	.w5(32'h398d305f),
	.w6(32'hb9a77449),
	.w7(32'hb954bdce),
	.w8(32'hb8ef1586),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2b45e),
	.w1(32'h39364206),
	.w2(32'hbb89cbcf),
	.w3(32'hba83002f),
	.w4(32'hbb8839ec),
	.w5(32'hbbf2e64c),
	.w6(32'h3b0ecf04),
	.w7(32'hbaa81a98),
	.w8(32'hbbd52a2e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc7c6c),
	.w1(32'hbb4570e8),
	.w2(32'hbbf7fc6a),
	.w3(32'hbbbc8201),
	.w4(32'hbb188b4f),
	.w5(32'hbbc8bb77),
	.w6(32'hbb91b7a3),
	.w7(32'hbb59f92f),
	.w8(32'hbba758be),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbdbbc),
	.w1(32'h39fe95b4),
	.w2(32'hbab21da8),
	.w3(32'hbb0e8f93),
	.w4(32'hba24ac84),
	.w5(32'hba9d9759),
	.w6(32'h3aff8fbd),
	.w7(32'h3a2f0929),
	.w8(32'hbb314280),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1f8eb),
	.w1(32'h3b86f56d),
	.w2(32'h3b30414b),
	.w3(32'hbab437d6),
	.w4(32'h3b652fc7),
	.w5(32'h3ad061aa),
	.w6(32'hbac3491f),
	.w7(32'h3b7832f6),
	.w8(32'h3ad4d737),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27ad37),
	.w1(32'h39b19a51),
	.w2(32'hbb4ca986),
	.w3(32'hbb1441e9),
	.w4(32'h3af0ec23),
	.w5(32'hbab8eb9b),
	.w6(32'hbb0c7df1),
	.w7(32'h3b37b58d),
	.w8(32'h38426357),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fdec8),
	.w1(32'hb8f770bc),
	.w2(32'hb900b8f2),
	.w3(32'h3813d969),
	.w4(32'hb5cd3fe5),
	.w5(32'hb8e936fe),
	.w6(32'h38a79cf5),
	.w7(32'hb8bf863b),
	.w8(32'hb9642d57),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997604b),
	.w1(32'hb97a7424),
	.w2(32'hb9aca390),
	.w3(32'hb9572dc1),
	.w4(32'hb9e56a87),
	.w5(32'hb82366fa),
	.w6(32'hb989d327),
	.w7(32'hb8c9b031),
	.w8(32'hb913083f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba6772),
	.w1(32'hb937582d),
	.w2(32'hb991d922),
	.w3(32'hb93c6e5b),
	.w4(32'hba32609c),
	.w5(32'hbaa55da3),
	.w6(32'hb81234da),
	.w7(32'hba357208),
	.w8(32'h3a398b7a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b16f2),
	.w1(32'hba00fd6e),
	.w2(32'h39dc42b4),
	.w3(32'h39f32945),
	.w4(32'hba088f8d),
	.w5(32'hb8064b7c),
	.w6(32'hb9d26423),
	.w7(32'h3987649a),
	.w8(32'h369b0a96),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab4954),
	.w1(32'hba6e7d1e),
	.w2(32'hba76217c),
	.w3(32'h3a08c551),
	.w4(32'hba98337f),
	.w5(32'hbabe3dde),
	.w6(32'hb64039b2),
	.w7(32'hba0f8826),
	.w8(32'hbaacaea5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7f05),
	.w1(32'h39ac7095),
	.w2(32'hbb40a2ab),
	.w3(32'hbb2d333f),
	.w4(32'h3aac4de2),
	.w5(32'hbb2ab1fe),
	.w6(32'hb9727124),
	.w7(32'h3b04e316),
	.w8(32'hbae32bd2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404686),
	.w1(32'hbac60ec8),
	.w2(32'hbb513c00),
	.w3(32'hbb1d413e),
	.w4(32'hb9a1b171),
	.w5(32'hbb648558),
	.w6(32'hbb5b0635),
	.w7(32'hbaf2ec91),
	.w8(32'hbb5402e8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbcbb5),
	.w1(32'hba67489d),
	.w2(32'hbac147a9),
	.w3(32'hba45a671),
	.w4(32'hba937998),
	.w5(32'hbaa734c4),
	.w6(32'hba543248),
	.w7(32'hba8c60f6),
	.w8(32'hb8bc18f9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64ac70),
	.w1(32'hbaabeeea),
	.w2(32'hbbd0e640),
	.w3(32'hbb57c293),
	.w4(32'hbb0d74cd),
	.w5(32'hbbbbe6a3),
	.w6(32'hb9850cad),
	.w7(32'hba4b0e5b),
	.w8(32'hbbe24468),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb172352),
	.w1(32'hba91ee8b),
	.w2(32'hbb49f30e),
	.w3(32'hbaf0c2f4),
	.w4(32'hba90329c),
	.w5(32'hbb3a7bfd),
	.w6(32'hba3bf850),
	.w7(32'hba0811f2),
	.w8(32'hbae4b76f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f7dd9),
	.w1(32'hba3f21c1),
	.w2(32'hba10e85d),
	.w3(32'hba198a45),
	.w4(32'hb9fc932f),
	.w5(32'hb9d2100d),
	.w6(32'hba377043),
	.w7(32'hba6fc022),
	.w8(32'hb9d8d753),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba440d5e),
	.w1(32'hba06cb49),
	.w2(32'hbaeaf925),
	.w3(32'hbaa0c5d8),
	.w4(32'hba767df7),
	.w5(32'hbafd82a2),
	.w6(32'hba77ca56),
	.w7(32'hba99d643),
	.w8(32'hbb13f72b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c71d21),
	.w1(32'h38845f8b),
	.w2(32'h3978a0f0),
	.w3(32'h39961590),
	.w4(32'hb8be4c0f),
	.w5(32'hb97acb46),
	.w6(32'h39ee7765),
	.w7(32'h39bc153b),
	.w8(32'h37eee1cb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a190d9),
	.w1(32'hb884b528),
	.w2(32'hb8c52b73),
	.w3(32'hba373e2a),
	.w4(32'h39010887),
	.w5(32'hb8964308),
	.w6(32'h37a2232f),
	.w7(32'h3484e3c2),
	.w8(32'hb8b05d68),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1e501),
	.w1(32'hba2b1362),
	.w2(32'hba33aa19),
	.w3(32'h3894ea24),
	.w4(32'hb9b542f4),
	.w5(32'hb9fd4603),
	.w6(32'hba12edf8),
	.w7(32'hba4ea105),
	.w8(32'hb9eff3b5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce5937),
	.w1(32'h3920e163),
	.w2(32'h3965b4aa),
	.w3(32'hb936d3c2),
	.w4(32'hb886fff9),
	.w5(32'hb939ad9b),
	.w6(32'h3a361404),
	.w7(32'h3a1c9fef),
	.w8(32'hba117d77),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba770d94),
	.w1(32'hb9d2c063),
	.w2(32'hba27206d),
	.w3(32'hbb0bb774),
	.w4(32'hba7bb191),
	.w5(32'hbaa1f50b),
	.w6(32'hbb473266),
	.w7(32'hba66f910),
	.w8(32'hba773846),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bce45),
	.w1(32'hbb0278e6),
	.w2(32'hbbf15523),
	.w3(32'hbb7ad412),
	.w4(32'hba9bd1c4),
	.w5(32'hbbc5fc23),
	.w6(32'hbb013401),
	.w7(32'h3aa1c41c),
	.w8(32'hbb956ef5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd470),
	.w1(32'hbad635ef),
	.w2(32'hbba56d8b),
	.w3(32'hba47b357),
	.w4(32'hba37a5cd),
	.w5(32'hbb649da8),
	.w6(32'hbad91aa4),
	.w7(32'hb9a9b6ad),
	.w8(32'hbb12a9f6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb768c19),
	.w1(32'hbb05fde4),
	.w2(32'hbbd5f516),
	.w3(32'hbb952645),
	.w4(32'hbb210ff7),
	.w5(32'hbbc0025a),
	.w6(32'hbb0d82ec),
	.w7(32'hbb0b3678),
	.w8(32'hbbac32d7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3adde9),
	.w1(32'h381f702b),
	.w2(32'h398452b1),
	.w3(32'hba47562a),
	.w4(32'h38d1927e),
	.w5(32'h39c92aee),
	.w6(32'hb9a4987a),
	.w7(32'hb951d3cf),
	.w8(32'hb9dee14f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de158),
	.w1(32'hbaa673e7),
	.w2(32'hba8b8fc6),
	.w3(32'hb9e0c660),
	.w4(32'hba421772),
	.w5(32'hba3774d2),
	.w6(32'hba77f86b),
	.w7(32'hbab52416),
	.w8(32'hba4c62ea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a9468),
	.w1(32'hba17922b),
	.w2(32'hb9e6b408),
	.w3(32'hb9822777),
	.w4(32'hb9cd1c56),
	.w5(32'hb9d0c948),
	.w6(32'hba1060cc),
	.w7(32'hba20bccd),
	.w8(32'hb9fd871b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2ad8b),
	.w1(32'hba2ef4b0),
	.w2(32'hb9fdd377),
	.w3(32'hb951db68),
	.w4(32'hb9c64f21),
	.w5(32'hb9bd4cc3),
	.w6(32'hba343943),
	.w7(32'hba3daad3),
	.w8(32'hb9e7e732),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d06ee),
	.w1(32'hbad4d848),
	.w2(32'hbb5f3dee),
	.w3(32'hbb1b9e80),
	.w4(32'h394c887b),
	.w5(32'hba8ab9d5),
	.w6(32'hbb2d2e2f),
	.w7(32'hb92ba637),
	.w8(32'hbb028886),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910e6dd),
	.w1(32'hb9b22914),
	.w2(32'hba061302),
	.w3(32'hb9f8cd04),
	.w4(32'hb9e9e182),
	.w5(32'hba1ae5a2),
	.w6(32'hba57b069),
	.w7(32'hbab08fdc),
	.w8(32'hba5b2269),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba720231),
	.w1(32'h3962b7cf),
	.w2(32'hb9700af8),
	.w3(32'hba676170),
	.w4(32'h3a4f97ab),
	.w5(32'hba075bab),
	.w6(32'hba6ded44),
	.w7(32'hb98d0e3a),
	.w8(32'hba627f72),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48d805),
	.w1(32'hb91b8b96),
	.w2(32'h37199658),
	.w3(32'hba169026),
	.w4(32'h39123770),
	.w5(32'h39c4a234),
	.w6(32'hba8de82e),
	.w7(32'h38283556),
	.w8(32'h39f1d48e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f413a),
	.w1(32'hba825a03),
	.w2(32'hba6a040e),
	.w3(32'h3a3a1234),
	.w4(32'hba491264),
	.w5(32'hba3e63ad),
	.w6(32'hba6988b2),
	.w7(32'hba775382),
	.w8(32'hba5ddf7c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee20e6),
	.w1(32'hba713db9),
	.w2(32'hbb0e8c80),
	.w3(32'hbac6565c),
	.w4(32'hba6d721a),
	.w5(32'hbab4c27e),
	.w6(32'hb9c86f7c),
	.w7(32'hb98119ef),
	.w8(32'hbaac0b92),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7559ec),
	.w1(32'hba54d851),
	.w2(32'hba32e2be),
	.w3(32'hba832fd1),
	.w4(32'hb9d0b326),
	.w5(32'hb9321025),
	.w6(32'hba40783b),
	.w7(32'hb9ed174b),
	.w8(32'h38f85502),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817b6f),
	.w1(32'hbb560a85),
	.w2(32'hbbf7fb88),
	.w3(32'hbb3d47fa),
	.w4(32'hba6611e4),
	.w5(32'hbb1fb51e),
	.w6(32'hbb8064f0),
	.w7(32'hbabc1795),
	.w8(32'hbaec7c7c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a958c),
	.w1(32'hb9cdf900),
	.w2(32'hb8eb3087),
	.w3(32'h38262970),
	.w4(32'hba5dd99d),
	.w5(32'hba1589cd),
	.w6(32'hb9effd07),
	.w7(32'hb964831b),
	.w8(32'hba3b7b49),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73ff4a),
	.w1(32'h3b083fb7),
	.w2(32'h3b3a516e),
	.w3(32'hbb23388b),
	.w4(32'h3b4c59f5),
	.w5(32'h3b4fd478),
	.w6(32'hbb67b8ad),
	.w7(32'h3ab9fdcc),
	.w8(32'h3aea69e0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule