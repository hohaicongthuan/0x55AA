module layer_6_featuremap_118(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0182bf),
	.w1(32'hbbe7fb67),
	.w2(32'h3b18e8bb),
	.w3(32'hbb10387e),
	.w4(32'h3ba14e0d),
	.w5(32'hba57ff6d),
	.w6(32'h3ae94316),
	.w7(32'h3c3e400b),
	.w8(32'h3be3b0ce),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f3c61),
	.w1(32'h3c601896),
	.w2(32'h3c5945ab),
	.w3(32'h3b13a77a),
	.w4(32'h3b8165f1),
	.w5(32'h3b95969d),
	.w6(32'hbca107cb),
	.w7(32'hbcb84b66),
	.w8(32'hbcb948b6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85bd09),
	.w1(32'hbbcb2468),
	.w2(32'hbc8e6550),
	.w3(32'hbafe0b9d),
	.w4(32'h3bbae032),
	.w5(32'h3c0b9647),
	.w6(32'h3b4097bc),
	.w7(32'hbc0043c7),
	.w8(32'hbb3a4056),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58ea50),
	.w1(32'h3a87f0ad),
	.w2(32'hbbebbcfd),
	.w3(32'hbbe324f0),
	.w4(32'hbc60a220),
	.w5(32'hbc6bde37),
	.w6(32'hbc0ce829),
	.w7(32'hbc953598),
	.w8(32'hbc9b22a6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7bc2b),
	.w1(32'h3b7e4502),
	.w2(32'h3c9094a0),
	.w3(32'hbbbefa65),
	.w4(32'hbc343777),
	.w5(32'hbc534515),
	.w6(32'h3b93e0c0),
	.w7(32'hbb0cbf72),
	.w8(32'hbaaf346e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c884b30),
	.w1(32'h3c864435),
	.w2(32'h3ce12a97),
	.w3(32'h3cdcd927),
	.w4(32'h3d1f5b56),
	.w5(32'h3d25bba0),
	.w6(32'h3cea9f7c),
	.w7(32'h3d2e4348),
	.w8(32'h3d34c1f6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce80959),
	.w1(32'hbc404c24),
	.w2(32'hbccdafc1),
	.w3(32'hbd0d6e0e),
	.w4(32'hbd5250d7),
	.w5(32'hbd31161c),
	.w6(32'hbd1788e2),
	.w7(32'hbd6174ee),
	.w8(32'hbd3d9d67),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83ce16),
	.w1(32'h3b59bf4a),
	.w2(32'hbc44d858),
	.w3(32'h3c462d0f),
	.w4(32'h3c87eb24),
	.w5(32'h3cbdb15d),
	.w6(32'h3b92c072),
	.w7(32'h3c2c4d67),
	.w8(32'h3bb7261e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadc81b),
	.w1(32'h3c32b305),
	.w2(32'h3c767adb),
	.w3(32'hbb096305),
	.w4(32'h3bd3b1c2),
	.w5(32'h3bd4728d),
	.w6(32'h3b9202e7),
	.w7(32'hbb6a9e89),
	.w8(32'h3b3eaca8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c530b41),
	.w1(32'h3bdfb802),
	.w2(32'h3c793f28),
	.w3(32'h3cb27681),
	.w4(32'h3d0afe14),
	.w5(32'h3cf0e141),
	.w6(32'h3cab878d),
	.w7(32'h3d0535bd),
	.w8(32'h3cd9b57e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ddb5f),
	.w1(32'hbb1e081a),
	.w2(32'h3a1257c7),
	.w3(32'h3b940ebd),
	.w4(32'h3bd8c685),
	.w5(32'hba25ca6f),
	.w6(32'h3b7aec2e),
	.w7(32'h3c057c07),
	.w8(32'h3b56771f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a704293),
	.w1(32'hbb37e0fa),
	.w2(32'h3ac74ded),
	.w3(32'hb9bd9347),
	.w4(32'h39631e23),
	.w5(32'h3b9f31ae),
	.w6(32'h3b853159),
	.w7(32'h3b9a79db),
	.w8(32'h3c315bf6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b69b),
	.w1(32'hbb8fac78),
	.w2(32'hbb639591),
	.w3(32'hbb8e2252),
	.w4(32'hbbd173e9),
	.w5(32'hbbf919e6),
	.w6(32'hbba724d0),
	.w7(32'hbba4070c),
	.w8(32'hbbfeb6d1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c312),
	.w1(32'hbbe56e9d),
	.w2(32'hbbd6ae16),
	.w3(32'h3a08fa90),
	.w4(32'h3b2e6214),
	.w5(32'h3bab5ec9),
	.w6(32'hbafda3bf),
	.w7(32'hbb7268e5),
	.w8(32'hbb448a0a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfc74b),
	.w1(32'h3bbea74c),
	.w2(32'h3c2c1735),
	.w3(32'hbb9a57d3),
	.w4(32'hbaec2957),
	.w5(32'hbb2fd91e),
	.w6(32'hba9689ac),
	.w7(32'h3a66c35e),
	.w8(32'h397c123f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf07f1d),
	.w1(32'hbacc679d),
	.w2(32'h3bd49ddb),
	.w3(32'h3ba174f2),
	.w4(32'h3c1cfe9c),
	.w5(32'h3c3e4bcc),
	.w6(32'h3b2e7a9d),
	.w7(32'h3bf53c3d),
	.w8(32'h3c37d974),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2120cd),
	.w1(32'hbb8992b9),
	.w2(32'hbbb5fa4d),
	.w3(32'hbc14b00f),
	.w4(32'hbc1c8869),
	.w5(32'hbba3dfd6),
	.w6(32'hbb6bb5fb),
	.w7(32'hbb9bda41),
	.w8(32'hbb5b0ea5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac1f7e),
	.w1(32'hbb568ded),
	.w2(32'h3c0d3e21),
	.w3(32'h3a8275f5),
	.w4(32'h3c60a6e3),
	.w5(32'h3c19516e),
	.w6(32'h3b2a2b03),
	.w7(32'h3c6b51ce),
	.w8(32'h3c25190c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e171),
	.w1(32'hbbc0ee34),
	.w2(32'hbc3caba6),
	.w3(32'hbbc66229),
	.w4(32'hbc25dd54),
	.w5(32'hbbf5f5b5),
	.w6(32'hbbc2174d),
	.w7(32'hbc3d2845),
	.w8(32'hbc3814e6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5004),
	.w1(32'h3b262812),
	.w2(32'hbb0d8cc7),
	.w3(32'hbc1afbb0),
	.w4(32'hbc2ca9cf),
	.w5(32'hbc247c19),
	.w6(32'h3a33c6e6),
	.w7(32'hbb692eac),
	.w8(32'h3b15c754),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b5513),
	.w1(32'hba8dbf21),
	.w2(32'hbaf614dc),
	.w3(32'hbba633df),
	.w4(32'hbbafdf41),
	.w5(32'hbb25cd69),
	.w6(32'hbbe385d4),
	.w7(32'hbc146d14),
	.w8(32'hbbbd5f95),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b389f7),
	.w1(32'h3bee0d77),
	.w2(32'h3c8cac70),
	.w3(32'h3b9c581b),
	.w4(32'h3b847a68),
	.w5(32'h3bbf8760),
	.w6(32'h3b3e767b),
	.w7(32'h3c0b3c54),
	.w8(32'h3be86438),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7902ce),
	.w1(32'h3c445e62),
	.w2(32'h3c9d5d01),
	.w3(32'hbbcc4e9e),
	.w4(32'h3b055af9),
	.w5(32'hba1a9497),
	.w6(32'h3bec8031),
	.w7(32'h3c3dac72),
	.w8(32'hba71bd6e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ca1d),
	.w1(32'h3bc76f9d),
	.w2(32'hbc0591c6),
	.w3(32'h3a322473),
	.w4(32'h3b3a063f),
	.w5(32'hbc3bbb2e),
	.w6(32'hbaa7b11a),
	.w7(32'hbbea8f9b),
	.w8(32'hbc242bc4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1b1a),
	.w1(32'hbaeb2b96),
	.w2(32'hbb19e691),
	.w3(32'hbb93fee8),
	.w4(32'h3a1a73b6),
	.w5(32'h39e4323d),
	.w6(32'h38ec909f),
	.w7(32'hbb032ed3),
	.w8(32'h3bc9affd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab701f7),
	.w1(32'hbb847d96),
	.w2(32'h3b3a1b2b),
	.w3(32'hbbe74e6b),
	.w4(32'hbbbe646c),
	.w5(32'hbae442cc),
	.w6(32'hbb99633d),
	.w7(32'hbaf97e9d),
	.w8(32'h3afb156a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e5f8),
	.w1(32'hbbb0af3f),
	.w2(32'hbb50dd2a),
	.w3(32'hbb6922d1),
	.w4(32'hbb9052b9),
	.w5(32'hbbee1fdd),
	.w6(32'hbb7d07ea),
	.w7(32'hba563509),
	.w8(32'hbacd9206),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf6db9),
	.w1(32'hbc0fa299),
	.w2(32'hbcab3654),
	.w3(32'hbcc7f558),
	.w4(32'hbd11af0b),
	.w5(32'hbcd0bd88),
	.w6(32'hbcc51a93),
	.w7(32'hbd1d412b),
	.w8(32'hbcec86b6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f0080),
	.w1(32'hbb51dc32),
	.w2(32'hbb913d82),
	.w3(32'hba8e1b1b),
	.w4(32'hbad0a5a3),
	.w5(32'h39bde545),
	.w6(32'hbb56a00c),
	.w7(32'hbb852245),
	.w8(32'hbb117645),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38329e),
	.w1(32'hbc117a34),
	.w2(32'h3b894bb0),
	.w3(32'hbc4a39d7),
	.w4(32'hbc157cb2),
	.w5(32'h3b6d4532),
	.w6(32'hbc67423c),
	.w7(32'hbc0b59c9),
	.w8(32'hbb96c13d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d52d),
	.w1(32'h39be8b29),
	.w2(32'h3c4afa07),
	.w3(32'h3bb1fa1e),
	.w4(32'h3c3b401d),
	.w5(32'h3c4ae4ce),
	.w6(32'h3c1dcced),
	.w7(32'h3c9be898),
	.w8(32'h3ccaf3e0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce50aa5),
	.w1(32'hbb91eb7d),
	.w2(32'h3c85c836),
	.w3(32'hb8dc5165),
	.w4(32'hbb421c9f),
	.w5(32'hbb6a73bc),
	.w6(32'hbc50e6fd),
	.w7(32'hbaa3b2ba),
	.w8(32'hbaea9b67),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b0b1e),
	.w1(32'h3bfd0548),
	.w2(32'h3ba210f5),
	.w3(32'hbba49f1c),
	.w4(32'hbc06156b),
	.w5(32'hbc040505),
	.w6(32'hbbca3710),
	.w7(32'hbc2a8a1b),
	.w8(32'h3abc95de),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2442a4),
	.w1(32'h3ae76329),
	.w2(32'hbb703a92),
	.w3(32'hbb51f58e),
	.w4(32'h3c1b8242),
	.w5(32'h3bad6b6f),
	.w6(32'h3b872a0b),
	.w7(32'hbb89449a),
	.w8(32'h3b12de89),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb67d),
	.w1(32'h3c16101b),
	.w2(32'h3c4f5a5c),
	.w3(32'h3c50593d),
	.w4(32'h3c8d7b6f),
	.w5(32'h3c877307),
	.w6(32'h3c4907c5),
	.w7(32'h3c8492c8),
	.w8(32'h3c77f9a8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c401b47),
	.w1(32'h3bd0c7e4),
	.w2(32'hbb56360d),
	.w3(32'h38bb6cbc),
	.w4(32'hbc2dd403),
	.w5(32'hbc53eba5),
	.w6(32'hbb5d2061),
	.w7(32'hbbf73961),
	.w8(32'hb9481ed7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba849d),
	.w1(32'hbadb7770),
	.w2(32'h3c42d876),
	.w3(32'hbb6b18a1),
	.w4(32'h3ba2ba3a),
	.w5(32'hbaa668c5),
	.w6(32'h3b430101),
	.w7(32'h3c91f679),
	.w8(32'h3c3195ce),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba32faf),
	.w1(32'hbba704f1),
	.w2(32'hbc0318c9),
	.w3(32'hbbfbccf2),
	.w4(32'hbc377588),
	.w5(32'hbc13f49f),
	.w6(32'hbc0fb28c),
	.w7(32'hbc451725),
	.w8(32'hbc294caa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd22f8c),
	.w1(32'hbc3fc569),
	.w2(32'hbbef860c),
	.w3(32'hbb29f221),
	.w4(32'h3b43ca7d),
	.w5(32'h3b034ae3),
	.w6(32'hbba2a162),
	.w7(32'h38a370f7),
	.w8(32'hbb801dd6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b555e),
	.w1(32'hbcc0e228),
	.w2(32'hbbbc33a9),
	.w3(32'h3c2f1630),
	.w4(32'hba06d450),
	.w5(32'hbc49880e),
	.w6(32'hbc3795ae),
	.w7(32'hbb642662),
	.w8(32'hba8c6e43),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fd937),
	.w1(32'h3c114d84),
	.w2(32'h3bdd6685),
	.w3(32'h3c00f8ec),
	.w4(32'hba840404),
	.w5(32'hbb8b26b9),
	.w6(32'h3c55e4f8),
	.w7(32'h3bad6b00),
	.w8(32'hbc13fca2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eada4),
	.w1(32'h3b463226),
	.w2(32'hbb84e27a),
	.w3(32'hbb921ad1),
	.w4(32'hbc466711),
	.w5(32'hbc2641fa),
	.w6(32'hbbc9167d),
	.w7(32'hbc7e1cd0),
	.w8(32'hbc52c5e7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee917),
	.w1(32'h3b4f0668),
	.w2(32'h3c871e50),
	.w3(32'h3a0c0ba0),
	.w4(32'h3c2e8bd3),
	.w5(32'h3c14206d),
	.w6(32'h3ba9a3f4),
	.w7(32'h3c92b6a8),
	.w8(32'h3c754c96),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ea108),
	.w1(32'hbbb2a7c0),
	.w2(32'hb9c50f6d),
	.w3(32'h3c16abfd),
	.w4(32'h3b509d00),
	.w5(32'h3bc6201f),
	.w6(32'hb9434584),
	.w7(32'h3a5d236a),
	.w8(32'h3ad1bf35),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e54d3),
	.w1(32'hbaeb26fe),
	.w2(32'hbbaf3cd0),
	.w3(32'hbc0a977e),
	.w4(32'hbc1d3c28),
	.w5(32'hbc26d2d8),
	.w6(32'hbb8df1bd),
	.w7(32'hbbdcb71c),
	.w8(32'hbc0c815a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe043c7),
	.w1(32'hbbf08ce0),
	.w2(32'hba55312b),
	.w3(32'h3b99af57),
	.w4(32'h3b33aef9),
	.w5(32'hbc03b8bb),
	.w6(32'h3b0ba262),
	.w7(32'hb9cb9fdc),
	.w8(32'hba183702),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c662037),
	.w1(32'h3c7cb171),
	.w2(32'h3c05072a),
	.w3(32'hba0f16b6),
	.w4(32'h3b5e6fe6),
	.w5(32'hbbe86bd3),
	.w6(32'hbae62fa4),
	.w7(32'hbbc1d7a8),
	.w8(32'hbc4ad043),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80b88a),
	.w1(32'h3bde7633),
	.w2(32'h3bd27fa3),
	.w3(32'hbc2abd77),
	.w4(32'hbc1bb66a),
	.w5(32'hbc24fd4a),
	.w6(32'h3a35b8d5),
	.w7(32'h3a59ff0a),
	.w8(32'h3ba5488a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2983f3),
	.w1(32'h3bbb2cfd),
	.w2(32'h3b42a43b),
	.w3(32'h3b535e69),
	.w4(32'h3b452be5),
	.w5(32'h3b801710),
	.w6(32'h3b132273),
	.w7(32'h39fb944c),
	.w8(32'h3b034897),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962e99),
	.w1(32'h39d10dae),
	.w2(32'h3c11f2d1),
	.w3(32'h3b04af83),
	.w4(32'hb972e2e5),
	.w5(32'hbbfc6019),
	.w6(32'hba4c1e01),
	.w7(32'h3bc536e5),
	.w8(32'h3bf557a6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e60c1),
	.w1(32'h3b47e1ba),
	.w2(32'hbbba71ef),
	.w3(32'hbb1190ff),
	.w4(32'hbc41b705),
	.w5(32'hbbdf1877),
	.w6(32'hbc0ea186),
	.w7(32'hbcaeecc5),
	.w8(32'hbc93c206),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb379a2),
	.w1(32'h3bc532d7),
	.w2(32'hbc1dbe1f),
	.w3(32'hbb0a04c0),
	.w4(32'hbc956257),
	.w5(32'hbc4fa222),
	.w6(32'hbae7f56e),
	.w7(32'hbca5a3f8),
	.w8(32'hbc4d2719),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31a10d),
	.w1(32'h3c1c09eb),
	.w2(32'hbc34f53d),
	.w3(32'hbb91434f),
	.w4(32'hbcb502e2),
	.w5(32'hbc8aeb97),
	.w6(32'hbbaed26b),
	.w7(32'hbcde9755),
	.w8(32'hbcc942b3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf70dbd),
	.w1(32'hbc19c47e),
	.w2(32'hbce8c099),
	.w3(32'hbd06701d),
	.w4(32'hbd4df218),
	.w5(32'hbd395126),
	.w6(32'hbd0167c3),
	.w7(32'hbd5f0d3e),
	.w8(32'hbd4db753),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5cb9b),
	.w1(32'h3ab46bdf),
	.w2(32'hbbbd833e),
	.w3(32'h3a5696e4),
	.w4(32'hbbd0ab0b),
	.w5(32'hbba14189),
	.w6(32'hbc5c669e),
	.w7(32'hbcbd5ccd),
	.w8(32'hbcc2aacd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0b2f),
	.w1(32'hba81afce),
	.w2(32'hba0f5621),
	.w3(32'h3a8493ee),
	.w4(32'h3974be32),
	.w5(32'hb9c4dfa6),
	.w6(32'hba067671),
	.w7(32'hba1a0f18),
	.w8(32'hba2996d3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25633b),
	.w1(32'hba469c68),
	.w2(32'hbaa42464),
	.w3(32'hbb51f2ce),
	.w4(32'hbb88a6fd),
	.w5(32'hbb6e8e49),
	.w6(32'hbb2f386c),
	.w7(32'hbb5d7768),
	.w8(32'hbb542826),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f5fe),
	.w1(32'h3aa79a29),
	.w2(32'h3a4d7bd0),
	.w3(32'h3912057f),
	.w4(32'hbaeb31d4),
	.w5(32'hbaae9785),
	.w6(32'h3a66cfa9),
	.w7(32'hbab11dda),
	.w8(32'h3a18f13d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af66cba),
	.w1(32'h37b2a774),
	.w2(32'h39347247),
	.w3(32'h3aa4c455),
	.w4(32'h3ad11d1d),
	.w5(32'h3aaef665),
	.w6(32'h3a4038d6),
	.w7(32'h3a791796),
	.w8(32'h3a369579),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d3a19e),
	.w1(32'hba0a2f91),
	.w2(32'h3addf29a),
	.w3(32'hba1120dc),
	.w4(32'h3ab56866),
	.w5(32'h3b190191),
	.w6(32'hbab5e6b5),
	.w7(32'h39294df9),
	.w8(32'h39920784),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fd5e7),
	.w1(32'hb99af7a2),
	.w2(32'hb9bd5e51),
	.w3(32'h3a2750e6),
	.w4(32'h3a67eb51),
	.w5(32'h39b875c4),
	.w6(32'h3a92543e),
	.w7(32'h3a900c91),
	.w8(32'h3a412616),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba084a6f),
	.w1(32'hbaeef175),
	.w2(32'hbac6a8e2),
	.w3(32'hbb201edd),
	.w4(32'hbafa37f6),
	.w5(32'hbb4a397d),
	.w6(32'hbb0ea318),
	.w7(32'hba378130),
	.w8(32'hbb27feb3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d2c0a),
	.w1(32'hbb4d1771),
	.w2(32'hbb00f672),
	.w3(32'h3ab584c7),
	.w4(32'h3b04994f),
	.w5(32'h3b4d8ad3),
	.w6(32'h3a3e7648),
	.w7(32'h3b40bb37),
	.w8(32'h3aa33dcf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6cdf2),
	.w1(32'h3a9a05d9),
	.w2(32'h390afefd),
	.w3(32'h3c183b96),
	.w4(32'h3c1f3e32),
	.w5(32'h3c0f7bd5),
	.w6(32'h3bb0d483),
	.w7(32'h3bae7feb),
	.w8(32'h3ba952fe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule