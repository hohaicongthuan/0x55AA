module layer_10_featuremap_411(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05c356),
	.w1(32'h3b86ac56),
	.w2(32'h381b2f30),
	.w3(32'hbc3a84dc),
	.w4(32'h3b3fdf2c),
	.w5(32'h39bf546f),
	.w6(32'h3a8c67eb),
	.w7(32'h3a8ccbc0),
	.w8(32'hbb83abb2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844c7e),
	.w1(32'hbc1e3437),
	.w2(32'hbc8060cc),
	.w3(32'hb99c0a29),
	.w4(32'hbb3d2be0),
	.w5(32'hbc3f2854),
	.w6(32'hba68ad8f),
	.w7(32'hbbac3923),
	.w8(32'hbc5818d2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0440d5),
	.w1(32'hbbc21d81),
	.w2(32'h3a13cd36),
	.w3(32'hbb87291e),
	.w4(32'hbc50cb33),
	.w5(32'hbc76ffe7),
	.w6(32'hbb19859f),
	.w7(32'hb91e7a50),
	.w8(32'hbc0b4e15),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27fa1a),
	.w1(32'hbbd2f77d),
	.w2(32'hbc676909),
	.w3(32'hbc69787a),
	.w4(32'hbc3f5b38),
	.w5(32'hbbefde88),
	.w6(32'hbbec6272),
	.w7(32'hbc509736),
	.w8(32'hbcab3912),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48f2d4),
	.w1(32'hbb617421),
	.w2(32'h3bf6d432),
	.w3(32'hbcb02fa7),
	.w4(32'hb94b6a9d),
	.w5(32'h3c278b0b),
	.w6(32'hbc4dd0de),
	.w7(32'hbb251776),
	.w8(32'h3b369761),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59dac),
	.w1(32'h3b2c7e55),
	.w2(32'h3bbba92c),
	.w3(32'h3b13f49b),
	.w4(32'h3b975c88),
	.w5(32'h3c149ddc),
	.w6(32'h3ae64b28),
	.w7(32'h3ba15176),
	.w8(32'h3b83b0e2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5458),
	.w1(32'hbbe4b52a),
	.w2(32'hbba9aa2f),
	.w3(32'h3be48422),
	.w4(32'h3b2ea616),
	.w5(32'h3d1e9523),
	.w6(32'h3b8076fe),
	.w7(32'hbb9c725f),
	.w8(32'h3be8699a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab08e09),
	.w1(32'hbb56a783),
	.w2(32'h3c382694),
	.w3(32'h3cb96a3b),
	.w4(32'h3b703c61),
	.w5(32'h3c960ed2),
	.w6(32'hbb342950),
	.w7(32'hba6e4ab1),
	.w8(32'h3b41b323),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0682),
	.w1(32'h3888938a),
	.w2(32'h3b5db79e),
	.w3(32'h38cac1e8),
	.w4(32'h3ab28270),
	.w5(32'h3ca28fd1),
	.w6(32'hbb9bbfa9),
	.w7(32'h3be6ea10),
	.w8(32'h3c57734f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1248cc),
	.w1(32'h3ba5961c),
	.w2(32'h3b217c6d),
	.w3(32'h3c801cd6),
	.w4(32'hbbab3ebb),
	.w5(32'hbb5a913f),
	.w6(32'h3c3c175c),
	.w7(32'h3b1b9608),
	.w8(32'h3b5f0148),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81be5d),
	.w1(32'hbb858e7a),
	.w2(32'hbb49ca45),
	.w3(32'h3b5b3cac),
	.w4(32'hbb170aa0),
	.w5(32'hbb8d965d),
	.w6(32'h3bb685d8),
	.w7(32'h3bf1d9f6),
	.w8(32'h3c70d974),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213c2b),
	.w1(32'h38b5b442),
	.w2(32'h3abda1bd),
	.w3(32'h3a63f308),
	.w4(32'hbb9e4c25),
	.w5(32'h3b12e8f8),
	.w6(32'h3bff377f),
	.w7(32'h3c07243f),
	.w8(32'h3c178ae9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e1a7),
	.w1(32'h3ab6e0c9),
	.w2(32'hbc4f24b1),
	.w3(32'h3c386ae6),
	.w4(32'hbc21c997),
	.w5(32'hbbdcd715),
	.w6(32'h3b843a4b),
	.w7(32'hbc140c7b),
	.w8(32'hbc119a6f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eeaed),
	.w1(32'hbc06fa45),
	.w2(32'h3baec506),
	.w3(32'hbc0b90c7),
	.w4(32'hbc87c471),
	.w5(32'hbc4bd4c8),
	.w6(32'hba18b9d1),
	.w7(32'hbb46ac37),
	.w8(32'h3aa3c0ec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b7819),
	.w1(32'h3b567ce5),
	.w2(32'hba5e7ef7),
	.w3(32'hbbf7df00),
	.w4(32'h3b9453c4),
	.w5(32'h3b0cb37d),
	.w6(32'hba3aa58a),
	.w7(32'h3b827b0c),
	.w8(32'h3c175d92),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb533aca),
	.w1(32'h394fc152),
	.w2(32'h3ab23706),
	.w3(32'hbc04b509),
	.w4(32'h3badfa35),
	.w5(32'h3b93e7c5),
	.w6(32'hbb76fe17),
	.w7(32'h3be6f755),
	.w8(32'h3bc26f0b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00c6d7),
	.w1(32'h3b11c2c1),
	.w2(32'h3c15e0ea),
	.w3(32'hbaaec628),
	.w4(32'hb9f58bf9),
	.w5(32'h3a021d71),
	.w6(32'hbba608f9),
	.w7(32'hbb67be46),
	.w8(32'h3b8f4761),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cad21),
	.w1(32'hba17e4b3),
	.w2(32'hba97e9d9),
	.w3(32'hb90aa7a0),
	.w4(32'hbaa9cfee),
	.w5(32'hbbb732be),
	.w6(32'h3a582050),
	.w7(32'h3b79a89a),
	.w8(32'h39770bf6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39015779),
	.w1(32'hbbcd4806),
	.w2(32'hbab55db9),
	.w3(32'hbc0bb520),
	.w4(32'hbbdbc9ae),
	.w5(32'h3b9642ee),
	.w6(32'h3b851ba4),
	.w7(32'h38bbe2d6),
	.w8(32'h3c415284),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c8df),
	.w1(32'hbb91f6da),
	.w2(32'hbbd1273e),
	.w3(32'h3bc024a7),
	.w4(32'h3b045906),
	.w5(32'hbbb116c0),
	.w6(32'h3a72ba12),
	.w7(32'h3b86ad95),
	.w8(32'h3adaaf8b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e6afa),
	.w1(32'h3bffb2c9),
	.w2(32'h3c186d64),
	.w3(32'h3ac5efed),
	.w4(32'h3c186a3f),
	.w5(32'h3acdaa34),
	.w6(32'hbad9d97b),
	.w7(32'h3a5f59f6),
	.w8(32'hbb6766e6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fff25),
	.w1(32'h3b8ac791),
	.w2(32'h3b05cd34),
	.w3(32'hb9702ec9),
	.w4(32'h3bb82f85),
	.w5(32'hbade9bdf),
	.w6(32'hbb63ad3f),
	.w7(32'hbbb72255),
	.w8(32'hbb1330a9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba574661),
	.w1(32'hba396b41),
	.w2(32'hbbc92090),
	.w3(32'hbc1d5873),
	.w4(32'hbc00dccf),
	.w5(32'hbab4817d),
	.w6(32'h3b6f60c5),
	.w7(32'hbb3a6819),
	.w8(32'h3ba89829),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fbe60),
	.w1(32'h3bb1cecc),
	.w2(32'h3c02ad65),
	.w3(32'h3bfa566a),
	.w4(32'hbb05510d),
	.w5(32'h3b714555),
	.w6(32'hba327f01),
	.w7(32'h3bbe1063),
	.w8(32'h3b8624c2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9c84),
	.w1(32'h3b8677e5),
	.w2(32'hbbe86403),
	.w3(32'hbb1c08fc),
	.w4(32'h3b80e313),
	.w5(32'hb92a1c9e),
	.w6(32'h3ba25886),
	.w7(32'hbb7e7800),
	.w8(32'h3b2e79a5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9155),
	.w1(32'h3c161ab8),
	.w2(32'h3bc97f20),
	.w3(32'h3c1e60a7),
	.w4(32'h3bf5c347),
	.w5(32'hbba3f616),
	.w6(32'hbaee5319),
	.w7(32'h3afa838a),
	.w8(32'hbadb19cc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6564),
	.w1(32'hbba990d9),
	.w2(32'hbac0ef09),
	.w3(32'hbb2b6c0e),
	.w4(32'h3a91f7c9),
	.w5(32'h3c058978),
	.w6(32'hba46dabd),
	.w7(32'hbb56e6d9),
	.w8(32'h3aacd52d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c7b27),
	.w1(32'h3bb0999e),
	.w2(32'h3aa2a401),
	.w3(32'h3b9d6dbc),
	.w4(32'h3bee10bf),
	.w5(32'hba81a2e2),
	.w6(32'h3be235ab),
	.w7(32'hbae009c5),
	.w8(32'hbb719b6a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a407f),
	.w1(32'hbbb62fbc),
	.w2(32'h3aa6e676),
	.w3(32'h3a92e586),
	.w4(32'h3b86d7e1),
	.w5(32'hbc1365d1),
	.w6(32'hbc0ddcd7),
	.w7(32'hbc077395),
	.w8(32'hbb86671c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeb94f),
	.w1(32'h3af29736),
	.w2(32'hba43f5f3),
	.w3(32'hbbb78567),
	.w4(32'hba95a8ca),
	.w5(32'h3af029ee),
	.w6(32'h3bc473d0),
	.w7(32'h3b7210fc),
	.w8(32'hbb41036f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107117),
	.w1(32'hbb903ad6),
	.w2(32'hbc1c87ff),
	.w3(32'h3acc9eb1),
	.w4(32'hbc12ad68),
	.w5(32'hbbffba4f),
	.w6(32'hbbdcce26),
	.w7(32'h3b8d8779),
	.w8(32'h3bdfd6ef),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe22f0e),
	.w1(32'hbbe4d29d),
	.w2(32'hbc0530f2),
	.w3(32'hbb8d31ea),
	.w4(32'hbb0b422a),
	.w5(32'hbbb963d4),
	.w6(32'h3b31426a),
	.w7(32'hbb52c567),
	.w8(32'hba315fab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04d8a),
	.w1(32'h3b1a088b),
	.w2(32'hbb41ae2c),
	.w3(32'hbb81d9c9),
	.w4(32'h3bc5f7be),
	.w5(32'h3a5ac83a),
	.w6(32'hbc02873c),
	.w7(32'hbb275176),
	.w8(32'hbb377101),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f0352),
	.w1(32'h3b8151f1),
	.w2(32'hba9860b8),
	.w3(32'h3b72a208),
	.w4(32'h3c58e436),
	.w5(32'h3cb0aa8f),
	.w6(32'h3b080d7b),
	.w7(32'h3c0fb6bf),
	.w8(32'h3c656ee6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a552),
	.w1(32'hba171265),
	.w2(32'hbb8b1afc),
	.w3(32'h3bf2fbe2),
	.w4(32'hbbb38818),
	.w5(32'hbc3e964e),
	.w6(32'h3a431e91),
	.w7(32'h39f627aa),
	.w8(32'hbbad932d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3657),
	.w1(32'h3befbe17),
	.w2(32'hbc5deb36),
	.w3(32'hbbaa22fb),
	.w4(32'hbc2f6ff1),
	.w5(32'hbc9a6ac7),
	.w6(32'h3b592c26),
	.w7(32'hbc02a4db),
	.w8(32'hbc1c713f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd557e8),
	.w1(32'hbc0addab),
	.w2(32'hbb9212f7),
	.w3(32'hbc720b6b),
	.w4(32'hbc06395f),
	.w5(32'h3baed38c),
	.w6(32'hbaaad0cd),
	.w7(32'h3b57d377),
	.w8(32'h3cb7ed8e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ccd2e),
	.w1(32'hbbd5d48e),
	.w2(32'hbc72fb90),
	.w3(32'h3c23b985),
	.w4(32'hbb8822c7),
	.w5(32'hbc96aeb5),
	.w6(32'h3b71af56),
	.w7(32'h394b7813),
	.w8(32'hbbd2818e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efcfc),
	.w1(32'h3b8a275f),
	.w2(32'h3add0aad),
	.w3(32'h3b90b2e3),
	.w4(32'hbc5001cf),
	.w5(32'hbbdb23f8),
	.w6(32'h3ba82478),
	.w7(32'hbb0e2097),
	.w8(32'h3bfca467),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10bf4f),
	.w1(32'hbb55b32d),
	.w2(32'hbb4b1491),
	.w3(32'h3acaffff),
	.w4(32'hbb273f6d),
	.w5(32'hbbe5bf6a),
	.w6(32'hb9cfe7f6),
	.w7(32'hbb6f3abf),
	.w8(32'hbba3ba05),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebef3),
	.w1(32'h3a50ff38),
	.w2(32'hbae0af6b),
	.w3(32'hbb4f0269),
	.w4(32'hbbd69170),
	.w5(32'hbba1a577),
	.w6(32'hbc060fdf),
	.w7(32'h3acf1735),
	.w8(32'hbb91627b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52046d),
	.w1(32'hbc7ee937),
	.w2(32'hbc519b1c),
	.w3(32'hbbca6d87),
	.w4(32'hbbcec0aa),
	.w5(32'h3b8e1735),
	.w6(32'h3ae12794),
	.w7(32'hbb9c1ef3),
	.w8(32'h3c1f4891),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c4741),
	.w1(32'hbc4ec913),
	.w2(32'hbc9fe489),
	.w3(32'h3c352162),
	.w4(32'hbc4f59e7),
	.w5(32'hbc3bc395),
	.w6(32'h3bc7a60a),
	.w7(32'hbbb42152),
	.w8(32'hbc5721fa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f8a6),
	.w1(32'h3c089147),
	.w2(32'h3b94b2a9),
	.w3(32'hbc95298b),
	.w4(32'h3bb46cc2),
	.w5(32'hbc310b8a),
	.w6(32'hbc20e452),
	.w7(32'hb9b3ec8b),
	.w8(32'hbc050362),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023254),
	.w1(32'hbb9e3320),
	.w2(32'h3b88bfa3),
	.w3(32'h3b4a7910),
	.w4(32'h3a8753ac),
	.w5(32'h3cc4e232),
	.w6(32'h3bc27e44),
	.w7(32'hba28deaa),
	.w8(32'h3b89bd90),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa478a),
	.w1(32'h3a5dfb64),
	.w2(32'hba291b6e),
	.w3(32'hba8711ee),
	.w4(32'h3b8ba9b1),
	.w5(32'h3abf9e7f),
	.w6(32'hbbf3d3b1),
	.w7(32'h3a9a83d7),
	.w8(32'h39e056b8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d657),
	.w1(32'hbb1f234c),
	.w2(32'hbc06e607),
	.w3(32'hbaf9f25f),
	.w4(32'hbbec5b93),
	.w5(32'hbbf0ec81),
	.w6(32'hbb87497d),
	.w7(32'h3a419ce5),
	.w8(32'hbae4c039),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35a099),
	.w1(32'h3b6a3517),
	.w2(32'h3b25a4ad),
	.w3(32'hbbb315e7),
	.w4(32'hbaded88d),
	.w5(32'h3b9c9c8d),
	.w6(32'hbb084210),
	.w7(32'hba99c820),
	.w8(32'h3ac9bfa3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc61d3f),
	.w1(32'hbb009e1a),
	.w2(32'h3c0bcae8),
	.w3(32'h3b8864f4),
	.w4(32'hbb193cc9),
	.w5(32'h3c84721e),
	.w6(32'hbb2cd351),
	.w7(32'hbafbce56),
	.w8(32'hbac40332),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab5a22),
	.w1(32'h3c474a82),
	.w2(32'h3ab9b80c),
	.w3(32'h3b37a29b),
	.w4(32'h3b041bba),
	.w5(32'hbbd3c28a),
	.w6(32'hbaef22c9),
	.w7(32'hbadbb2ac),
	.w8(32'hbc15a20e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb59b94),
	.w1(32'hbb679de8),
	.w2(32'hbb742817),
	.w3(32'hbc21911c),
	.w4(32'hbbf37d4e),
	.w5(32'hbb4edfeb),
	.w6(32'hbc3c5159),
	.w7(32'hbae3db10),
	.w8(32'hbb9e1594),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd4d0),
	.w1(32'hbb466b78),
	.w2(32'hbadfc577),
	.w3(32'hbb182e1a),
	.w4(32'h3ac8982c),
	.w5(32'hbb9f882e),
	.w6(32'h3b03bd28),
	.w7(32'h3ac0e024),
	.w8(32'hb92875aa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bece7),
	.w1(32'hbbffc932),
	.w2(32'h3c0a68fc),
	.w3(32'hbb20c95c),
	.w4(32'h3bf9ff07),
	.w5(32'h3ce64661),
	.w6(32'h3b747522),
	.w7(32'h3b9f1b3f),
	.w8(32'h3ca25f41),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ad256),
	.w1(32'h3ab6e6df),
	.w2(32'h3c83f7ac),
	.w3(32'h3c8b8956),
	.w4(32'h3c541705),
	.w5(32'h3c60b9f0),
	.w6(32'h3b93d57f),
	.w7(32'h3aa50441),
	.w8(32'h3bcb05dc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced912),
	.w1(32'hbc29667a),
	.w2(32'hbc9229d7),
	.w3(32'h3c7627ab),
	.w4(32'hbba08f3a),
	.w5(32'hbc399cfc),
	.w6(32'h3b8ac734),
	.w7(32'hbb6d8ac7),
	.w8(32'hbbc823b2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaead2ff),
	.w1(32'hbc756885),
	.w2(32'hbc9dfa88),
	.w3(32'h3ac942d3),
	.w4(32'hbc3d32b4),
	.w5(32'hbccfcd5c),
	.w6(32'hbb026c13),
	.w7(32'hbc4b5765),
	.w8(32'hbca19d87),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e725),
	.w1(32'hbb238ef0),
	.w2(32'hbb763f6f),
	.w3(32'hbc038d25),
	.w4(32'hbb7f1d95),
	.w5(32'hbb64260d),
	.w6(32'hbc092050),
	.w7(32'hbbc8e4d9),
	.w8(32'hbbab46d6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb063f5f),
	.w1(32'h3b8547a2),
	.w2(32'hbb4d8e29),
	.w3(32'h3bc81651),
	.w4(32'h3b77c4f2),
	.w5(32'h3a45b589),
	.w6(32'h3b1a2c17),
	.w7(32'h37f853ba),
	.w8(32'h3bf2f7f8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b44cb),
	.w1(32'h3ba04f33),
	.w2(32'hbbcc6f96),
	.w3(32'h3b33c89e),
	.w4(32'h3bdfe67d),
	.w5(32'hbc7a6fbc),
	.w6(32'h3c33b515),
	.w7(32'hbaf09c24),
	.w8(32'hbbef4fde),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2178),
	.w1(32'h3b20a2d3),
	.w2(32'h3ab9ae0b),
	.w3(32'h3b1f9a8e),
	.w4(32'h3b27e5f7),
	.w5(32'h3b604b0e),
	.w6(32'h3ba2dd53),
	.w7(32'h3c134ed5),
	.w8(32'h3b3736a3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c9d27),
	.w1(32'h3b9287c3),
	.w2(32'h39072a70),
	.w3(32'h3c4aa08b),
	.w4(32'h3b842b2e),
	.w5(32'hbc51fa1e),
	.w6(32'hbb48859b),
	.w7(32'hba86a1c4),
	.w8(32'h3a0c0442),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93826),
	.w1(32'hbc634b8e),
	.w2(32'hbbcc9665),
	.w3(32'hbb9095a4),
	.w4(32'hbbe2ed21),
	.w5(32'h3a433971),
	.w6(32'h3bf39e37),
	.w7(32'hba6e9172),
	.w8(32'h3b66f613),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be13c3d),
	.w1(32'h3bac7c98),
	.w2(32'hbb9d9633),
	.w3(32'h3ae62794),
	.w4(32'h3b466356),
	.w5(32'hbb1e0c04),
	.w6(32'hbbae4b3f),
	.w7(32'h3b05a3d4),
	.w8(32'hbbcc19ad),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32cd67),
	.w1(32'hbc0d0d3c),
	.w2(32'hbaed517d),
	.w3(32'hbc965da0),
	.w4(32'hbc00f9aa),
	.w5(32'hbb85757d),
	.w6(32'hbc4bf414),
	.w7(32'h3a3c0ab9),
	.w8(32'h3b1fc403),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66a041),
	.w1(32'h3c48767e),
	.w2(32'h3c0530fc),
	.w3(32'hbab8d55b),
	.w4(32'h3bad6d0b),
	.w5(32'hbc0ea283),
	.w6(32'hb97c532c),
	.w7(32'h3b8409f0),
	.w8(32'hbc0d5c3e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1369bf),
	.w1(32'hbb1a536e),
	.w2(32'h3c2060ba),
	.w3(32'hbbc4f9c1),
	.w4(32'h3aadd00e),
	.w5(32'h3ccac1d1),
	.w6(32'h3ae6a973),
	.w7(32'h3bfe99ee),
	.w8(32'h3c89a1d4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee5c0d),
	.w1(32'h3bbd8401),
	.w2(32'h3b9e639b),
	.w3(32'h3c33c4e6),
	.w4(32'h3c1249ff),
	.w5(32'h3bf01b88),
	.w6(32'h3b9df7d9),
	.w7(32'h3b2683cd),
	.w8(32'h3a5a8c19),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86ef10),
	.w1(32'hbb2ce3d9),
	.w2(32'h3bab27c4),
	.w3(32'hb9b0501f),
	.w4(32'h3c697f5a),
	.w5(32'h3ba9edbd),
	.w6(32'hbbdf05ab),
	.w7(32'h3c2733ce),
	.w8(32'hbb92e05d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811d988),
	.w1(32'h3c09496b),
	.w2(32'hbb578082),
	.w3(32'hbc615d8b),
	.w4(32'h3bf4c886),
	.w5(32'hb9b8bd25),
	.w6(32'hbc8a71f7),
	.w7(32'hbafd6696),
	.w8(32'h3b05f5a8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b59f),
	.w1(32'h3bcd42b9),
	.w2(32'hbb29d010),
	.w3(32'h39a8606b),
	.w4(32'hbb1c07c7),
	.w5(32'hbb5c8029),
	.w6(32'hbaed5d07),
	.w7(32'h3b78ff42),
	.w8(32'h3b2fca59),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f99c1),
	.w1(32'h3ab8cc96),
	.w2(32'hbaed342b),
	.w3(32'h3acab54c),
	.w4(32'hbb44f7ef),
	.w5(32'h3bd55f1d),
	.w6(32'h3ba3719e),
	.w7(32'h3bec4755),
	.w8(32'h3b7fb79e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9760a23),
	.w1(32'hbb60f853),
	.w2(32'hbbe5714e),
	.w3(32'hbb9c4987),
	.w4(32'hbc65e1cf),
	.w5(32'hbc2ab913),
	.w6(32'h3b929a6c),
	.w7(32'h394ea801),
	.w8(32'hbb74418c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e8a0),
	.w1(32'hbb8b7e7b),
	.w2(32'hb6fc0129),
	.w3(32'hbc2e29f2),
	.w4(32'hbc025f58),
	.w5(32'h3c1f7c2d),
	.w6(32'hbbeed04d),
	.w7(32'hbb19f90e),
	.w8(32'h3b82567d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc4978),
	.w1(32'hba8c3653),
	.w2(32'hba362608),
	.w3(32'hbc2f021a),
	.w4(32'h3c3dbd99),
	.w5(32'hbc3f1d2f),
	.w6(32'hbba1b96c),
	.w7(32'h3abcf6aa),
	.w8(32'hb952b235),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9717),
	.w1(32'hba152e61),
	.w2(32'h3b9e9bd1),
	.w3(32'h3a1b943e),
	.w4(32'h3b07aa85),
	.w5(32'hbb011ca0),
	.w6(32'hbaec6bce),
	.w7(32'h3ae36e94),
	.w8(32'h3b1585ca),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f642),
	.w1(32'h3b0a71c0),
	.w2(32'hbbc28f55),
	.w3(32'h3b05a89e),
	.w4(32'h3c0178fc),
	.w5(32'hbb3b83b1),
	.w6(32'hbbbbb826),
	.w7(32'hbc5e9f50),
	.w8(32'hbbcde40d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdfdb5),
	.w1(32'h3b3c9934),
	.w2(32'h3b88de92),
	.w3(32'hbc11c67c),
	.w4(32'h3b303acd),
	.w5(32'hbbf21aa9),
	.w6(32'hbb28c2ef),
	.w7(32'hbab01932),
	.w8(32'hbb3e7c9e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d6b89),
	.w1(32'hbba47456),
	.w2(32'hbb66de8b),
	.w3(32'h3bb0253e),
	.w4(32'hbb3aac9b),
	.w5(32'h3d090514),
	.w6(32'h3b1ddfaf),
	.w7(32'hbb5fc282),
	.w8(32'h3b83fe5a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79c437),
	.w1(32'hbb9f05c1),
	.w2(32'hbb569ce1),
	.w3(32'hbbe52e83),
	.w4(32'hbbfca5ee),
	.w5(32'h3cc61369),
	.w6(32'hbb024374),
	.w7(32'hbc299e7b),
	.w8(32'h3b5958fb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb678a81),
	.w1(32'hbad54091),
	.w2(32'hbc08cc2f),
	.w3(32'hbbedb6bf),
	.w4(32'hbb7b3647),
	.w5(32'hbca274ef),
	.w6(32'hba935a46),
	.w7(32'h3c063657),
	.w8(32'hbb3bbb95),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e04ea),
	.w1(32'h3aed9077),
	.w2(32'h397cd876),
	.w3(32'hb889ed3f),
	.w4(32'hbbbbf48a),
	.w5(32'h3b854385),
	.w6(32'hbb8d80e6),
	.w7(32'hbbc90053),
	.w8(32'hba3651fe),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae2a13),
	.w1(32'h3b1f5f27),
	.w2(32'h3ab82fd2),
	.w3(32'h3c27c843),
	.w4(32'h3b623ebc),
	.w5(32'hbb6810b9),
	.w6(32'h3bcf7d56),
	.w7(32'hba89f2ab),
	.w8(32'hbac8510b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcdc9d),
	.w1(32'hba3f8a9a),
	.w2(32'hbb1d7b18),
	.w3(32'h3b9116e0),
	.w4(32'hbc02b90b),
	.w5(32'h3b56ef97),
	.w6(32'h3b97bedf),
	.w7(32'h3bd09e51),
	.w8(32'h3b90cbaf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f05f),
	.w1(32'hbb7349f5),
	.w2(32'hba013f42),
	.w3(32'hbbcea48e),
	.w4(32'hbc247f7d),
	.w5(32'hbab32d6c),
	.w6(32'hbbabe9ad),
	.w7(32'hba1da33a),
	.w8(32'hb8ceb612),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad669c0),
	.w1(32'hbba9e9c6),
	.w2(32'h3b8ddbcf),
	.w3(32'hbc14df2c),
	.w4(32'h3a851b46),
	.w5(32'hbbc09258),
	.w6(32'h3b68f9d0),
	.w7(32'h3a8378bc),
	.w8(32'hb911b60c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9768c2),
	.w1(32'hbbca865e),
	.w2(32'hbc3848fd),
	.w3(32'h3b9e383c),
	.w4(32'hba8aa27d),
	.w5(32'hbc38dcad),
	.w6(32'h390ab33c),
	.w7(32'hbb95ee9a),
	.w8(32'hb9ecc8e5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc174098),
	.w1(32'hbbdd10e1),
	.w2(32'hbc39b16b),
	.w3(32'hbb6a26c4),
	.w4(32'h39f5e3f5),
	.w5(32'h3cfcad09),
	.w6(32'hba06ab03),
	.w7(32'h3bebe181),
	.w8(32'h3c166de3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b911d),
	.w1(32'hba9c1ba3),
	.w2(32'hbb00b7ab),
	.w3(32'hbc8a80e3),
	.w4(32'h3c8b5574),
	.w5(32'h3c612896),
	.w6(32'hbbed147a),
	.w7(32'h3c9a102e),
	.w8(32'h3c9eb5de),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e838f),
	.w1(32'hbc22f58f),
	.w2(32'hbbea7d5b),
	.w3(32'hbb38f620),
	.w4(32'hbbf6a794),
	.w5(32'hbbd514b9),
	.w6(32'h3b73466e),
	.w7(32'hbc01b6b3),
	.w8(32'hbc1dfd17),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2b96),
	.w1(32'hbc3aad78),
	.w2(32'hbbe005f3),
	.w3(32'hbc065de8),
	.w4(32'hbc4c9de4),
	.w5(32'h3bff4c5a),
	.w6(32'hbc10cc63),
	.w7(32'hbc5099b1),
	.w8(32'hbc1d2624),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc36123),
	.w1(32'hbc180e08),
	.w2(32'hbb941c32),
	.w3(32'hbbff514c),
	.w4(32'hbb0c6e57),
	.w5(32'h3b7146f6),
	.w6(32'hbc1ce7d0),
	.w7(32'h3606775c),
	.w8(32'h3b2a0333),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbe862),
	.w1(32'h3b4db795),
	.w2(32'h3b3a88f2),
	.w3(32'hbc1e1654),
	.w4(32'h3c09d29a),
	.w5(32'h3bb2fb73),
	.w6(32'hba9d1dde),
	.w7(32'hbb127827),
	.w8(32'hbb09c59f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7224),
	.w1(32'hbb91b335),
	.w2(32'hbbac1b5d),
	.w3(32'h3ad9f5be),
	.w4(32'hbbc7a229),
	.w5(32'hbc498048),
	.w6(32'hbb80101d),
	.w7(32'h3b79afd8),
	.w8(32'h3b05eec3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2448),
	.w1(32'hbbbec8bb),
	.w2(32'hbb32be00),
	.w3(32'hbab09b3a),
	.w4(32'hba182072),
	.w5(32'h3b38947f),
	.w6(32'h38e394d7),
	.w7(32'hbb1dc74c),
	.w8(32'h3b3b7673),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b1ba7),
	.w1(32'hb9c5654c),
	.w2(32'hbaf4b5f6),
	.w3(32'hba2d1474),
	.w4(32'hbbbe0d33),
	.w5(32'hbc16272b),
	.w6(32'h3bc7784a),
	.w7(32'h3a23a5b9),
	.w8(32'hbbdafe02),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd58ca1),
	.w1(32'hbc0179a2),
	.w2(32'hba880901),
	.w3(32'h3b96d445),
	.w4(32'hb9db4c5e),
	.w5(32'hbcd2b431),
	.w6(32'hbb3af685),
	.w7(32'hbbb33a99),
	.w8(32'hbbadd19f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0697d6),
	.w1(32'hbb43aee4),
	.w2(32'h3bf20b70),
	.w3(32'h3c69e36b),
	.w4(32'h3c92d431),
	.w5(32'hbc1b29fe),
	.w6(32'h3babb46b),
	.w7(32'h3c5f6a5e),
	.w8(32'h3bd8c51a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac4aac),
	.w1(32'hbb0f71cc),
	.w2(32'h3c2ee6f9),
	.w3(32'h3c6b5fa1),
	.w4(32'hbc065190),
	.w5(32'h3af3f33a),
	.w6(32'h3c6da31c),
	.w7(32'hbc151ef2),
	.w8(32'h39690aab),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b500240),
	.w1(32'h3b1421e5),
	.w2(32'hbb713e38),
	.w3(32'h3bba9fea),
	.w4(32'hbbf4be81),
	.w5(32'h3a49a85b),
	.w6(32'hb8345a75),
	.w7(32'hbbb6b500),
	.w8(32'hbb0a2a96),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f81c),
	.w1(32'h3a2ed6a1),
	.w2(32'hbba8af36),
	.w3(32'hbbae451a),
	.w4(32'h3abc0272),
	.w5(32'hbba9955e),
	.w6(32'hbbaa247f),
	.w7(32'hb946d9fa),
	.w8(32'hbb1260bd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa148de),
	.w1(32'hbc05a459),
	.w2(32'hbaf18138),
	.w3(32'hbbb85e11),
	.w4(32'hbb3e3119),
	.w5(32'hbae07e5d),
	.w6(32'hbb62e2a9),
	.w7(32'hbbd0ff58),
	.w8(32'hbb2b2f0a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a850041),
	.w1(32'hbb39e04c),
	.w2(32'h3c212d7e),
	.w3(32'hbb785023),
	.w4(32'h3bcae408),
	.w5(32'h3bfcc43b),
	.w6(32'h3b6b1d62),
	.w7(32'hba8ac45c),
	.w8(32'h3c0c0d56),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc36d46),
	.w1(32'hbb09b76d),
	.w2(32'hbbac2376),
	.w3(32'h3cac5163),
	.w4(32'hbc85e3ce),
	.w5(32'hbc8b2467),
	.w6(32'h3bd926c6),
	.w7(32'hbbfcc238),
	.w8(32'hbc2408f7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183340),
	.w1(32'h3b54002d),
	.w2(32'h3bb05e19),
	.w3(32'hbc0cce9f),
	.w4(32'hba4f554c),
	.w5(32'h3c062081),
	.w6(32'hbb84cea1),
	.w7(32'h3ac0fae0),
	.w8(32'h3bc24186),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ece04),
	.w1(32'h3c046c08),
	.w2(32'h3c1118b7),
	.w3(32'h3b68a7b8),
	.w4(32'h38ab9e50),
	.w5(32'h3bbfa92b),
	.w6(32'hbbbcd5e4),
	.w7(32'h3c1c25b6),
	.w8(32'h3c556428),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a4f7c),
	.w1(32'h3b7d39d9),
	.w2(32'hba88b319),
	.w3(32'h3ba2d0e5),
	.w4(32'h3b6836fd),
	.w5(32'hbb3e4884),
	.w6(32'h39c29ce6),
	.w7(32'hbad0be87),
	.w8(32'hbba08565),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b21e),
	.w1(32'h3b6c4232),
	.w2(32'hbb24cbc9),
	.w3(32'h3b3bb9f0),
	.w4(32'h3b410139),
	.w5(32'h3c664174),
	.w6(32'h3b1d78aa),
	.w7(32'hbb5f6735),
	.w8(32'h3baa504e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb397219),
	.w1(32'hbbf4c8db),
	.w2(32'hbbf3477d),
	.w3(32'hbc5b0fc4),
	.w4(32'hbc422ffc),
	.w5(32'hbb9e214f),
	.w6(32'hbbbbeb9a),
	.w7(32'hbb035530),
	.w8(32'hbc15d263),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134a51),
	.w1(32'h3bd1af09),
	.w2(32'h3c55620f),
	.w3(32'hbbf9f4c7),
	.w4(32'h3c27251d),
	.w5(32'hbbe64788),
	.w6(32'hbc025fd7),
	.w7(32'h3c84b850),
	.w8(32'h3c007bea),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36dac1),
	.w1(32'h3bc09dcc),
	.w2(32'h3be722c3),
	.w3(32'h3c47f0cc),
	.w4(32'h3b36cda0),
	.w5(32'hbc11ae7b),
	.w6(32'hbac83962),
	.w7(32'hbb9c259e),
	.w8(32'hbbc02335),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc162c1b),
	.w1(32'h3ae52b53),
	.w2(32'hbb27d52c),
	.w3(32'h3be22290),
	.w4(32'hb9e1ddc0),
	.w5(32'h38473048),
	.w6(32'hbc09356f),
	.w7(32'h3b096f86),
	.w8(32'hb94679a0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934d228),
	.w1(32'h3aaf32cb),
	.w2(32'h3a013b7c),
	.w3(32'hbaee8c62),
	.w4(32'h3afb1179),
	.w5(32'hbc13873f),
	.w6(32'h39b5de26),
	.w7(32'h3c047861),
	.w8(32'h3b59585e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cc00),
	.w1(32'h3b03d8fe),
	.w2(32'hbbb25099),
	.w3(32'h3b63a9bd),
	.w4(32'h3c8dcff7),
	.w5(32'hbcb274a8),
	.w6(32'h3bd9624f),
	.w7(32'h3c3034b5),
	.w8(32'hbb94d8f9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c086575),
	.w1(32'hbb338a4f),
	.w2(32'hbc082ccc),
	.w3(32'h3c57bfb5),
	.w4(32'h3b81a81a),
	.w5(32'hba5402eb),
	.w6(32'h3b0f1cfd),
	.w7(32'hbac3c879),
	.w8(32'h3b166bae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1dcd),
	.w1(32'hbbaf327c),
	.w2(32'hba8d4181),
	.w3(32'h3b97841e),
	.w4(32'hbc20659f),
	.w5(32'h3ca42401),
	.w6(32'h3b7967da),
	.w7(32'hb9f5223b),
	.w8(32'h3c635e67),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977564),
	.w1(32'hbbacd63a),
	.w2(32'h3aeb2da5),
	.w3(32'h375b0530),
	.w4(32'hbc023bc4),
	.w5(32'h3b8bf325),
	.w6(32'h3a811b2f),
	.w7(32'hbb82a09f),
	.w8(32'hbaae0def),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90e157),
	.w1(32'h3b127d06),
	.w2(32'hbb783d4c),
	.w3(32'h3bc3026c),
	.w4(32'h3c76fb81),
	.w5(32'hbb947e69),
	.w6(32'h3b9be0e9),
	.w7(32'h3b30e3e8),
	.w8(32'h3ba07bb0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cca6ee),
	.w1(32'hbbaed08d),
	.w2(32'hbbaff943),
	.w3(32'h3b892aef),
	.w4(32'hbb21ed30),
	.w5(32'hbbeb014e),
	.w6(32'h3b6d5ff6),
	.w7(32'h3bacf9ad),
	.w8(32'h3a2138e6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5ffe),
	.w1(32'h3b595f51),
	.w2(32'h3bf16030),
	.w3(32'hba8f0eeb),
	.w4(32'h3b8e7de9),
	.w5(32'hbc019de8),
	.w6(32'h3bccf62d),
	.w7(32'h3b5842a1),
	.w8(32'h3b36c2bc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bb35),
	.w1(32'hbb944624),
	.w2(32'h3bf6fc33),
	.w3(32'hbba5a263),
	.w4(32'hbc7af70f),
	.w5(32'h3cd65903),
	.w6(32'hbad0b0ae),
	.w7(32'hbc0ec3df),
	.w8(32'h3bf7dca1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31648),
	.w1(32'hbb802899),
	.w2(32'hb986baf9),
	.w3(32'hbbc13778),
	.w4(32'hbbb1ff60),
	.w5(32'h3a21d224),
	.w6(32'h3a2b92a1),
	.w7(32'hbc0fdb04),
	.w8(32'hbae059f7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7acb),
	.w1(32'hbbb27c8d),
	.w2(32'hbc0a5a69),
	.w3(32'hba74f3a7),
	.w4(32'hbaa27ce5),
	.w5(32'hbb95e2b0),
	.w6(32'hba1438dd),
	.w7(32'hba8a954b),
	.w8(32'h3a9dfe25),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38871f16),
	.w1(32'hbba43a11),
	.w2(32'hbb858f4f),
	.w3(32'hbb220121),
	.w4(32'hbb25d5a7),
	.w5(32'hbc029c1c),
	.w6(32'hbaa4b00c),
	.w7(32'h3a219389),
	.w8(32'hba307e43),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11333d),
	.w1(32'h3bc55411),
	.w2(32'hba961742),
	.w3(32'hbb0551bf),
	.w4(32'h3cabace7),
	.w5(32'hbd1a0d64),
	.w6(32'hbbe90b51),
	.w7(32'h3c5febed),
	.w8(32'hbc61673b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c9c2),
	.w1(32'h3ae6a081),
	.w2(32'hbb361daf),
	.w3(32'h3cc58a28),
	.w4(32'h3b73e0ae),
	.w5(32'hbc56a2cd),
	.w6(32'h3b484871),
	.w7(32'h3ba67e3d),
	.w8(32'h3ab676c6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1aa1e),
	.w1(32'h3bbe5a16),
	.w2(32'hbb00f0c6),
	.w3(32'hba545a59),
	.w4(32'hbbeb437e),
	.w5(32'h3a257199),
	.w6(32'hbbb32d8a),
	.w7(32'hbaff5e4f),
	.w8(32'h3b818a04),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe55a5f),
	.w1(32'h3b9e9fc0),
	.w2(32'hbbb5b632),
	.w3(32'hbc031d25),
	.w4(32'hba8094cb),
	.w5(32'hbbe650c4),
	.w6(32'hbbb1ad94),
	.w7(32'hba4b4675),
	.w8(32'hbaaf924b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba269e29),
	.w1(32'h3b6fb8ee),
	.w2(32'hbb3a29b5),
	.w3(32'hbb31eaa9),
	.w4(32'hba82e6e2),
	.w5(32'hbb30b729),
	.w6(32'h3b95c8ef),
	.w7(32'h3a947f3f),
	.w8(32'h3baff9b8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a363506),
	.w1(32'h3aed3b6b),
	.w2(32'h3b5f0c28),
	.w3(32'h3be89599),
	.w4(32'hba7bd7a9),
	.w5(32'h3be5eac8),
	.w6(32'h3bd34df9),
	.w7(32'hb9d514d4),
	.w8(32'h3b93432a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d81a),
	.w1(32'hbc9885d4),
	.w2(32'hbc94e4eb),
	.w3(32'hbb7db819),
	.w4(32'hbc87bb99),
	.w5(32'hbc68a9d7),
	.w6(32'hbb633703),
	.w7(32'hbc46e766),
	.w8(32'hbc86ecbe),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc391f29),
	.w1(32'hbb8b6a7f),
	.w2(32'hbc200bca),
	.w3(32'hbc837a68),
	.w4(32'h3bccd164),
	.w5(32'h3a705e11),
	.w6(32'hbc959aeb),
	.w7(32'hbc871f2f),
	.w8(32'h3be422b7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d00b1),
	.w1(32'hbacad6ef),
	.w2(32'hbb51782f),
	.w3(32'hbc2f573e),
	.w4(32'hbb0d293e),
	.w5(32'h3d0f3fa2),
	.w6(32'hbb0fb10f),
	.w7(32'h3b39a904),
	.w8(32'h3c5c3a71),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1620df),
	.w1(32'h3af06160),
	.w2(32'h3ba9d567),
	.w3(32'hbb12a2f0),
	.w4(32'h3bb1f4ac),
	.w5(32'hbbed8795),
	.w6(32'h3af7af10),
	.w7(32'h3bf618c6),
	.w8(32'h3a1c0e92),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f280),
	.w1(32'h3b31c130),
	.w2(32'hba672b3a),
	.w3(32'h3c956142),
	.w4(32'h3c075e12),
	.w5(32'hbc4c9be6),
	.w6(32'h3b27fc3c),
	.w7(32'h3c07098a),
	.w8(32'h3adc4884),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156e30),
	.w1(32'hba1944ca),
	.w2(32'h3b93548f),
	.w3(32'h3ab5acf2),
	.w4(32'h3c457d74),
	.w5(32'h3b0ac1d6),
	.w6(32'h3ab6be64),
	.w7(32'hbb28c321),
	.w8(32'h3c310c7b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb2640),
	.w1(32'h3beca409),
	.w2(32'h3b58a83c),
	.w3(32'h3c42ccb7),
	.w4(32'h3c4ad3f6),
	.w5(32'h3c518184),
	.w6(32'h3c8deca8),
	.w7(32'hba436c84),
	.w8(32'h3a1948de),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7288c),
	.w1(32'hbbe33d7e),
	.w2(32'h3b474141),
	.w3(32'hbbe51101),
	.w4(32'hbb60ae95),
	.w5(32'hbc339b6d),
	.w6(32'h3b2e6fff),
	.w7(32'hbb896b09),
	.w8(32'hbb484fc9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92eea4),
	.w1(32'h3c052ff9),
	.w2(32'h3b96b903),
	.w3(32'h3c41dd74),
	.w4(32'h3b9839f5),
	.w5(32'h3c27066b),
	.w6(32'h3a9105ea),
	.w7(32'h3c796d39),
	.w8(32'h3c980e69),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11397e),
	.w1(32'hba9c9f91),
	.w2(32'h3b32e840),
	.w3(32'hbbbd3191),
	.w4(32'h3b7cb574),
	.w5(32'hbc0f0d35),
	.w6(32'hbbaa5a88),
	.w7(32'h3bc73671),
	.w8(32'h38a726b0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17f4f1),
	.w1(32'hbb8cd744),
	.w2(32'h3bddf9a2),
	.w3(32'hbac813fc),
	.w4(32'hbb9174dc),
	.w5(32'hbc86ec8b),
	.w6(32'hbb3b4138),
	.w7(32'hbc32d4be),
	.w8(32'hbc6bcf0d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfefe80),
	.w1(32'h3ba7d8e7),
	.w2(32'hbc4ce890),
	.w3(32'h3c0b217f),
	.w4(32'hbc699c06),
	.w5(32'h3cd7d1d1),
	.w6(32'h3af43389),
	.w7(32'hbc5414a0),
	.w8(32'hbb1d9ecd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717426),
	.w1(32'h3a9f269d),
	.w2(32'h3ba66302),
	.w3(32'hbc485497),
	.w4(32'h3b8f3c43),
	.w5(32'hbc02f971),
	.w6(32'hbc092f55),
	.w7(32'h3bd6c89c),
	.w8(32'hbc2d00f4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd8d3),
	.w1(32'h3ab6220d),
	.w2(32'h3c298011),
	.w3(32'h3c121e3b),
	.w4(32'h3bc7af6e),
	.w5(32'h3b3b242a),
	.w6(32'hbb512ea8),
	.w7(32'h3af84626),
	.w8(32'h3b909765),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1eee),
	.w1(32'hbb17b831),
	.w2(32'hb99bf008),
	.w3(32'h3c292200),
	.w4(32'hbbd993c0),
	.w5(32'h3b619605),
	.w6(32'h3b2aa99f),
	.w7(32'hbc007257),
	.w8(32'hbbacc8c2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9675c6),
	.w1(32'hbba80f01),
	.w2(32'hbaa3464d),
	.w3(32'hbb4ec2a3),
	.w4(32'hbc1bc81d),
	.w5(32'hbbeeeea5),
	.w6(32'h3a980146),
	.w7(32'hbae8d924),
	.w8(32'hbbeb8b0c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133f1a),
	.w1(32'hbb173ffe),
	.w2(32'h3a8dec8b),
	.w3(32'h3b8c2ab7),
	.w4(32'hbb212bb9),
	.w5(32'h3c34d69e),
	.w6(32'hbaf68cc2),
	.w7(32'h39c434dd),
	.w8(32'h3c39cc77),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384057ad),
	.w1(32'h3b581615),
	.w2(32'h3ba1b721),
	.w3(32'hbbe17a05),
	.w4(32'h3bfa55f1),
	.w5(32'hbc918fc3),
	.w6(32'hba132cf2),
	.w7(32'h3bddde7e),
	.w8(32'hbbad8d4b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971412),
	.w1(32'hbc063c75),
	.w2(32'hbc1c4ef5),
	.w3(32'h3c407d34),
	.w4(32'hbc1cd2ac),
	.w5(32'hbc1b81a0),
	.w6(32'h3b557b04),
	.w7(32'h3bc0e3a4),
	.w8(32'hbc2d0b23),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae0489),
	.w1(32'h3a6b0864),
	.w2(32'h3a56b280),
	.w3(32'hbc3e4995),
	.w4(32'h3bda74a1),
	.w5(32'hbc4c756a),
	.w6(32'hbc066c0a),
	.w7(32'h3b8ffdf7),
	.w8(32'hbbf7800c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb7fd),
	.w1(32'hbb142346),
	.w2(32'hbb7b4f26),
	.w3(32'h3ab1eaec),
	.w4(32'hbb3f6b36),
	.w5(32'hbc2cdd41),
	.w6(32'hbb1734f8),
	.w7(32'hb9da3e57),
	.w8(32'h3b2c9971),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d559),
	.w1(32'h3bf8c479),
	.w2(32'h3c1ce83a),
	.w3(32'h3840394b),
	.w4(32'hbaa70a2c),
	.w5(32'h3adb69f5),
	.w6(32'h3a933613),
	.w7(32'hbb84d5ee),
	.w8(32'h3b0eb447),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf701e0),
	.w1(32'h3b5d4e93),
	.w2(32'hbbd244cf),
	.w3(32'hbbc03d09),
	.w4(32'h3bbe39d6),
	.w5(32'hbbacd5de),
	.w6(32'hbba7a942),
	.w7(32'h3bb85494),
	.w8(32'hbb87f3b2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa77f),
	.w1(32'hbb79383d),
	.w2(32'hbbb585b1),
	.w3(32'hbb8c4687),
	.w4(32'hba874d8a),
	.w5(32'h3befa51b),
	.w6(32'hbbde2b28),
	.w7(32'hbb77fe5f),
	.w8(32'hba0bc275),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9e4a),
	.w1(32'h3c1b8a4a),
	.w2(32'h3b345f07),
	.w3(32'hbbea7724),
	.w4(32'h3a86f8cb),
	.w5(32'hbb0c5800),
	.w6(32'h3baabd02),
	.w7(32'h3afe4201),
	.w8(32'h3a3823ef),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26160e),
	.w1(32'hbb5d9771),
	.w2(32'hbbbab808),
	.w3(32'hbc08136a),
	.w4(32'h3c9c14ed),
	.w5(32'hbc2f480a),
	.w6(32'hbbba5059),
	.w7(32'h3b4c40e6),
	.w8(32'hbb220901),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8235),
	.w1(32'hbb911b56),
	.w2(32'hbbc26499),
	.w3(32'h3c1da225),
	.w4(32'hbbdbbed4),
	.w5(32'hb781b1ba),
	.w6(32'h3c20ed12),
	.w7(32'hbb84a921),
	.w8(32'hb9eec8a8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc268720),
	.w1(32'h3bd6396c),
	.w2(32'h3b68a75d),
	.w3(32'hbc6284c6),
	.w4(32'hba3850fb),
	.w5(32'hbc19de6e),
	.w6(32'hbc433a87),
	.w7(32'hbbdddc26),
	.w8(32'hbb4de391),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2bbed),
	.w1(32'hbaaba362),
	.w2(32'hbb15f1fc),
	.w3(32'h3bf6eaa7),
	.w4(32'hbaf3deb9),
	.w5(32'hbc2c92e1),
	.w6(32'h3b8dd418),
	.w7(32'hbc0992a2),
	.w8(32'hbc57078c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d49e48),
	.w1(32'hbc257d7f),
	.w2(32'hbb3644ed),
	.w3(32'hba73aab4),
	.w4(32'hbac4902e),
	.w5(32'h3ad4580d),
	.w6(32'h3a1be24a),
	.w7(32'hbbbbd5e3),
	.w8(32'hbb65e66d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3271),
	.w1(32'hbbc6d951),
	.w2(32'hbb5b02e4),
	.w3(32'hb8a0230b),
	.w4(32'hbc0d2e2d),
	.w5(32'h3d005e28),
	.w6(32'hbae68f78),
	.w7(32'hbc3f4c3e),
	.w8(32'h3bab3bf7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95cc0a),
	.w1(32'hbb59d224),
	.w2(32'hb926039e),
	.w3(32'hbc4c72c9),
	.w4(32'hbbbf7d5b),
	.w5(32'h3bcdda34),
	.w6(32'hbb9bb8ec),
	.w7(32'hbc120451),
	.w8(32'hbc475a5a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9045227),
	.w1(32'hbc66f2a4),
	.w2(32'hbc3daae3),
	.w3(32'hbbe2ee2c),
	.w4(32'hbc4fffc8),
	.w5(32'hbc87e196),
	.w6(32'hbb31c4d8),
	.w7(32'hbbce122f),
	.w8(32'hbbf6f233),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b3e6),
	.w1(32'hbb4f243a),
	.w2(32'hbbc86883),
	.w3(32'hbbe9ebd5),
	.w4(32'hbc16958b),
	.w5(32'hbc0026d2),
	.w6(32'hbbe375db),
	.w7(32'h3b5200c4),
	.w8(32'hbc21ff5f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb97312),
	.w1(32'hbb73c600),
	.w2(32'hbb4b67d5),
	.w3(32'h3adc7051),
	.w4(32'hbc4b8c3d),
	.w5(32'h3c915360),
	.w6(32'hb92a00ee),
	.w7(32'hbbb11b6b),
	.w8(32'h3c29a5ef),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b107f8e),
	.w1(32'hbba594ae),
	.w2(32'hbc20179c),
	.w3(32'h3954e1e0),
	.w4(32'hbb93f906),
	.w5(32'hbc6ed624),
	.w6(32'hb9642d66),
	.w7(32'h3a09b285),
	.w8(32'hbc0838fb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba435c5),
	.w1(32'hbbf83790),
	.w2(32'hbb024695),
	.w3(32'hbb6572ac),
	.w4(32'hbc4fb7b3),
	.w5(32'h3d382e35),
	.w6(32'h3a8323e1),
	.w7(32'hbc43d725),
	.w8(32'h3bce7fab),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4022c5),
	.w1(32'h3b95c68a),
	.w2(32'h3c0aae83),
	.w3(32'hbc658793),
	.w4(32'h3c3bfdb0),
	.w5(32'hbc99e29d),
	.w6(32'hbb29d49f),
	.w7(32'h3bc828f1),
	.w8(32'hbb708199),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb9f46),
	.w1(32'h3bd6e6a2),
	.w2(32'h3b537601),
	.w3(32'h3cae0758),
	.w4(32'hbb2270e3),
	.w5(32'h3d599515),
	.w6(32'h3be85662),
	.w7(32'h3b40dc39),
	.w8(32'h3cafe07f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc317),
	.w1(32'hbb383c60),
	.w2(32'h3b77f8fb),
	.w3(32'hbc2880b7),
	.w4(32'hbc8aefd6),
	.w5(32'h3c613faf),
	.w6(32'hba82d209),
	.w7(32'h398fb760),
	.w8(32'h3aee140c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49950e),
	.w1(32'hbb696f61),
	.w2(32'h3bf79cc4),
	.w3(32'hb9e1731d),
	.w4(32'h3b4c8660),
	.w5(32'h3b751d77),
	.w6(32'hbac180a6),
	.w7(32'h3b22f942),
	.w8(32'h3beb1466),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82551a),
	.w1(32'h3b79f160),
	.w2(32'hba7c7bcc),
	.w3(32'h3c1a75c7),
	.w4(32'hbc483475),
	.w5(32'h3d2d5548),
	.w6(32'h3c206a08),
	.w7(32'hbbb72a6d),
	.w8(32'h3c835dae),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb2a4),
	.w1(32'h3ab22081),
	.w2(32'h3aa84afa),
	.w3(32'hbb9e0a5f),
	.w4(32'h3a4541f0),
	.w5(32'h36a11417),
	.w6(32'h3bcef616),
	.w7(32'h3b8f1144),
	.w8(32'h3b140368),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170759),
	.w1(32'hbb0af4a7),
	.w2(32'h38efc6cf),
	.w3(32'hbbbe8d83),
	.w4(32'hbb55b9c4),
	.w5(32'hbba95e0e),
	.w6(32'hbaf2baf6),
	.w7(32'h3b30cd08),
	.w8(32'hbab1fba0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c03d),
	.w1(32'hbb263191),
	.w2(32'hbb111e09),
	.w3(32'hb9bfb0b0),
	.w4(32'hbc204901),
	.w5(32'h3aaf0985),
	.w6(32'hb9897181),
	.w7(32'hbbcbd25e),
	.w8(32'hbb9fc10a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4218bc),
	.w1(32'hbb67fa56),
	.w2(32'hbc5cf15a),
	.w3(32'hbb326809),
	.w4(32'hbc1ba3f7),
	.w5(32'hbc8740ee),
	.w6(32'h3c1899c8),
	.w7(32'hb9dba916),
	.w8(32'hba9e6572),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc514210),
	.w1(32'hb989813c),
	.w2(32'h3be76b5d),
	.w3(32'hbc57c726),
	.w4(32'hbbbdfc65),
	.w5(32'h3b69e7f3),
	.w6(32'hbc4dddd2),
	.w7(32'hbb109691),
	.w8(32'h3b9d7b74),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74fc4c),
	.w1(32'h3a800ef4),
	.w2(32'hbb793aea),
	.w3(32'h3a61c099),
	.w4(32'h3c06a767),
	.w5(32'hbcc3b718),
	.w6(32'h39a67517),
	.w7(32'h3c6f166f),
	.w8(32'hbba16ed6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee6f40),
	.w1(32'h3a69957b),
	.w2(32'hb9d7e4f6),
	.w3(32'h3c26468a),
	.w4(32'hbba46154),
	.w5(32'h3c8719ea),
	.w6(32'hb8eb343e),
	.w7(32'hbbde9c92),
	.w8(32'h3bd7bb15),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d3db1),
	.w1(32'h3a9cf6e9),
	.w2(32'hbaeab971),
	.w3(32'hbc09a36e),
	.w4(32'hba0b0590),
	.w5(32'hbc594511),
	.w6(32'hb97d69c4),
	.w7(32'h3aab2a76),
	.w8(32'hbb357db6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a196ee7),
	.w1(32'hbabb8846),
	.w2(32'hbbdff7e9),
	.w3(32'h3c4087dc),
	.w4(32'h3b5e2501),
	.w5(32'hbc9e4a3f),
	.w6(32'hbb3e4e4d),
	.w7(32'h3ae42a8a),
	.w8(32'hbbd964c8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8151d9),
	.w1(32'h3b2582ea),
	.w2(32'h3bc77aa5),
	.w3(32'h3bcd7835),
	.w4(32'h3a14a76f),
	.w5(32'hba22f462),
	.w6(32'h3ba76ead),
	.w7(32'hbb369705),
	.w8(32'hbae88d6f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba693712),
	.w1(32'h3b4e80e2),
	.w2(32'h3b98743e),
	.w3(32'hbc088a46),
	.w4(32'h3b70ebd5),
	.w5(32'h3cfa4511),
	.w6(32'hbaff0ebb),
	.w7(32'hbc3e4ebe),
	.w8(32'hbb8f0493),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392762bb),
	.w1(32'h3bd82f8b),
	.w2(32'hbbb2b0c1),
	.w3(32'hbbad2607),
	.w4(32'h3acfba2f),
	.w5(32'h3d49d5ff),
	.w6(32'hbb170260),
	.w7(32'h3c47d432),
	.w8(32'h3c2bbb05),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3876d090),
	.w1(32'hbb914196),
	.w2(32'hb7fcc5fe),
	.w3(32'hbc28cfd8),
	.w4(32'hbc0329b1),
	.w5(32'h3d325142),
	.w6(32'h3a4ff184),
	.w7(32'hbb27028a),
	.w8(32'h3b84c146),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c1694),
	.w1(32'h3b692a19),
	.w2(32'hba8a81c1),
	.w3(32'hbc351641),
	.w4(32'h3b922795),
	.w5(32'hbc087d1a),
	.w6(32'hbc0e7c9b),
	.w7(32'hbb3f35ae),
	.w8(32'hbb347b04),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38509d0a),
	.w1(32'h3a3749a5),
	.w2(32'h3aca4e14),
	.w3(32'h3b598214),
	.w4(32'h3a471c1f),
	.w5(32'hbb402805),
	.w6(32'h3ae6ff7a),
	.w7(32'h3acc480d),
	.w8(32'hbb3e83a1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb17e4),
	.w1(32'h3c3559ab),
	.w2(32'hbb8af8ca),
	.w3(32'hbb18ff67),
	.w4(32'h3b8c4ebb),
	.w5(32'hbac8bb56),
	.w6(32'hbb680a64),
	.w7(32'h3bd21dfd),
	.w8(32'hbb71d0b0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71f98f),
	.w1(32'hbba2225f),
	.w2(32'hbc5df6c3),
	.w3(32'h3b95c432),
	.w4(32'hbb9ca5c8),
	.w5(32'h39bd713e),
	.w6(32'h3b9a430f),
	.w7(32'hbb88ce12),
	.w8(32'hbafcc1b1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ef46e),
	.w1(32'hbb1fed7e),
	.w2(32'hbc0da790),
	.w3(32'hbc112472),
	.w4(32'h3c0ec3fd),
	.w5(32'h3b56dcd2),
	.w6(32'hbc20183c),
	.w7(32'h3aa75037),
	.w8(32'hbc1f5f12),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd58c4),
	.w1(32'hbb9592ff),
	.w2(32'hbb860b8e),
	.w3(32'hbbd12938),
	.w4(32'h3913ea75),
	.w5(32'hbc1f543d),
	.w6(32'hbb7ee2f6),
	.w7(32'h3a286f07),
	.w8(32'hbb3cb45b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d44f),
	.w1(32'h3c6cc448),
	.w2(32'hbc26b276),
	.w3(32'h3af405ea),
	.w4(32'h3c3bdd55),
	.w5(32'h3c83ad28),
	.w6(32'hbb05358e),
	.w7(32'h3c9831d8),
	.w8(32'hb986f890),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9ffd5),
	.w1(32'h3b551384),
	.w2(32'hb63cc17c),
	.w3(32'hbb7d4a49),
	.w4(32'hbb592486),
	.w5(32'hbc412aa5),
	.w6(32'h3b3c6a3e),
	.w7(32'hbb52011c),
	.w8(32'hbc42617a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ead4),
	.w1(32'h3c3fbb7c),
	.w2(32'hb9d9a340),
	.w3(32'h3bf64dda),
	.w4(32'h3bcf5ba8),
	.w5(32'h3c3c70ac),
	.w6(32'h3adc9916),
	.w7(32'h3bb56e41),
	.w8(32'h3ba6067e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5a1f8),
	.w1(32'hbb22a321),
	.w2(32'hb97c7b37),
	.w3(32'hbaea62bf),
	.w4(32'h3c0fe4cc),
	.w5(32'hbcd24727),
	.w6(32'h3a8ac7a2),
	.w7(32'h3a12eacc),
	.w8(32'hbc0e6a0e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7722ba),
	.w1(32'hbc21251e),
	.w2(32'hbb600478),
	.w3(32'h3c2f461f),
	.w4(32'hbc1dd450),
	.w5(32'hbc24b237),
	.w6(32'h3abe9496),
	.w7(32'hbc0e121a),
	.w8(32'hbb8b9590),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac768a2),
	.w1(32'h39c1321c),
	.w2(32'hb99544bb),
	.w3(32'hbbadbac8),
	.w4(32'hbc45b60a),
	.w5(32'hba15e057),
	.w6(32'hba95c032),
	.w7(32'hbb36140a),
	.w8(32'hbbeb647f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d610),
	.w1(32'hbbf82af6),
	.w2(32'hbb2821b2),
	.w3(32'h3c300c55),
	.w4(32'hbc206583),
	.w5(32'hbc0b9289),
	.w6(32'h3c0ba5ed),
	.w7(32'hbbc1b6ef),
	.w8(32'hbb813ecd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7afce),
	.w1(32'hbaf4b9f4),
	.w2(32'h3b9f17ff),
	.w3(32'hba8f6856),
	.w4(32'hbc299484),
	.w5(32'h3c293ec2),
	.w6(32'hbb1389ff),
	.w7(32'h3bd32790),
	.w8(32'h3c2dde46),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8978d3),
	.w1(32'hbc47105a),
	.w2(32'hbc703bfc),
	.w3(32'hbc035e9f),
	.w4(32'hbc2d618b),
	.w5(32'hbc065b3c),
	.w6(32'h3b2a84f4),
	.w7(32'hbbdae11c),
	.w8(32'h3c133016),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc623099),
	.w1(32'hbc202a8b),
	.w2(32'hbbb1bed0),
	.w3(32'hbba5af6f),
	.w4(32'hbbbf1473),
	.w5(32'h3b99ff7e),
	.w6(32'h39c14e6f),
	.w7(32'hbbfed3ce),
	.w8(32'hbbe8b55d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94999b),
	.w1(32'hba72342a),
	.w2(32'h3b4c65f6),
	.w3(32'hbb819bb0),
	.w4(32'h3bc96454),
	.w5(32'h3be2ba05),
	.w6(32'hbbb1b231),
	.w7(32'h3be42dec),
	.w8(32'h3b9ab2a6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5a236),
	.w1(32'hbae5b304),
	.w2(32'h395217ee),
	.w3(32'hbbccd2ec),
	.w4(32'h3b52a4b2),
	.w5(32'h3bbbb8cd),
	.w6(32'hbbe966d5),
	.w7(32'hb9dc8e6b),
	.w8(32'hb99801ff),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3db53c),
	.w1(32'hbc4d934d),
	.w2(32'hba84fbf4),
	.w3(32'h3a3dae94),
	.w4(32'h3b80c7d8),
	.w5(32'h3b92319c),
	.w6(32'h3af93ff1),
	.w7(32'h3b091f1e),
	.w8(32'hbbdd6c8e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c2691),
	.w1(32'hbbbcb519),
	.w2(32'hbb8df932),
	.w3(32'hbbfda25e),
	.w4(32'h3a9cb88e),
	.w5(32'h3c3f8602),
	.w6(32'hbb4e0343),
	.w7(32'hba73b80e),
	.w8(32'hbb928872),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6caf87),
	.w1(32'h3b47643c),
	.w2(32'h3a518d0b),
	.w3(32'h3aeeb861),
	.w4(32'h3b53a4a5),
	.w5(32'hb9d2c0fa),
	.w6(32'hbb116ca9),
	.w7(32'hba89a5e4),
	.w8(32'h3bb5c8d0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a71ed),
	.w1(32'hbbdb44c6),
	.w2(32'hbc3bb58d),
	.w3(32'h3b4e6543),
	.w4(32'hbbedb87c),
	.w5(32'h3c16173d),
	.w6(32'h3be39c96),
	.w7(32'h3b613c78),
	.w8(32'h3904a45c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2376d),
	.w1(32'hbb1f030f),
	.w2(32'hba2c934a),
	.w3(32'h3b0c5779),
	.w4(32'hbb825d31),
	.w5(32'h3a987372),
	.w6(32'hbb3b1d31),
	.w7(32'h3a4ffd5e),
	.w8(32'h3911b9ac),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0378dd),
	.w1(32'hbb4d2b83),
	.w2(32'hbbd2da26),
	.w3(32'h3b7469f7),
	.w4(32'hba21acf8),
	.w5(32'hbb9ea245),
	.w6(32'hbad6b8b7),
	.w7(32'hbad8a377),
	.w8(32'hbacaf74a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab982c2),
	.w1(32'h3b203f7a),
	.w2(32'h3b87994c),
	.w3(32'hbbd39b1d),
	.w4(32'h3a05f168),
	.w5(32'hbbccdc97),
	.w6(32'hbba771da),
	.w7(32'h3bfcddcc),
	.w8(32'h3c82a1c1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b357d7b),
	.w1(32'hbb2d1539),
	.w2(32'hbb8a9857),
	.w3(32'h3c26aeea),
	.w4(32'hbbf8956c),
	.w5(32'hbc02d803),
	.w6(32'h3c3f1532),
	.w7(32'hbb607c26),
	.w8(32'hbb0b5f3d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8103e6),
	.w1(32'h38f9fd54),
	.w2(32'h3ba347ba),
	.w3(32'h39d9d8de),
	.w4(32'hb9eb1dd2),
	.w5(32'hbb7b5a01),
	.w6(32'hbb202d32),
	.w7(32'hbaa7c080),
	.w8(32'h3baa57c2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc362f),
	.w1(32'h3b9ad408),
	.w2(32'hbb4459f2),
	.w3(32'h3a4362e0),
	.w4(32'hbb74e1d7),
	.w5(32'hbb27a2f3),
	.w6(32'h3b86275a),
	.w7(32'hbbcd3dbf),
	.w8(32'hbb033a6d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc410e9c),
	.w1(32'hbc0008e5),
	.w2(32'hbbc0cc76),
	.w3(32'hbb8b4b57),
	.w4(32'hbb8339e6),
	.w5(32'hbbf4ebb9),
	.w6(32'hbb8985ef),
	.w7(32'hbbc50f9c),
	.w8(32'hbb548eca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3b36),
	.w1(32'hbb561fbd),
	.w2(32'hbc63d43e),
	.w3(32'hbb2d3cb7),
	.w4(32'h3c0b0cb8),
	.w5(32'hbc08c0ef),
	.w6(32'hbb3e7867),
	.w7(32'h3bcd8479),
	.w8(32'hb955600f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2adcc5),
	.w1(32'hbb91fc97),
	.w2(32'hbc001ab3),
	.w3(32'h3b0766e9),
	.w4(32'hbb5b0642),
	.w5(32'hbbc127c2),
	.w6(32'hbbd78abb),
	.w7(32'hbba69dd6),
	.w8(32'hbc53e8e8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc549ee2),
	.w1(32'h3c0f5f53),
	.w2(32'h3c3ad361),
	.w3(32'hbc11b6e1),
	.w4(32'h39f9a19a),
	.w5(32'hbb37fe7a),
	.w6(32'hbc3b264f),
	.w7(32'hb9a3d393),
	.w8(32'h3a658f1b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcec789),
	.w1(32'hbb00446a),
	.w2(32'hbb90f167),
	.w3(32'hbc2d6230),
	.w4(32'hbbca7077),
	.w5(32'hbb636cf8),
	.w6(32'hbbc92a70),
	.w7(32'hbbb4c8eb),
	.w8(32'h3a89d76a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e6d6),
	.w1(32'h3b9c14ff),
	.w2(32'hbb45cc4e),
	.w3(32'hbba7f05d),
	.w4(32'h3bfe4176),
	.w5(32'h3c8b95fe),
	.w6(32'hbbd639bf),
	.w7(32'hbb8a6a92),
	.w8(32'h3bb0ce66),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb859c64),
	.w1(32'hbb7ef8cb),
	.w2(32'hba8f576c),
	.w3(32'h3c245240),
	.w4(32'hbbf36382),
	.w5(32'hbac491a8),
	.w6(32'h3c2a0046),
	.w7(32'hbb65b6f6),
	.w8(32'h3b96f759),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d6d0a),
	.w1(32'hba558fd5),
	.w2(32'h3b84031f),
	.w3(32'hbbb7c0ed),
	.w4(32'h3b775a9f),
	.w5(32'hbbf639ff),
	.w6(32'h391b54be),
	.w7(32'h3b9771d5),
	.w8(32'h3bc8b62f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac41d),
	.w1(32'hbbad2e15),
	.w2(32'h3c039a6b),
	.w3(32'hbb1e86b4),
	.w4(32'hbb9a308d),
	.w5(32'hbc0ac002),
	.w6(32'h3bb82ffb),
	.w7(32'hbc043bf5),
	.w8(32'hbaff333f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db7996),
	.w1(32'h3b2b5647),
	.w2(32'h3b285018),
	.w3(32'hbaf00229),
	.w4(32'h3b48834b),
	.w5(32'hbaa61ba4),
	.w6(32'hbb92c2b1),
	.w7(32'h3a29c293),
	.w8(32'h3b1cbc55),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885cf5c),
	.w1(32'hbc1aed8a),
	.w2(32'hbc1a2be8),
	.w3(32'h3b0b5e8f),
	.w4(32'hbaa2b034),
	.w5(32'hbb5ba415),
	.w6(32'h3b094dee),
	.w7(32'hb9b92629),
	.w8(32'h3b95ec64),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc341f67),
	.w1(32'h3a7e2a4e),
	.w2(32'h3b1a73af),
	.w3(32'hbc5a3f4a),
	.w4(32'hba31081f),
	.w5(32'h3c223cfb),
	.w6(32'hbbaae584),
	.w7(32'hba91e833),
	.w8(32'h3b5bd669),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b82a9),
	.w1(32'h3a9aa2d3),
	.w2(32'h39a0f6f7),
	.w3(32'h3b81ab37),
	.w4(32'hbad29cf8),
	.w5(32'hbb893271),
	.w6(32'h3b8ae00a),
	.w7(32'hbb367cd0),
	.w8(32'h3ab79c5c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec3ef6),
	.w1(32'h3baaed7e),
	.w2(32'h3c1140f6),
	.w3(32'hbb8175b8),
	.w4(32'hbadf06c1),
	.w5(32'h3bee416d),
	.w6(32'hbbc0af5a),
	.w7(32'h39835997),
	.w8(32'h3b5416b8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7053bd),
	.w1(32'h3c10cf04),
	.w2(32'h3a185517),
	.w3(32'h3b2973ca),
	.w4(32'h3b8a7e35),
	.w5(32'h3cc9c469),
	.w6(32'h3beb02ee),
	.w7(32'hbb2d6424),
	.w8(32'hbb8b9d88),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befe1a9),
	.w1(32'h3c489cd2),
	.w2(32'hba1f5601),
	.w3(32'h3b99baea),
	.w4(32'h3c8af54f),
	.w5(32'h3d3b286c),
	.w6(32'hbc062c07),
	.w7(32'h3b7138de),
	.w8(32'hbc1e2d0e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b883d99),
	.w1(32'hbb3aab1f),
	.w2(32'hbbad8c0c),
	.w3(32'h3c9840b5),
	.w4(32'hbb7a95e6),
	.w5(32'hbb722741),
	.w6(32'h3af8a5ef),
	.w7(32'hbbb7b6dd),
	.w8(32'hbbae25de),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba015e),
	.w1(32'hbaf192cd),
	.w2(32'hbbfb42fb),
	.w3(32'hbbe46eb4),
	.w4(32'hbbff7658),
	.w5(32'hbb9df11a),
	.w6(32'hbbb35ef4),
	.w7(32'hbc07c111),
	.w8(32'hbba869ce),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a11fc),
	.w1(32'h3ae49890),
	.w2(32'h3ae0bbe8),
	.w3(32'hbb1027c2),
	.w4(32'h3b64ad42),
	.w5(32'h3ca8464f),
	.w6(32'hbc0efcaa),
	.w7(32'hbb8dd1a8),
	.w8(32'h3b2d96cd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee7d3),
	.w1(32'h3af330e5),
	.w2(32'h3b38a8f0),
	.w3(32'h3ba2cfc1),
	.w4(32'hbbc4ddf0),
	.w5(32'hbb1777f0),
	.w6(32'h3acfe03a),
	.w7(32'hbb7e5c83),
	.w8(32'h3a59c391),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b168),
	.w1(32'hbb3fd6c1),
	.w2(32'h3b43479c),
	.w3(32'h39292a04),
	.w4(32'hbbeb1c4e),
	.w5(32'hbbd62042),
	.w6(32'h3a4b9724),
	.w7(32'hbc0a1d66),
	.w8(32'h3b478b0c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd671a9),
	.w1(32'hb9af73d9),
	.w2(32'hbbac3cb7),
	.w3(32'hbb41c2ce),
	.w4(32'hb97e01bc),
	.w5(32'hb9596fd6),
	.w6(32'hba8f2ea3),
	.w7(32'hba85f6de),
	.w8(32'hbae1b038),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ffe7b),
	.w1(32'h3bf30983),
	.w2(32'h3ad8c007),
	.w3(32'hbab95a1f),
	.w4(32'h3bdeea74),
	.w5(32'hbb212488),
	.w6(32'hbab7a9df),
	.w7(32'hbb22376d),
	.w8(32'h3b71152d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9affc47),
	.w1(32'hbb8924e1),
	.w2(32'h3ac132ad),
	.w3(32'h3bcfc39a),
	.w4(32'h3af8ba6d),
	.w5(32'h3c361818),
	.w6(32'h3bcd2664),
	.w7(32'h3bbb8425),
	.w8(32'h3c482c9f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1e1b),
	.w1(32'hb98a573f),
	.w2(32'h3b8319aa),
	.w3(32'hbba46598),
	.w4(32'h3ba88793),
	.w5(32'h3bc9fe82),
	.w6(32'h3b801bb8),
	.w7(32'h398c8bd3),
	.w8(32'hbb032c89),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38402cca),
	.w1(32'hba4979b1),
	.w2(32'h3b819e9d),
	.w3(32'h3ba103bd),
	.w4(32'hbbeb97de),
	.w5(32'hbbb100c0),
	.w6(32'hbb929ba2),
	.w7(32'hbba93931),
	.w8(32'hb9850368),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886685),
	.w1(32'h3a2a72e4),
	.w2(32'hbbbc1391),
	.w3(32'hbbeb9ed7),
	.w4(32'hb8cf1f91),
	.w5(32'hb98456fe),
	.w6(32'hbbbe6960),
	.w7(32'h39f8403c),
	.w8(32'h3c227260),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc74bd),
	.w1(32'h3c333748),
	.w2(32'h3b95dbf0),
	.w3(32'hbba6eb25),
	.w4(32'hbb10b13f),
	.w5(32'h3b4fa51e),
	.w6(32'h3ade4352),
	.w7(32'hbae86f27),
	.w8(32'h3aad8ae9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94857d),
	.w1(32'h3bbef284),
	.w2(32'h3b00accb),
	.w3(32'h3b312d24),
	.w4(32'h3b888586),
	.w5(32'h3b05ac57),
	.w6(32'h3ac539c4),
	.w7(32'hbac6f7dc),
	.w8(32'hbbaea1f1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970bc5),
	.w1(32'h3b707fe0),
	.w2(32'h3bcc1074),
	.w3(32'h3ab351f8),
	.w4(32'hbb7a5d3c),
	.w5(32'hbbd5ece4),
	.w6(32'hbb95e873),
	.w7(32'hba3198a3),
	.w8(32'hbbb6dedd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b014821),
	.w1(32'hbad8376b),
	.w2(32'h3b720747),
	.w3(32'h3aa6d160),
	.w4(32'h3be1e569),
	.w5(32'h3ad7a483),
	.w6(32'h38df5cb1),
	.w7(32'h3c2dad16),
	.w8(32'hbb0cc783),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b828357),
	.w1(32'hbb6a975a),
	.w2(32'hbb8cd219),
	.w3(32'h3b6736a8),
	.w4(32'hbb0cbf52),
	.w5(32'hb7036dab),
	.w6(32'h3b957ab9),
	.w7(32'h3a5ceb29),
	.w8(32'h3b9bbd78),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c8c6b),
	.w1(32'h3bebf636),
	.w2(32'h3c4b1492),
	.w3(32'hb8ad2a75),
	.w4(32'h3b34f5c7),
	.w5(32'h3906a54b),
	.w6(32'h3bc83344),
	.w7(32'h3bdaee99),
	.w8(32'hbb07481f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ede3e),
	.w1(32'hbb034d9d),
	.w2(32'hbaa24e67),
	.w3(32'h3c3ce6ec),
	.w4(32'h3b9daf5e),
	.w5(32'h3b4d07bc),
	.w6(32'h3b834b4c),
	.w7(32'h3bbaaab5),
	.w8(32'h3b925bf2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed153),
	.w1(32'h3a51f0ae),
	.w2(32'h3b897f89),
	.w3(32'h3c052a17),
	.w4(32'hbb7dcc33),
	.w5(32'h3ba01db7),
	.w6(32'h3acc905e),
	.w7(32'hbaa7b021),
	.w8(32'h39865eea),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa379b),
	.w1(32'hbaabce86),
	.w2(32'hbb8ffc93),
	.w3(32'hbaf09a82),
	.w4(32'hbab1864c),
	.w5(32'hb99f3a0a),
	.w6(32'hba8f458e),
	.w7(32'hbb1d8fae),
	.w8(32'hbb8f155c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f997e2),
	.w1(32'h39e8aedb),
	.w2(32'hb9bd7a59),
	.w3(32'hbb3d672c),
	.w4(32'hbbf2ab48),
	.w5(32'hbba4e9bf),
	.w6(32'hbaf1e2d9),
	.w7(32'hbbe92e9a),
	.w8(32'h3aa50206),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd66d0),
	.w1(32'hbb9d97a3),
	.w2(32'hbbb2d414),
	.w3(32'hbba2af1b),
	.w4(32'h3c681778),
	.w5(32'h3cf3d319),
	.w6(32'hbaaa07f2),
	.w7(32'h3ccb46c6),
	.w8(32'h3cd8c533),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfd6f0),
	.w1(32'hbb60c9ac),
	.w2(32'hbbb0b86a),
	.w3(32'h3c95f801),
	.w4(32'hbb4650c9),
	.w5(32'hba1afb1f),
	.w6(32'hbb577f3e),
	.w7(32'hbbbebe83),
	.w8(32'h3b105e50),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcad51b),
	.w1(32'hbb391fa5),
	.w2(32'hbc03b450),
	.w3(32'hbb0a628f),
	.w4(32'h3ba597e1),
	.w5(32'h3a8cb5c9),
	.w6(32'h3a52166c),
	.w7(32'h3bbbdc48),
	.w8(32'h3bcbab21),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2eee66),
	.w1(32'hbb2ed408),
	.w2(32'h3b8d85c0),
	.w3(32'h3c1dae82),
	.w4(32'h3932a77a),
	.w5(32'h3c560135),
	.w6(32'hba1668a4),
	.w7(32'hbbc68807),
	.w8(32'hba967ce9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95fb71),
	.w1(32'h3afda615),
	.w2(32'h3be74349),
	.w3(32'h3b8cba78),
	.w4(32'h3be751df),
	.w5(32'h3a30b416),
	.w6(32'hbb34d304),
	.w7(32'hbb27dff4),
	.w8(32'hbb17a4fb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c6644),
	.w1(32'h3b9d173a),
	.w2(32'h3abe6d48),
	.w3(32'h3a6ef41a),
	.w4(32'hb9f2a027),
	.w5(32'hbb9476cd),
	.w6(32'hbad59344),
	.w7(32'h3c354a7e),
	.w8(32'h3c12e4f1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74bec3),
	.w1(32'h3b0912e3),
	.w2(32'h3ad8db04),
	.w3(32'h3bb73004),
	.w4(32'h3a9c8d02),
	.w5(32'h3b13227d),
	.w6(32'h3bcb419e),
	.w7(32'hbb0dd2a6),
	.w8(32'hbae0f0f9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule