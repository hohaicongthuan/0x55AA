module layer_10_featuremap_57(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7c10e),
	.w1(32'hbca14821),
	.w2(32'hbbff4c9b),
	.w3(32'h3d355465),
	.w4(32'h3b679758),
	.w5(32'h3ce219d8),
	.w6(32'h3c9a307a),
	.w7(32'h3ca2c56d),
	.w8(32'hbb185069),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7ce10),
	.w1(32'hbc5c5228),
	.w2(32'hbb57a729),
	.w3(32'h3c89039e),
	.w4(32'hbb9f638e),
	.w5(32'h3c6861c4),
	.w6(32'h3c9a7efb),
	.w7(32'h3c88a682),
	.w8(32'h3c6e70c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60252c),
	.w1(32'h3b157d50),
	.w2(32'h3bce7efa),
	.w3(32'h3c7d65ca),
	.w4(32'h3c5900d1),
	.w5(32'h3b1fdba4),
	.w6(32'h3d086748),
	.w7(32'h3cd47dfc),
	.w8(32'hba1378e1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc30bc1),
	.w1(32'hbb69281b),
	.w2(32'h3a871ac2),
	.w3(32'h3c8a666c),
	.w4(32'h3c19151d),
	.w5(32'hbceca6ac),
	.w6(32'h3b93f5fc),
	.w7(32'h3a5aa712),
	.w8(32'h3a6c6e22),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b5b3),
	.w1(32'h3bb27e0f),
	.w2(32'h3c580dbd),
	.w3(32'hbca9b406),
	.w4(32'hbc332dd7),
	.w5(32'hbb8cb60a),
	.w6(32'hbc2e8990),
	.w7(32'hbc737a00),
	.w8(32'hbc16ac48),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ea880),
	.w1(32'hbbabafbc),
	.w2(32'h3bae03d5),
	.w3(32'h3bbb6ab3),
	.w4(32'h3b5ae221),
	.w5(32'hb8170bd3),
	.w6(32'hbc3c4f1c),
	.w7(32'h3b917c63),
	.w8(32'h3a4eb6f5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a077c),
	.w1(32'h3b9c52be),
	.w2(32'h39a0462c),
	.w3(32'hbb8985f0),
	.w4(32'hbb0a4575),
	.w5(32'hbc4322d6),
	.w6(32'hbb5dda2b),
	.w7(32'h3a725aa2),
	.w8(32'hbb0eb794),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c072c71),
	.w1(32'h3a2cf488),
	.w2(32'hbc1165af),
	.w3(32'hbc89708f),
	.w4(32'hbaf589a4),
	.w5(32'h3b9e91c6),
	.w6(32'hbc5371a5),
	.w7(32'hbc840400),
	.w8(32'hbb44fa22),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a616c),
	.w1(32'hbc5c560f),
	.w2(32'hba9c5de1),
	.w3(32'h3b2077a9),
	.w4(32'h3ae18987),
	.w5(32'h3a86eadb),
	.w6(32'h3b04ccab),
	.w7(32'h3b86edc3),
	.w8(32'h3ab5bedf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c363fc8),
	.w1(32'h3c580867),
	.w2(32'h3a93ad81),
	.w3(32'hbb884a00),
	.w4(32'h3b67b115),
	.w5(32'h3b2a54e6),
	.w6(32'hbba09e7b),
	.w7(32'hb9b22c75),
	.w8(32'hbb48cb8a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf14ddb),
	.w1(32'h384d06c9),
	.w2(32'h3be2e747),
	.w3(32'h3a6a0b44),
	.w4(32'h3ab8f098),
	.w5(32'hbb5baaf4),
	.w6(32'h3aed58e2),
	.w7(32'h3adc7973),
	.w8(32'h39110392),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c1d50a),
	.w1(32'h3a4d516c),
	.w2(32'h3bcbb79e),
	.w3(32'hbaabc16d),
	.w4(32'hbacadfe7),
	.w5(32'h3bb5e50a),
	.w6(32'h3c02628b),
	.w7(32'h3bef609b),
	.w8(32'hbb0ac794),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb3e03),
	.w1(32'h3c3bbe7e),
	.w2(32'h3c3a4c7c),
	.w3(32'h3c2d034f),
	.w4(32'h3c3d7c41),
	.w5(32'h3b487e89),
	.w6(32'hbb00c23c),
	.w7(32'h3b3e078f),
	.w8(32'h3c25708a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f22f8),
	.w1(32'h3bb2ec5c),
	.w2(32'hbb8da5d8),
	.w3(32'h38f8e0b1),
	.w4(32'hba8fea1b),
	.w5(32'hbb670a20),
	.w6(32'h3ad643df),
	.w7(32'h3b86a6a5),
	.w8(32'hbb6fda17),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccf4d8),
	.w1(32'hbb0b3714),
	.w2(32'hbb88764c),
	.w3(32'h3c96c29f),
	.w4(32'h3cdad4ad),
	.w5(32'hb9306210),
	.w6(32'hbc8ad277),
	.w7(32'hbb29c74f),
	.w8(32'h3c290b64),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ef666),
	.w1(32'h3ba302b9),
	.w2(32'h3ae78351),
	.w3(32'hbc825a30),
	.w4(32'hbb8c095e),
	.w5(32'h3b442e92),
	.w6(32'h3b2244bb),
	.w7(32'hbaad3504),
	.w8(32'hbaaba8e3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3adb1d),
	.w1(32'hba1ff1a7),
	.w2(32'hbb9f9a54),
	.w3(32'h3a2144b8),
	.w4(32'h3b08a680),
	.w5(32'hbaf2f100),
	.w6(32'h3b293772),
	.w7(32'h3b4ac3d5),
	.w8(32'h3ae39255),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b4143),
	.w1(32'hbc1de914),
	.w2(32'h3b2f2d72),
	.w3(32'hbc1aec90),
	.w4(32'hbbca1b92),
	.w5(32'h3c04ef10),
	.w6(32'hba9f3297),
	.w7(32'h3aeadff0),
	.w8(32'hb99e9738),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba674),
	.w1(32'h3b1a6bf4),
	.w2(32'h3c0c32a8),
	.w3(32'hbb7a7582),
	.w4(32'hbb97023b),
	.w5(32'h3c81fc48),
	.w6(32'hb9cd9d66),
	.w7(32'hbadc4066),
	.w8(32'hbb00f96b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8e94),
	.w1(32'hbbdd386b),
	.w2(32'h3afad954),
	.w3(32'h3d0440f1),
	.w4(32'h3d0083ea),
	.w5(32'hbb61846f),
	.w6(32'h3bab1168),
	.w7(32'h3c6faf48),
	.w8(32'hbbb4eaf1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7288df),
	.w1(32'hba9483bd),
	.w2(32'h3bc5e91a),
	.w3(32'hba14e054),
	.w4(32'h3b85595f),
	.w5(32'h3bc5be8e),
	.w6(32'hbb7b969f),
	.w7(32'h3ba99e2b),
	.w8(32'h3ba5bc06),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c2c8),
	.w1(32'h3aeaa3c3),
	.w2(32'h3b60b13d),
	.w3(32'h3c98a952),
	.w4(32'h3bd25a1e),
	.w5(32'hbbdad68b),
	.w6(32'h3a965d43),
	.w7(32'hbbaff276),
	.w8(32'hbac138fe),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5839e3),
	.w1(32'hbb5eb637),
	.w2(32'h3acb775e),
	.w3(32'h3c26ffff),
	.w4(32'hba1dffb0),
	.w5(32'hbb9c1284),
	.w6(32'hbcaebd68),
	.w7(32'hbc929cc9),
	.w8(32'hbc7de814),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b475341),
	.w1(32'h3b8afa7e),
	.w2(32'h3bb45deb),
	.w3(32'h3bae96c5),
	.w4(32'h3bb739af),
	.w5(32'h3c32e220),
	.w6(32'hbbc75936),
	.w7(32'hbb21db83),
	.w8(32'h3a502506),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2f0bc),
	.w1(32'h3ace78c8),
	.w2(32'hb99a8be0),
	.w3(32'hba64001a),
	.w4(32'h3ba13c9b),
	.w5(32'h3a67df91),
	.w6(32'hbb616c19),
	.w7(32'h3b6aa914),
	.w8(32'hbcb59a59),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9614d),
	.w1(32'hbc3622e5),
	.w2(32'h3c2838ff),
	.w3(32'hba91046f),
	.w4(32'hbba3290d),
	.w5(32'h3bbd6863),
	.w6(32'hbca397f9),
	.w7(32'hbc25ba89),
	.w8(32'h3b2d5423),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c43c),
	.w1(32'h3aa75c77),
	.w2(32'h3a27f644),
	.w3(32'h3cbda68f),
	.w4(32'h3c34b0b0),
	.w5(32'hb9860200),
	.w6(32'hbc1cf689),
	.w7(32'h3bf0e916),
	.w8(32'h39d0f7f6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a374e0d),
	.w1(32'h3b05f7af),
	.w2(32'hbbd24b51),
	.w3(32'hba70476e),
	.w4(32'h3b254133),
	.w5(32'h3a3ef5ac),
	.w6(32'h3a61b8a6),
	.w7(32'h3aa89da0),
	.w8(32'h3be1f635),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb551a3),
	.w1(32'hbbd10a12),
	.w2(32'hbb69928a),
	.w3(32'h3b960a94),
	.w4(32'h3b12a6a5),
	.w5(32'hbb9c39af),
	.w6(32'h3c6afb49),
	.w7(32'h3c2a970f),
	.w8(32'hba94408b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23cab6),
	.w1(32'hbaab3f65),
	.w2(32'hbbe3ed3a),
	.w3(32'hbc402046),
	.w4(32'hbb0a201a),
	.w5(32'h3a906eb2),
	.w6(32'h3c81b837),
	.w7(32'h3c616089),
	.w8(32'hbab116f6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab69e0),
	.w1(32'hbbd66b59),
	.w2(32'h3c65ddb4),
	.w3(32'h3b2c0d36),
	.w4(32'hb9c33bb1),
	.w5(32'h3ae1b194),
	.w6(32'h37c6ed99),
	.w7(32'hbac64952),
	.w8(32'h3c0ad4ba),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bf26c),
	.w1(32'h3c4d3ead),
	.w2(32'h3b51742c),
	.w3(32'hbafcd6e2),
	.w4(32'hbbb8b21a),
	.w5(32'hbc4212dd),
	.w6(32'h3c3c9edb),
	.w7(32'h3ba9404c),
	.w8(32'h3c8e555d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0099f5),
	.w1(32'h3b0e4c44),
	.w2(32'hbb1fbd4c),
	.w3(32'hbbd45c5a),
	.w4(32'h39d13e10),
	.w5(32'hb8c3360e),
	.w6(32'h3c638553),
	.w7(32'hbb4989c1),
	.w8(32'h3ad9d292),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f61c),
	.w1(32'hbbb8fadf),
	.w2(32'h3b94ccb3),
	.w3(32'hba91d026),
	.w4(32'hbba3a5dd),
	.w5(32'h3bfed02a),
	.w6(32'h39cb69ee),
	.w7(32'h3a4de229),
	.w8(32'hbb9e1ac9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5078b),
	.w1(32'h3c899270),
	.w2(32'hbaec826a),
	.w3(32'h3c4d89e4),
	.w4(32'hbbdf2510),
	.w5(32'hbb29b409),
	.w6(32'hbb9d82dd),
	.w7(32'hbaaa470a),
	.w8(32'hbb5ae34d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42dcdc),
	.w1(32'h39969bb9),
	.w2(32'h3c144cc7),
	.w3(32'h3a60d84a),
	.w4(32'h366c2a8e),
	.w5(32'h3b3a3dc9),
	.w6(32'hba1ce103),
	.w7(32'h3ab3ef93),
	.w8(32'h3b3c1d28),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41adce),
	.w1(32'h3b03f037),
	.w2(32'hbbe74877),
	.w3(32'hbc681923),
	.w4(32'hbcca8f0c),
	.w5(32'hb9c8bda0),
	.w6(32'h3c40ddd9),
	.w7(32'h3ca00bdd),
	.w8(32'h3b9f1093),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9a14f),
	.w1(32'hbc287fc0),
	.w2(32'hbc4397af),
	.w3(32'h3a7acdbf),
	.w4(32'hbb80ee98),
	.w5(32'h3c2a53fc),
	.w6(32'h3b916e15),
	.w7(32'h3bd11adf),
	.w8(32'hbc2a9581),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe056b),
	.w1(32'hbb8156e3),
	.w2(32'hba8cf50c),
	.w3(32'h3bdc3214),
	.w4(32'hbb4a7072),
	.w5(32'hbc19fe28),
	.w6(32'hbca193a0),
	.w7(32'hbb309465),
	.w8(32'hbbe8ae00),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2965d2),
	.w1(32'hb939b42a),
	.w2(32'h3b08abb2),
	.w3(32'h3c7acb68),
	.w4(32'h3c98b25b),
	.w5(32'hbb0a4bba),
	.w6(32'hbbc7f660),
	.w7(32'hbbf618aa),
	.w8(32'hbbe5501d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a1df7),
	.w1(32'h3b9c5a5a),
	.w2(32'hbc1b642b),
	.w3(32'h3c190f24),
	.w4(32'h3b833448),
	.w5(32'h3c03af3c),
	.w6(32'h3bfd9c83),
	.w7(32'h3b4b34d0),
	.w8(32'h3c340647),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909049),
	.w1(32'h3ac65767),
	.w2(32'h3ac9213a),
	.w3(32'h3c68d4b2),
	.w4(32'h3c0e7e50),
	.w5(32'hbbe4c672),
	.w6(32'h3b98fead),
	.w7(32'h3c090975),
	.w8(32'h3b3ee739),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35b5fe),
	.w1(32'h3c22dd55),
	.w2(32'hbae299d4),
	.w3(32'hbc822d8c),
	.w4(32'hbc74d07d),
	.w5(32'hbb98493f),
	.w6(32'h3be108f7),
	.w7(32'h3c8b6c4a),
	.w8(32'hbaee77d1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52489),
	.w1(32'h3bab1616),
	.w2(32'hbc001b51),
	.w3(32'hbbf97f59),
	.w4(32'hba8ef4af),
	.w5(32'hbc4c99d4),
	.w6(32'hbb7e9f8b),
	.w7(32'hba99fc97),
	.w8(32'hbace2e79),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86aa6c),
	.w1(32'h3b22492a),
	.w2(32'h3b6b2475),
	.w3(32'hbb8aaba9),
	.w4(32'h39766d96),
	.w5(32'hbba02fb7),
	.w6(32'h3ba79d80),
	.w7(32'hbb304bb8),
	.w8(32'h3b2fdde5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f512),
	.w1(32'hbc18c9d5),
	.w2(32'hba392d9d),
	.w3(32'hbb0cf168),
	.w4(32'h3b762741),
	.w5(32'h3baf6d3c),
	.w6(32'hbb8e3b49),
	.w7(32'hbb74cd0b),
	.w8(32'h3b98c245),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacf3a8),
	.w1(32'h38b459a2),
	.w2(32'hbbebba37),
	.w3(32'hbc127eed),
	.w4(32'hbc09319d),
	.w5(32'h3c16822e),
	.w6(32'h3b85ea4f),
	.w7(32'h3bc9aa34),
	.w8(32'h39882237),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8385c),
	.w1(32'hb992cd2f),
	.w2(32'hb683cc12),
	.w3(32'hbc970a7c),
	.w4(32'hbcda293b),
	.w5(32'hbb8b671c),
	.w6(32'hbba4930a),
	.w7(32'hbac738af),
	.w8(32'hbc028b6b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00951e),
	.w1(32'h39a68950),
	.w2(32'h3975ddf7),
	.w3(32'hbb9f99f9),
	.w4(32'h3a18f6b2),
	.w5(32'hbbcb9ad2),
	.w6(32'hbb52d1d5),
	.w7(32'hbaaa1df1),
	.w8(32'h398cabb4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf652ef),
	.w1(32'h3c07bde8),
	.w2(32'hba8e4ca6),
	.w3(32'h3a21934e),
	.w4(32'h3c27e6be),
	.w5(32'hbb012760),
	.w6(32'hbbbb062e),
	.w7(32'hbb215d55),
	.w8(32'h3b96db8d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6060ca),
	.w1(32'hbb8518ca),
	.w2(32'hbc113afb),
	.w3(32'hbbeafb30),
	.w4(32'h3b317a09),
	.w5(32'hbc887303),
	.w6(32'h3beebcdc),
	.w7(32'h3c688981),
	.w8(32'h3c301496),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca40333),
	.w1(32'hbc38edc3),
	.w2(32'h3a6f3188),
	.w3(32'hbc9b0293),
	.w4(32'hbb0406fa),
	.w5(32'hb903e099),
	.w6(32'h3c41bf8f),
	.w7(32'h3b543b2b),
	.w8(32'h3c57b080),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c8f1),
	.w1(32'hbb8f4cab),
	.w2(32'h39fa54f2),
	.w3(32'hbabc9e77),
	.w4(32'hbbc2cb19),
	.w5(32'h3ba1cd59),
	.w6(32'h3aaa0813),
	.w7(32'h3bd99b1a),
	.w8(32'h3a17f529),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f580f),
	.w1(32'h3987298c),
	.w2(32'hbc607a0c),
	.w3(32'h3b5e4503),
	.w4(32'h3bbcd150),
	.w5(32'h3c97eb90),
	.w6(32'h3c73a1b6),
	.w7(32'h3c292ecd),
	.w8(32'hbbd06254),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aabfd),
	.w1(32'hbc6f7e6d),
	.w2(32'h3be5607b),
	.w3(32'h3cdadbf5),
	.w4(32'h3cca4df5),
	.w5(32'hbbb22d8c),
	.w6(32'hba036a10),
	.w7(32'h3b3d3487),
	.w8(32'h3b8b948e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a5f9),
	.w1(32'h3b61189c),
	.w2(32'h3a98febd),
	.w3(32'h3c692429),
	.w4(32'h3c8ebc87),
	.w5(32'h399f67b6),
	.w6(32'h3bd27ab4),
	.w7(32'h3c10957a),
	.w8(32'h3b97dde4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b88c),
	.w1(32'hbc097d38),
	.w2(32'h3888eefb),
	.w3(32'hbcb265ee),
	.w4(32'hbc8e0b1a),
	.w5(32'h3a9e3e87),
	.w6(32'h3c0e7d45),
	.w7(32'hbbb7276e),
	.w8(32'hbbd15748),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04703f),
	.w1(32'hbb22de37),
	.w2(32'h38ee53fa),
	.w3(32'hbc13f1f7),
	.w4(32'hbbd67b39),
	.w5(32'hb9e6b966),
	.w6(32'hbc6b97a5),
	.w7(32'hb9f91c3e),
	.w8(32'h3b21ef1b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d04de),
	.w1(32'h3bc15942),
	.w2(32'h3ba33384),
	.w3(32'hbac3a1dc),
	.w4(32'h3bf982f8),
	.w5(32'h3ba840fe),
	.w6(32'h3aeaa551),
	.w7(32'h3c2a96b4),
	.w8(32'hbb20e7b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cf3b5),
	.w1(32'h3c4c0483),
	.w2(32'h3afb4496),
	.w3(32'hbac5ee42),
	.w4(32'h3ac98a20),
	.w5(32'h3bfae4d6),
	.w6(32'hbc8fec1a),
	.w7(32'hbc6cf968),
	.w8(32'hba188fb3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fcf98),
	.w1(32'h3b5d59f1),
	.w2(32'hbbbb5d19),
	.w3(32'hbb9f8c8d),
	.w4(32'hbad7126e),
	.w5(32'hbbf02109),
	.w6(32'hbc1582bf),
	.w7(32'hbb9bcdd5),
	.w8(32'h3ac7b1fc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a8968),
	.w1(32'h3bfc3305),
	.w2(32'h3883e7e2),
	.w3(32'hbc9757ab),
	.w4(32'hbbc99567),
	.w5(32'h3aedf17f),
	.w6(32'hbb1e1894),
	.w7(32'hba0cbad6),
	.w8(32'h3966d3e1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41423d),
	.w1(32'h3b83de0e),
	.w2(32'h3b7de951),
	.w3(32'hbbc333cd),
	.w4(32'hbba4d0b1),
	.w5(32'h3bbf7785),
	.w6(32'h3b699a0c),
	.w7(32'h3b897002),
	.w8(32'h3bd1187e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb501),
	.w1(32'hbaabf709),
	.w2(32'h3a802f42),
	.w3(32'hbb16da1b),
	.w4(32'h3a703685),
	.w5(32'hbbc7490a),
	.w6(32'h3bcf613d),
	.w7(32'h3bdcb92c),
	.w8(32'hbb869c17),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5c6b),
	.w1(32'h3be73e72),
	.w2(32'h3b0e0dbc),
	.w3(32'h39c1e8ff),
	.w4(32'hbb657357),
	.w5(32'hba4c0f79),
	.w6(32'hb9fd250c),
	.w7(32'h39da8b05),
	.w8(32'hbb52edfc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b581454),
	.w1(32'h3ac5649d),
	.w2(32'h3b07a345),
	.w3(32'h3b21c826),
	.w4(32'h3b7ec958),
	.w5(32'h3b135a5d),
	.w6(32'hba86ff46),
	.w7(32'hb9c174d1),
	.w8(32'h3be3d36a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d8126),
	.w1(32'h3ba18b5b),
	.w2(32'hbbfbaabd),
	.w3(32'hbb2249f6),
	.w4(32'h3b00581d),
	.w5(32'h3a27d311),
	.w6(32'hba6f7f35),
	.w7(32'h3b253fc3),
	.w8(32'h3bb29272),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb995),
	.w1(32'h3c0208db),
	.w2(32'hbaaec828),
	.w3(32'h3b862677),
	.w4(32'h3ba6caf6),
	.w5(32'hba1f62d1),
	.w6(32'h3ab0fa2c),
	.w7(32'h3b94e84e),
	.w8(32'h3b5f59f0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d3c98),
	.w1(32'hb9817d5e),
	.w2(32'h3b5337fb),
	.w3(32'hbb687719),
	.w4(32'hbabd1d1d),
	.w5(32'hbb0c60e7),
	.w6(32'hba38333c),
	.w7(32'hb9ab7ba4),
	.w8(32'hbba3b87b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63aa33),
	.w1(32'h3bf0e5ad),
	.w2(32'hbb105cba),
	.w3(32'hba0d17ba),
	.w4(32'h3ba112dc),
	.w5(32'hbb21492d),
	.w6(32'hbb37d2d8),
	.w7(32'hb9b1d1c4),
	.w8(32'h396b269d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae430),
	.w1(32'h3b86ad43),
	.w2(32'hba86d7b5),
	.w3(32'hbb8a2dc4),
	.w4(32'h3c4ea267),
	.w5(32'h3b648006),
	.w6(32'hbbc00461),
	.w7(32'hbb4b3db6),
	.w8(32'hbbb637e6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8f00),
	.w1(32'h3a95137a),
	.w2(32'hbba9c64b),
	.w3(32'h3bc9f7d3),
	.w4(32'h3bd21321),
	.w5(32'h37f254f5),
	.w6(32'h3bc91380),
	.w7(32'h3bce0cbf),
	.w8(32'hb9c530e9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93ee09),
	.w1(32'h3aa83ae3),
	.w2(32'hbb7424aa),
	.w3(32'h3b62c8bd),
	.w4(32'hbb84e8c7),
	.w5(32'hbbb6c81a),
	.w6(32'h3bde25d1),
	.w7(32'h3c2e2232),
	.w8(32'hbc0d7fca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2298),
	.w1(32'hba4f75c8),
	.w2(32'hbbca6978),
	.w3(32'hbc90d607),
	.w4(32'hbb510048),
	.w5(32'hbb8f0ef5),
	.w6(32'hbc8a503b),
	.w7(32'hbc1c9a03),
	.w8(32'hbc38ff57),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324ec8),
	.w1(32'hb82d0da9),
	.w2(32'hbb2134f1),
	.w3(32'h3c0e1ef2),
	.w4(32'h3bef32ef),
	.w5(32'hbb303812),
	.w6(32'hba9ebaaa),
	.w7(32'hbb811eff),
	.w8(32'hba630603),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba374b0),
	.w1(32'h3bb7d2f2),
	.w2(32'hbb58375d),
	.w3(32'hbc3e039f),
	.w4(32'hbba5ced9),
	.w5(32'hbc1bc5e7),
	.w6(32'hbb4bea3e),
	.w7(32'hbbd10bb1),
	.w8(32'h3bbe34b0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaabf13),
	.w1(32'hbaa5bb3f),
	.w2(32'hbb0fff47),
	.w3(32'hbc767c75),
	.w4(32'hbc3abb58),
	.w5(32'hbbcadc29),
	.w6(32'h3a8070d2),
	.w7(32'hbbd8ac26),
	.w8(32'h3c4fce98),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b634ca9),
	.w1(32'h3b926a91),
	.w2(32'h3b258a6f),
	.w3(32'hbcc95192),
	.w4(32'hbc8d1cb7),
	.w5(32'h3c831d7b),
	.w6(32'h3bffef02),
	.w7(32'h3b4948f7),
	.w8(32'hba463c5b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44ae4f),
	.w1(32'hbb94ae56),
	.w2(32'h3b5d500a),
	.w3(32'h3c188bdc),
	.w4(32'hbc0954c0),
	.w5(32'h39a8fdaf),
	.w6(32'h3c47c9d9),
	.w7(32'h3c467273),
	.w8(32'h3a950292),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0deffd),
	.w1(32'h3b63fa64),
	.w2(32'h3b06d403),
	.w3(32'h3ba13556),
	.w4(32'hb93832cd),
	.w5(32'h3ae653e9),
	.w6(32'h3bb328b6),
	.w7(32'h39acb0aa),
	.w8(32'hbb275694),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739a581),
	.w1(32'hb986a099),
	.w2(32'hbb82649d),
	.w3(32'hbbcc449b),
	.w4(32'hbb1ce5e4),
	.w5(32'h3b6e0630),
	.w6(32'hbaf1996b),
	.w7(32'hbab2b3bb),
	.w8(32'hbac6f346),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4db83),
	.w1(32'hbacba7b0),
	.w2(32'h3bdff0cc),
	.w3(32'h3b248c41),
	.w4(32'h3ab19c56),
	.w5(32'h3bdfd1fb),
	.w6(32'hbb1e7f1c),
	.w7(32'hbb672d3f),
	.w8(32'hbbaa7d01),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4beaa8),
	.w1(32'hbbcf77cf),
	.w2(32'hbc9df642),
	.w3(32'hbb909947),
	.w4(32'h3a9bd428),
	.w5(32'hbc848125),
	.w6(32'hbc264d9b),
	.w7(32'hbc5dca9a),
	.w8(32'h3a5240da),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9e3aa),
	.w1(32'hba63ddb2),
	.w2(32'h3b04bc54),
	.w3(32'hbc99690f),
	.w4(32'hbc504cd4),
	.w5(32'h3b86d518),
	.w6(32'hbbbbf077),
	.w7(32'hbb926c13),
	.w8(32'h3ba4c6ce),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40af97),
	.w1(32'h3b87598a),
	.w2(32'h3c15c1a7),
	.w3(32'hbc3b6732),
	.w4(32'hbba54453),
	.w5(32'h3b080d14),
	.w6(32'h3c21c1b5),
	.w7(32'h3bb33b7c),
	.w8(32'h3c066658),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f689),
	.w1(32'h3b89f511),
	.w2(32'hbb35522a),
	.w3(32'hbbae8208),
	.w4(32'hbc35dad5),
	.w5(32'hbb5603bc),
	.w6(32'h3c3404f4),
	.w7(32'hbabbb7f5),
	.w8(32'hbbc2904c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8380d9),
	.w1(32'h3bf52bf3),
	.w2(32'h3a988a89),
	.w3(32'h3b18c13d),
	.w4(32'h3c634304),
	.w5(32'h3b1e5bbd),
	.w6(32'hbaa1fb96),
	.w7(32'h3c0a8329),
	.w8(32'h3b2fedec),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971c463),
	.w1(32'h3b3300dd),
	.w2(32'hbc18a48c),
	.w3(32'h3b7924d4),
	.w4(32'h3b5eaee5),
	.w5(32'hbc2395ad),
	.w6(32'h39a020ae),
	.w7(32'h3ae5a3b2),
	.w8(32'h3bec4f3c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1739bd),
	.w1(32'hbb673262),
	.w2(32'h3bc79dcf),
	.w3(32'hbc81f520),
	.w4(32'hbb9e8f60),
	.w5(32'h3aa0b99d),
	.w6(32'h3b4571b2),
	.w7(32'h3bd01204),
	.w8(32'hbb4ee589),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c768e94),
	.w1(32'h3c7751ef),
	.w2(32'h3beeb8cf),
	.w3(32'hbbbcecf9),
	.w4(32'hbbe99129),
	.w5(32'h39e4e588),
	.w6(32'hbb888d91),
	.w7(32'h3b103e89),
	.w8(32'hbc73521d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877696),
	.w1(32'h3bf099d6),
	.w2(32'h3c096f10),
	.w3(32'hbadfc3c2),
	.w4(32'h3b896b8c),
	.w5(32'h3c9546cb),
	.w6(32'hbc0bdc1a),
	.w7(32'hbba5f27c),
	.w8(32'h3ba3c106),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1db0b),
	.w1(32'hba9aacfa),
	.w2(32'hb9481a08),
	.w3(32'h3ca91b3f),
	.w4(32'h3c3f0439),
	.w5(32'hbb3ea53b),
	.w6(32'hbbee9035),
	.w7(32'hbc153a13),
	.w8(32'hbbcb0200),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4de64),
	.w1(32'h3b6735c3),
	.w2(32'h3b6757b6),
	.w3(32'hbb1e9d56),
	.w4(32'h39d03dff),
	.w5(32'h3b87c7cb),
	.w6(32'h3ae11073),
	.w7(32'h3b974e41),
	.w8(32'h3a94b406),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b9d81),
	.w1(32'h3c16f275),
	.w2(32'h3ad74505),
	.w3(32'h3b558560),
	.w4(32'h3bcbb006),
	.w5(32'hba6651d3),
	.w6(32'hbb3500b6),
	.w7(32'hba22d434),
	.w8(32'h3ac4d56f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189b82),
	.w1(32'h3ac8e526),
	.w2(32'hbb2ac1f3),
	.w3(32'hba8fcb6c),
	.w4(32'h3a6aa458),
	.w5(32'hbc0965ad),
	.w6(32'h3badade8),
	.w7(32'h3bab1d40),
	.w8(32'h3b789f3d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8290da),
	.w1(32'h3c070bc5),
	.w2(32'hb932b3e0),
	.w3(32'hbc754b67),
	.w4(32'hbbaeb274),
	.w5(32'h3a4b69f8),
	.w6(32'h3c6f2f6c),
	.w7(32'h3be25ccc),
	.w8(32'h3a7e4e4e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72f0d2),
	.w1(32'h3bbe62bd),
	.w2(32'hbc388992),
	.w3(32'hbb2a155c),
	.w4(32'h3a58a855),
	.w5(32'hba8d188f),
	.w6(32'h3b8fa47f),
	.w7(32'h3c3bfb9c),
	.w8(32'h3b96d1ec),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eaf58),
	.w1(32'h3bb99dc7),
	.w2(32'h3be7eda9),
	.w3(32'hbc9992d0),
	.w4(32'hbc87aacd),
	.w5(32'hbc6f3a1a),
	.w6(32'h3c3c1b74),
	.w7(32'h3c352e4b),
	.w8(32'h3bd638de),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc15bec),
	.w1(32'h3a8f5213),
	.w2(32'h3bcaac1c),
	.w3(32'hbcf27b66),
	.w4(32'hbcc8ffb1),
	.w5(32'h3c3bfb23),
	.w6(32'h3bf5f3c8),
	.w7(32'h3b89af44),
	.w8(32'h3c544935),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c831),
	.w1(32'hbbf7b98e),
	.w2(32'hbaef221d),
	.w3(32'h3aa0a6da),
	.w4(32'h3ba742e5),
	.w5(32'hbc0a4f73),
	.w6(32'h3aaba6e9),
	.w7(32'h3c10488e),
	.w8(32'hbb93cc6a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca26814),
	.w1(32'h3c99549a),
	.w2(32'h3b118ba4),
	.w3(32'hbc415ebf),
	.w4(32'hbc944223),
	.w5(32'hbbf7d88a),
	.w6(32'h3c63aadb),
	.w7(32'h3c81835a),
	.w8(32'h392a374f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8643b3),
	.w1(32'h3c99046d),
	.w2(32'h3a774635),
	.w3(32'hbc461a75),
	.w4(32'hbc2cabbb),
	.w5(32'h3ab051ad),
	.w6(32'h3c74eaea),
	.w7(32'h3c5a4fc0),
	.w8(32'hbb07a86e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c146d),
	.w1(32'h3b3080ab),
	.w2(32'hb9bbf23e),
	.w3(32'hbc22f381),
	.w4(32'hbc8da952),
	.w5(32'hbb87830f),
	.w6(32'hbc384409),
	.w7(32'hbc47dd49),
	.w8(32'hbbc302bd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c2268),
	.w1(32'hbabbefda),
	.w2(32'h3b8bda2f),
	.w3(32'hbba869b9),
	.w4(32'hba84318e),
	.w5(32'h3aee9e66),
	.w6(32'hbaabd09f),
	.w7(32'h3b9759d9),
	.w8(32'h3b9a4072),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2c7d2),
	.w1(32'hbbc86137),
	.w2(32'hbb6b455b),
	.w3(32'hbc361ae8),
	.w4(32'hbc2fdeb6),
	.w5(32'hbb51fc09),
	.w6(32'h3b8099fa),
	.w7(32'hba9340f9),
	.w8(32'hbbd0b3c9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dae56),
	.w1(32'hba871995),
	.w2(32'hbbd806ca),
	.w3(32'h3a1a5226),
	.w4(32'hba609d17),
	.w5(32'hbbe3ac7f),
	.w6(32'h39eea451),
	.w7(32'h3b5b4461),
	.w8(32'hbbb2c3d0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a661efa),
	.w1(32'hbb76ca10),
	.w2(32'hbb9d8668),
	.w3(32'hbaf948aa),
	.w4(32'hbb470393),
	.w5(32'hbbee3778),
	.w6(32'h3b108eee),
	.w7(32'h3b9875f1),
	.w8(32'hbb7e090f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3e1e9),
	.w1(32'h3bd7eac1),
	.w2(32'hbc275ff2),
	.w3(32'hbc1cd3c5),
	.w4(32'hb9b09f99),
	.w5(32'hbc01a79e),
	.w6(32'h3a4100f1),
	.w7(32'h3a7f60cf),
	.w8(32'hbc063ca4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c93f9),
	.w1(32'h3b9a05cd),
	.w2(32'hbba99033),
	.w3(32'hbc87259e),
	.w4(32'hba41242c),
	.w5(32'hbbdcc74a),
	.w6(32'hbbc108a4),
	.w7(32'hbb937b30),
	.w8(32'h3ba9c5de),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8158),
	.w1(32'h3c862195),
	.w2(32'hbb11f57e),
	.w3(32'hbc8d7969),
	.w4(32'hbc06172d),
	.w5(32'h3aebff9c),
	.w6(32'h3c854c4c),
	.w7(32'h3c66f362),
	.w8(32'h3958d8b3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23ad3f),
	.w1(32'h3bb75127),
	.w2(32'h3b79f7fb),
	.w3(32'hbc8c1523),
	.w4(32'hbc1af9bc),
	.w5(32'h3c0e8ec7),
	.w6(32'h3ae609b1),
	.w7(32'h3c003a1c),
	.w8(32'h3be4feb7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e48aa),
	.w1(32'h3c324296),
	.w2(32'hbb996917),
	.w3(32'h3bcad8aa),
	.w4(32'hbb4ba321),
	.w5(32'hbc28677c),
	.w6(32'h3c0523a8),
	.w7(32'h3a1d0d13),
	.w8(32'h3c225725),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ce1ac),
	.w1(32'h3b523c86),
	.w2(32'h3b9226f4),
	.w3(32'hbc30ee6d),
	.w4(32'hbc1e35c5),
	.w5(32'hbcbe78de),
	.w6(32'h3b2a0ff9),
	.w7(32'hba953bee),
	.w8(32'hbb6fac2e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c138aee),
	.w1(32'h3bb89564),
	.w2(32'h3b5dc980),
	.w3(32'hbd03bfac),
	.w4(32'hbc74b2ef),
	.w5(32'hbc026245),
	.w6(32'hbb3bce84),
	.w7(32'h3a4625ae),
	.w8(32'hbb851ece),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad42c),
	.w1(32'h3c77a237),
	.w2(32'h3aeef13e),
	.w3(32'hb97c74a9),
	.w4(32'hba03f284),
	.w5(32'h3877758f),
	.w6(32'hbbd958d0),
	.w7(32'hbc2432c1),
	.w8(32'h3c4fdee8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b52246),
	.w1(32'h3b8da4e6),
	.w2(32'hbb96d4cd),
	.w3(32'hbb6881df),
	.w4(32'h3b2d7348),
	.w5(32'h3aaf8746),
	.w6(32'h3c13b270),
	.w7(32'h3c4036c2),
	.w8(32'hbc460fcc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d492c),
	.w1(32'hbc1c6ded),
	.w2(32'h3b676d4f),
	.w3(32'h3bf68ced),
	.w4(32'h3bc681fb),
	.w5(32'hbaf85974),
	.w6(32'hbb397582),
	.w7(32'hba6f55a8),
	.w8(32'h3b92fd18),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa2122),
	.w1(32'h3b97e466),
	.w2(32'h3af6a322),
	.w3(32'hbbcbfb1e),
	.w4(32'hbba17f13),
	.w5(32'hbb63f258),
	.w6(32'h3c02df13),
	.w7(32'h3bd93104),
	.w8(32'h3c144ec7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9dfa8),
	.w1(32'h3b952e61),
	.w2(32'h3b164a5b),
	.w3(32'hbca8f96b),
	.w4(32'hbc931d94),
	.w5(32'hbb582726),
	.w6(32'h3c984e1a),
	.w7(32'h3c96e464),
	.w8(32'hbb0f964e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb526a),
	.w1(32'h3b725f5c),
	.w2(32'hbaf44ad5),
	.w3(32'hbba8c495),
	.w4(32'hbb05765c),
	.w5(32'hbb82a54c),
	.w6(32'h3b5f2a81),
	.w7(32'h3b8a3713),
	.w8(32'h3bbc2515),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22971),
	.w1(32'hbb2930b1),
	.w2(32'hbbef87ff),
	.w3(32'hba36deb3),
	.w4(32'h3a102177),
	.w5(32'hbab9ae6d),
	.w6(32'h3bc7b9c8),
	.w7(32'hbae1b019),
	.w8(32'hbb6e7f7d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2be0e),
	.w1(32'hbb9e4b7b),
	.w2(32'hbb5eeb5e),
	.w3(32'h3adc27fd),
	.w4(32'h3b15248b),
	.w5(32'hba55c375),
	.w6(32'hbb672ac6),
	.w7(32'hbadec864),
	.w8(32'hbad35e9c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8970be),
	.w1(32'hbad50d8b),
	.w2(32'h3a93b7a3),
	.w3(32'hb96a0916),
	.w4(32'h38561b05),
	.w5(32'hbc0c5dae),
	.w6(32'h3a18d114),
	.w7(32'h3a438257),
	.w8(32'h3b93c28d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45cfc2),
	.w1(32'hbb8e7886),
	.w2(32'h38153265),
	.w3(32'hbbcc11bb),
	.w4(32'hbc28bad7),
	.w5(32'hb9f65ed1),
	.w6(32'h3bc2636e),
	.w7(32'h3bc1d2f5),
	.w8(32'h3ad0aaab),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37fd37),
	.w1(32'hbb6164e6),
	.w2(32'hbc246331),
	.w3(32'hba091784),
	.w4(32'hbb2796dc),
	.w5(32'hbc3602ee),
	.w6(32'h3ad3f5bd),
	.w7(32'hb9aaa1fd),
	.w8(32'h3b8992d8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084874),
	.w1(32'hbc82bedb),
	.w2(32'hbb7880a2),
	.w3(32'hbc436588),
	.w4(32'hbc2d1d3d),
	.w5(32'hbb4faf50),
	.w6(32'h3c010894),
	.w7(32'h3a9a4603),
	.w8(32'h3b54a024),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe71a7),
	.w1(32'hba2ab8bc),
	.w2(32'h3be9e437),
	.w3(32'hbaf46aa4),
	.w4(32'h3b6e7cb2),
	.w5(32'h3bdb2786),
	.w6(32'h3aa5d307),
	.w7(32'h3c267693),
	.w8(32'h3b17aa61),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa99eb6),
	.w1(32'h38924605),
	.w2(32'h3c20ba1e),
	.w3(32'h3b98ad6b),
	.w4(32'h3b95f5ed),
	.w5(32'hbbeb2eb3),
	.w6(32'h3c1a3867),
	.w7(32'h3c329ad1),
	.w8(32'h3c362071),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed4746),
	.w1(32'h3c66dfc9),
	.w2(32'hbad2d334),
	.w3(32'hbcc4c34d),
	.w4(32'hbb6936cf),
	.w5(32'hbbe00d95),
	.w6(32'hba5e651f),
	.w7(32'hbbbd6ee5),
	.w8(32'h3a840f6e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe80bb),
	.w1(32'h3b7b065d),
	.w2(32'hbb53d385),
	.w3(32'hbc48610a),
	.w4(32'hbc0ecc06),
	.w5(32'h3c535481),
	.w6(32'h3bfe4065),
	.w7(32'h3c1b0616),
	.w8(32'hbb4c5320),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b563e92),
	.w1(32'h3b08fdf7),
	.w2(32'hba494ca9),
	.w3(32'h3d119083),
	.w4(32'h3d08780f),
	.w5(32'h3af6f181),
	.w6(32'hbc42034d),
	.w7(32'hbc41e870),
	.w8(32'h3b8fbab7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c429b94),
	.w1(32'h3a04bfeb),
	.w2(32'h3b9fee4e),
	.w3(32'hbc08fe72),
	.w4(32'hbc43a080),
	.w5(32'hbcb2422a),
	.w6(32'h3c976350),
	.w7(32'h3c1e1161),
	.w8(32'hbc303032),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b479),
	.w1(32'hbc5dd7ec),
	.w2(32'hbbad7d8e),
	.w3(32'hbcc06e0e),
	.w4(32'hbca0548f),
	.w5(32'h3baf9dc1),
	.w6(32'hbc89fa7a),
	.w7(32'hbc62f72e),
	.w8(32'hb97201bc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba97589),
	.w1(32'hbabe899e),
	.w2(32'hbb3db474),
	.w3(32'hba5179d7),
	.w4(32'h3c756b33),
	.w5(32'hbac7ab94),
	.w6(32'hb9c688c1),
	.w7(32'hbbd7dd8c),
	.w8(32'hbb7b79fc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89f091),
	.w1(32'h3b671cec),
	.w2(32'hbb162958),
	.w3(32'h3abcd003),
	.w4(32'h3be81a04),
	.w5(32'hbba7b378),
	.w6(32'hbb9028c0),
	.w7(32'hbb40cf72),
	.w8(32'h3b8b9fd5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c045a5f),
	.w1(32'h3a8e7d49),
	.w2(32'hbc10dea8),
	.w3(32'hbc289cd5),
	.w4(32'hbc7be2dc),
	.w5(32'hbc02afea),
	.w6(32'h3bcfc954),
	.w7(32'h3c0a63d4),
	.w8(32'hbb67c343),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8830d6),
	.w1(32'hbba92c54),
	.w2(32'h3c252b88),
	.w3(32'hbc059447),
	.w4(32'hbc08ced1),
	.w5(32'h3b9c0c05),
	.w6(32'h3c20b6ea),
	.w7(32'h3c119895),
	.w8(32'h3a8c5272),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d26c),
	.w1(32'h3c153492),
	.w2(32'h3874d32d),
	.w3(32'h3c038733),
	.w4(32'h3bbb098f),
	.w5(32'h3b67e84a),
	.w6(32'h39f173b0),
	.w7(32'h3c30a944),
	.w8(32'hba27c7c9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55aab4),
	.w1(32'hbac744c3),
	.w2(32'h3bc5e594),
	.w3(32'h3b9001cf),
	.w4(32'h3b678fcb),
	.w5(32'hbba1ee6b),
	.w6(32'hbb18e6ad),
	.w7(32'hba9cc619),
	.w8(32'h3c0fbab5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0673e),
	.w1(32'h3a99ddf6),
	.w2(32'h3b812a16),
	.w3(32'hbc2a8dc2),
	.w4(32'hbb02adea),
	.w5(32'h3ab04d00),
	.w6(32'h3c336f13),
	.w7(32'hb9be5941),
	.w8(32'hbb375061),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbba1bf),
	.w1(32'h3bc798c8),
	.w2(32'h3c0f4103),
	.w3(32'h3b9267bf),
	.w4(32'h3b9e6201),
	.w5(32'h3c69d596),
	.w6(32'h3b960bbb),
	.w7(32'h3b914ab3),
	.w8(32'h3c18788c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae1083),
	.w1(32'h3bf5bd1c),
	.w2(32'hbb844719),
	.w3(32'h3cbd3ccb),
	.w4(32'h3c5959e5),
	.w5(32'h3cf27d8e),
	.w6(32'h3ca4527a),
	.w7(32'h3c16c480),
	.w8(32'h3b945a1f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc890fa8),
	.w1(32'hbb4e4249),
	.w2(32'h3b784e10),
	.w3(32'h3d02880a),
	.w4(32'h3d02999e),
	.w5(32'h3a2163fe),
	.w6(32'h3c0ff50a),
	.w7(32'h3c6d559a),
	.w8(32'hbbc85fa4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116132),
	.w1(32'h3c35a3ea),
	.w2(32'hba89ec46),
	.w3(32'h3b137240),
	.w4(32'h3c22e694),
	.w5(32'h3b11ed5c),
	.w6(32'hbc32aa8e),
	.w7(32'hbbc73f5e),
	.w8(32'hba0e2060),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773700),
	.w1(32'hba8d73a6),
	.w2(32'h3b388ac9),
	.w3(32'h3a3ca905),
	.w4(32'h3acbdad1),
	.w5(32'hbb75e8d4),
	.w6(32'hbb79bb75),
	.w7(32'hbb1bc32d),
	.w8(32'h3c0a3f97),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa24b3b),
	.w1(32'h3a6b5eaf),
	.w2(32'h3c13127d),
	.w3(32'hbc0cda31),
	.w4(32'hbbaf9859),
	.w5(32'h3b5b6057),
	.w6(32'h3b14881f),
	.w7(32'h3bc19dfe),
	.w8(32'h3c00bf77),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ead48),
	.w1(32'hb798d7fa),
	.w2(32'hbc28ae31),
	.w3(32'h3c467b72),
	.w4(32'h3c30ed4c),
	.w5(32'h3c9c4a35),
	.w6(32'h3bd40320),
	.w7(32'h3b622c17),
	.w8(32'hb5b60d74),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f336d),
	.w1(32'hbb302af7),
	.w2(32'hbb9e9ea6),
	.w3(32'hbbb51506),
	.w4(32'hbbef3b9d),
	.w5(32'hbb936fbe),
	.w6(32'h3cd9c4b9),
	.w7(32'h3d0a63e5),
	.w8(32'hb9f60dfa),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a3ecc),
	.w1(32'hbb31cce3),
	.w2(32'hbbcd5bc7),
	.w3(32'hbc336a9a),
	.w4(32'h39b37f04),
	.w5(32'h3bd0dcba),
	.w6(32'hbb41d4a2),
	.w7(32'h3b9dd052),
	.w8(32'h3c584d5c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983024d),
	.w1(32'h3c06f162),
	.w2(32'h3b933f79),
	.w3(32'hbc64b215),
	.w4(32'hbb85e0c4),
	.w5(32'hbc548634),
	.w6(32'h3c0960f4),
	.w7(32'h3c0b38e1),
	.w8(32'h3a65c1fb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd49aca),
	.w1(32'h3c22a8be),
	.w2(32'hbb82e473),
	.w3(32'hbce794dd),
	.w4(32'hbc4c9929),
	.w5(32'h3a824deb),
	.w6(32'h3bcb7ec6),
	.w7(32'h3b73ec9c),
	.w8(32'h3a4480bd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6267),
	.w1(32'hbb5f9973),
	.w2(32'h3c3f863e),
	.w3(32'h397dfa61),
	.w4(32'hba64496b),
	.w5(32'h3c423c08),
	.w6(32'h3aa61def),
	.w7(32'h3ab9b4d5),
	.w8(32'h3bf17ff4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4efbcd),
	.w1(32'h3b09c219),
	.w2(32'hbc9c90d5),
	.w3(32'h3c8e272f),
	.w4(32'h3c962aa3),
	.w5(32'h3b278389),
	.w6(32'h3c39dc95),
	.w7(32'h3b1e301c),
	.w8(32'hbc8e7740),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8070e),
	.w1(32'hbc0915a3),
	.w2(32'hbb89b800),
	.w3(32'hbc14244a),
	.w4(32'hbcbc69a1),
	.w5(32'hbbf97b78),
	.w6(32'hbc7c70b9),
	.w7(32'hbbb746f6),
	.w8(32'h3c8de988),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaf446),
	.w1(32'h3ab66f84),
	.w2(32'h37cd1031),
	.w3(32'hbc796d64),
	.w4(32'hbc00502b),
	.w5(32'h3ac8460a),
	.w6(32'h3c49fb90),
	.w7(32'h3c92af9c),
	.w8(32'hb97d2dc8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2e1ca),
	.w1(32'h3aaae59a),
	.w2(32'hbb940a8c),
	.w3(32'h3c59940a),
	.w4(32'h3b404923),
	.w5(32'h3b301170),
	.w6(32'h3bcfd590),
	.w7(32'hba639613),
	.w8(32'h3b32a26d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22036b),
	.w1(32'h3ac791dc),
	.w2(32'h3bb913c4),
	.w3(32'h3bb1f8f9),
	.w4(32'h3b99d4d3),
	.w5(32'h39445a29),
	.w6(32'hba96ee22),
	.w7(32'hbb889d77),
	.w8(32'hba66ed78),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42ce76),
	.w1(32'h3c36a2d4),
	.w2(32'h399f80be),
	.w3(32'h3b78624e),
	.w4(32'h3bcfb618),
	.w5(32'hb9ed0a83),
	.w6(32'h3b8ff76d),
	.w7(32'h3c10c35e),
	.w8(32'hbaa015ff),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2064d7),
	.w1(32'h39ff5c8f),
	.w2(32'hb887dfe4),
	.w3(32'hba3cfbbb),
	.w4(32'h3a4043a9),
	.w5(32'hbb59c4a4),
	.w6(32'hb9e7c540),
	.w7(32'hb9ce6492),
	.w8(32'hb9431ad2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a335045),
	.w1(32'hbb508795),
	.w2(32'hbbb04b2b),
	.w3(32'h3a0920ac),
	.w4(32'hbad04eca),
	.w5(32'hbb6f270b),
	.w6(32'h3be50141),
	.w7(32'hbafee32a),
	.w8(32'hbc0ce69b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d4c85),
	.w1(32'hbbe04c54),
	.w2(32'h3aa11d94),
	.w3(32'h3b0c553b),
	.w4(32'hbb557a9f),
	.w5(32'hbaf4f82e),
	.w6(32'hbb58e028),
	.w7(32'hbb0a5c31),
	.w8(32'hbaca1383),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a250938),
	.w1(32'h38f1a3f9),
	.w2(32'h3a78635d),
	.w3(32'hbb0fad12),
	.w4(32'hba621386),
	.w5(32'h3bf3352e),
	.w6(32'hbb1c2e08),
	.w7(32'hbaa3942e),
	.w8(32'hbba184bf),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9d7e3),
	.w1(32'hbad4aa13),
	.w2(32'hbba0eb26),
	.w3(32'h3b0402ae),
	.w4(32'h3ba000af),
	.w5(32'hbb3dc28a),
	.w6(32'h3be7f42a),
	.w7(32'h3c1b2492),
	.w8(32'hbb3930e7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea49b6),
	.w1(32'hbbe8f5a3),
	.w2(32'h3b2dd492),
	.w3(32'hbb95f188),
	.w4(32'hbbbc35a4),
	.w5(32'hb9ae7c94),
	.w6(32'hbbc94437),
	.w7(32'hbbbb37f7),
	.w8(32'hbb1252f3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06f3a5),
	.w1(32'hbb5a70f3),
	.w2(32'hba730950),
	.w3(32'h3bf8accf),
	.w4(32'h3b4c0b6e),
	.w5(32'hb96b44c0),
	.w6(32'h3c257d6a),
	.w7(32'h3b9054dc),
	.w8(32'h39964b9f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb406d),
	.w1(32'hbb66eda3),
	.w2(32'hba9f0f6e),
	.w3(32'hb9fd5b93),
	.w4(32'h3b1bec8e),
	.w5(32'h3ae4cf27),
	.w6(32'h3b2d7453),
	.w7(32'h3b8bf239),
	.w8(32'h3b1b75ad),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873f82),
	.w1(32'hbb3700fa),
	.w2(32'hba797f33),
	.w3(32'h3add8884),
	.w4(32'hbb12b831),
	.w5(32'hbb89ed8a),
	.w6(32'hbb6d4dfa),
	.w7(32'hbbcf5736),
	.w8(32'hbc0df74b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c661),
	.w1(32'hba795e6b),
	.w2(32'h3868a435),
	.w3(32'h3c3f0d66),
	.w4(32'h3b5cea20),
	.w5(32'h3b13908e),
	.w6(32'h3c134f34),
	.w7(32'hbaf9d2f9),
	.w8(32'hbaaecef0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24164c),
	.w1(32'hba8058b8),
	.w2(32'h3b0c5ea2),
	.w3(32'h3c22bf74),
	.w4(32'h3a5ec93e),
	.w5(32'h3ad1fb27),
	.w6(32'h3bc5d83d),
	.w7(32'hbb68cbb0),
	.w8(32'h3b886f5c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbf314),
	.w1(32'hbc384576),
	.w2(32'hbb5546f6),
	.w3(32'h3af04cf4),
	.w4(32'h3b2f8b24),
	.w5(32'hbc4a9a3e),
	.w6(32'h3b60c06b),
	.w7(32'h39cb9639),
	.w8(32'hbc3db454),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c53ea),
	.w1(32'hbb8d2c8b),
	.w2(32'hb9f397eb),
	.w3(32'hbc950ce3),
	.w4(32'hbb754afa),
	.w5(32'h3b2cd0d1),
	.w6(32'hbc3b44fb),
	.w7(32'hbbb4d313),
	.w8(32'h3a394e23),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb321c33),
	.w1(32'hbb1386e1),
	.w2(32'hba89bba6),
	.w3(32'h3b78365c),
	.w4(32'h3ad97152),
	.w5(32'hbc2d6662),
	.w6(32'h3b37caf6),
	.w7(32'h3ad4221e),
	.w8(32'hbc59af90),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3378),
	.w1(32'h3c83a901),
	.w2(32'h3aafd3bd),
	.w3(32'hbc23e306),
	.w4(32'h3bb24408),
	.w5(32'hbba9706a),
	.w6(32'hba88cf9e),
	.w7(32'h3baf71bd),
	.w8(32'h39915b8a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a55f4),
	.w1(32'hbb4c168b),
	.w2(32'hbaf0b56c),
	.w3(32'hbb604b65),
	.w4(32'h3b33ff3d),
	.w5(32'hbb1d47c6),
	.w6(32'hb9ee81f7),
	.w7(32'h3b2c1777),
	.w8(32'hbc29c8a7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50d3eb),
	.w1(32'hbbaabda1),
	.w2(32'h3bdc708e),
	.w3(32'hbbf122c7),
	.w4(32'hbad736ec),
	.w5(32'h3bc89bed),
	.w6(32'hbc003a56),
	.w7(32'hbb97c9f3),
	.w8(32'h3b8c1b95),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73ea87),
	.w1(32'h3bbe8132),
	.w2(32'hbb089320),
	.w3(32'h3bc4518c),
	.w4(32'hbb48779c),
	.w5(32'hba905547),
	.w6(32'hba5a69f5),
	.w7(32'hb91c05ce),
	.w8(32'hbac43c35),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9c6c),
	.w1(32'hbb013505),
	.w2(32'hbb961522),
	.w3(32'h39b8f054),
	.w4(32'h3b31d3df),
	.w5(32'h3bc4b793),
	.w6(32'h3aab9c08),
	.w7(32'h3b4fd800),
	.w8(32'hba2e930c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1972a2),
	.w1(32'hbc5910af),
	.w2(32'h3bee6140),
	.w3(32'hbb90a3af),
	.w4(32'hbc14e5c1),
	.w5(32'h3bebaa19),
	.w6(32'hbc083edc),
	.w7(32'hbb7839b6),
	.w8(32'h3b89e79e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d3204),
	.w1(32'hbba65026),
	.w2(32'h3b00e655),
	.w3(32'hb96578a7),
	.w4(32'hbc248b70),
	.w5(32'hbc11a243),
	.w6(32'h3b21c59b),
	.w7(32'hbb126d68),
	.w8(32'hbc65f4ae),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b321),
	.w1(32'hba98de6d),
	.w2(32'h3c896ef7),
	.w3(32'hbc3c556d),
	.w4(32'hbbdb4dec),
	.w5(32'h3c58db7a),
	.w6(32'hbc24aff7),
	.w7(32'hbc1e5c1f),
	.w8(32'h3c5a408c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d9a4),
	.w1(32'hbb87016e),
	.w2(32'h3b517cea),
	.w3(32'h3bfc833b),
	.w4(32'hbb62c516),
	.w5(32'h3b47e7d4),
	.w6(32'h39d16f88),
	.w7(32'hbb89210f),
	.w8(32'h39ccd792),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c9261),
	.w1(32'hbba01627),
	.w2(32'h3b327dbb),
	.w3(32'h3ace4f67),
	.w4(32'hbb857e44),
	.w5(32'hbbda7889),
	.w6(32'hb9f127d3),
	.w7(32'hbbd6db7e),
	.w8(32'hbabd1886),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7ab46),
	.w1(32'h3a1d9755),
	.w2(32'hbb6411d8),
	.w3(32'hbaf0aeeb),
	.w4(32'hbb011e06),
	.w5(32'h3a5f9ea6),
	.w6(32'hbb57464c),
	.w7(32'hbb2f8d84),
	.w8(32'hb930553a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5b35e),
	.w1(32'h3b4a7589),
	.w2(32'hba97ff7b),
	.w3(32'h3bd32969),
	.w4(32'h3c0a1582),
	.w5(32'hbb8e4466),
	.w6(32'h3c4a8485),
	.w7(32'h3c55431f),
	.w8(32'hbbd85eb3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330870),
	.w1(32'h3ba610fb),
	.w2(32'h37f1e466),
	.w3(32'h385d729a),
	.w4(32'h3baf7ee6),
	.w5(32'hbb1f65c7),
	.w6(32'hbb35bbfe),
	.w7(32'hbac15f6e),
	.w8(32'hba9852ed),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa2863),
	.w1(32'hbb25a1f3),
	.w2(32'hba689d3a),
	.w3(32'hbb28e9c9),
	.w4(32'h3b333424),
	.w5(32'hbbbc59e7),
	.w6(32'hbabf0811),
	.w7(32'h3b85c7f0),
	.w8(32'h3b6aa4b6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64c56),
	.w1(32'hbbf12439),
	.w2(32'h3ad403e1),
	.w3(32'hbb061c93),
	.w4(32'hbbeb1113),
	.w5(32'hbb22d4b7),
	.w6(32'h3b17e0d6),
	.w7(32'h3abaa5f1),
	.w8(32'hbb29adac),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9879d6),
	.w1(32'h3a19fcfc),
	.w2(32'h3bc0f4a8),
	.w3(32'hb980778e),
	.w4(32'hbaa2e374),
	.w5(32'h3c130ed5),
	.w6(32'hbae890af),
	.w7(32'hbb7a9c09),
	.w8(32'h3bcee486),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa31d7),
	.w1(32'hbbcfd013),
	.w2(32'hbb8d7f51),
	.w3(32'h3ac451c1),
	.w4(32'hbb1abb7a),
	.w5(32'hbbd9df2e),
	.w6(32'h3970b7e2),
	.w7(32'hbbf48fb7),
	.w8(32'hbc30a59a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f6b7a),
	.w1(32'hbb7930da),
	.w2(32'hbc0d1ace),
	.w3(32'hb7525eee),
	.w4(32'hbb0e6e80),
	.w5(32'hbc82455b),
	.w6(32'h39fe728e),
	.w7(32'h3ba0a0b6),
	.w8(32'hbbd73680),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55c179),
	.w1(32'h399c6363),
	.w2(32'hbb16552f),
	.w3(32'hbc9de0f5),
	.w4(32'hbb9d44aa),
	.w5(32'hbbfc9065),
	.w6(32'hbc1b75d5),
	.w7(32'h3b8676d3),
	.w8(32'hbad9c192),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a548),
	.w1(32'h3a8a5e90),
	.w2(32'h3bb392d4),
	.w3(32'hbbad7626),
	.w4(32'h3ae30294),
	.w5(32'h3bd5543a),
	.w6(32'hbafc67ac),
	.w7(32'h38a0b0b5),
	.w8(32'h3a82b9b1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7cd92),
	.w1(32'h3c050b59),
	.w2(32'h3b2f8f62),
	.w3(32'h3c652538),
	.w4(32'h3c922db6),
	.w5(32'h3ae3508b),
	.w6(32'h3bd820a0),
	.w7(32'h3ab35092),
	.w8(32'h394479fc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1cace),
	.w1(32'h3b212f73),
	.w2(32'hbb1f72fc),
	.w3(32'h3ba0f66b),
	.w4(32'h3ab52330),
	.w5(32'hbb2d63d6),
	.w6(32'h3b4a1016),
	.w7(32'h373c398c),
	.w8(32'hbb453338),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1bf1),
	.w1(32'hbae355d8),
	.w2(32'h3bd951fa),
	.w3(32'h3a0201b4),
	.w4(32'hba877138),
	.w5(32'h3be968b7),
	.w6(32'hba906c5f),
	.w7(32'hbb1430e4),
	.w8(32'h3ad6d452),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97b58),
	.w1(32'hba475ac8),
	.w2(32'h3c06d2ef),
	.w3(32'h3be5f56e),
	.w4(32'hbb0e31ce),
	.w5(32'h3c3fb23c),
	.w6(32'h3b0e0dc3),
	.w7(32'hbbc9207f),
	.w8(32'h3b1f24ba),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cf4ba),
	.w1(32'hbb9fdd57),
	.w2(32'h3b897f68),
	.w3(32'h3c61bba0),
	.w4(32'hba961358),
	.w5(32'h3b1a30ff),
	.w6(32'h3be523f0),
	.w7(32'hbbfa1f87),
	.w8(32'h3b7bfa5e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e2d6),
	.w1(32'h3b08a2cb),
	.w2(32'hb9799f00),
	.w3(32'h3aa8d9d8),
	.w4(32'hba23a63c),
	.w5(32'h3ab09d3d),
	.w6(32'h3b236e1d),
	.w7(32'hb9d10e31),
	.w8(32'hb8506daa),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed3161),
	.w1(32'h38e704f8),
	.w2(32'hbb125a04),
	.w3(32'h3b5de3ab),
	.w4(32'h3af62a1d),
	.w5(32'h3b237ca4),
	.w6(32'h3b780807),
	.w7(32'h3bbb1c6a),
	.w8(32'h379a2e45),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2d129),
	.w1(32'hbb77fad0),
	.w2(32'h3ad3ff66),
	.w3(32'h3c03d483),
	.w4(32'hbb535394),
	.w5(32'hbb00a941),
	.w6(32'h3bc49dda),
	.w7(32'hbb2a268a),
	.w8(32'hbb83c414),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912b4b),
	.w1(32'hbbb73926),
	.w2(32'hbc2f7050),
	.w3(32'hbbab1229),
	.w4(32'hbc271a75),
	.w5(32'hbc8fe0bb),
	.w6(32'hbc10614a),
	.w7(32'hbbd42a63),
	.w8(32'hbc927711),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bfd21),
	.w1(32'h3c4d6320),
	.w2(32'h3a603044),
	.w3(32'h3be8aac7),
	.w4(32'h3c99294d),
	.w5(32'h3b005869),
	.w6(32'h3b74a6aa),
	.w7(32'h3c55f1ee),
	.w8(32'h3a26ae0c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808e56),
	.w1(32'hba4a8695),
	.w2(32'hbb759114),
	.w3(32'h3b29b7fa),
	.w4(32'h3b84cddd),
	.w5(32'hbb6cecec),
	.w6(32'h3a8293c7),
	.w7(32'h3a2cd367),
	.w8(32'hbbaa89f2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c912),
	.w1(32'hbbfaaeae),
	.w2(32'h3bb65c6e),
	.w3(32'hbb9fefcb),
	.w4(32'hbb5dd5fa),
	.w5(32'h3bf5b8fb),
	.w6(32'hbc0962a5),
	.w7(32'hbb87b732),
	.w8(32'h3bc5da65),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a3791),
	.w1(32'h3c229fcc),
	.w2(32'h3c194d8f),
	.w3(32'h3cb07dd2),
	.w4(32'h3c51c406),
	.w5(32'h3b6a759b),
	.w6(32'h3c5e45b4),
	.w7(32'h3bbf5353),
	.w8(32'hba4375ff),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103170),
	.w1(32'h3b52374f),
	.w2(32'h3bb2ced2),
	.w3(32'h3c2c5d9b),
	.w4(32'h3ba59aed),
	.w5(32'h3b852f92),
	.w6(32'h3c555f2d),
	.w7(32'h3b89a6c8),
	.w8(32'hbb059810),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3970a6),
	.w1(32'hbba69b5f),
	.w2(32'h3a6015fb),
	.w3(32'hbaa7a0ee),
	.w4(32'hbbb23112),
	.w5(32'h3c528d37),
	.w6(32'hbaf01dbe),
	.w7(32'hbbc62d48),
	.w8(32'h3aaab78b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f3d5d),
	.w1(32'h3b7ae7fd),
	.w2(32'hba1da330),
	.w3(32'h3cd5a4f1),
	.w4(32'h3c4258d6),
	.w5(32'hbb054321),
	.w6(32'h3c01b0c0),
	.w7(32'h3a1f6779),
	.w8(32'hbb56afa3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2212be),
	.w1(32'h3b840649),
	.w2(32'h3b3a54ec),
	.w3(32'hbb1a5f36),
	.w4(32'h3b212cb4),
	.w5(32'h3b126cf5),
	.w6(32'hbb7aa5ed),
	.w7(32'h3ad16fca),
	.w8(32'hb98a8e5d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8ae0),
	.w1(32'hbb0b861d),
	.w2(32'h3c47431d),
	.w3(32'h3ac4bb2c),
	.w4(32'hbadefd42),
	.w5(32'h3c55183b),
	.w6(32'hb8cecef5),
	.w7(32'hbbadce6a),
	.w8(32'h3c42a6c9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cb7ed),
	.w1(32'h3b96cfe8),
	.w2(32'h3a26b4a3),
	.w3(32'h3c614476),
	.w4(32'h3a859f59),
	.w5(32'h3b86e28c),
	.w6(32'h3ba0a94b),
	.w7(32'hbbaf956a),
	.w8(32'hbb835a9d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122a1c),
	.w1(32'hbad0a0d0),
	.w2(32'hbba9f99a),
	.w3(32'h3bd998e0),
	.w4(32'hbbd6b736),
	.w5(32'hbc1f6b26),
	.w6(32'hba8f6d84),
	.w7(32'hbb95f2e6),
	.w8(32'hbc1d86dd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33bed6),
	.w1(32'hbc4cc6f5),
	.w2(32'h3acd8a0f),
	.w3(32'hbc979396),
	.w4(32'hbc30eccf),
	.w5(32'hbc075907),
	.w6(32'hbc760fe8),
	.w7(32'hbbe05538),
	.w8(32'hbc1e2eb7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac46c7c),
	.w1(32'h3b2d080d),
	.w2(32'h3b764f7f),
	.w3(32'hbb82ca63),
	.w4(32'h3a768fb1),
	.w5(32'h3b38211c),
	.w6(32'hbc058560),
	.w7(32'hba842bcd),
	.w8(32'h3b61ae86),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d79ec),
	.w1(32'hb9a35564),
	.w2(32'h38ad333e),
	.w3(32'h3b5211b4),
	.w4(32'hbaeae989),
	.w5(32'h3add24a2),
	.w6(32'h3b4a36dd),
	.w7(32'hbb48c2d6),
	.w8(32'h3a06863f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c04513),
	.w1(32'h390e0f3e),
	.w2(32'h3c80e0d9),
	.w3(32'h3b40e5ec),
	.w4(32'h3af3e4ee),
	.w5(32'h3c418cd6),
	.w6(32'h3b50870e),
	.w7(32'h3b5678e8),
	.w8(32'h3bba822c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be106c7),
	.w1(32'hbb4dfdae),
	.w2(32'hbc113dae),
	.w3(32'h3ae855b4),
	.w4(32'hbba32b09),
	.w5(32'hbbe47c53),
	.w6(32'h3bdac2f0),
	.w7(32'hb952f1e0),
	.w8(32'hbb219662),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc112d6e),
	.w1(32'hbc2c717f),
	.w2(32'h3b96de75),
	.w3(32'hbaabb32d),
	.w4(32'hbb1a4ed7),
	.w5(32'hbb96bb54),
	.w6(32'h3ba6b2ee),
	.w7(32'h3b76a216),
	.w8(32'hbaf1b01b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a642079),
	.w1(32'h39eec22b),
	.w2(32'h3b62d4bf),
	.w3(32'hbbacda6b),
	.w4(32'hbbda07af),
	.w5(32'h3a181378),
	.w6(32'h3a9a764c),
	.w7(32'hb990f030),
	.w8(32'h3b835358),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96452c),
	.w1(32'hbc18b5ba),
	.w2(32'hbac3f8a1),
	.w3(32'hbad7d73e),
	.w4(32'hbc3ec65d),
	.w5(32'h3b36d589),
	.w6(32'hbabdae92),
	.w7(32'hbc23696e),
	.w8(32'h3a318322),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a0fe),
	.w1(32'hbb6e5b49),
	.w2(32'h3a472d68),
	.w3(32'h3b2e57a3),
	.w4(32'h38b007d3),
	.w5(32'h3b386eea),
	.w6(32'h39d329da),
	.w7(32'hba281532),
	.w8(32'h3b40a727),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f72ba),
	.w1(32'h3af83c30),
	.w2(32'h3c025477),
	.w3(32'h3bfdfcb5),
	.w4(32'h3b903f24),
	.w5(32'h3c4c4f34),
	.w6(32'h3bf021b5),
	.w7(32'h3ba49063),
	.w8(32'h3c264448),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad19f64),
	.w1(32'hbb57c7a2),
	.w2(32'h399e9f90),
	.w3(32'h3c1e394d),
	.w4(32'hbc05fe74),
	.w5(32'hba26397d),
	.w6(32'h3b5cfbe6),
	.w7(32'hbb8d1eb6),
	.w8(32'h3ad8bebe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a306),
	.w1(32'hbbffc84e),
	.w2(32'hbbcd2e43),
	.w3(32'hbbb17a9b),
	.w4(32'hbc2d7199),
	.w5(32'h3b0778ae),
	.w6(32'hbbb258fe),
	.w7(32'hbb99cb4d),
	.w8(32'hbbc084f7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc300855),
	.w1(32'hbc21a9fe),
	.w2(32'hbc1958ac),
	.w3(32'hb8097af3),
	.w4(32'h3a5c545e),
	.w5(32'hbca1cfca),
	.w6(32'hbb7e0bda),
	.w7(32'hbbb2ca84),
	.w8(32'hbc642ef8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4bd08),
	.w1(32'hbc5999a4),
	.w2(32'hba97508c),
	.w3(32'hbcea54fa),
	.w4(32'hbc2c4887),
	.w5(32'hbc441f58),
	.w6(32'hbc1fd490),
	.w7(32'hbba57d78),
	.w8(32'hbb13da97),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3dc8a),
	.w1(32'hba61f1c1),
	.w2(32'h3b0b98c6),
	.w3(32'hbbc3afa4),
	.w4(32'h3b5594c5),
	.w5(32'h3c07e66c),
	.w6(32'hb921d9ac),
	.w7(32'h3bc26593),
	.w8(32'h3bcec777),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0431fa),
	.w1(32'hbb47985e),
	.w2(32'hbbcd8ec7),
	.w3(32'hbad0f30e),
	.w4(32'h3b5ffbc3),
	.w5(32'hbc0a866e),
	.w6(32'hbb4f5ca1),
	.w7(32'h3bb5a2df),
	.w8(32'hbc68b8db),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf4de2),
	.w1(32'h3aef14aa),
	.w2(32'hbb9a2d83),
	.w3(32'hb9cfb24c),
	.w4(32'h3bc9c1f9),
	.w5(32'hbb249c57),
	.w6(32'hbc1c561d),
	.w7(32'hbbe188a1),
	.w8(32'hbb7b08b0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbca977),
	.w1(32'h3c089bcc),
	.w2(32'hb9d69ad5),
	.w3(32'h3bd36efb),
	.w4(32'h3bb5da38),
	.w5(32'h3aede296),
	.w6(32'h3baeb790),
	.w7(32'hbb3b872f),
	.w8(32'hbaeb4f07),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d6b54),
	.w1(32'h3b24b09e),
	.w2(32'h3bab73da),
	.w3(32'h3af77bbf),
	.w4(32'h3b45b1f7),
	.w5(32'h3ad6729c),
	.w6(32'hbb7af7ff),
	.w7(32'hbb2d76bc),
	.w8(32'hbaa9da85),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b247731),
	.w1(32'h3bd6e97c),
	.w2(32'h3b3290e7),
	.w3(32'h3ac7d0cd),
	.w4(32'h3b60527a),
	.w5(32'hbb1826be),
	.w6(32'hbaf7ad3a),
	.w7(32'h3b5a89c9),
	.w8(32'hbb566858),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a7142),
	.w1(32'h3b6e5a5f),
	.w2(32'hbb1de07c),
	.w3(32'h3c0585b8),
	.w4(32'hbaed4db0),
	.w5(32'hbb90b515),
	.w6(32'h3babe63c),
	.w7(32'hbb0c1a3e),
	.w8(32'hbbb5951f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b699f3d),
	.w1(32'h3ae20e87),
	.w2(32'hbaf25b8c),
	.w3(32'h3a4fa073),
	.w4(32'hbab726df),
	.w5(32'hbaa8319c),
	.w6(32'hbb923a91),
	.w7(32'hbb9027f8),
	.w8(32'hbb197069),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928054d),
	.w1(32'h39acde60),
	.w2(32'h3b5278a1),
	.w3(32'h39b4d08e),
	.w4(32'hb9f2ded0),
	.w5(32'h3b91abab),
	.w6(32'hbb457491),
	.w7(32'hbaecb868),
	.w8(32'hbafa48d1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22b780),
	.w1(32'hba736c5d),
	.w2(32'hbc4f2b84),
	.w3(32'hbad9ba44),
	.w4(32'h3ba881e7),
	.w5(32'hbc8ec57f),
	.w6(32'hbb40c243),
	.w7(32'h3af2cfde),
	.w8(32'hbc924295),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a774a),
	.w1(32'hbbc69517),
	.w2(32'hbbaad630),
	.w3(32'hbc8631cc),
	.w4(32'hbbb2e1bf),
	.w5(32'h3a7d53c7),
	.w6(32'hbc47d228),
	.w7(32'hbb3ddb28),
	.w8(32'hbb9be406),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46284d),
	.w1(32'h3a1369b6),
	.w2(32'hbc0e1c85),
	.w3(32'h3b97c60a),
	.w4(32'h3bcceff5),
	.w5(32'hbc906448),
	.w6(32'h3984cb22),
	.w7(32'h3a783635),
	.w8(32'hbc28ec5e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fa1e2),
	.w1(32'hbbde8eda),
	.w2(32'h3a582a58),
	.w3(32'hbcb264b5),
	.w4(32'hbc2b4fdb),
	.w5(32'h3c04c476),
	.w6(32'hbc213909),
	.w7(32'hbb159446),
	.w8(32'hbac56145),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1160cb),
	.w1(32'h3c04e109),
	.w2(32'hbb88451a),
	.w3(32'h3b74a5f8),
	.w4(32'h3c1ad93e),
	.w5(32'h3b8527d6),
	.w6(32'hbb154fa6),
	.w7(32'h3b9cb870),
	.w8(32'hbab1571d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85812b),
	.w1(32'h3b087447),
	.w2(32'hbaf79884),
	.w3(32'h3b990b49),
	.w4(32'h3ba6cff0),
	.w5(32'hbbfbd34c),
	.w6(32'h3bd4dc60),
	.w7(32'h3bf400f8),
	.w8(32'hbbd71cc9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd136),
	.w1(32'hbaffe9b5),
	.w2(32'hb983ab04),
	.w3(32'hbc195b8f),
	.w4(32'hbc008a55),
	.w5(32'hbb036ddb),
	.w6(32'hbb1fcf20),
	.w7(32'hbb95a3a9),
	.w8(32'hbbc621de),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b003a34),
	.w1(32'hb9c0e8af),
	.w2(32'h3b9b9e62),
	.w3(32'hbad7c454),
	.w4(32'h3bbcf317),
	.w5(32'h3c2151a4),
	.w6(32'h3b21758e),
	.w7(32'h3c45262d),
	.w8(32'h3bec6d0d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0859c9),
	.w1(32'hbabbb50c),
	.w2(32'hbb33e0e6),
	.w3(32'h3bdf3115),
	.w4(32'h3b53473d),
	.w5(32'hba87172b),
	.w6(32'h3b50e164),
	.w7(32'hbacddeea),
	.w8(32'hbb4528a8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38733e),
	.w1(32'hba4c3c49),
	.w2(32'hba9044fc),
	.w3(32'h3bdeed47),
	.w4(32'h3c06d0de),
	.w5(32'hba4558ac),
	.w6(32'h3a80aba5),
	.w7(32'h3b7f0e5d),
	.w8(32'hb9c9e878),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80aa8c),
	.w1(32'hbb2b8ebb),
	.w2(32'h3a04d95f),
	.w3(32'hba9c46b8),
	.w4(32'hba90061d),
	.w5(32'hbc21ea75),
	.w6(32'hbb54e98b),
	.w7(32'hbbafa04e),
	.w8(32'hbb35e936),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba923d99),
	.w1(32'hbae8f829),
	.w2(32'hbbdaa05d),
	.w3(32'h3b2748a7),
	.w4(32'h3c1b73c2),
	.w5(32'hbaa84404),
	.w6(32'h3a17ec1e),
	.w7(32'h39e3d500),
	.w8(32'hbbd8defa),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936b3a),
	.w1(32'h3be196d5),
	.w2(32'hbc2150b2),
	.w3(32'h3c12e0e6),
	.w4(32'h3c0b73b3),
	.w5(32'hbc69d04e),
	.w6(32'hbb83f7a7),
	.w7(32'h3ab1ca8b),
	.w8(32'hbc4033c7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a2997),
	.w1(32'hbbc83069),
	.w2(32'hb982031c),
	.w3(32'hbcaf77e6),
	.w4(32'hbc6e9c46),
	.w5(32'h3908f805),
	.w6(32'hbc99f217),
	.w7(32'hbc37e9a0),
	.w8(32'h3af95ac5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3daa0),
	.w1(32'hbb0d7dff),
	.w2(32'hb94a49d2),
	.w3(32'h396b57dc),
	.w4(32'hbaecb973),
	.w5(32'hba5eec33),
	.w6(32'h3aa10407),
	.w7(32'h39c76017),
	.w8(32'hba91e3d9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bcccf),
	.w1(32'hbb20be04),
	.w2(32'h3b4e43fc),
	.w3(32'hbb5cc143),
	.w4(32'hbb0e205f),
	.w5(32'h3b429195),
	.w6(32'hbb2c7fb4),
	.w7(32'hb9918e8c),
	.w8(32'hbb3f0f91),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d590),
	.w1(32'h3c101f99),
	.w2(32'hbb18d426),
	.w3(32'h3bda9a5e),
	.w4(32'h3c512e33),
	.w5(32'hba623875),
	.w6(32'h3a606180),
	.w7(32'h3b809e22),
	.w8(32'hbb0d2380),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a18839),
	.w1(32'h3b13f1fb),
	.w2(32'h3bc20a0b),
	.w3(32'h3af0feef),
	.w4(32'h3b0f1f74),
	.w5(32'hbbd95264),
	.w6(32'hbac81821),
	.w7(32'hba9f223c),
	.w8(32'h3b47aa56),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e4ea7),
	.w1(32'h3bb7a3ce),
	.w2(32'h3bddebd7),
	.w3(32'h3a4ea93f),
	.w4(32'h3b7effab),
	.w5(32'h3c128ede),
	.w6(32'hbbf98f59),
	.w7(32'hb99cb625),
	.w8(32'h3af12981),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becc269),
	.w1(32'h3bdda233),
	.w2(32'h3b224341),
	.w3(32'h3c005df8),
	.w4(32'hbb0e2446),
	.w5(32'h3c15b7b8),
	.w6(32'hbbddb248),
	.w7(32'hbb7c99b3),
	.w8(32'h3be10125),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda5de1),
	.w1(32'h39459652),
	.w2(32'h3b88d6d2),
	.w3(32'h3a9313a0),
	.w4(32'hbaaee7b8),
	.w5(32'h393d717e),
	.w6(32'hb9e989a3),
	.w7(32'hbb42728b),
	.w8(32'hbab28961),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule