module layer_10_featuremap_338(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dc047),
	.w1(32'hba1aa8b2),
	.w2(32'hbab1b1f7),
	.w3(32'h3a9189c9),
	.w4(32'h3a9f6765),
	.w5(32'hbacf3334),
	.w6(32'h3b112020),
	.w7(32'hba62d1ac),
	.w8(32'hbac41d26),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37214b),
	.w1(32'h397cf979),
	.w2(32'hbb513430),
	.w3(32'h3b34b461),
	.w4(32'h39ef535a),
	.w5(32'hbb971a2e),
	.w6(32'hb9948a81),
	.w7(32'hbbaf86cd),
	.w8(32'hb94d89e0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b875cdc),
	.w1(32'hba7c30b0),
	.w2(32'h3b9af5f4),
	.w3(32'hbb182363),
	.w4(32'hba79d233),
	.w5(32'h3a8cbb40),
	.w6(32'h3c220799),
	.w7(32'h3a84cbcf),
	.w8(32'hba562418),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44a2e6),
	.w1(32'hbb058ece),
	.w2(32'h38d400d1),
	.w3(32'h3b856ee3),
	.w4(32'h3a4f895c),
	.w5(32'hbb6c63ba),
	.w6(32'hbaa9f699),
	.w7(32'hbabc585d),
	.w8(32'hbc398208),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f4da),
	.w1(32'hbb7bf071),
	.w2(32'h3bba0693),
	.w3(32'hbbc8dddf),
	.w4(32'hbb655a99),
	.w5(32'h3a7f84be),
	.w6(32'hbc32eb86),
	.w7(32'hbba32190),
	.w8(32'hba5160e7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba384f33),
	.w1(32'hbaae3572),
	.w2(32'hba02b1bc),
	.w3(32'h3b4d7b95),
	.w4(32'h3ab4cc02),
	.w5(32'h39c71669),
	.w6(32'hbaf29ddb),
	.w7(32'hbb54a888),
	.w8(32'hbab3ace2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9610),
	.w1(32'hbb9bfc86),
	.w2(32'h3ac67205),
	.w3(32'h3bc02d70),
	.w4(32'h3b237255),
	.w5(32'h3a467718),
	.w6(32'h3b7b6bfe),
	.w7(32'h3acda062),
	.w8(32'hbb2e6df1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b19e),
	.w1(32'hbc098026),
	.w2(32'hba88fdf4),
	.w3(32'h3bd56fde),
	.w4(32'h3aeee9d2),
	.w5(32'hbbb35a09),
	.w6(32'h3cbeeec2),
	.w7(32'h3bee3158),
	.w8(32'hba10d92b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6663d3),
	.w1(32'hbaa158a3),
	.w2(32'hba9f347e),
	.w3(32'hb99d5a73),
	.w4(32'h39012ede),
	.w5(32'h3ac99102),
	.w6(32'hbaeb3d99),
	.w7(32'hbaaeef7a),
	.w8(32'h37c159ee),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05badf),
	.w1(32'hba6f45ab),
	.w2(32'h3b17527a),
	.w3(32'hba0c3038),
	.w4(32'hb9138f49),
	.w5(32'h3b308daf),
	.w6(32'h3acd4a68),
	.w7(32'h3a10592b),
	.w8(32'hba8a7351),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656690),
	.w1(32'hbb9c3191),
	.w2(32'h378d51e8),
	.w3(32'h3b384683),
	.w4(32'hba248dcd),
	.w5(32'hbb2d9878),
	.w6(32'hbb878535),
	.w7(32'hbb977aea),
	.w8(32'h3b2ad4c9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f2a09c),
	.w1(32'hbc0aa8b1),
	.w2(32'hbb3025f7),
	.w3(32'h3aa7ec2d),
	.w4(32'h3ba92136),
	.w5(32'hbbaa4f79),
	.w6(32'h3cf86645),
	.w7(32'h3c98a5e1),
	.w8(32'h37e1837b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99c6a0),
	.w1(32'h3a81a12b),
	.w2(32'h3b9a3686),
	.w3(32'hba7dfca6),
	.w4(32'h3a07794f),
	.w5(32'h3a07e0ca),
	.w6(32'h3b611775),
	.w7(32'h3bbe990c),
	.w8(32'hbb3e0348),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e14fe),
	.w1(32'h3ab30895),
	.w2(32'h3b106abf),
	.w3(32'hbbb555a9),
	.w4(32'hbb8d6751),
	.w5(32'hbae5b289),
	.w6(32'hbb42a186),
	.w7(32'hbb352092),
	.w8(32'hbb930c3f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a818d3c),
	.w1(32'h39bb7fd1),
	.w2(32'h39d10f68),
	.w3(32'h3b7aa53b),
	.w4(32'h3ad82e1d),
	.w5(32'h3aa81672),
	.w6(32'hbb2266a4),
	.w7(32'hbb44550f),
	.w8(32'hb95158ce),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffed50),
	.w1(32'h3bc4ef88),
	.w2(32'hbb3817e3),
	.w3(32'h3aa11215),
	.w4(32'h3bc846ba),
	.w5(32'h3a10458e),
	.w6(32'h389001c9),
	.w7(32'h3a6d2f5d),
	.w8(32'hba1fc398),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accb38c),
	.w1(32'hba0131e2),
	.w2(32'h39b02024),
	.w3(32'h3bd6b565),
	.w4(32'h3b2bae7e),
	.w5(32'hbb103fed),
	.w6(32'hb97800fa),
	.w7(32'hbb8805c5),
	.w8(32'h3aae0f5b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb344e),
	.w1(32'h3b29e4f9),
	.w2(32'h3b9d6a9e),
	.w3(32'h3a0969d3),
	.w4(32'hbae2a402),
	.w5(32'hbb327248),
	.w6(32'h3c2aad67),
	.w7(32'h3ba07bf5),
	.w8(32'hbc4c49ef),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f62e),
	.w1(32'h3aeb9168),
	.w2(32'hba98f0bd),
	.w3(32'hbb3957b3),
	.w4(32'hbb6a7044),
	.w5(32'hbb09468f),
	.w6(32'h39d5ce91),
	.w7(32'h3a1aa53c),
	.w8(32'hbaf70765),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc1481),
	.w1(32'hbbd3fbab),
	.w2(32'hbb389eed),
	.w3(32'hbbe83abe),
	.w4(32'hbbbc7df1),
	.w5(32'h3ab7335b),
	.w6(32'hbbb03d1a),
	.w7(32'hbac806c9),
	.w8(32'hbb536643),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69a61),
	.w1(32'h3a004c6b),
	.w2(32'h3ad13a4a),
	.w3(32'h3b4244dc),
	.w4(32'h3b828c0e),
	.w5(32'h3abd81bf),
	.w6(32'hbace253a),
	.w7(32'hbb2d4d85),
	.w8(32'h3a4035ef),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162c1f),
	.w1(32'hbb2c164c),
	.w2(32'hbb6c1dd3),
	.w3(32'hb9f51114),
	.w4(32'h3a234c0b),
	.w5(32'hbbbee6e6),
	.w6(32'hba4ca4da),
	.w7(32'h39bfd787),
	.w8(32'hbb753ab6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47195b),
	.w1(32'h3b00e6f6),
	.w2(32'hbb96325c),
	.w3(32'hbb913253),
	.w4(32'h3b7f9a5d),
	.w5(32'h3af4d537),
	.w6(32'h3ceead36),
	.w7(32'h3c15828b),
	.w8(32'hbc164bf1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e52c5),
	.w1(32'h3af98cdd),
	.w2(32'h3a8d59f6),
	.w3(32'h3b1f04c1),
	.w4(32'h3bf98c2f),
	.w5(32'h3b04de74),
	.w6(32'hbab68935),
	.w7(32'h3bd69aa0),
	.w8(32'hba3b4669),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb44ad2),
	.w1(32'h3b09d9ec),
	.w2(32'h3a35736f),
	.w3(32'hbb27dbe4),
	.w4(32'hbbabe535),
	.w5(32'h3b5f7de6),
	.w6(32'hbc20c53d),
	.w7(32'hbb67eac5),
	.w8(32'h3bbdc1d9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42dabc),
	.w1(32'hbb48c251),
	.w2(32'h3a33c15c),
	.w3(32'h3b354046),
	.w4(32'h3b2977f9),
	.w5(32'h3b856307),
	.w6(32'hbabf875c),
	.w7(32'hb94bd855),
	.w8(32'h39acccb5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30007b),
	.w1(32'hbaf90f78),
	.w2(32'h3adbe2be),
	.w3(32'h3b31fb6f),
	.w4(32'h3ab8b42c),
	.w5(32'h3909fb15),
	.w6(32'hbb1d1167),
	.w7(32'hba9f337c),
	.w8(32'hbb0eb12f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba640fd4),
	.w1(32'h3a868ca2),
	.w2(32'hbb83e0fc),
	.w3(32'hbc1cf4f9),
	.w4(32'hba0dc98d),
	.w5(32'h3b9e9ab9),
	.w6(32'hbc8385b0),
	.w7(32'hbbebfe3c),
	.w8(32'hbc285d98),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f54c1),
	.w1(32'hbb2b3634),
	.w2(32'hbaa0773c),
	.w3(32'hbb8bca82),
	.w4(32'hbbcd608c),
	.w5(32'hb9411015),
	.w6(32'hbbd8eb37),
	.w7(32'hbba16110),
	.w8(32'h3b06dc41),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf09695),
	.w1(32'hbb6bf25f),
	.w2(32'h3a20ad07),
	.w3(32'hb9201ed9),
	.w4(32'hba38af23),
	.w5(32'h3b8ed12f),
	.w6(32'hbc50fe5a),
	.w7(32'hbc10f114),
	.w8(32'hbb40bef4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6346),
	.w1(32'hbbd3276d),
	.w2(32'hbc11b24f),
	.w3(32'hbbbd9ba0),
	.w4(32'hbabd3a78),
	.w5(32'h3ab5fa1b),
	.w6(32'h3c5139c3),
	.w7(32'h3b073f9c),
	.w8(32'h3b6d4130),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da5e95),
	.w1(32'hbb1ed8e1),
	.w2(32'hb9942764),
	.w3(32'hb9213ec9),
	.w4(32'h3b1e4551),
	.w5(32'hbb754bfa),
	.w6(32'h3b9b33a0),
	.w7(32'h3bb93233),
	.w8(32'hbbf07229),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb273e22),
	.w1(32'h3afde42a),
	.w2(32'hbb4656b7),
	.w3(32'hbb788859),
	.w4(32'hbb6ff088),
	.w5(32'hba43d65e),
	.w6(32'hbb56909a),
	.w7(32'hbb748ad6),
	.w8(32'hb9c3806f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92819d),
	.w1(32'h3a177382),
	.w2(32'hb9d0e86e),
	.w3(32'hba9a1591),
	.w4(32'hba6692db),
	.w5(32'h3b683647),
	.w6(32'hbba3ad01),
	.w7(32'hbb684a73),
	.w8(32'hbbc06685),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cdb5d),
	.w1(32'h3b6ea134),
	.w2(32'h3a8310c6),
	.w3(32'h3a55bf7d),
	.w4(32'h3a88002b),
	.w5(32'hba7fa45a),
	.w6(32'hbbefdb80),
	.w7(32'hbbb3c918),
	.w8(32'h3b2027ff),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c085d),
	.w1(32'hbb741739),
	.w2(32'hb8d7eca7),
	.w3(32'h3b9e7b0f),
	.w4(32'h3b14f393),
	.w5(32'h3a72262c),
	.w6(32'h3b1631c6),
	.w7(32'hbb1d1fcd),
	.w8(32'hbc115896),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ac103),
	.w1(32'hbc3e008b),
	.w2(32'h3c22e8c0),
	.w3(32'hbbdf4c8d),
	.w4(32'hbbb4453f),
	.w5(32'h3c1cccc8),
	.w6(32'h3c8a3e25),
	.w7(32'hbaf9e6e9),
	.w8(32'h3bc3c521),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6989d),
	.w1(32'hbb14b36f),
	.w2(32'hbb75b342),
	.w3(32'hbb4e2757),
	.w4(32'hbb38b54d),
	.w5(32'h38b4daed),
	.w6(32'hbc0fea50),
	.w7(32'hbbac479a),
	.w8(32'h3c0d543e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf89ed),
	.w1(32'hbba2ab64),
	.w2(32'hbba964bc),
	.w3(32'hbb80c527),
	.w4(32'hbb8a02cd),
	.w5(32'h3b0fb58e),
	.w6(32'hbbc72e99),
	.w7(32'h3abfe3a5),
	.w8(32'h3b657194),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ac8b2),
	.w1(32'h3b23184f),
	.w2(32'h3ac0d59a),
	.w3(32'hbb6a2dd4),
	.w4(32'hbb00048b),
	.w5(32'hbb30cbbe),
	.w6(32'hbbda5744),
	.w7(32'hbb473f27),
	.w8(32'hbb041efd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df601),
	.w1(32'h3c094f77),
	.w2(32'h3b590262),
	.w3(32'hbbd52ea5),
	.w4(32'hba91050a),
	.w5(32'h3aa136df),
	.w6(32'h3c496e74),
	.w7(32'h3bc439b6),
	.w8(32'h3a4c8131),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30c02),
	.w1(32'hbb098bb8),
	.w2(32'h3b1ae0df),
	.w3(32'h3ace74eb),
	.w4(32'h3b347a60),
	.w5(32'hbac00a41),
	.w6(32'hbb83a17d),
	.w7(32'h39b5b324),
	.w8(32'h3b1ae8ff),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7f611),
	.w1(32'h3b4d05f2),
	.w2(32'h3a492359),
	.w3(32'hbb85780d),
	.w4(32'hbb85474b),
	.w5(32'hb927215f),
	.w6(32'hba423dce),
	.w7(32'hbaf53c12),
	.w8(32'h3ac14ba2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1e0b),
	.w1(32'hbba6a000),
	.w2(32'hbb16ffa4),
	.w3(32'h3baad133),
	.w4(32'h3be75e0e),
	.w5(32'hbb01c13f),
	.w6(32'hbb191249),
	.w7(32'hbc111d11),
	.w8(32'hbb7167bb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf35cf),
	.w1(32'hbbadee32),
	.w2(32'hbb9c497e),
	.w3(32'hbbd78cd2),
	.w4(32'hbb1afa92),
	.w5(32'h3bdbdff1),
	.w6(32'hbc80170c),
	.w7(32'hbaf8dae6),
	.w8(32'h3c4780e7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8c9df),
	.w1(32'hbba9632c),
	.w2(32'hba125e0f),
	.w3(32'h3a9792a3),
	.w4(32'hbaaca604),
	.w5(32'h3af0ba58),
	.w6(32'hbb154d5d),
	.w7(32'hbadd4056),
	.w8(32'h3c063be0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d53c3),
	.w1(32'hbb4fb388),
	.w2(32'h3b58385c),
	.w3(32'hbb6da0ac),
	.w4(32'h3a0dc17c),
	.w5(32'hba720e39),
	.w6(32'hbb919410),
	.w7(32'hbb257f45),
	.w8(32'hbb46d39d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104524),
	.w1(32'hbb6258dc),
	.w2(32'h3a9854f7),
	.w3(32'h3a7bac03),
	.w4(32'hbac52016),
	.w5(32'hbbfbf543),
	.w6(32'h3c5f3561),
	.w7(32'h3ba937ed),
	.w8(32'hbbf7fc23),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52da1d),
	.w1(32'hbb3e1ad1),
	.w2(32'hbb3bac1d),
	.w3(32'hbb52bd61),
	.w4(32'hbabdc247),
	.w5(32'h38efb279),
	.w6(32'hbb8298eb),
	.w7(32'hbaf9b135),
	.w8(32'hbaaaa049),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee2cb),
	.w1(32'hbb52d2fe),
	.w2(32'hba99f7fe),
	.w3(32'h3a99a5ce),
	.w4(32'h3a84661b),
	.w5(32'h3bc7de5a),
	.w6(32'hba6b0213),
	.w7(32'hba8850c4),
	.w8(32'h3ab45d53),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c99ff),
	.w1(32'h3a1295d1),
	.w2(32'hb8e75836),
	.w3(32'h3b85a3e3),
	.w4(32'h3a91c628),
	.w5(32'hb903d998),
	.w6(32'hbb178b5d),
	.w7(32'h3a378a91),
	.w8(32'h3ac7321b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5f636),
	.w1(32'hbb3f9a82),
	.w2(32'hbaefe0ec),
	.w3(32'hbaabbb78),
	.w4(32'h3aa709bb),
	.w5(32'hb9032923),
	.w6(32'hba3312b5),
	.w7(32'h3ba054fd),
	.w8(32'hbb02f0a1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c41c87),
	.w1(32'hb9d84aef),
	.w2(32'hbb0d0eec),
	.w3(32'hba90cd97),
	.w4(32'h3ae539cd),
	.w5(32'hbac831dd),
	.w6(32'h3c3161f9),
	.w7(32'h3acee98a),
	.w8(32'hbbbc9070),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4f4f7),
	.w1(32'h3b3ab54e),
	.w2(32'h3a206d16),
	.w3(32'hbb5adce3),
	.w4(32'h3b0a44bf),
	.w5(32'hbba6ecf7),
	.w6(32'h3ca3c654),
	.w7(32'h3bf64724),
	.w8(32'hbc004f17),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe5c55),
	.w1(32'hbbb7e60c),
	.w2(32'hbb1013af),
	.w3(32'hbba8cbf5),
	.w4(32'hbb31dfcf),
	.w5(32'hbb0f9c4b),
	.w6(32'hbb7ed034),
	.w7(32'h3acc1d49),
	.w8(32'hbbd550a5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39442306),
	.w1(32'h3c4cfcd3),
	.w2(32'h3bf0efd1),
	.w3(32'hba3eb908),
	.w4(32'h3b518ad1),
	.w5(32'h39076b5a),
	.w6(32'hbbc52519),
	.w7(32'hbb075cc6),
	.w8(32'hbb0ace66),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a5f39a),
	.w1(32'h3c1987ed),
	.w2(32'h3b44f243),
	.w3(32'hbb065dcc),
	.w4(32'h3bb12834),
	.w5(32'hbb6afdaf),
	.w6(32'hba08f17b),
	.w7(32'h3b143f28),
	.w8(32'hbadacdb3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3102f3),
	.w1(32'h3b663016),
	.w2(32'h39979498),
	.w3(32'h3b2852c2),
	.w4(32'hbadf17ee),
	.w5(32'h3a6bbfb5),
	.w6(32'h3baf1ddd),
	.w7(32'hba852ce7),
	.w8(32'hbb0a124f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51b04d),
	.w1(32'hbb93fdcf),
	.w2(32'hbaeb51a8),
	.w3(32'h3a666323),
	.w4(32'h3ad06735),
	.w5(32'h3b50361f),
	.w6(32'hbb13af3d),
	.w7(32'hbabc5e52),
	.w8(32'h3b9fddc6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b399924),
	.w1(32'hbb3e216c),
	.w2(32'hbb1e9499),
	.w3(32'hbb75a3bd),
	.w4(32'hbba862a1),
	.w5(32'hba8efcc8),
	.w6(32'h3b6bdaf6),
	.w7(32'hbb14dac3),
	.w8(32'hbb68d85c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3e630),
	.w1(32'hbb0a1707),
	.w2(32'hba329546),
	.w3(32'hba6aa54d),
	.w4(32'hbb14b421),
	.w5(32'hba239b24),
	.w6(32'h3aa214b8),
	.w7(32'h39d5be02),
	.w8(32'hbb2486c5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1bbe6),
	.w1(32'h3b704d07),
	.w2(32'h3ae3f5cd),
	.w3(32'h3b6b4fd2),
	.w4(32'h3afef6e9),
	.w5(32'h3ba98412),
	.w6(32'hbba1c4fe),
	.w7(32'hbbac5e67),
	.w8(32'hbc2d13e7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79546d),
	.w1(32'hbb6085be),
	.w2(32'hb9e6b1e4),
	.w3(32'hb9c7fa2c),
	.w4(32'hbb720b06),
	.w5(32'hbb1e0dad),
	.w6(32'hbb9265af),
	.w7(32'h3a16f4bf),
	.w8(32'hbbe1f014),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e11c4),
	.w1(32'h3c54c2ce),
	.w2(32'h3bd814ec),
	.w3(32'hbac7bc07),
	.w4(32'h3bed0fbe),
	.w5(32'hbaa42634),
	.w6(32'hbb9ce9da),
	.w7(32'h383e3237),
	.w8(32'hbba83560),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0644ee),
	.w1(32'hbabd5d0a),
	.w2(32'hbaf18b00),
	.w3(32'hb9e86b3d),
	.w4(32'hb9b87973),
	.w5(32'hbbfd4a4b),
	.w6(32'hbc06e8d2),
	.w7(32'hbb7e4bfb),
	.w8(32'hbc316ee4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010263),
	.w1(32'hbbf2b6d3),
	.w2(32'hbb9e8192),
	.w3(32'hbc0fd584),
	.w4(32'hbb3e1ee4),
	.w5(32'h39b05594),
	.w6(32'h3bad9540),
	.w7(32'h3b817f6e),
	.w8(32'hbb5bbacf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966ab3),
	.w1(32'hbbb18e46),
	.w2(32'hbb883a93),
	.w3(32'hbb6216f1),
	.w4(32'hbb2e3612),
	.w5(32'h3b60885a),
	.w6(32'h3c52f617),
	.w7(32'hbb8c41d6),
	.w8(32'hbc39f0bf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a729),
	.w1(32'hbb448470),
	.w2(32'hbb5bdc7d),
	.w3(32'h3c6426f2),
	.w4(32'h3b9ccc54),
	.w5(32'hbb90dac4),
	.w6(32'h3b280968),
	.w7(32'h3affc305),
	.w8(32'hbb062768),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13f4ba),
	.w1(32'hbbf44f7b),
	.w2(32'hbba2fe2c),
	.w3(32'hba9f7c96),
	.w4(32'hbbb688c2),
	.w5(32'h3b6436f5),
	.w6(32'hbbce9f9c),
	.w7(32'hbbdf7d60),
	.w8(32'h3c5a745b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7c041),
	.w1(32'hb984bec7),
	.w2(32'hba506e46),
	.w3(32'h3a6dc300),
	.w4(32'h3b91a834),
	.w5(32'h3bbd6df0),
	.w6(32'hbbecaf73),
	.w7(32'h3b866484),
	.w8(32'h3c30c992),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a954f),
	.w1(32'h3b737caf),
	.w2(32'hbaf77f6a),
	.w3(32'hbb777b05),
	.w4(32'hbb03558c),
	.w5(32'hbb015001),
	.w6(32'hbaab61ac),
	.w7(32'hbba03d6a),
	.w8(32'hbaed8ba5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec116),
	.w1(32'hba45543b),
	.w2(32'hba5db19f),
	.w3(32'h36f98545),
	.w4(32'h3b1c40cd),
	.w5(32'hba56782c),
	.w6(32'h3b38506d),
	.w7(32'hbab960bc),
	.w8(32'h3b821fbb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f2576),
	.w1(32'h3acec3ac),
	.w2(32'h3a8c79d3),
	.w3(32'hba2a7ad8),
	.w4(32'h3b04b6f0),
	.w5(32'hbbb1afa5),
	.w6(32'h3b5a9142),
	.w7(32'hba9b0d22),
	.w8(32'hbbb43553),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae34e2c),
	.w1(32'h3b836f2a),
	.w2(32'h3bb80fe1),
	.w3(32'hbb25ebce),
	.w4(32'hbb4bc1fa),
	.w5(32'h3a32a12c),
	.w6(32'hbaf69799),
	.w7(32'h3b11ef05),
	.w8(32'hbb84b0fe),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5a4e3),
	.w1(32'hba8dd48e),
	.w2(32'hbac30590),
	.w3(32'h3b89b182),
	.w4(32'hb9be209f),
	.w5(32'hbb915f7b),
	.w6(32'hba2af9fc),
	.w7(32'hbba5709b),
	.w8(32'hb9c86d7b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9411b1),
	.w1(32'h3bc397b6),
	.w2(32'h3bcb3690),
	.w3(32'hbbec5bc6),
	.w4(32'hbb2fc856),
	.w5(32'hbba94efb),
	.w6(32'h3bff89a5),
	.w7(32'h3c1bdce3),
	.w8(32'hbbb34a44),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade281d),
	.w1(32'hbb311154),
	.w2(32'hbb539593),
	.w3(32'hbbe3af4e),
	.w4(32'hbb947d0c),
	.w5(32'hbb8b7b67),
	.w6(32'h3d22388d),
	.w7(32'h3c8340c6),
	.w8(32'hba8872f8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a417d),
	.w1(32'hbb41a953),
	.w2(32'hbb88ac25),
	.w3(32'hbb97a04a),
	.w4(32'h3b1b6aff),
	.w5(32'h3abd57d3),
	.w6(32'hbb8dc388),
	.w7(32'h3b51e1d8),
	.w8(32'h3ad353c1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e369),
	.w1(32'hba64ec3e),
	.w2(32'hba82dcc5),
	.w3(32'h39dd88c6),
	.w4(32'hbb560d1e),
	.w5(32'h3b0aa7a9),
	.w6(32'h3ba86376),
	.w7(32'hbabfa019),
	.w8(32'hbad7a3b4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f13b),
	.w1(32'hbaef4d09),
	.w2(32'hbb8bb1c2),
	.w3(32'h3b341a1d),
	.w4(32'h3b1dacda),
	.w5(32'hba852a74),
	.w6(32'h3b6f02e5),
	.w7(32'hbb6d2f32),
	.w8(32'hbc0a9873),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ad1ee),
	.w1(32'h3b5373d7),
	.w2(32'hbb3bcee1),
	.w3(32'hbc452971),
	.w4(32'hb97d8203),
	.w5(32'hbb6f7e66),
	.w6(32'hbba503a8),
	.w7(32'h3a79d72a),
	.w8(32'hbba07909),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152c7a),
	.w1(32'h3af8c448),
	.w2(32'h3b803041),
	.w3(32'hbc0731e3),
	.w4(32'hbb967654),
	.w5(32'hbb16803e),
	.w6(32'h3acd167e),
	.w7(32'h3afbddcd),
	.w8(32'hbb1be2a4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebf6c7),
	.w1(32'hbb793900),
	.w2(32'hbc31e493),
	.w3(32'hbbd51e39),
	.w4(32'hbb61657b),
	.w5(32'h3b994393),
	.w6(32'h3c3de196),
	.w7(32'hbb55c1aa),
	.w8(32'hba5e8a11),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba042b42),
	.w1(32'hbb1f3191),
	.w2(32'h3bb5ef7e),
	.w3(32'h3b131797),
	.w4(32'hbb770f63),
	.w5(32'hbb32ffdf),
	.w6(32'hbbb73241),
	.w7(32'hbad71190),
	.w8(32'h3ab51b69),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091da9),
	.w1(32'h3c1621b4),
	.w2(32'hbb6ef7a1),
	.w3(32'hbba7a007),
	.w4(32'hba1c8a58),
	.w5(32'hba1718cb),
	.w6(32'h3c96daaf),
	.w7(32'h3c0ff876),
	.w8(32'h3a3c3d6a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a11e0),
	.w1(32'hbc108a67),
	.w2(32'hbbb0be48),
	.w3(32'hbb2589d4),
	.w4(32'h3ba5838e),
	.w5(32'h3adcbc3e),
	.w6(32'hba8ad515),
	.w7(32'hbb8cea40),
	.w8(32'hb9183f3c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62c269),
	.w1(32'h3b233e75),
	.w2(32'h3b077884),
	.w3(32'h3bb3f75c),
	.w4(32'h3b81925a),
	.w5(32'hb880fd7f),
	.w6(32'hb8d6a662),
	.w7(32'hbb046ab5),
	.w8(32'h3b734931),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c5efd),
	.w1(32'hbba0bc9b),
	.w2(32'hbb44209f),
	.w3(32'hba34ee85),
	.w4(32'h3955df8f),
	.w5(32'hba64506e),
	.w6(32'h3c588ca5),
	.w7(32'h3c12a753),
	.w8(32'hbb240c42),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e4c3f),
	.w1(32'hbb513587),
	.w2(32'hbb3eecc7),
	.w3(32'h3b99a3b1),
	.w4(32'h3b1540bd),
	.w5(32'hba1da91e),
	.w6(32'hbb8ce7c1),
	.w7(32'hb999bb49),
	.w8(32'h3b09ec4c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14e10b),
	.w1(32'hbb859a88),
	.w2(32'h3bf9804f),
	.w3(32'hbb5af483),
	.w4(32'hbb2bd9ad),
	.w5(32'hbb3dad80),
	.w6(32'h3b68d5aa),
	.w7(32'h3b83292f),
	.w8(32'hbbbf7238),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc47e),
	.w1(32'hba35fe2d),
	.w2(32'hbae22a25),
	.w3(32'hbb08264d),
	.w4(32'h3a30fe00),
	.w5(32'hbb3459d8),
	.w6(32'hbc20a770),
	.w7(32'h3a171718),
	.w8(32'hbafdf6c8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63ca43),
	.w1(32'hbbfbb17a),
	.w2(32'hbab814b7),
	.w3(32'hbbb4ccf9),
	.w4(32'hbb521a2c),
	.w5(32'h3ba36338),
	.w6(32'h3b824d30),
	.w7(32'hbae00c85),
	.w8(32'hbc2025f7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7317f),
	.w1(32'h3a5df927),
	.w2(32'hbb0e6fc8),
	.w3(32'h3becc358),
	.w4(32'h3bf9b009),
	.w5(32'h3b719fdf),
	.w6(32'hbbdf946f),
	.w7(32'h3b374cc0),
	.w8(32'h3b842f84),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27111d),
	.w1(32'h3bc4b796),
	.w2(32'h3bc0e589),
	.w3(32'h3b0971a2),
	.w4(32'h3b320365),
	.w5(32'hbb3630d4),
	.w6(32'h3c0b6396),
	.w7(32'h3baefd9d),
	.w8(32'hbba08e1c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9176a1),
	.w1(32'hbb175910),
	.w2(32'hbb699535),
	.w3(32'hbb3b80ea),
	.w4(32'h3b85bd22),
	.w5(32'h3a3df5ac),
	.w6(32'hbb77fe5b),
	.w7(32'hbad36efa),
	.w8(32'h3bd5a065),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac29fa4),
	.w1(32'hbbac78e3),
	.w2(32'hbb699053),
	.w3(32'h390f53b8),
	.w4(32'h3afa3047),
	.w5(32'h3b253fd3),
	.w6(32'h3b54f8aa),
	.w7(32'h3c01a056),
	.w8(32'h3a382fab),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3a882),
	.w1(32'h3b05a154),
	.w2(32'h3a5cbf4c),
	.w3(32'hbb4b1142),
	.w4(32'hbb4498f2),
	.w5(32'h3b986d72),
	.w6(32'h3ad8faa6),
	.w7(32'h3bc77259),
	.w8(32'hb896bd13),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1e038),
	.w1(32'h3bc0232b),
	.w2(32'hbb43e611),
	.w3(32'hbb89018f),
	.w4(32'h3b1b962e),
	.w5(32'h392f959b),
	.w6(32'h3c9e9796),
	.w7(32'h3c8cfffc),
	.w8(32'hbab9f088),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021b5e),
	.w1(32'hbb5b5a09),
	.w2(32'hbb04af49),
	.w3(32'hbbdd2f9c),
	.w4(32'hbb4b3295),
	.w5(32'h3bb611b5),
	.w6(32'h3bf8e739),
	.w7(32'h3b4e2bb3),
	.w8(32'h3a4c7c8e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f068),
	.w1(32'hbc57eab8),
	.w2(32'h3c0717f4),
	.w3(32'h3c38e893),
	.w4(32'hbbbf82f9),
	.w5(32'hbb5a771b),
	.w6(32'h3c6ff95b),
	.w7(32'h3bebbf74),
	.w8(32'h3c1f9aeb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c369a),
	.w1(32'hba96bdb2),
	.w2(32'hbaadbd33),
	.w3(32'h3ad6cee2),
	.w4(32'hbb13a2ba),
	.w5(32'hbaeede4e),
	.w6(32'hbba55bdd),
	.w7(32'h39f29774),
	.w8(32'h3903d1ea),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068802),
	.w1(32'h3960a13a),
	.w2(32'h3aadce9c),
	.w3(32'hb9a20a5f),
	.w4(32'h3af86511),
	.w5(32'h3b474a31),
	.w6(32'hbb6f214f),
	.w7(32'h3b1b86e0),
	.w8(32'h3bb6beb0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81b0dd),
	.w1(32'hbb752aa9),
	.w2(32'h3b6b70df),
	.w3(32'hbb42a86f),
	.w4(32'hbb263a96),
	.w5(32'h3add3635),
	.w6(32'h3c7c8434),
	.w7(32'h3b4511cb),
	.w8(32'hbabab092),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cfcd7),
	.w1(32'hbaa077b0),
	.w2(32'hb828f9c1),
	.w3(32'hb9f430f0),
	.w4(32'hb93fd482),
	.w5(32'h3a18bd38),
	.w6(32'hba2dd52e),
	.w7(32'hb9385d2b),
	.w8(32'h37c2208e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6071a),
	.w1(32'hbc3075e9),
	.w2(32'h3c32f427),
	.w3(32'h3c088769),
	.w4(32'hbbd87648),
	.w5(32'h3b193224),
	.w6(32'h3c8f78dd),
	.w7(32'h3c37ff7a),
	.w8(32'h3c1adbd3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f07a0),
	.w1(32'hbb3b5efd),
	.w2(32'h3aebd0e9),
	.w3(32'h3acb4255),
	.w4(32'hbb689aea),
	.w5(32'h39950a68),
	.w6(32'h3ba63a18),
	.w7(32'h3ae8a464),
	.w8(32'h3b399b6d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87cafc1),
	.w1(32'h38c32b3c),
	.w2(32'h36ffc6f4),
	.w3(32'hb983ac2e),
	.w4(32'h37bcf7f8),
	.w5(32'h384e246d),
	.w6(32'hba01246f),
	.w7(32'hb8cb1bd7),
	.w8(32'hb7e3b905),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a943a1a),
	.w1(32'h3a32bd30),
	.w2(32'hbada455c),
	.w3(32'hb96c04c9),
	.w4(32'h3a82c46c),
	.w5(32'hba3be009),
	.w6(32'hba8cb84e),
	.w7(32'hb9993f7e),
	.w8(32'hbabf6cf3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb475659),
	.w1(32'hbac1e505),
	.w2(32'h3a92cd67),
	.w3(32'hba7825cd),
	.w4(32'hbaa467bc),
	.w5(32'hb9d34e7f),
	.w6(32'h3b59bb4f),
	.w7(32'h3aaf5652),
	.w8(32'hb8805f8b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fdde9),
	.w1(32'h3a1ce40b),
	.w2(32'h3a378587),
	.w3(32'hbadae417),
	.w4(32'h3aa54670),
	.w5(32'h3b13fc80),
	.w6(32'hbb7395a5),
	.w7(32'h395a8fea),
	.w8(32'h3b92434b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93553fe),
	.w1(32'h3a3e4b64),
	.w2(32'hba75c9ae),
	.w3(32'hba9b0dcb),
	.w4(32'h399a0187),
	.w5(32'h39a098f7),
	.w6(32'hbb4eb277),
	.w7(32'hbb43562f),
	.w8(32'hba116c12),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dac6e),
	.w1(32'h3a594918),
	.w2(32'h3a14584f),
	.w3(32'hba9d8644),
	.w4(32'h39ad00bc),
	.w5(32'h393334c9),
	.w6(32'hbaddffbb),
	.w7(32'h39ee4a05),
	.w8(32'h3ae0b3c7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6c96b),
	.w1(32'hbb5c0b5a),
	.w2(32'hbb9cb94f),
	.w3(32'h3b121e47),
	.w4(32'hba95b80f),
	.w5(32'hbbd44862),
	.w6(32'h3b568ce6),
	.w7(32'h3bc5d131),
	.w8(32'h3ac58e3f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fa2d7),
	.w1(32'h396f39e8),
	.w2(32'hbb74cb64),
	.w3(32'hbbab9003),
	.w4(32'hbb363da0),
	.w5(32'hbb32639f),
	.w6(32'hb9c44264),
	.w7(32'hbb70d7dc),
	.w8(32'hbb8d307c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae887),
	.w1(32'h399f6bda),
	.w2(32'h3839f99c),
	.w3(32'hba62107e),
	.w4(32'h3a060aed),
	.w5(32'h3a030d1d),
	.w6(32'hba582bc6),
	.w7(32'h3a1533b9),
	.w8(32'h3afad581),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997c1ef),
	.w1(32'h394362dc),
	.w2(32'h39691aa7),
	.w3(32'h395aaa6e),
	.w4(32'h396135c8),
	.w5(32'h395f4380),
	.w6(32'h3923585f),
	.w7(32'h38ba8cef),
	.w8(32'h380ecd5a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab3389),
	.w1(32'h39807381),
	.w2(32'hba091d44),
	.w3(32'h37dd0bc6),
	.w4(32'hb7aae1f8),
	.w5(32'hba829cb9),
	.w6(32'h3904c637),
	.w7(32'hba44c3f6),
	.w8(32'hba3f921f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878252b),
	.w1(32'hb890e5ba),
	.w2(32'hb87909dc),
	.w3(32'hb87ec075),
	.w4(32'hb84729b1),
	.w5(32'hb7e0bb1a),
	.w6(32'h366fc9b3),
	.w7(32'hb6dff6ef),
	.w8(32'h3631e4fc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96689f5),
	.w1(32'hb8b87999),
	.w2(32'hb9b34aa7),
	.w3(32'hb9a15c85),
	.w4(32'hb9be1320),
	.w5(32'hb9a6f7c5),
	.w6(32'hb93a3e88),
	.w7(32'h37923abf),
	.w8(32'h37aa61c4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09dfa3),
	.w1(32'hb9b618e2),
	.w2(32'h397e4ebd),
	.w3(32'hbafbe503),
	.w4(32'h3988b1d3),
	.w5(32'h3974a021),
	.w6(32'hbb1656c7),
	.w7(32'hb8d0a8a5),
	.w8(32'h3ac83c0b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eb5e2),
	.w1(32'h3a151296),
	.w2(32'h3959a013),
	.w3(32'h39fd86ba),
	.w4(32'h3987e8b7),
	.w5(32'h391b7189),
	.w6(32'hb800a2b0),
	.w7(32'hb89251c2),
	.w8(32'h38c0f935),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951773d),
	.w1(32'h39425f5d),
	.w2(32'h3aa66f21),
	.w3(32'hb8506b11),
	.w4(32'hba62fe5f),
	.w5(32'h39ca5251),
	.w6(32'h3b967bc7),
	.w7(32'h3ab4c8e5),
	.w8(32'hba43a722),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e5a83),
	.w1(32'h3ac8d5c4),
	.w2(32'hba57197c),
	.w3(32'hba7f7b60),
	.w4(32'h396597d1),
	.w5(32'h3a275717),
	.w6(32'hbbb4ae13),
	.w7(32'h38bf3fe0),
	.w8(32'h3b6edcc2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d454d),
	.w1(32'h3805cada),
	.w2(32'h38143afc),
	.w3(32'hb5dce62b),
	.w4(32'h375abc54),
	.w5(32'h38216555),
	.w6(32'hb8412db7),
	.w7(32'h372e335a),
	.w8(32'h378dd567),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8946446),
	.w1(32'hb859260e),
	.w2(32'h3873e117),
	.w3(32'hb8eebf65),
	.w4(32'hb8d6a7f8),
	.w5(32'h370f7adc),
	.w6(32'hb7ac934e),
	.w7(32'hb846b3c7),
	.w8(32'h385c549f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c8232),
	.w1(32'hb81eb345),
	.w2(32'h3781422e),
	.w3(32'hb80f6d0c),
	.w4(32'hb8890238),
	.w5(32'hb7d01709),
	.w6(32'h37958927),
	.w7(32'hb828734f),
	.w8(32'hb803a301),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe1bf9),
	.w1(32'hb8ac2988),
	.w2(32'h398d08ec),
	.w3(32'hb9cdeabc),
	.w4(32'hb9709a0a),
	.w5(32'h392497e3),
	.w6(32'hb9c3aebc),
	.w7(32'hb8c05628),
	.w8(32'h399b8d7d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39979375),
	.w1(32'hbb9638d8),
	.w2(32'hba6dc597),
	.w3(32'h3be9775b),
	.w4(32'hb9d33cd6),
	.w5(32'hbbea5a2d),
	.w6(32'h3bbc8e92),
	.w7(32'h3b16bcd2),
	.w8(32'h3b6664e9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a249b),
	.w1(32'h3aba781d),
	.w2(32'h3aa31e73),
	.w3(32'hbb0bcca8),
	.w4(32'hbadb211f),
	.w5(32'hba964f93),
	.w6(32'h3beb57c3),
	.w7(32'h3b007e2b),
	.w8(32'hbb63039c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399df55a),
	.w1(32'hb839bf72),
	.w2(32'hb99d009f),
	.w3(32'h383eea3d),
	.w4(32'hba227230),
	.w5(32'hb9f653e2),
	.w6(32'h3ad036d4),
	.w7(32'h39781133),
	.w8(32'hba281f96),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c099c),
	.w1(32'hba4a408b),
	.w2(32'h39560f3f),
	.w3(32'h3a1ff5b1),
	.w4(32'hba6d0930),
	.w5(32'hbaecaf2b),
	.w6(32'h3b275937),
	.w7(32'h39cb0726),
	.w8(32'hba4b3ced),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d6353),
	.w1(32'hb9037bb4),
	.w2(32'hb9b170f8),
	.w3(32'hbac3bd30),
	.w4(32'h39bc4434),
	.w5(32'h398cec77),
	.w6(32'hba968ffa),
	.w7(32'h3a1be90d),
	.w8(32'h3a7fcfa7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995a48),
	.w1(32'h397d5a94),
	.w2(32'h3a8b0ef8),
	.w3(32'hba578446),
	.w4(32'hb918d7ca),
	.w5(32'hb8e67140),
	.w6(32'h3a5134e1),
	.w7(32'h36b97cdc),
	.w8(32'hba6a86e4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab802ea),
	.w1(32'h3b29be6e),
	.w2(32'h3a44937f),
	.w3(32'hbbc6ebd4),
	.w4(32'h3a85cc09),
	.w5(32'hba5e877b),
	.w6(32'hbb765ee8),
	.w7(32'h39f97283),
	.w8(32'hb9031524),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef39a3),
	.w1(32'hba4e099a),
	.w2(32'h3aeceb11),
	.w3(32'hbb22a594),
	.w4(32'hbab9640c),
	.w5(32'h392c9f4a),
	.w6(32'h3c32c8a2),
	.w7(32'h3b1c71c6),
	.w8(32'hbbb22282),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84c327),
	.w1(32'h3a6bcc83),
	.w2(32'hb7cbc73c),
	.w3(32'hba192743),
	.w4(32'h3a549838),
	.w5(32'h3a40a184),
	.w6(32'hbb3a45c9),
	.w7(32'h39827ee6),
	.w8(32'h3b0aeed2),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3a224),
	.w1(32'hb71e7580),
	.w2(32'hbae06c74),
	.w3(32'hb9e23f3e),
	.w4(32'hb9c064c4),
	.w5(32'h39ec1c0d),
	.w6(32'h3afaf744),
	.w7(32'h3a7aa9b1),
	.w8(32'hba540bc8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15afd0),
	.w1(32'hba0e7c01),
	.w2(32'h3a86e3cf),
	.w3(32'hbadcc0b4),
	.w4(32'h3addaa61),
	.w5(32'hbb25f52b),
	.w6(32'h3bec57f5),
	.w7(32'h3b0de9f9),
	.w8(32'hbb650d83),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399babf5),
	.w1(32'hba1d98fa),
	.w2(32'hbb3abcd3),
	.w3(32'h3a8d8c5a),
	.w4(32'hb87ac9cf),
	.w5(32'hbb4d37d5),
	.w6(32'h3a221031),
	.w7(32'h3b48d9d1),
	.w8(32'h3b16d86b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e8d4),
	.w1(32'h3a88bb82),
	.w2(32'h3a72e5a2),
	.w3(32'hba854c48),
	.w4(32'hb97ebe6a),
	.w5(32'h3a15ee2a),
	.w6(32'h3ba9422c),
	.w7(32'h399933eb),
	.w8(32'hbb43b861),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ffaf),
	.w1(32'hb8ac124f),
	.w2(32'h3916d36e),
	.w3(32'hb9f236f1),
	.w4(32'h36921f1c),
	.w5(32'h3980026c),
	.w6(32'hb93dd982),
	.w7(32'h39f21213),
	.w8(32'h3a5b3529),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb90aa),
	.w1(32'h3b029aca),
	.w2(32'hb9fe8e37),
	.w3(32'hbb10e649),
	.w4(32'h3ab79e1b),
	.w5(32'h3b4d6cef),
	.w6(32'hbc0a13f9),
	.w7(32'h39f8cc08),
	.w8(32'h3b575fe9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78285b0),
	.w1(32'hb8edd15a),
	.w2(32'h38877c51),
	.w3(32'h38fedc63),
	.w4(32'h39b6a6f9),
	.w5(32'hba836b85),
	.w6(32'h3ac8b7a0),
	.w7(32'h3a092c98),
	.w8(32'hba604563),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b25db),
	.w1(32'hb876b915),
	.w2(32'hb78071c1),
	.w3(32'h394ebdde),
	.w4(32'h38641fef),
	.w5(32'hb8f838f9),
	.w6(32'h390da589),
	.w7(32'hb6f4c1bf),
	.w8(32'hb7fd7898),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38044329),
	.w1(32'h37fe1e97),
	.w2(32'h3853e5e3),
	.w3(32'h384029c7),
	.w4(32'h3923cf6c),
	.w5(32'h38f458e1),
	.w6(32'hb855774d),
	.w7(32'h384fba3c),
	.w8(32'h3814ca12),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae79797),
	.w1(32'hba37c5b0),
	.w2(32'h399f4d61),
	.w3(32'h3a411d66),
	.w4(32'hbab765bf),
	.w5(32'hb987dbef),
	.w6(32'h3b08b384),
	.w7(32'h39d2f113),
	.w8(32'h3838287b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa59fb),
	.w1(32'hba044b69),
	.w2(32'h39e930eb),
	.w3(32'hb9193e66),
	.w4(32'hba4428bc),
	.w5(32'h3a585dfa),
	.w6(32'hba61a0ef),
	.w7(32'h3b543bb6),
	.w8(32'h3b8b46df),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7c063),
	.w1(32'hb9d4d366),
	.w2(32'h3960e45a),
	.w3(32'hba55770f),
	.w4(32'hb91fdb0b),
	.w5(32'hb9f8df76),
	.w6(32'h3b0c056e),
	.w7(32'h3b25e58e),
	.w8(32'h3ad377ed),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37731771),
	.w1(32'h38296835),
	.w2(32'h37488594),
	.w3(32'h3644ae15),
	.w4(32'h3783946c),
	.w5(32'h37cc81fd),
	.w6(32'hb63b841b),
	.w7(32'h34d425d9),
	.w8(32'hb7043371),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd9824),
	.w1(32'h3a21882f),
	.w2(32'h3a83f80b),
	.w3(32'hbb314c00),
	.w4(32'hbaaec6cc),
	.w5(32'h39911ce5),
	.w6(32'h3b6e4745),
	.w7(32'h3adaae54),
	.w8(32'hb7b5f318),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb020ce6),
	.w1(32'h386a45e4),
	.w2(32'h3a8f4b24),
	.w3(32'hbad568b5),
	.w4(32'h3a763361),
	.w5(32'h3b15c04b),
	.w6(32'hb7d3dced),
	.w7(32'h3b17ef9a),
	.w8(32'h3b68c910),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a683f1e),
	.w1(32'hb9c8f196),
	.w2(32'h3abafb1f),
	.w3(32'hba8efed8),
	.w4(32'hb99a9cf8),
	.w5(32'h3aa27175),
	.w6(32'h3c0b73f6),
	.w7(32'h3b0e2fad),
	.w8(32'hba3fdb5a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e4e5),
	.w1(32'hbb106da8),
	.w2(32'hbb46a98e),
	.w3(32'hbbcc07b5),
	.w4(32'h3aadfb75),
	.w5(32'h3b55dd7d),
	.w6(32'hbc1a7493),
	.w7(32'hbb0ff5de),
	.w8(32'h3b0737e0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9b31c),
	.w1(32'h3a1dfe29),
	.w2(32'hba3b996a),
	.w3(32'hb9014981),
	.w4(32'hba11a532),
	.w5(32'hbab1521d),
	.w6(32'hbacc39e0),
	.w7(32'hbaa426b6),
	.w8(32'hba6c0010),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a6838),
	.w1(32'hba6d3e17),
	.w2(32'hb9d93226),
	.w3(32'hbab842e4),
	.w4(32'hbaa07c2f),
	.w5(32'hb9fddf50),
	.w6(32'hba17c04b),
	.w7(32'hb99958fa),
	.w8(32'hb9950e16),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d789c),
	.w1(32'h39c96500),
	.w2(32'h394d9441),
	.w3(32'hba96c4b3),
	.w4(32'h3a0c26ca),
	.w5(32'h3a739d83),
	.w6(32'hba9f4da4),
	.w7(32'h3a4717f1),
	.w8(32'h3b1ef53c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11f6a1),
	.w1(32'h3ac56dbf),
	.w2(32'hba060f2e),
	.w3(32'hbb1648aa),
	.w4(32'h39b91214),
	.w5(32'h380901ac),
	.w6(32'hbb4f3128),
	.w7(32'h3a298e2d),
	.w8(32'h3ac8d91b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dca02),
	.w1(32'hba846c1e),
	.w2(32'hbabc02c6),
	.w3(32'hbaa54135),
	.w4(32'hba4cc1fa),
	.w5(32'hb9d2729c),
	.w6(32'hbb243d9b),
	.w7(32'hba4d2964),
	.w8(32'h3aa1137b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0247a1),
	.w1(32'hb9e68128),
	.w2(32'hb80257cd),
	.w3(32'hb9643a2f),
	.w4(32'hba2ad002),
	.w5(32'hb992028e),
	.w6(32'h3b0c4230),
	.w7(32'h3a1ba344),
	.w8(32'hb9be67ab),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c77fd),
	.w1(32'hb8c670d3),
	.w2(32'hb90d6292),
	.w3(32'h3815d404),
	.w4(32'hb96727f9),
	.w5(32'hb88d1547),
	.w6(32'hb89ad1d0),
	.w7(32'hb9708130),
	.w8(32'hb9e21efa),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74a16bb),
	.w1(32'hb994d6d6),
	.w2(32'hb882cc5b),
	.w3(32'h34742880),
	.w4(32'hba2270d4),
	.w5(32'hba930f05),
	.w6(32'h3ba7bf0a),
	.w7(32'h3aad3d42),
	.w8(32'hbb0a88b7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9756045),
	.w1(32'hb95fbffe),
	.w2(32'hb9bdf221),
	.w3(32'h39826b4d),
	.w4(32'hb902e0e7),
	.w5(32'h3a2056ec),
	.w6(32'h3a7328cc),
	.w7(32'h39d33111),
	.w8(32'h38cd8496),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38eb10),
	.w1(32'h3aa16305),
	.w2(32'h3ae16ae1),
	.w3(32'hba6ef17c),
	.w4(32'h3a90e617),
	.w5(32'h3afe9ef6),
	.w6(32'hbb13a6f7),
	.w7(32'h3ab9eff3),
	.w8(32'h3b6086a4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934a22e),
	.w1(32'hb903ecdf),
	.w2(32'h39c1ddf4),
	.w3(32'h38d27931),
	.w4(32'hb99a6f66),
	.w5(32'h39b6aa64),
	.w6(32'h390eb889),
	.w7(32'hb9575efb),
	.w8(32'h39ee6d76),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec789),
	.w1(32'hbb1535e3),
	.w2(32'h3a376126),
	.w3(32'hba9e45a6),
	.w4(32'hbb140b38),
	.w5(32'hb9e98648),
	.w6(32'h3a471f2f),
	.w7(32'h3ab2d81d),
	.w8(32'h3a34107f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38685442),
	.w1(32'hb894171d),
	.w2(32'hb63fc6a1),
	.w3(32'h37bdf123),
	.w4(32'hb787028d),
	.w5(32'h389d6c3b),
	.w6(32'hb8c458f2),
	.w7(32'hb8729b66),
	.w8(32'h37b0451f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c1654),
	.w1(32'h39c9641e),
	.w2(32'h39272810),
	.w3(32'hb89eeefb),
	.w4(32'hb78478b4),
	.w5(32'hb890c4ad),
	.w6(32'h392d0496),
	.w7(32'h3999a97e),
	.w8(32'h39bfd91c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8645cd),
	.w1(32'h39c9b45f),
	.w2(32'h3a2829db),
	.w3(32'h37a7626f),
	.w4(32'hb8d27413),
	.w5(32'h3a53db8a),
	.w6(32'hbb0fdbc7),
	.w7(32'hbab92776),
	.w8(32'h3a43e125),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad15053),
	.w1(32'hbbadca23),
	.w2(32'h3a55cce2),
	.w3(32'h3bd7773a),
	.w4(32'h39b84329),
	.w5(32'hbac4ee88),
	.w6(32'h3c1cd5cf),
	.w7(32'h3ba21927),
	.w8(32'h3b12f5de),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2f5ed),
	.w1(32'hb9d45016),
	.w2(32'h38ace5eb),
	.w3(32'hba7b58be),
	.w4(32'hba388d4a),
	.w5(32'h390bc396),
	.w6(32'hba2ee353),
	.w7(32'hba03a79c),
	.w8(32'h39493fe9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c6fa0),
	.w1(32'h39cdfc0c),
	.w2(32'h3a0f6d0b),
	.w3(32'hbaabbbf6),
	.w4(32'h3a213b4f),
	.w5(32'h3ad26ab1),
	.w6(32'hbb7a1549),
	.w7(32'hba0f1b22),
	.w8(32'h3b52f7b3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba137d22),
	.w1(32'h3a1cfb67),
	.w2(32'h3a42f5c0),
	.w3(32'hbaafd5ad),
	.w4(32'h39e6058e),
	.w5(32'h3b0ee0e9),
	.w6(32'hbae6fc2c),
	.w7(32'hba9fb5f8),
	.w8(32'hba7b766e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d7ced),
	.w1(32'h3a931e8a),
	.w2(32'h3ac838d1),
	.w3(32'hbb99e255),
	.w4(32'hb8f9ba15),
	.w5(32'h3aa1fd8a),
	.w6(32'h39949b70),
	.w7(32'h3ac1c2b6),
	.w8(32'hbaf9fd18),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dc261),
	.w1(32'h3a16c12a),
	.w2(32'h3a248676),
	.w3(32'hba756ede),
	.w4(32'hba58d3a1),
	.w5(32'h39dfbd2f),
	.w6(32'h3b47e635),
	.w7(32'h3a242055),
	.w8(32'h39ed15b6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf986e1),
	.w1(32'hba9d0c59),
	.w2(32'h3a9837fd),
	.w3(32'hbb38d866),
	.w4(32'hbb1a55cd),
	.w5(32'hbad6e78d),
	.w6(32'h3b899d88),
	.w7(32'h3a0e4d97),
	.w8(32'hbb279bfa),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2d60e),
	.w1(32'hb996b54f),
	.w2(32'hb724c840),
	.w3(32'hb9be821a),
	.w4(32'hba156874),
	.w5(32'hb9fd7c7d),
	.w6(32'hba09c9a6),
	.w7(32'hba73734b),
	.w8(32'hb9c50085),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ca94f),
	.w1(32'h3a86284b),
	.w2(32'hbab165d2),
	.w3(32'hbb4403b4),
	.w4(32'hb9bac462),
	.w5(32'hbaaf263e),
	.w6(32'hb9ebfda7),
	.w7(32'hbb07e5ac),
	.w8(32'hbb43e9d4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4028375),
	.w1(32'hb7c8ae19),
	.w2(32'hb876ddea),
	.w3(32'h36f3ac86),
	.w4(32'hb798b640),
	.w5(32'hb7ed49fd),
	.w6(32'hb810a0e8),
	.w7(32'hb84262bd),
	.w8(32'hb80cdd75),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c07dd2),
	.w1(32'hb8b46728),
	.w2(32'hba0f047d),
	.w3(32'hba064910),
	.w4(32'hb9b9cd42),
	.w5(32'hb8fd13b7),
	.w6(32'h3a5896cb),
	.w7(32'h3a9a1808),
	.w8(32'h3a359934),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b7608),
	.w1(32'h3a37f8ad),
	.w2(32'hb9af2f90),
	.w3(32'hb976fbf4),
	.w4(32'h38bfe3cb),
	.w5(32'hb9bc2566),
	.w6(32'hba2b0c66),
	.w7(32'hb91baa87),
	.w8(32'h39a18db1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83a522),
	.w1(32'h3ab6514b),
	.w2(32'hba97eeca),
	.w3(32'hbb8654ed),
	.w4(32'hbaafa848),
	.w5(32'hba269efb),
	.w6(32'hba3e3392),
	.w7(32'hbaa222fe),
	.w8(32'hbb028f48),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37346758),
	.w1(32'hb6e9cb99),
	.w2(32'hb6fa6e4a),
	.w3(32'hb751aa2a),
	.w4(32'hb70f7a9c),
	.w5(32'hb7d2790c),
	.w6(32'hb84752ae),
	.w7(32'hb770bf10),
	.w8(32'hb75575d1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924dd7d),
	.w1(32'h391a2106),
	.w2(32'h3808d884),
	.w3(32'h38cf2dec),
	.w4(32'h37b4d08d),
	.w5(32'h3616503c),
	.w6(32'h381aed1b),
	.w7(32'h384ac2f3),
	.w8(32'h38cae21c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ace053),
	.w1(32'h3a723250),
	.w2(32'hb9cdfc1d),
	.w3(32'hba9cff3d),
	.w4(32'h3a4be7d9),
	.w5(32'hba2f75cb),
	.w6(32'hba03b370),
	.w7(32'h39b9b002),
	.w8(32'h3a2534f0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba54c),
	.w1(32'hbb91c880),
	.w2(32'hbb4b88fd),
	.w3(32'hbb60a6bd),
	.w4(32'hbb8a8066),
	.w5(32'hbaa3d6be),
	.w6(32'h3a8bcf17),
	.w7(32'hbbaa6e75),
	.w8(32'hbb57d0d4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc5847),
	.w1(32'hbb8c6625),
	.w2(32'h3bae1e84),
	.w3(32'h3b961b66),
	.w4(32'h3a726f61),
	.w5(32'h3b784805),
	.w6(32'h3c266c4b),
	.w7(32'h3b315840),
	.w8(32'h3b49e4cc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d1081),
	.w1(32'h382cdccc),
	.w2(32'h3966b8b1),
	.w3(32'hb9e14900),
	.w4(32'h36a91b8d),
	.w5(32'h396e5c22),
	.w6(32'hb90637e3),
	.w7(32'h393633d4),
	.w8(32'h37e57618),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cf274),
	.w1(32'hb9379a6d),
	.w2(32'h3b61b228),
	.w3(32'h3ac6f3ed),
	.w4(32'h3963f0be),
	.w5(32'hbaa1d345),
	.w6(32'h3c1212f8),
	.w7(32'h3b9b2654),
	.w8(32'hbafbcd29),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0734c8),
	.w1(32'hba0aded8),
	.w2(32'hbab0a4b4),
	.w3(32'hbc46415a),
	.w4(32'hba07f5e7),
	.w5(32'h3b0d18d1),
	.w6(32'hbbb04b29),
	.w7(32'hbb7ac06e),
	.w8(32'h3a5cd175),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1807b),
	.w1(32'h398ad13d),
	.w2(32'hb746a380),
	.w3(32'h3adad641),
	.w4(32'h3a10b8d6),
	.w5(32'h3adde571),
	.w6(32'h3b7169b3),
	.w7(32'h3ae4feb1),
	.w8(32'h37a94192),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382bfa01),
	.w1(32'hb768f31f),
	.w2(32'hb7362cd1),
	.w3(32'h37a09d95),
	.w4(32'hb817b227),
	.w5(32'h378599e3),
	.w6(32'h37cbf876),
	.w7(32'h36b69da4),
	.w8(32'hb7e9be17),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915b354),
	.w1(32'hb8a98b5f),
	.w2(32'h396e5f7d),
	.w3(32'h39499400),
	.w4(32'hb8a932d9),
	.w5(32'h395a9db0),
	.w6(32'h399232f0),
	.w7(32'hb81c1402),
	.w8(32'h391e7453),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57d701e),
	.w1(32'h36376483),
	.w2(32'h37100818),
	.w3(32'hb6c5fe58),
	.w4(32'hb77b4762),
	.w5(32'hb8452948),
	.w6(32'h37953e9a),
	.w7(32'hb7213f11),
	.w8(32'hb808645d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa136ec),
	.w1(32'hbaa0a05e),
	.w2(32'h3b00a834),
	.w3(32'h3b2e150f),
	.w4(32'h39a0e017),
	.w5(32'h3a1e88e5),
	.w6(32'h3ba8aa7e),
	.w7(32'h3b2a6f86),
	.w8(32'hb8b157e7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0693c7),
	.w1(32'hb96d8818),
	.w2(32'h39f6c7eb),
	.w3(32'h3a41c67c),
	.w4(32'hb8387c27),
	.w5(32'hba87d527),
	.w6(32'h3a96aad5),
	.w7(32'h3a7cb37a),
	.w8(32'hb7cde211),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8008),
	.w1(32'h3aa81f6c),
	.w2(32'h3a577ba1),
	.w3(32'hbac6c3b5),
	.w4(32'h3a020a44),
	.w5(32'h394ade7a),
	.w6(32'hbb954e5e),
	.w7(32'h3a7362ae),
	.w8(32'h3b426972),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b7c8a8),
	.w1(32'h3999a804),
	.w2(32'hb959dac5),
	.w3(32'h3910fcab),
	.w4(32'h39beec4c),
	.w5(32'hb9b49837),
	.w6(32'hba1046f1),
	.w7(32'h39e6851b),
	.w8(32'h3a01fe05),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127cde),
	.w1(32'hb99b9bbb),
	.w2(32'h3b177011),
	.w3(32'hb8ee6f78),
	.w4(32'h3946a487),
	.w5(32'h3aad3ca4),
	.w6(32'h3baa6fab),
	.w7(32'h3b458785),
	.w8(32'h3ae16c0f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a166b0a),
	.w1(32'hba8ae0fc),
	.w2(32'h3a05915e),
	.w3(32'h3ac3f64c),
	.w4(32'hbadc757d),
	.w5(32'h392ebdd6),
	.w6(32'h3ac4db90),
	.w7(32'hba67fe4d),
	.w8(32'h39352c57),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ca16ea),
	.w1(32'hb7c511c2),
	.w2(32'hb88ecf3c),
	.w3(32'hb6f7bbcb),
	.w4(32'hb7a80cc5),
	.w5(32'hb81a580f),
	.w6(32'hb84f52e0),
	.w7(32'hb8530022),
	.w8(32'hb88286bb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5963bc),
	.w1(32'hba7a51eb),
	.w2(32'hba5305bd),
	.w3(32'h3a99ebe1),
	.w4(32'hbac1f49d),
	.w5(32'hbb202d2b),
	.w6(32'h3b2fa978),
	.w7(32'h3a230062),
	.w8(32'hbb089db0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57babc9),
	.w1(32'h369205d9),
	.w2(32'hb8daebae),
	.w3(32'hb7e5cef9),
	.w4(32'h3771c676),
	.w5(32'hb891f279),
	.w6(32'hb8e77e7e),
	.w7(32'hb84e8aff),
	.w8(32'hb904c138),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0e26),
	.w1(32'hba98cd19),
	.w2(32'hb74a8686),
	.w3(32'hbaab0d0b),
	.w4(32'hbaa91617),
	.w5(32'hba5ef777),
	.w6(32'h3a9b656b),
	.w7(32'h3a343382),
	.w8(32'h38ac5adf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39787877),
	.w1(32'h3a3c523f),
	.w2(32'hb9f31bf6),
	.w3(32'hbb2f7404),
	.w4(32'hba039b3f),
	.w5(32'hb76d7078),
	.w6(32'hbb96e95a),
	.w7(32'hba3b5775),
	.w8(32'h3b0c14c8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19ee8f),
	.w1(32'h3a4670b9),
	.w2(32'h3ab50969),
	.w3(32'hbab5c5bb),
	.w4(32'h3a287b10),
	.w5(32'h3aafa089),
	.w6(32'hba9f83a6),
	.w7(32'h3afb5fd6),
	.w8(32'h3b6ca504),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9862128),
	.w1(32'hb9a7c88e),
	.w2(32'hb9d5a485),
	.w3(32'hb9988539),
	.w4(32'hb9e45110),
	.w5(32'hb9c982a3),
	.w6(32'hb921d8e0),
	.w7(32'hb942f304),
	.w8(32'hb8d74805),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949fcd8),
	.w1(32'h3b2bb222),
	.w2(32'h3afb22b8),
	.w3(32'hbb97ec75),
	.w4(32'h3af0108f),
	.w5(32'h3acd9273),
	.w6(32'hbb93bb1e),
	.w7(32'hb98f7647),
	.w8(32'h3b53c676),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a338131),
	.w1(32'h3ad8ca9c),
	.w2(32'h3aafb5bf),
	.w3(32'hb938451d),
	.w4(32'hb9c89c06),
	.w5(32'h3a326644),
	.w6(32'h3b71bc83),
	.w7(32'h3a6a6c0e),
	.w8(32'hb96cfc56),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb071030),
	.w1(32'h38e64b72),
	.w2(32'h3aa28463),
	.w3(32'hbaf7321f),
	.w4(32'h39c5c847),
	.w5(32'h3a4a2321),
	.w6(32'h3a638883),
	.w7(32'h3b5bea6e),
	.w8(32'h3b46cedf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a3dc69),
	.w1(32'h37cde17e),
	.w2(32'hb6dcf231),
	.w3(32'hb6e43750),
	.w4(32'hb79e060a),
	.w5(32'hb721f4b1),
	.w6(32'h38672e49),
	.w7(32'h37bc96ca),
	.w8(32'hb8abcd83),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9245466),
	.w1(32'hb8a5b44b),
	.w2(32'h3892e84e),
	.w3(32'h380d39fb),
	.w4(32'h39b09268),
	.w5(32'h39af7376),
	.w6(32'hb91b96b1),
	.w7(32'hb8697380),
	.w8(32'h37fb187e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b728),
	.w1(32'hbba74ebf),
	.w2(32'hbb0002dd),
	.w3(32'h3bd06e93),
	.w4(32'hb6b830ac),
	.w5(32'hbb026f64),
	.w6(32'h3bd6c6f3),
	.w7(32'h3acc9dc6),
	.w8(32'h3a8ae3bf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67650),
	.w1(32'hbb599c93),
	.w2(32'h39b7b713),
	.w3(32'h3b61b25c),
	.w4(32'hba7be1dd),
	.w5(32'hba8fd9ae),
	.w6(32'h3b3cfbf1),
	.w7(32'hb92a224c),
	.w8(32'hbafa2b17),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2bf5a),
	.w1(32'h3a5d6ac6),
	.w2(32'h3a5d1573),
	.w3(32'hbad687fd),
	.w4(32'h3acbd484),
	.w5(32'hba0334a5),
	.w6(32'hbb03ca1d),
	.w7(32'h3a743fd5),
	.w8(32'h3b1476c2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaecf64),
	.w1(32'hbb0da9a6),
	.w2(32'hbb7fe405),
	.w3(32'hbbdabbb7),
	.w4(32'h39584973),
	.w5(32'h3b3f6772),
	.w6(32'h3bc7e5db),
	.w7(32'hbb052377),
	.w8(32'hbbec6d68),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c3b1f),
	.w1(32'h39c8851c),
	.w2(32'hb8553dc2),
	.w3(32'h393f3877),
	.w4(32'h38916619),
	.w5(32'hb9970638),
	.w6(32'h3a78ceae),
	.w7(32'h3a2381f5),
	.w8(32'hba8839d2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62bda5),
	.w1(32'hba086952),
	.w2(32'hba171c0b),
	.w3(32'h3ac974f3),
	.w4(32'hb945e347),
	.w5(32'hba9e20db),
	.w6(32'h3a389fc7),
	.w7(32'hb9cc3946),
	.w8(32'hba84e457),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa70b0),
	.w1(32'hbbddd2f0),
	.w2(32'h3b03a756),
	.w3(32'h3c486657),
	.w4(32'hbaa150e9),
	.w5(32'hbae6685e),
	.w6(32'h3c8086d5),
	.w7(32'h3c343883),
	.w8(32'h3b95f109),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b1cc),
	.w1(32'h3a87d90d),
	.w2(32'h3b4829e7),
	.w3(32'h3b0f1706),
	.w4(32'h385a9e6a),
	.w5(32'hbaf03921),
	.w6(32'h3c1611dc),
	.w7(32'h3b9a659d),
	.w8(32'hbb320ead),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2be2d6),
	.w1(32'hbb69fd2b),
	.w2(32'h3b12fade),
	.w3(32'h3ba95663),
	.w4(32'h3995e4b7),
	.w5(32'hba56ea5e),
	.w6(32'h3c4727ff),
	.w7(32'h3bb3a417),
	.w8(32'h3aabc137),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababb83),
	.w1(32'hb887d9f7),
	.w2(32'hbaf3427d),
	.w3(32'hbaa10402),
	.w4(32'h3954fb86),
	.w5(32'h39b6a5fe),
	.w6(32'hbb3f86bd),
	.w7(32'h3a1098aa),
	.w8(32'h3b483363),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a583e8),
	.w1(32'h3aa42de0),
	.w2(32'hba91f253),
	.w3(32'hbb4a239d),
	.w4(32'h39e185c7),
	.w5(32'h3a5b8985),
	.w6(32'hbbc21bf5),
	.w7(32'hba748b84),
	.w8(32'h3b6a050d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f7b515),
	.w1(32'hb7ba6f0a),
	.w2(32'hb81cafa0),
	.w3(32'hb7a902ed),
	.w4(32'hb7b4303a),
	.w5(32'hb75ee08f),
	.w6(32'hb8144ace),
	.w7(32'hb7bba5bc),
	.w8(32'hb83b057f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bea411),
	.w1(32'h37e8cee6),
	.w2(32'hb6e25d84),
	.w3(32'h37c7e965),
	.w4(32'h36822b27),
	.w5(32'hb7b3b1fc),
	.w6(32'hb807e5a6),
	.w7(32'hb84aa2e2),
	.w8(32'hb7f7457f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e264f),
	.w1(32'hba2c7ea3),
	.w2(32'hba218b04),
	.w3(32'hb9e0a032),
	.w4(32'hbabdebb7),
	.w5(32'hbaa21bf0),
	.w6(32'h3a9a84a8),
	.w7(32'h3a898427),
	.w8(32'h3aa61ecc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3630bead),
	.w1(32'hb810550b),
	.w2(32'hb8835683),
	.w3(32'hb6c72996),
	.w4(32'hb7b7403b),
	.w5(32'h3b16fd80),
	.w6(32'hb7072397),
	.w7(32'hb802c127),
	.w8(32'h3aed4cac),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b356bd6),
	.w1(32'h3adfd524),
	.w2(32'h3a9fde1f),
	.w3(32'h3b9fc132),
	.w4(32'h38a93e22),
	.w5(32'h3aee5ae3),
	.w6(32'h3b8df0c2),
	.w7(32'h397866b9),
	.w8(32'hb9940b2f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a48e8),
	.w1(32'hba90bd4e),
	.w2(32'h3ac1ee92),
	.w3(32'h3bc88628),
	.w4(32'h3b23ca80),
	.w5(32'hbbb0a90b),
	.w6(32'h3b3bed9f),
	.w7(32'hba7b1475),
	.w8(32'hbb9a45ca),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4fff3),
	.w1(32'hbb3d60af),
	.w2(32'hbb29120f),
	.w3(32'hbb2c240b),
	.w4(32'hbb922a8e),
	.w5(32'hbb7f9fb6),
	.w6(32'hb989d76f),
	.w7(32'hbb022e2d),
	.w8(32'h3a4f4cbe),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0d7c3),
	.w1(32'h3b4e896e),
	.w2(32'h3b566a2e),
	.w3(32'hbbb46a62),
	.w4(32'hbba90929),
	.w5(32'hb98dbf3f),
	.w6(32'h3a464d35),
	.w7(32'hbb2fb812),
	.w8(32'hb989cf0a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068f56),
	.w1(32'hbc0ff4d6),
	.w2(32'h3b147559),
	.w3(32'h3b760b49),
	.w4(32'hbae51595),
	.w5(32'hbb8419fb),
	.w6(32'h3caa1e27),
	.w7(32'h3befc387),
	.w8(32'hbadd315f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb681862),
	.w1(32'hba9b0aaa),
	.w2(32'hb9731b11),
	.w3(32'hbb655d46),
	.w4(32'hbb132b2a),
	.w5(32'h3a02891a),
	.w6(32'h3a8a2cee),
	.w7(32'h3ad6d020),
	.w8(32'hbb39bce7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126500),
	.w1(32'hbabdfdf8),
	.w2(32'hbbb8dc90),
	.w3(32'hbb2d728b),
	.w4(32'hbbab072d),
	.w5(32'h3b8e3a5e),
	.w6(32'hbb94a99e),
	.w7(32'hbbe84814),
	.w8(32'h3b4b7d0f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07871a),
	.w1(32'hba5d96dc),
	.w2(32'h39360a25),
	.w3(32'h3ba2239b),
	.w4(32'h3b2a1685),
	.w5(32'hbb171808),
	.w6(32'h3be87fa1),
	.w7(32'h3b63200c),
	.w8(32'hba5cbb8f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5b4b1),
	.w1(32'h3ba1dd96),
	.w2(32'h3a3ba233),
	.w3(32'hbb25b9d4),
	.w4(32'hb8e3edc3),
	.w5(32'hbae7f53d),
	.w6(32'h392d87d0),
	.w7(32'hba83b5b0),
	.w8(32'hbac296ae),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79085),
	.w1(32'hbb9bb503),
	.w2(32'h3ad36890),
	.w3(32'hb9cc8785),
	.w4(32'hba004e8d),
	.w5(32'h3b0f528d),
	.w6(32'h3a1200f5),
	.w7(32'hba2b842f),
	.w8(32'hb990967f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cb791),
	.w1(32'hb916f9d0),
	.w2(32'hbb60ccaa),
	.w3(32'h3b345951),
	.w4(32'hbadfb399),
	.w5(32'hbb45fc4b),
	.w6(32'hba0afe87),
	.w7(32'hbb59dcc9),
	.w8(32'h3b083ea3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ae5f8),
	.w1(32'h3be52cd2),
	.w2(32'h3b9ba0b6),
	.w3(32'h3b304fc2),
	.w4(32'h3b080a91),
	.w5(32'h3b8585cd),
	.w6(32'h3c016bed),
	.w7(32'h3bdadc47),
	.w8(32'h3bd24e28),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c324748),
	.w1(32'h3b9c5cff),
	.w2(32'h3bfb5e56),
	.w3(32'h3b6a670a),
	.w4(32'h3ba2e4b6),
	.w5(32'hb9b24215),
	.w6(32'h3b16305f),
	.w7(32'h3ba294bb),
	.w8(32'h3b8ec2c8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d58b1),
	.w1(32'h3b30ab5c),
	.w2(32'hbb266a12),
	.w3(32'hbb661540),
	.w4(32'h3b88b9fc),
	.w5(32'h3c0c027b),
	.w6(32'h3c2a9162),
	.w7(32'hbac04279),
	.w8(32'h3af3664f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6780),
	.w1(32'h3ba9e03b),
	.w2(32'h395e5271),
	.w3(32'h3b344eeb),
	.w4(32'h3b3fc936),
	.w5(32'hbb1ccacd),
	.w6(32'h3bde314e),
	.w7(32'h398660d3),
	.w8(32'hbbc0f664),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4841),
	.w1(32'hbb6dedce),
	.w2(32'hba93e252),
	.w3(32'hbb406371),
	.w4(32'hba20edd4),
	.w5(32'h3a347156),
	.w6(32'h390a12b7),
	.w7(32'h38836797),
	.w8(32'hbb826ebf),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb634d32),
	.w1(32'hbbd283b0),
	.w2(32'hbbef5803),
	.w3(32'hba83d2d9),
	.w4(32'hbb66622a),
	.w5(32'hbb3f198d),
	.w6(32'hbb68ce1c),
	.w7(32'hbbf79746),
	.w8(32'h3a8f3c9c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40e402),
	.w1(32'h3b2a3fec),
	.w2(32'hbb001ba6),
	.w3(32'hb9c42609),
	.w4(32'h3a464940),
	.w5(32'h3ac96deb),
	.w6(32'h3bf640af),
	.w7(32'h3911509d),
	.w8(32'hb9c8a60f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39453bd7),
	.w1(32'hba49e675),
	.w2(32'h3a95cc84),
	.w3(32'h3ba347f4),
	.w4(32'h3b42ac08),
	.w5(32'h3b95ddce),
	.w6(32'h3abbfe56),
	.w7(32'h3b996c8e),
	.w8(32'hb9a54e7f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6193b4),
	.w1(32'hbb7ef770),
	.w2(32'hbba08bd6),
	.w3(32'hb9985cc0),
	.w4(32'hbb213db9),
	.w5(32'h3ae60dd6),
	.w6(32'hbb96faf7),
	.w7(32'hbbce62d1),
	.w8(32'hba1a424b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82fe71),
	.w1(32'h3b3d47de),
	.w2(32'h3a10fb25),
	.w3(32'hbae361c6),
	.w4(32'hbb521faf),
	.w5(32'hbbf63c0f),
	.w6(32'h3ae0e7fb),
	.w7(32'hbad7aa62),
	.w8(32'hbc054375),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa0d0),
	.w1(32'hbb481ff8),
	.w2(32'hbbd63749),
	.w3(32'hbb9dfb44),
	.w4(32'hbbf86292),
	.w5(32'hbb83d56d),
	.w6(32'hbb6ebb68),
	.w7(32'hbbc77d31),
	.w8(32'h39d70dac),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951cc9b),
	.w1(32'h3b28f8a9),
	.w2(32'hbb14350e),
	.w3(32'hba7784a6),
	.w4(32'h3b33b9d7),
	.w5(32'h3b03fedf),
	.w6(32'h3bba0ae0),
	.w7(32'h3b2b29b4),
	.w8(32'hbb4fe11b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b48a4),
	.w1(32'h39d2e235),
	.w2(32'hbb568c12),
	.w3(32'hbadad51a),
	.w4(32'h38c7e493),
	.w5(32'h3aff3772),
	.w6(32'hbaf89786),
	.w7(32'hbb7a75f6),
	.w8(32'h3b560259),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ecdeb),
	.w1(32'h3afcdbad),
	.w2(32'h38a1f39b),
	.w3(32'hba7dd64e),
	.w4(32'h3b9c0a0a),
	.w5(32'h3bc9a29c),
	.w6(32'h3c31cc77),
	.w7(32'hbac10eb6),
	.w8(32'h3a4ae760),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244742),
	.w1(32'hbae3eae6),
	.w2(32'hbb12a8cb),
	.w3(32'h3ba8770e),
	.w4(32'h3b8a1a31),
	.w5(32'h3b6a9aec),
	.w6(32'hbad8e27b),
	.w7(32'hbaa3d455),
	.w8(32'h3b137e0a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2434ce),
	.w1(32'h3af6b6b4),
	.w2(32'h3b29084f),
	.w3(32'h3b516af1),
	.w4(32'h3bc1cfb9),
	.w5(32'hbb707bac),
	.w6(32'h3c00cb9b),
	.w7(32'h3ac2d949),
	.w8(32'hbb4016d5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d032a1),
	.w1(32'h3b10c0d9),
	.w2(32'hbac4b317),
	.w3(32'hbc2e8393),
	.w4(32'hb8e02720),
	.w5(32'hba888dc9),
	.w6(32'hbb9bb2c4),
	.w7(32'hbb8cf801),
	.w8(32'hbc449694),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fef52),
	.w1(32'hbb072207),
	.w2(32'h399800a6),
	.w3(32'hb8e3f0f7),
	.w4(32'hb9b02428),
	.w5(32'hbaf01dbd),
	.w6(32'h3b3f683c),
	.w7(32'h3b366017),
	.w8(32'hbb34372f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80473cb),
	.w1(32'hbab5ec78),
	.w2(32'hbb25d2a6),
	.w3(32'h3b79aea3),
	.w4(32'hbb0dcd69),
	.w5(32'hbab07dcd),
	.w6(32'hbb713bd8),
	.w7(32'hbb7d9b63),
	.w8(32'h3b1bbc62),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule