module layer_8_featuremap_240(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb019e5),
	.w1(32'hbb4d170c),
	.w2(32'hbbc7f2c1),
	.w3(32'h3a9af40a),
	.w4(32'hbb9d0236),
	.w5(32'hbc0c7e3b),
	.w6(32'h3b00f54c),
	.w7(32'hbabb295f),
	.w8(32'h3b78135d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8d5f9),
	.w1(32'hbabdc734),
	.w2(32'hbafeacf3),
	.w3(32'hbbf6f061),
	.w4(32'hbaf0f23a),
	.w5(32'hba71d0fe),
	.w6(32'h3bde9e88),
	.w7(32'h3b138935),
	.w8(32'hb9df5f96),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba351f43),
	.w1(32'h3b6e01e1),
	.w2(32'hbc1c8d4d),
	.w3(32'h3b0793dd),
	.w4(32'hbbf2b42c),
	.w5(32'hbc008aa7),
	.w6(32'h3c859c74),
	.w7(32'h3b2ad538),
	.w8(32'hbc5d78d5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fccd1),
	.w1(32'hbb500c91),
	.w2(32'hbc5c451a),
	.w3(32'hbb844971),
	.w4(32'hbc28cc8e),
	.w5(32'hbc61134e),
	.w6(32'h3c126be6),
	.w7(32'h383b9b06),
	.w8(32'hbc126f1f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc841443),
	.w1(32'hbb8d32b2),
	.w2(32'hbb841162),
	.w3(32'h3bed0e78),
	.w4(32'hb9237e04),
	.w5(32'hbb25a301),
	.w6(32'h3b97a4a6),
	.w7(32'h3afcaae3),
	.w8(32'hb8960081),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e702c),
	.w1(32'h3c84988e),
	.w2(32'h3ba46532),
	.w3(32'hb9b9b74d),
	.w4(32'h3c517b78),
	.w5(32'h3a7e5bea),
	.w6(32'hba9ac961),
	.w7(32'h3ab422b3),
	.w8(32'hbbabb664),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b997b13),
	.w1(32'h3aa16d02),
	.w2(32'h3b80c205),
	.w3(32'h3b1b6155),
	.w4(32'h3b1ed9d8),
	.w5(32'h3ab6c678),
	.w6(32'h3a125733),
	.w7(32'h3b503dba),
	.w8(32'h3ac5a2fb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa876d4),
	.w1(32'hbc74f246),
	.w2(32'hbb7f96f1),
	.w3(32'hb99c3be3),
	.w4(32'hbc8c0ff4),
	.w5(32'hbb589ffd),
	.w6(32'hbc8563cb),
	.w7(32'hbc566e6d),
	.w8(32'hbb690119),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6756be),
	.w1(32'hbc7dd731),
	.w2(32'hbb3d674f),
	.w3(32'hbb2c1f79),
	.w4(32'hbc5f9f22),
	.w5(32'hbbd2cb28),
	.w6(32'hbc14f0a8),
	.w7(32'hba14266e),
	.w8(32'hbb29e638),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7a41),
	.w1(32'hbc5b76d0),
	.w2(32'hbc596928),
	.w3(32'hbbdbb7d8),
	.w4(32'hbc4109fe),
	.w5(32'hbc204c82),
	.w6(32'h3aea768b),
	.w7(32'hbc2478ff),
	.w8(32'hbaa05a84),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b872ddc),
	.w1(32'h3a2b191b),
	.w2(32'h3a255fa0),
	.w3(32'h3c0ad6ea),
	.w4(32'h3a119fc2),
	.w5(32'hbb8bc83d),
	.w6(32'h3b0092be),
	.w7(32'h3b3057bd),
	.w8(32'h3bc66e2e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d118b),
	.w1(32'hbaed8dec),
	.w2(32'h39f81eb9),
	.w3(32'hba63fe89),
	.w4(32'h3b29cc23),
	.w5(32'hb90c946a),
	.w6(32'h3b3907e4),
	.w7(32'h3be850b1),
	.w8(32'h3c0a3a69),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c567fed),
	.w1(32'h3b21db10),
	.w2(32'h3b026e8d),
	.w3(32'h3c47b9d6),
	.w4(32'h3b96d420),
	.w5(32'h3a2a64ef),
	.w6(32'h3be2defc),
	.w7(32'h3ba50c66),
	.w8(32'h3b91f3d3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c56c6),
	.w1(32'hbcc78f30),
	.w2(32'hbd2f68e7),
	.w3(32'h3c000c06),
	.w4(32'hbc9296e2),
	.w5(32'hbcb2f0e7),
	.w6(32'hbb505e40),
	.w7(32'hbc55804a),
	.w8(32'hbcb60a79),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca348cf),
	.w1(32'hbba35e4e),
	.w2(32'h3b16d643),
	.w3(32'hbb2ebffe),
	.w4(32'hbb2efa29),
	.w5(32'h3b79af6f),
	.w6(32'hbc00b26b),
	.w7(32'h3a399349),
	.w8(32'hbaba804c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e1b5),
	.w1(32'hbbcab194),
	.w2(32'hba02628c),
	.w3(32'h3b049d59),
	.w4(32'hbc064fca),
	.w5(32'h3b2cc1b8),
	.w6(32'hbb4a6aa0),
	.w7(32'h3c09b7b1),
	.w8(32'h3a60feba),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24e14c),
	.w1(32'h3b1831d9),
	.w2(32'h3b9099ad),
	.w3(32'h3bd8ab6f),
	.w4(32'h3b852f48),
	.w5(32'hba346dac),
	.w6(32'hbba7c0a0),
	.w7(32'hbb5a243e),
	.w8(32'h3bff2c12),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093e72),
	.w1(32'hbd02bd5f),
	.w2(32'hbd5b875e),
	.w3(32'hbb4c54bc),
	.w4(32'hbd0cd57c),
	.w5(32'hbd35dfd9),
	.w6(32'hbc280de4),
	.w7(32'hbcc403ec),
	.w8(32'hbd062c58),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2beda8),
	.w1(32'hbc8d1786),
	.w2(32'h3af9a358),
	.w3(32'hbcb1ee09),
	.w4(32'hbcb54e39),
	.w5(32'hbbbd4215),
	.w6(32'h3bd0abe3),
	.w7(32'h3ae7f6c2),
	.w8(32'h3b9ebb13),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96759f),
	.w1(32'hbc105134),
	.w2(32'hbbd98def),
	.w3(32'h3bb203ff),
	.w4(32'hbbac22e5),
	.w5(32'hbbbedb25),
	.w6(32'hbbb76e5d),
	.w7(32'hbb74b727),
	.w8(32'hbbe518a9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ac47b),
	.w1(32'hbaf9d0e4),
	.w2(32'hbc27cf60),
	.w3(32'h3b595f4e),
	.w4(32'h3b96481c),
	.w5(32'hbc034cf5),
	.w6(32'h3b675f2c),
	.w7(32'h3bf81e56),
	.w8(32'hbab48217),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3b33),
	.w1(32'h3cb76317),
	.w2(32'h3d2a3c69),
	.w3(32'hbbac2668),
	.w4(32'h3ccbec8a),
	.w5(32'h3c942b04),
	.w6(32'h3c4a877e),
	.w7(32'h3cd3c187),
	.w8(32'h3c7ef4bd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17abf9),
	.w1(32'h3c399f2d),
	.w2(32'h3c761f16),
	.w3(32'h3c9057b6),
	.w4(32'hbba0607a),
	.w5(32'hb9000be2),
	.w6(32'h3c0a9863),
	.w7(32'h3c1f7024),
	.w8(32'h3c3e1332),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c697528),
	.w1(32'h3ca6209a),
	.w2(32'h3cd59f6a),
	.w3(32'hbb817338),
	.w4(32'h3c85a5ee),
	.w5(32'h3c8393e9),
	.w6(32'h3c6ec8c4),
	.w7(32'h3ca5b010),
	.w8(32'h3c6322c6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ecb23),
	.w1(32'h3bce6580),
	.w2(32'h3c14bb94),
	.w3(32'h3c2999f0),
	.w4(32'h3c09c71a),
	.w5(32'h3ba2b4a2),
	.w6(32'hb9749466),
	.w7(32'h3ab087f4),
	.w8(32'hbaa751fc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be77051),
	.w1(32'hbb8107cf),
	.w2(32'hbb85dd7f),
	.w3(32'hb993dcaa),
	.w4(32'hbb965d82),
	.w5(32'hbc5c5625),
	.w6(32'h3c803670),
	.w7(32'hbb950534),
	.w8(32'hbb3bda90),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5e99),
	.w1(32'h3b807004),
	.w2(32'h3ae25f41),
	.w3(32'hbc30d3bd),
	.w4(32'hbbe71401),
	.w5(32'hbbce9730),
	.w6(32'h3bc38f2f),
	.w7(32'h3bdfa90b),
	.w8(32'hba9bafd1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbac230),
	.w1(32'hbcdb53ec),
	.w2(32'hbc9eb9ff),
	.w3(32'hbc225f89),
	.w4(32'hbd122845),
	.w5(32'hbd102d88),
	.w6(32'h3bcd9244),
	.w7(32'hbc1ac913),
	.w8(32'hbb4cc009),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8fd0),
	.w1(32'hbc49f243),
	.w2(32'h3a8b60c7),
	.w3(32'hbc40e6e4),
	.w4(32'hbc0c8dba),
	.w5(32'hba277ddd),
	.w6(32'hbbf34e7e),
	.w7(32'hbb2731b2),
	.w8(32'h3a770584),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8005),
	.w1(32'h3b4401c0),
	.w2(32'h3c03b102),
	.w3(32'hb9d93bd3),
	.w4(32'h3b08719f),
	.w5(32'h3bb1da0d),
	.w6(32'h392816d5),
	.w7(32'h3ae03b7d),
	.w8(32'h3c8086e2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fb58b),
	.w1(32'hbbd90d20),
	.w2(32'h3a620a0f),
	.w3(32'h3c4c59de),
	.w4(32'h3b0dae4a),
	.w5(32'h3b550075),
	.w6(32'hbb9ceb73),
	.w7(32'h3b7bc557),
	.w8(32'h3b614b84),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f5200),
	.w1(32'hbb49f909),
	.w2(32'h3b1b1f59),
	.w3(32'hba1fa8de),
	.w4(32'h3b59a150),
	.w5(32'h3b92e658),
	.w6(32'hb6f330ec),
	.w7(32'h3ad0388f),
	.w8(32'hb939a741),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc63f75),
	.w1(32'hbc9a5413),
	.w2(32'hbcfe3a94),
	.w3(32'h3a1f823f),
	.w4(32'hbc79660f),
	.w5(32'hbc75aed4),
	.w6(32'hba23c4aa),
	.w7(32'hbc6f95ac),
	.w8(32'hbc469c96),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4c973),
	.w1(32'h3ba64a87),
	.w2(32'h3c59bc66),
	.w3(32'hbb8cbbcd),
	.w4(32'h3c244990),
	.w5(32'h3bf744a0),
	.w6(32'h3b093368),
	.w7(32'h3bf51c77),
	.w8(32'h3c90122e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b9824),
	.w1(32'h3c2a4a9e),
	.w2(32'h3c8b44be),
	.w3(32'h3c88998d),
	.w4(32'h3cb47cca),
	.w5(32'h3cb9dd40),
	.w6(32'h3c096621),
	.w7(32'h3c8e3204),
	.w8(32'h3c546b99),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e38ce),
	.w1(32'hbae1cc1d),
	.w2(32'hbc6cbab6),
	.w3(32'h3ab5da00),
	.w4(32'hbb8accf5),
	.w5(32'hbbdd8833),
	.w6(32'h3bc7a848),
	.w7(32'h3b975a3d),
	.w8(32'hb9a52286),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d66e),
	.w1(32'h3b83e12c),
	.w2(32'h3b977330),
	.w3(32'h3b167796),
	.w4(32'h3b58e77e),
	.w5(32'h3b8f1a23),
	.w6(32'h3bac3011),
	.w7(32'h3b9a61b4),
	.w8(32'h3b01ff61),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545d8b),
	.w1(32'hbbeef938),
	.w2(32'hbb2b87b4),
	.w3(32'h3bf9df4c),
	.w4(32'hbbc7472b),
	.w5(32'hba9aae3e),
	.w6(32'hbb90e0cb),
	.w7(32'hba3aee21),
	.w8(32'hbb6bab60),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b0053),
	.w1(32'hbc7a04da),
	.w2(32'hbcdfe8f6),
	.w3(32'hbada6bd6),
	.w4(32'hbc62b0b7),
	.w5(32'hbca83747),
	.w6(32'h3bc3f169),
	.w7(32'hbbf4ef46),
	.w8(32'hbc1eddd1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78f92a),
	.w1(32'hbb9efcd7),
	.w2(32'hbc0f2530),
	.w3(32'hbc0f7b88),
	.w4(32'hbb8baa7a),
	.w5(32'hbc0a6368),
	.w6(32'h3afb0f27),
	.w7(32'hbc2bdd94),
	.w8(32'hbc20d821),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e810a),
	.w1(32'hbc03cb9a),
	.w2(32'hbaa52a2c),
	.w3(32'hbc9990d3),
	.w4(32'hbc089f8b),
	.w5(32'hbacb7e12),
	.w6(32'hbbc7164c),
	.w7(32'h3bd9a301),
	.w8(32'hbbdf386a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad85110),
	.w1(32'hbc2addca),
	.w2(32'h3b498a3d),
	.w3(32'hba9dedb3),
	.w4(32'hbc4b4f2c),
	.w5(32'h3ab0f3e1),
	.w6(32'hbba56fc6),
	.w7(32'h3aa1ac7c),
	.w8(32'hbc003742),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb302c0f),
	.w1(32'h3bb02dd2),
	.w2(32'h3aff4a50),
	.w3(32'hba6d1894),
	.w4(32'h3b9141b1),
	.w5(32'h3b9effc0),
	.w6(32'h3bae13f2),
	.w7(32'h3b98a753),
	.w8(32'hbacadc10),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373f22a2),
	.w1(32'hbcd331e4),
	.w2(32'hbd3d8dcd),
	.w3(32'h3b9cba41),
	.w4(32'hbcf5d75d),
	.w5(32'hbd1e3654),
	.w6(32'hbc31f301),
	.w7(32'hbccb3a81),
	.w8(32'hbcca521f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcebbf29),
	.w1(32'hbb73b983),
	.w2(32'h3c60057c),
	.w3(32'hbbc88832),
	.w4(32'hbc2e9a7a),
	.w5(32'h3b01a825),
	.w6(32'h3b2a5e11),
	.w7(32'h3bc45dc7),
	.w8(32'hbb0db1c0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b81de4),
	.w1(32'hbc001648),
	.w2(32'h3a064527),
	.w3(32'hbbf7066b),
	.w4(32'hbbf0d4c6),
	.w5(32'hb8a53eda),
	.w6(32'hba16a2ab),
	.w7(32'h3b197968),
	.w8(32'h3b8c7b16),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbf6b9),
	.w1(32'hb9f365ac),
	.w2(32'h3b89dc4e),
	.w3(32'h3b1f6aa1),
	.w4(32'h3b36037b),
	.w5(32'h3b56fb82),
	.w6(32'hbb741b80),
	.w7(32'h3b44fcca),
	.w8(32'h3b2fc32b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bded076),
	.w1(32'hbc0e9e7d),
	.w2(32'hbc915e2f),
	.w3(32'h3b1ba2b0),
	.w4(32'hbc7e10a6),
	.w5(32'hbc71d830),
	.w6(32'hbb43b7da),
	.w7(32'hbc0b1610),
	.w8(32'hbc1e4471),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86bcd0),
	.w1(32'hbbb53961),
	.w2(32'hbc39d620),
	.w3(32'hbbae2f36),
	.w4(32'hbbfa2adc),
	.w5(32'hbc2b5eb2),
	.w6(32'hbbaea29f),
	.w7(32'hbbf94554),
	.w8(32'hbb976f9f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16b0e0),
	.w1(32'hbc8f9e58),
	.w2(32'hbd14fdd0),
	.w3(32'hbb50e1fa),
	.w4(32'hbcbf0fad),
	.w5(32'hbd064da2),
	.w6(32'hbb385a69),
	.w7(32'hbc84ac81),
	.w8(32'hbc642e31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4bd6),
	.w1(32'h3bf2a328),
	.w2(32'h3baff2a7),
	.w3(32'h3b4fca00),
	.w4(32'h3c379479),
	.w5(32'h3bc148b6),
	.w6(32'h3c1881af),
	.w7(32'h3c647c08),
	.w8(32'h3c0589ea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97b37),
	.w1(32'h3c2eca6a),
	.w2(32'h3caccf2c),
	.w3(32'hbb32b516),
	.w4(32'hbc31fb42),
	.w5(32'h3c0024ce),
	.w6(32'h3c02a976),
	.w7(32'hbb2317e9),
	.w8(32'h3b5ed7d8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c793ce0),
	.w1(32'h3acdc093),
	.w2(32'h3ba12228),
	.w3(32'h3a73338d),
	.w4(32'hbb4cbd9e),
	.w5(32'h3ba47ad5),
	.w6(32'h3bf9d493),
	.w7(32'h3b0e7f9f),
	.w8(32'hbb8b5ec2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95cb40),
	.w1(32'hbcc44bd5),
	.w2(32'hbccc4bdb),
	.w3(32'hb862ecbe),
	.w4(32'hbc241413),
	.w5(32'hbb8ac59c),
	.w6(32'hbaadfd13),
	.w7(32'hbbc919ee),
	.w8(32'hbb594cdd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1397b0),
	.w1(32'hbca327e3),
	.w2(32'hbd12a93c),
	.w3(32'h3bba9138),
	.w4(32'hbce9488a),
	.w5(32'hbcf71d4f),
	.w6(32'hbc067bf3),
	.w7(32'hbc92c315),
	.w8(32'hbcb9afae),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ac5d4),
	.w1(32'hbcbe4c78),
	.w2(32'hbd22a48e),
	.w3(32'hbc488f09),
	.w4(32'hbcd78d30),
	.w5(32'hbd163b63),
	.w6(32'h3b3b5426),
	.w7(32'hbc66b1b3),
	.w8(32'hbc8ad65a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb5e0c),
	.w1(32'h3aa5ca08),
	.w2(32'h3ba0c223),
	.w3(32'hbcac0e6e),
	.w4(32'hba493729),
	.w5(32'h3c1c9c5c),
	.w6(32'h3bb41a12),
	.w7(32'hbb44912a),
	.w8(32'h3bd2d93b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86b1d),
	.w1(32'h3b155b5b),
	.w2(32'h3c0de2f9),
	.w3(32'h3c04304c),
	.w4(32'hbb61e0a7),
	.w5(32'h3baaa133),
	.w6(32'h3b2cbfa2),
	.w7(32'h3ab17e4c),
	.w8(32'h3bb4bf37),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea40d4),
	.w1(32'h3af38ee4),
	.w2(32'h3b11cbe2),
	.w3(32'h3c541b24),
	.w4(32'hb97c4f30),
	.w5(32'hbb077f8f),
	.w6(32'h3b127aad),
	.w7(32'h3b459f97),
	.w8(32'h3b94f10d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdc2fe),
	.w1(32'h3c7bf3c8),
	.w2(32'h3cf03c8c),
	.w3(32'hb9cf98e9),
	.w4(32'h3bcb2672),
	.w5(32'h3c3e2fb3),
	.w6(32'h3bc0f0c6),
	.w7(32'h3c551808),
	.w8(32'h3c8f6e2f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc56fa0),
	.w1(32'h3bcb3883),
	.w2(32'hbb1c6a88),
	.w3(32'h3c903515),
	.w4(32'hbc4209c3),
	.w5(32'hbbae9095),
	.w6(32'h3a69afb9),
	.w7(32'hbb09bbe0),
	.w8(32'h3b2820ca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ba29e),
	.w1(32'hbbcd02bf),
	.w2(32'h3bb7408e),
	.w3(32'h3b102b09),
	.w4(32'hbae9873e),
	.w5(32'h3b81862a),
	.w6(32'hbbc81b46),
	.w7(32'hbb067fce),
	.w8(32'hba8c8afd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978f78),
	.w1(32'hbcb9cef7),
	.w2(32'hbc38029b),
	.w3(32'hbc5ab770),
	.w4(32'hbcbc8fda),
	.w5(32'hbc6734fe),
	.w6(32'hbc1ccb61),
	.w7(32'hbc014076),
	.w8(32'hbbf71d90),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22c978),
	.w1(32'hbaa9f06e),
	.w2(32'h3b0317c4),
	.w3(32'hbc14c227),
	.w4(32'hba8ce8a7),
	.w5(32'hbb370d19),
	.w6(32'hbb91fee7),
	.w7(32'hba8448f7),
	.w8(32'h3b2910d7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388508c9),
	.w1(32'hbb211cf6),
	.w2(32'h3b2811e4),
	.w3(32'hbab70e79),
	.w4(32'hbb9530ef),
	.w5(32'h3a7def05),
	.w6(32'hbb029b0c),
	.w7(32'h3a761100),
	.w8(32'h3ae8b839),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fd5a9),
	.w1(32'hbb833286),
	.w2(32'hbb1db31b),
	.w3(32'hba7b75e9),
	.w4(32'hbbb2dbd0),
	.w5(32'hbc1cacfc),
	.w6(32'h3aca9aff),
	.w7(32'h390c704d),
	.w8(32'hbb08cab3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcce40c),
	.w1(32'hbc26a31c),
	.w2(32'hbc8a7f10),
	.w3(32'hbb84d31a),
	.w4(32'hbc0a63fc),
	.w5(32'hbc20a1c5),
	.w6(32'hbb3ea9e5),
	.w7(32'hbb30d6b3),
	.w8(32'hbc3ea9bf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f773),
	.w1(32'h3c636e73),
	.w2(32'h3be55a4f),
	.w3(32'h3c177560),
	.w4(32'h3c2feb46),
	.w5(32'h3c08aa51),
	.w6(32'h3c28274c),
	.w7(32'h3c29fb74),
	.w8(32'h3c3df3a2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2e678),
	.w1(32'hbca1c21f),
	.w2(32'hbd1372e7),
	.w3(32'h3b36542a),
	.w4(32'hbca7ea77),
	.w5(32'hbd038a1d),
	.w6(32'hbc2da775),
	.w7(32'hbcbc3ca9),
	.w8(32'hbccce6ee),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc011f5),
	.w1(32'h3c84ccf1),
	.w2(32'h3d1c0f3c),
	.w3(32'hbcacb75d),
	.w4(32'h3c790fd4),
	.w5(32'h3ca5fb9e),
	.w6(32'hbb68211e),
	.w7(32'h3c91d1eb),
	.w8(32'h3c4ed431),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9aaedf),
	.w1(32'h3ac66170),
	.w2(32'h39305ff7),
	.w3(32'hba050e76),
	.w4(32'h3adfe1d7),
	.w5(32'h3a61b869),
	.w6(32'hbabe1483),
	.w7(32'hbb6beca3),
	.w8(32'h3b94c313),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbacbc),
	.w1(32'h3a0599f0),
	.w2(32'hbc0c880b),
	.w3(32'h3b15dfb4),
	.w4(32'h3ba93d7e),
	.w5(32'h3b970f4a),
	.w6(32'h3c883719),
	.w7(32'h3c0635df),
	.w8(32'hbaedc801),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba23b5),
	.w1(32'hbaca6132),
	.w2(32'hbc223574),
	.w3(32'h3c84fd3a),
	.w4(32'hbc247e7b),
	.w5(32'h3b5cebb8),
	.w6(32'h3c233154),
	.w7(32'h3b720a5f),
	.w8(32'h3b4b6646),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cb9e9),
	.w1(32'hbc2b1b07),
	.w2(32'h3b9e0f9a),
	.w3(32'h3b8d2021),
	.w4(32'hbc05c7a3),
	.w5(32'hbbbfdeb8),
	.w6(32'hbc039090),
	.w7(32'hbb520a1c),
	.w8(32'h39e07108),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b416187),
	.w1(32'h3ab97006),
	.w2(32'h3a982e29),
	.w3(32'h3b69c4c0),
	.w4(32'h3bf55209),
	.w5(32'h3b17bdf4),
	.w6(32'hbb12f55a),
	.w7(32'hbbfdbafe),
	.w8(32'hbb4d04db),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad694c8),
	.w1(32'h3b952e8a),
	.w2(32'h3c4fad26),
	.w3(32'hbb82829a),
	.w4(32'h3b3edc2c),
	.w5(32'h3a9d0517),
	.w6(32'h3c400890),
	.w7(32'h3c5af8b2),
	.w8(32'h3bec8767),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c288a61),
	.w1(32'h3ba52b09),
	.w2(32'h3c19b546),
	.w3(32'h3bb215b5),
	.w4(32'h3bc770a4),
	.w5(32'h3c234fbd),
	.w6(32'hba3957fc),
	.w7(32'h3b144284),
	.w8(32'h3ba151c8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d8ec),
	.w1(32'hba3b374a),
	.w2(32'h3bbc6905),
	.w3(32'hbb862d16),
	.w4(32'hbb901202),
	.w5(32'h3aea4158),
	.w6(32'h3b3c0744),
	.w7(32'h3abd8609),
	.w8(32'h3b253724),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6b542),
	.w1(32'hbb9e7feb),
	.w2(32'hbc4a7c86),
	.w3(32'h3bb4977d),
	.w4(32'hbb964823),
	.w5(32'hbb01e24e),
	.w6(32'h3b8408d8),
	.w7(32'hbbc7c8b9),
	.w8(32'h3b823712),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e3f36),
	.w1(32'hbc91f755),
	.w2(32'hbcbf7a4c),
	.w3(32'h3c612717),
	.w4(32'hbc6b96fe),
	.w5(32'hbc8cb6d1),
	.w6(32'hbb923fb4),
	.w7(32'hbcb5e441),
	.w8(32'hbc302776),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc672a93),
	.w1(32'hbb6b8d6e),
	.w2(32'hbcc500d6),
	.w3(32'hbc17ec49),
	.w4(32'hbbb82758),
	.w5(32'hbbeeddf3),
	.w6(32'h394882d0),
	.w7(32'hbb9eb13b),
	.w8(32'hbc518acd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ba654),
	.w1(32'hbca6d619),
	.w2(32'hbcec979c),
	.w3(32'h3c087114),
	.w4(32'hbc3cf23a),
	.w5(32'hbc8e6f0d),
	.w6(32'hbc8136e8),
	.w7(32'hbca847b1),
	.w8(32'hbca92410),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc718ad4),
	.w1(32'hbc344c96),
	.w2(32'hbc2c2d9e),
	.w3(32'hbcc433ad),
	.w4(32'hbc82ff3d),
	.w5(32'hbc549ba5),
	.w6(32'h3a8f93b6),
	.w7(32'hbbd28781),
	.w8(32'hbb9e3ded),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5851),
	.w1(32'hbbc4603b),
	.w2(32'hbc3b2e05),
	.w3(32'hbc32797f),
	.w4(32'hbbfaf2b9),
	.w5(32'hbc81cf2e),
	.w6(32'hbc034903),
	.w7(32'hbad7f0a3),
	.w8(32'hbc264d34),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2033e),
	.w1(32'hbce94934),
	.w2(32'hbd373077),
	.w3(32'hbbd65e0b),
	.w4(32'hbd1a0527),
	.w5(32'hbd2a853d),
	.w6(32'h3b3f7c8e),
	.w7(32'hbc96d8f7),
	.w8(32'hbc9bb972),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcffdc65),
	.w1(32'h3bde43db),
	.w2(32'h3be6ca46),
	.w3(32'hbbddd00e),
	.w4(32'h3abdfd30),
	.w5(32'hbbb13bce),
	.w6(32'h3c16fe62),
	.w7(32'h3be7f4ee),
	.w8(32'hbb1c14b6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa25b50),
	.w1(32'hba063eb2),
	.w2(32'h3a61ba71),
	.w3(32'hbb468913),
	.w4(32'h3ae2c2dc),
	.w5(32'h3b84cc90),
	.w6(32'hba73aa4e),
	.w7(32'h39b7eef3),
	.w8(32'h3b17316f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b2d2f),
	.w1(32'hbb0d600f),
	.w2(32'h39614df4),
	.w3(32'h3be9ad9a),
	.w4(32'hbbb167a9),
	.w5(32'hbb2f1edd),
	.w6(32'hbb8cfa6b),
	.w7(32'hbb529068),
	.w8(32'hbb12737f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd2da5),
	.w1(32'hbbacf912),
	.w2(32'hbac0e9a2),
	.w3(32'hbb9a238d),
	.w4(32'h3b441729),
	.w5(32'h3b93eae2),
	.w6(32'hbb0f63ce),
	.w7(32'hbb15897c),
	.w8(32'hbaca14b3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801710),
	.w1(32'h3baf6cd1),
	.w2(32'hb99a3b69),
	.w3(32'h3bed9789),
	.w4(32'hbb639509),
	.w5(32'h3b178f19),
	.w6(32'hbb3bfb27),
	.w7(32'h3c014618),
	.w8(32'h3bbe9793),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2d6e),
	.w1(32'h3b302b26),
	.w2(32'hbbf66643),
	.w3(32'h3c2e82c5),
	.w4(32'hbb096389),
	.w5(32'hba4c329d),
	.w6(32'h3c6214e2),
	.w7(32'h3c13fa9f),
	.w8(32'h3c1002ca),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d751),
	.w1(32'h3c2f1849),
	.w2(32'h3c033642),
	.w3(32'h3c4ae172),
	.w4(32'h3bc1fbfd),
	.w5(32'h3c3edec2),
	.w6(32'h3b57f829),
	.w7(32'h3b0cdadd),
	.w8(32'h3ba2e6e6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc1fb),
	.w1(32'h3b60baf8),
	.w2(32'h3b3f0a55),
	.w3(32'h3b425347),
	.w4(32'h3b638138),
	.w5(32'h3ab14526),
	.w6(32'h3a60f119),
	.w7(32'hbac5f92f),
	.w8(32'h3b232fae),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8989),
	.w1(32'hbb932430),
	.w2(32'hbb881562),
	.w3(32'h3b876c65),
	.w4(32'hbbf96c4c),
	.w5(32'hbbc10fe1),
	.w6(32'hb9c1d5d8),
	.w7(32'hbb8f1d86),
	.w8(32'hbb884048),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396bdb61),
	.w1(32'h394157b3),
	.w2(32'h3b7cd347),
	.w3(32'h3b0b2d6c),
	.w4(32'h3b14f9d2),
	.w5(32'hbbacc3e4),
	.w6(32'hbb3d13de),
	.w7(32'h3b538d88),
	.w8(32'hbb164868),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7107a2),
	.w1(32'hbbdff417),
	.w2(32'hbb9c3a95),
	.w3(32'hbc426631),
	.w4(32'hbb15523e),
	.w5(32'hbad0d364),
	.w6(32'h3a3f491d),
	.w7(32'h390bdf99),
	.w8(32'hba54e53c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6072),
	.w1(32'h3c500017),
	.w2(32'h3cc701a4),
	.w3(32'h3ae641ff),
	.w4(32'h3aad08a9),
	.w5(32'hb9576b1c),
	.w6(32'h3b8572f0),
	.w7(32'h3c49fe9f),
	.w8(32'h3aa3aaba),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7d538),
	.w1(32'hbc9b494e),
	.w2(32'hbcd04f75),
	.w3(32'hbb0e8fd9),
	.w4(32'hbcd20d1b),
	.w5(32'hbcf80921),
	.w6(32'hb6614cd8),
	.w7(32'hbc696010),
	.w8(32'hbc8a526d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a2ca1),
	.w1(32'hbcbe9fc0),
	.w2(32'hbd24792d),
	.w3(32'hbbe21faf),
	.w4(32'hbcf36986),
	.w5(32'hbce7e7ee),
	.w6(32'hbb255a79),
	.w7(32'hbc912895),
	.w8(32'hbc6218f9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4d55),
	.w1(32'hbc0c12fe),
	.w2(32'hbc1d4fc6),
	.w3(32'hbb86235d),
	.w4(32'hbc092cbf),
	.w5(32'h3b7f0c1f),
	.w6(32'h3b3f3e1e),
	.w7(32'hbc3efd89),
	.w8(32'hbc223287),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aae05),
	.w1(32'hbc1fe343),
	.w2(32'hbc0bdc81),
	.w3(32'h3bae126b),
	.w4(32'hbb9146fb),
	.w5(32'h3abe3d14),
	.w6(32'hbbb3bfe1),
	.w7(32'hbc0c5ddd),
	.w8(32'hbc29c9ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeabb20),
	.w1(32'hbba2dc8b),
	.w2(32'h3817722c),
	.w3(32'h3be3e6ca),
	.w4(32'hbb618e56),
	.w5(32'h3ad39e4c),
	.w6(32'h3a458492),
	.w7(32'hbaae26a9),
	.w8(32'hba902cf4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0ff46),
	.w1(32'hbc0e18e6),
	.w2(32'hbc04d94b),
	.w3(32'h3c7610c3),
	.w4(32'h3b237552),
	.w5(32'h3ade70e4),
	.w6(32'h3a08754d),
	.w7(32'hbb2c5d3f),
	.w8(32'hba41373e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825d5c),
	.w1(32'hbb1f2892),
	.w2(32'h3aaec6ea),
	.w3(32'hbb4c12c5),
	.w4(32'hbba5006c),
	.w5(32'h39d834d3),
	.w6(32'h3b9bf858),
	.w7(32'hbb1b1421),
	.w8(32'hbc047703),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806ec1),
	.w1(32'hbc250bec),
	.w2(32'hbc62c4cd),
	.w3(32'hba9f4f71),
	.w4(32'hbc4e0da3),
	.w5(32'hbc65e5d7),
	.w6(32'hbb8c1b12),
	.w7(32'hbc1e85c6),
	.w8(32'hbbf5d579),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6514),
	.w1(32'hbb708319),
	.w2(32'h3bddb739),
	.w3(32'h3bab4c4f),
	.w4(32'hbc1c0615),
	.w5(32'hb9d12652),
	.w6(32'hbb5a78b0),
	.w7(32'h3931368d),
	.w8(32'hbb624f81),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96127a9),
	.w1(32'hbb7a0f4f),
	.w2(32'h3bdbe341),
	.w3(32'h3a85d5c1),
	.w4(32'h3baf0adb),
	.w5(32'h3aaf149b),
	.w6(32'hbc29c8bc),
	.w7(32'hbb8de662),
	.w8(32'hbb223af3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3706667e),
	.w1(32'h3ac03dc0),
	.w2(32'hbbc27643),
	.w3(32'hbb07ed02),
	.w4(32'h3ac1f9d2),
	.w5(32'h3afae6a0),
	.w6(32'h3c706f01),
	.w7(32'h3b5cc594),
	.w8(32'hbc1eee6c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4e6e),
	.w1(32'h3ba72a25),
	.w2(32'h3baa68ab),
	.w3(32'h3c5738a6),
	.w4(32'h3c07f647),
	.w5(32'h3bdd1653),
	.w6(32'hbb0a8ff7),
	.w7(32'h3b8ac864),
	.w8(32'h3c2fbda6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cc727),
	.w1(32'hbb4c2ffe),
	.w2(32'hba097d99),
	.w3(32'h3b9ee9d8),
	.w4(32'hbb1e92ad),
	.w5(32'h3a9f35a8),
	.w6(32'h3b866bb2),
	.w7(32'h38f3e697),
	.w8(32'hba8400e0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9892dbc),
	.w1(32'hbaa844cd),
	.w2(32'hba4347dc),
	.w3(32'h3acc83d5),
	.w4(32'h3b8e38bb),
	.w5(32'h3b20c67d),
	.w6(32'h3b1b4161),
	.w7(32'h3bd92881),
	.w8(32'h3b5f936d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc419652),
	.w1(32'h399a89e4),
	.w2(32'h3b9f83ae),
	.w3(32'hbaf7a8df),
	.w4(32'hbaeb2bb5),
	.w5(32'h3a398d02),
	.w6(32'hbb029118),
	.w7(32'h3aa321f4),
	.w8(32'h3b528aa5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca7f19),
	.w1(32'h3b8ffdf1),
	.w2(32'h3c6475ba),
	.w3(32'h3b943f32),
	.w4(32'hbb7026a4),
	.w5(32'h3c6fc0fb),
	.w6(32'h3a503da9),
	.w7(32'h3b2cb9d2),
	.w8(32'hbb02a2a1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25b7af),
	.w1(32'hbbdfb47e),
	.w2(32'hbbe1de0c),
	.w3(32'hbbaeb0b8),
	.w4(32'hb9d3d502),
	.w5(32'hba2ff8a8),
	.w6(32'h3a550455),
	.w7(32'hbb9f8e8c),
	.w8(32'hbc217fcb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f52f9),
	.w1(32'h3a4cb062),
	.w2(32'hb93d8911),
	.w3(32'h3a60cb15),
	.w4(32'h3a7b0725),
	.w5(32'h3a8e7363),
	.w6(32'h3b955e52),
	.w7(32'h3b9e2a67),
	.w8(32'h3a17c092),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfe276),
	.w1(32'hbb145fc1),
	.w2(32'h398fba37),
	.w3(32'h3b38c67a),
	.w4(32'hbaa482f8),
	.w5(32'h3b3405c6),
	.w6(32'h3afd0574),
	.w7(32'h3a38b9ae),
	.w8(32'h3ae27e21),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a919107),
	.w1(32'h3c21fe35),
	.w2(32'h3c80d217),
	.w3(32'h3b0a381a),
	.w4(32'h3c07bfce),
	.w5(32'h3c946739),
	.w6(32'h3a60d3bd),
	.w7(32'h3baf5bf0),
	.w8(32'h3c4c4350),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87c663),
	.w1(32'h3ba3c8ff),
	.w2(32'h3c109e9b),
	.w3(32'h3c312ed1),
	.w4(32'h3aacf365),
	.w5(32'h3b3c74b7),
	.w6(32'h3b3997d1),
	.w7(32'h3b90c8fc),
	.w8(32'h3c144c51),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154a69),
	.w1(32'hbca419f5),
	.w2(32'hbcf56cc6),
	.w3(32'h3bd909b5),
	.w4(32'hbc87fc4c),
	.w5(32'hbcb6e524),
	.w6(32'hbba402cc),
	.w7(32'hbc9d37e0),
	.w8(32'hbcd1a304),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c8444),
	.w1(32'h3c1d5773),
	.w2(32'h3bb34621),
	.w3(32'hbbd0a8ad),
	.w4(32'h3b0ac788),
	.w5(32'hba9cca39),
	.w6(32'h3b3fb925),
	.w7(32'h3b414162),
	.w8(32'h3aa6cfaf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdd4f8),
	.w1(32'hbc8c897a),
	.w2(32'hbcb65228),
	.w3(32'hbbadf0e8),
	.w4(32'hbc4d4039),
	.w5(32'hbc606b78),
	.w6(32'hbc491483),
	.w7(32'hbc3da0a4),
	.w8(32'hbc694aa1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c39aa),
	.w1(32'hbb575e07),
	.w2(32'hbafbbf0b),
	.w3(32'hbc88e14d),
	.w4(32'hbbbf049d),
	.w5(32'h3b63ec9c),
	.w6(32'hba09b63c),
	.w7(32'hbb2b985b),
	.w8(32'h3ad6a48b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d377),
	.w1(32'h3ac2e38e),
	.w2(32'h3b710174),
	.w3(32'h3ba5de00),
	.w4(32'h3b6da069),
	.w5(32'h3b841fc4),
	.w6(32'h3bbbb492),
	.w7(32'h3b9c6783),
	.w8(32'h3bb500a9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7e4cb),
	.w1(32'hbb9751e1),
	.w2(32'h3bd8d951),
	.w3(32'h3be52adb),
	.w4(32'hbae851a4),
	.w5(32'h3b89447f),
	.w6(32'h3b70abc8),
	.w7(32'h3c309cb7),
	.w8(32'h3b1f617c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720191),
	.w1(32'hbbe5ea3f),
	.w2(32'hbc52279a),
	.w3(32'hbab28d46),
	.w4(32'hba2a9392),
	.w5(32'h3b345be2),
	.w6(32'hba2e0ed4),
	.w7(32'hbc3f1719),
	.w8(32'hbc36c60d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4939f1),
	.w1(32'hbbc84886),
	.w2(32'hbc09abd8),
	.w3(32'h3bed0e11),
	.w4(32'hbc6dfaf6),
	.w5(32'hbbb44e49),
	.w6(32'h3b96aab4),
	.w7(32'hba7c34f5),
	.w8(32'hbc01657a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96610c),
	.w1(32'h3afc49c6),
	.w2(32'h3aee3fba),
	.w3(32'hbad5cb45),
	.w4(32'h3aa4d726),
	.w5(32'h3a4d9bfc),
	.w6(32'h3b160f7c),
	.w7(32'h3b2f4416),
	.w8(32'h3b2c63d2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b644ee1),
	.w1(32'h3b7358e0),
	.w2(32'h3be7346e),
	.w3(32'h3a49f9bd),
	.w4(32'hbb367247),
	.w5(32'hbb2b973d),
	.w6(32'hb91c0de2),
	.w7(32'hbb420ca0),
	.w8(32'h3a24d10e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule