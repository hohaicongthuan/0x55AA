module layer_8_featuremap_236(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06a29),
	.w1(32'hbb000c53),
	.w2(32'h3b1a8bb8),
	.w3(32'hbb9020c7),
	.w4(32'h3b0b41de),
	.w5(32'hbbc27010),
	.w6(32'h3a77f997),
	.w7(32'h3b8d0dc0),
	.w8(32'hbae33ecc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68dcf5),
	.w1(32'h3d07866c),
	.w2(32'h3d99650f),
	.w3(32'h3af6f66b),
	.w4(32'h3c8b6e68),
	.w5(32'h3d5a55e6),
	.w6(32'h3a1c796d),
	.w7(32'h3cff43b2),
	.w8(32'h3c835722),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5617fd),
	.w1(32'h3b393c4d),
	.w2(32'h3a60d72d),
	.w3(32'h3d0998c5),
	.w4(32'hbb85c987),
	.w5(32'hba8e4be7),
	.w6(32'hbba0c27b),
	.w7(32'hbb514d0e),
	.w8(32'hbb640708),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a879e6e),
	.w1(32'h3b1a0cb0),
	.w2(32'hba17aeb9),
	.w3(32'hbb78be31),
	.w4(32'h3b9f11b4),
	.w5(32'h3b8cd0f4),
	.w6(32'h3bbf365f),
	.w7(32'h3b8c6e0b),
	.w8(32'h3b92f130),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebb1f0),
	.w1(32'hbcea9e1b),
	.w2(32'hbbcc7e3f),
	.w3(32'h3ae87e5a),
	.w4(32'hbd36c30c),
	.w5(32'hbcdfd04a),
	.w6(32'hbd4233d0),
	.w7(32'hbd03fd17),
	.w8(32'hbd282095),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9efaf),
	.w1(32'h3c0d314b),
	.w2(32'h3bc97f7d),
	.w3(32'hbd28f3ce),
	.w4(32'h3b525d85),
	.w5(32'h3b345003),
	.w6(32'h3bb222ef),
	.w7(32'h3bcac67f),
	.w8(32'hba68286c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94b8a4),
	.w1(32'hbca798e6),
	.w2(32'hbd2af404),
	.w3(32'h3b90e2e0),
	.w4(32'hbc5ccaf9),
	.w5(32'hbd0348ee),
	.w6(32'hbb2df50e),
	.w7(32'hbc9bd4a0),
	.w8(32'hbc3aa0c6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf14a0d),
	.w1(32'h3a79044a),
	.w2(32'hb9a7c5e8),
	.w3(32'hbcb0f973),
	.w4(32'h3b41b626),
	.w5(32'h3a9e43c7),
	.w6(32'h3a106cdf),
	.w7(32'hbafd3255),
	.w8(32'hba95d907),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de354),
	.w1(32'h3c1d7406),
	.w2(32'h3ca44e77),
	.w3(32'hba714323),
	.w4(32'hbc0e1b36),
	.w5(32'hbb5a4f86),
	.w6(32'hba9ff87f),
	.w7(32'h3ae2275a),
	.w8(32'hbbd4dfdc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d7b5a),
	.w1(32'h3aac950a),
	.w2(32'hbbc8a9ac),
	.w3(32'hbc855826),
	.w4(32'hbb0a187f),
	.w5(32'hbb87066a),
	.w6(32'hba8b3c48),
	.w7(32'hbba64f22),
	.w8(32'hba2b4fd8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556d47),
	.w1(32'hb9ebce6f),
	.w2(32'h3aace9a3),
	.w3(32'hbbe563bb),
	.w4(32'hbb56cdf5),
	.w5(32'hb96fe468),
	.w6(32'h3bea6f64),
	.w7(32'h3c0ae703),
	.w8(32'h3c21373f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb90500),
	.w1(32'hb9f6fee1),
	.w2(32'hbb80ec25),
	.w3(32'h3ab9575f),
	.w4(32'h39ce6ef6),
	.w5(32'h3a92fb34),
	.w6(32'h3abec6ca),
	.w7(32'hbaa9a6fd),
	.w8(32'hbacb372d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8ddae),
	.w1(32'hbb4fd072),
	.w2(32'h3a286589),
	.w3(32'hbb4d33a1),
	.w4(32'h3abef688),
	.w5(32'hbb3eb9cb),
	.w6(32'hbbf07cc0),
	.w7(32'hbac0f4f5),
	.w8(32'hbbd84c1f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26880),
	.w1(32'h3aca0ea0),
	.w2(32'h3afc154d),
	.w3(32'hbb9b6814),
	.w4(32'hba802ee7),
	.w5(32'h3b4b48af),
	.w6(32'hbad7c1d3),
	.w7(32'hbb93a8df),
	.w8(32'h3a25b74b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3dc05),
	.w1(32'hbc50a578),
	.w2(32'hbd2bce74),
	.w3(32'h3a954510),
	.w4(32'h3a8f96b9),
	.w5(32'hbcc2669b),
	.w6(32'h3c4f7330),
	.w7(32'hbc6fdfa1),
	.w8(32'hb97f9bae),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9d42d),
	.w1(32'h3b57d045),
	.w2(32'h39577d25),
	.w3(32'hbbf07e8d),
	.w4(32'hb9cab50f),
	.w5(32'hbbaa5cca),
	.w6(32'hbb4b42b3),
	.w7(32'h3b49ef30),
	.w8(32'hb92bc460),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b569011),
	.w1(32'h3b20209b),
	.w2(32'h3a3522aa),
	.w3(32'hbacf661a),
	.w4(32'h3ae9ccb2),
	.w5(32'h3b171fc8),
	.w6(32'h3a7124c4),
	.w7(32'h3b39221a),
	.w8(32'hb9dc054f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bd782),
	.w1(32'h3a68252b),
	.w2(32'hbb13b4f5),
	.w3(32'h3b62f7f9),
	.w4(32'h3c263a2c),
	.w5(32'h3aceaa19),
	.w6(32'hbb9d52c3),
	.w7(32'h3aecfafc),
	.w8(32'h3b3a20fc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fdc62),
	.w1(32'h3c024753),
	.w2(32'hbb30b497),
	.w3(32'hbb38fb08),
	.w4(32'h3c10d317),
	.w5(32'h3a83734e),
	.w6(32'h3af090e2),
	.w7(32'hbb6e40ac),
	.w8(32'hbbc24d39),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe6996),
	.w1(32'hbd173126),
	.w2(32'hbd9c2738),
	.w3(32'hbb8b35bb),
	.w4(32'hbcbad6e9),
	.w5(32'hbd6d3b54),
	.w6(32'hbba4364c),
	.w7(32'hbd12e1ec),
	.w8(32'hbcb45d8b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd669010),
	.w1(32'hbb3d17ec),
	.w2(32'h3ad4ac7f),
	.w3(32'hbd24789c),
	.w4(32'hbbe18e40),
	.w5(32'hbbfc6e94),
	.w6(32'hbb7edb12),
	.w7(32'h39e11997),
	.w8(32'hbba49b77),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661997),
	.w1(32'h3b226e91),
	.w2(32'h3b1d072b),
	.w3(32'hbbd82cf5),
	.w4(32'h3af415c3),
	.w5(32'h3bb38a61),
	.w6(32'hba22fda3),
	.w7(32'h396fa96f),
	.w8(32'h3ac6b5e4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514ea8),
	.w1(32'h3b11b044),
	.w2(32'h3994620a),
	.w3(32'hba2c5f4a),
	.w4(32'h3b8ca315),
	.w5(32'h3bce597b),
	.w6(32'hbb055ec6),
	.w7(32'hbb74fadb),
	.w8(32'h3b0ab93b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80e03),
	.w1(32'h3b128b41),
	.w2(32'h3b5a1535),
	.w3(32'h3bb243be),
	.w4(32'hbb65f8db),
	.w5(32'h392e0d20),
	.w6(32'h3b67b791),
	.w7(32'hbb9c861b),
	.w8(32'hbbc4d15a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8dedf),
	.w1(32'hba29ce42),
	.w2(32'h3abe481c),
	.w3(32'hbb635c7d),
	.w4(32'h3adc2cbe),
	.w5(32'h3bcb2dee),
	.w6(32'hbb877f8d),
	.w7(32'hbb914fa5),
	.w8(32'hbbd4f14f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a5708),
	.w1(32'hbabf14b8),
	.w2(32'h3bc81255),
	.w3(32'h3b4c2444),
	.w4(32'hbb6e6ae0),
	.w5(32'hb9c1d307),
	.w6(32'hbacd4e9c),
	.w7(32'h3be8e838),
	.w8(32'hba2ed735),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113b2f),
	.w1(32'hbb1183de),
	.w2(32'h3b56ec67),
	.w3(32'hbab700d3),
	.w4(32'hbb8be8e1),
	.w5(32'hbad7b61e),
	.w6(32'h38957c38),
	.w7(32'h3b15776e),
	.w8(32'hbb5f2d0e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a520ac2),
	.w1(32'h3b7cc7ed),
	.w2(32'h3ab3aed0),
	.w3(32'hba0533ff),
	.w4(32'h3b59b5c0),
	.w5(32'h39fb3d89),
	.w6(32'hbbcf816b),
	.w7(32'hbab29de3),
	.w8(32'hbb0ec039),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a38fe),
	.w1(32'h3c50671f),
	.w2(32'h3c01a4ee),
	.w3(32'hbbd07371),
	.w4(32'h3bf620a7),
	.w5(32'h3b65e36b),
	.w6(32'h3c9a91ad),
	.w7(32'h3c6cf2cb),
	.w8(32'hbb02715d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51447e),
	.w1(32'h3ba06e49),
	.w2(32'h3c3661a8),
	.w3(32'hbc836e57),
	.w4(32'hba20a8ab),
	.w5(32'hb9185030),
	.w6(32'h3ba8ac7a),
	.w7(32'h3bc708d6),
	.w8(32'h3bd2c2a4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c034c02),
	.w1(32'h3b2949b0),
	.w2(32'h3b4836c1),
	.w3(32'h3a2cc037),
	.w4(32'hbbd1a955),
	.w5(32'hbb8e3e93),
	.w6(32'h3c477380),
	.w7(32'h3c8838f9),
	.w8(32'h3c41c3c3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9277e),
	.w1(32'h3b4c963b),
	.w2(32'h3b8d637a),
	.w3(32'hbbd5e75d),
	.w4(32'h3ac42f4a),
	.w5(32'h3b96b3c9),
	.w6(32'h3b416dcb),
	.w7(32'h3b651caf),
	.w8(32'h3925f98c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95962bb),
	.w1(32'h3bb29864),
	.w2(32'h3be47324),
	.w3(32'h3b13bb1c),
	.w4(32'h3b16c9ca),
	.w5(32'h3b50b08e),
	.w6(32'h3b7653ec),
	.w7(32'h3b3a03c2),
	.w8(32'h3c17abed),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d199),
	.w1(32'hba337c23),
	.w2(32'hbc052b7d),
	.w3(32'h3b59b7ed),
	.w4(32'hbb25a0a0),
	.w5(32'h3ac77d14),
	.w6(32'hba8ebc27),
	.w7(32'hb9499867),
	.w8(32'hbb662af4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3b4c),
	.w1(32'hbc0e940d),
	.w2(32'hbaff98a2),
	.w3(32'hbb38e55d),
	.w4(32'hbaec091c),
	.w5(32'h3ba56919),
	.w6(32'hbbe3f41e),
	.w7(32'hbb1473e7),
	.w8(32'hbb89f6ce),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa509e),
	.w1(32'h3b06912d),
	.w2(32'h3b9909af),
	.w3(32'h3b4bc1f7),
	.w4(32'hb991eb08),
	.w5(32'hbacb963a),
	.w6(32'h3ad75ba9),
	.w7(32'h3ac53bf1),
	.w8(32'h3b43aa79),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabb206),
	.w1(32'h3bab79eb),
	.w2(32'h3b0a8282),
	.w3(32'hbb312e01),
	.w4(32'h3bd12c9b),
	.w5(32'h3b23083b),
	.w6(32'h3b0d6b68),
	.w7(32'hbade0cf7),
	.w8(32'hbb7c25c4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67820a),
	.w1(32'hbbbf344e),
	.w2(32'hbb9da70e),
	.w3(32'hbb2cb633),
	.w4(32'hbbde863b),
	.w5(32'hbc240791),
	.w6(32'hbb6ea93b),
	.w7(32'hbc239a38),
	.w8(32'hbb89b229),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ca29),
	.w1(32'h3a60d1d9),
	.w2(32'hbb1521b5),
	.w3(32'hbbcd8c4b),
	.w4(32'hb9f79edf),
	.w5(32'h3b0cb7af),
	.w6(32'hba9d589d),
	.w7(32'hba76c9aa),
	.w8(32'h3a11344a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa51410),
	.w1(32'h389f4a0d),
	.w2(32'hbbbdbd16),
	.w3(32'hba94494c),
	.w4(32'h3a72bdf6),
	.w5(32'hbad3fae3),
	.w6(32'h3a67f3f7),
	.w7(32'hbb807c6e),
	.w8(32'hbb74c2d5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9acf5b),
	.w1(32'h3b621d69),
	.w2(32'h3b663fb7),
	.w3(32'hbaaaa310),
	.w4(32'h3b758b79),
	.w5(32'h3b5114b0),
	.w6(32'h3aa8c911),
	.w7(32'h3ad3bb5a),
	.w8(32'h3b39658d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9d39),
	.w1(32'hbc28ca2e),
	.w2(32'h3af3b359),
	.w3(32'h3b9c38ff),
	.w4(32'hbc0653b0),
	.w5(32'h3a85018c),
	.w6(32'hba6b4404),
	.w7(32'h3c07c24c),
	.w8(32'h3c2907ac),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0149c2),
	.w1(32'hbb9734ef),
	.w2(32'hbbdb5b81),
	.w3(32'h3bf8a9cd),
	.w4(32'hbb0042ba),
	.w5(32'hbb8624b7),
	.w6(32'hba3631c9),
	.w7(32'hbb77462a),
	.w8(32'h3a940ba1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1f98),
	.w1(32'hbbb2e397),
	.w2(32'hbb46c796),
	.w3(32'h3a1ea4f0),
	.w4(32'hbace661c),
	.w5(32'hbb229926),
	.w6(32'h3b20ed79),
	.w7(32'hbae66b05),
	.w8(32'h3b3e3b7b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69cad5),
	.w1(32'h3b09049b),
	.w2(32'h3bce8ecd),
	.w3(32'hbb5e3bf9),
	.w4(32'hbb14d67a),
	.w5(32'hb9da58ab),
	.w6(32'h3a004df8),
	.w7(32'h3b56939a),
	.w8(32'h396ad449),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897ba7),
	.w1(32'h3adfd2ad),
	.w2(32'h39b50fe6),
	.w3(32'h3aee625e),
	.w4(32'h3b16681d),
	.w5(32'h3b1f9d44),
	.w6(32'h3be9122e),
	.w7(32'h3ba8907d),
	.w8(32'hba9f9849),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a98a),
	.w1(32'hbc61f768),
	.w2(32'hbc9e8252),
	.w3(32'hbb82314b),
	.w4(32'hbc0c219c),
	.w5(32'hbc7a1f61),
	.w6(32'hbbb5c8d7),
	.w7(32'hbc3ba002),
	.w8(32'hbbff82cb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dc2ee),
	.w1(32'h3a7a0830),
	.w2(32'h3c00d8fb),
	.w3(32'hbc62b011),
	.w4(32'h3bded33e),
	.w5(32'h3a9f8710),
	.w6(32'h3bfdf12b),
	.w7(32'h3b91834e),
	.w8(32'hbb0af38c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15fbf),
	.w1(32'h3b7c295e),
	.w2(32'h3c020ccf),
	.w3(32'h3bc58a5d),
	.w4(32'h3afa7da5),
	.w5(32'h3bc43023),
	.w6(32'h3aca5ecf),
	.w7(32'h3c021094),
	.w8(32'h3b5900f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0473e),
	.w1(32'h3a874d17),
	.w2(32'h3bee9a51),
	.w3(32'h3b5342e4),
	.w4(32'h395886fd),
	.w5(32'h3af4fbb5),
	.w6(32'hb81e2898),
	.w7(32'h3b9050a2),
	.w8(32'hbb48e34f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfc5a),
	.w1(32'hbac7027d),
	.w2(32'h3bf19ee5),
	.w3(32'hbbd3e873),
	.w4(32'hbb9df0bf),
	.w5(32'hba9739a1),
	.w6(32'hbbac1fe9),
	.w7(32'hbaea9b52),
	.w8(32'hbbaf72aa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac76885),
	.w1(32'h3aafc98f),
	.w2(32'hbaccc024),
	.w3(32'hbb7d8371),
	.w4(32'hbafeb5d6),
	.w5(32'h3a5646d6),
	.w6(32'h3a447e8a),
	.w7(32'hba9a06ed),
	.w8(32'h3b59d1e5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc10c03),
	.w1(32'h3b907f6d),
	.w2(32'h3d3b05cb),
	.w3(32'h3ad9e3dd),
	.w4(32'hbc0bd1b3),
	.w5(32'h3cbf2bcc),
	.w6(32'hbc982637),
	.w7(32'h3bb80aa8),
	.w8(32'hbc3d936d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87523f),
	.w1(32'hbb7e6e2a),
	.w2(32'h3b0ed352),
	.w3(32'hb910d733),
	.w4(32'hbaab0f12),
	.w5(32'h3bd382a4),
	.w6(32'hbb86779f),
	.w7(32'hbb40e4e3),
	.w8(32'hbaf628e8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fdff6),
	.w1(32'hbc169ddf),
	.w2(32'h3a74e7f8),
	.w3(32'h3b83ca92),
	.w4(32'hbbad9f53),
	.w5(32'h3a6f5a32),
	.w6(32'hbb674a79),
	.w7(32'hbba13361),
	.w8(32'h3ba42348),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291576),
	.w1(32'h3bafd992),
	.w2(32'h3b49206b),
	.w3(32'h3b708561),
	.w4(32'h3aa6e73d),
	.w5(32'hbb8ec88a),
	.w6(32'hbae1c875),
	.w7(32'h3b48dc30),
	.w8(32'h3a9ca1e4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85d4ba),
	.w1(32'hba40808d),
	.w2(32'hbc54cfc6),
	.w3(32'hba8a7ac0),
	.w4(32'hbb198370),
	.w5(32'hbb4fd739),
	.w6(32'h3b24e75b),
	.w7(32'hbbb6fddc),
	.w8(32'h3abb3746),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242eff),
	.w1(32'h3b7ef081),
	.w2(32'hbbb55af0),
	.w3(32'h3b291a50),
	.w4(32'h3ae5d131),
	.w5(32'hbbdfc3c1),
	.w6(32'h3b231448),
	.w7(32'hbc0962ec),
	.w8(32'hbc213265),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bad6c),
	.w1(32'h3c45cf44),
	.w2(32'h3c7e03cb),
	.w3(32'hbc161110),
	.w4(32'h3c33edfe),
	.w5(32'h3c664aef),
	.w6(32'h3c3099b1),
	.w7(32'h3c59aacc),
	.w8(32'h3c48158a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e6e16),
	.w1(32'h3b89a46c),
	.w2(32'h398e3315),
	.w3(32'h3c574504),
	.w4(32'hba993d7f),
	.w5(32'h3b785b53),
	.w6(32'h3bf9a507),
	.w7(32'h3b4ba9a8),
	.w8(32'h39965f64),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf37418),
	.w1(32'h3b631ec6),
	.w2(32'hbb3a446a),
	.w3(32'h3b0f8437),
	.w4(32'hba503a28),
	.w5(32'hba3891c1),
	.w6(32'h3be6e175),
	.w7(32'h3a12227e),
	.w8(32'h3b201c7c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf76a3),
	.w1(32'hba8a3cfa),
	.w2(32'hbbd2efd1),
	.w3(32'h3ab0baab),
	.w4(32'h3a51dbe4),
	.w5(32'hbbabf420),
	.w6(32'h39da36bf),
	.w7(32'hbbbec3ee),
	.w8(32'hbc0a7052),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170356),
	.w1(32'hbbb9a955),
	.w2(32'hbc60d2a9),
	.w3(32'hbbda8cb9),
	.w4(32'hbba5a33e),
	.w5(32'hbc4c381e),
	.w6(32'h3b57f82c),
	.w7(32'hbb0aec60),
	.w8(32'hbb0e5f2e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81e514),
	.w1(32'hbc2719f9),
	.w2(32'hbc567595),
	.w3(32'hbc6eb470),
	.w4(32'hbc1c1d8c),
	.w5(32'hbc736670),
	.w6(32'hbc0ab48e),
	.w7(32'hbc372db9),
	.w8(32'hbc185471),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc208a28),
	.w1(32'h3bd40eb8),
	.w2(32'h3c170be2),
	.w3(32'hbc246010),
	.w4(32'h3c4326b2),
	.w5(32'h3c493b44),
	.w6(32'h3c15f4e3),
	.w7(32'h3bfb8d47),
	.w8(32'h3bfe956d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021a5d),
	.w1(32'hb950aeaa),
	.w2(32'hbac7051d),
	.w3(32'h3c52c49a),
	.w4(32'hbbbb45aa),
	.w5(32'h3a2750bb),
	.w6(32'h3aa2df4b),
	.w7(32'hbbd45926),
	.w8(32'hbb7ee5c5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fbfd0),
	.w1(32'h3c0f0aba),
	.w2(32'h3b329a1d),
	.w3(32'hbb93a4fa),
	.w4(32'hba14ff0d),
	.w5(32'h3ae19bac),
	.w6(32'h3b08d46d),
	.w7(32'h3ba42236),
	.w8(32'h3aedf747),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6cfb6),
	.w1(32'hbbd8dd98),
	.w2(32'hbb55f6dc),
	.w3(32'h3b4970ee),
	.w4(32'hbbd02053),
	.w5(32'hbb7b27d6),
	.w6(32'h3929f268),
	.w7(32'hb96d9964),
	.w8(32'hbb5ef4cf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c9f0),
	.w1(32'h3bbfb838),
	.w2(32'h3b50551b),
	.w3(32'hbc0c5774),
	.w4(32'h3bc7d0ec),
	.w5(32'h3aab91b8),
	.w6(32'h3b99aab0),
	.w7(32'h3b5fc220),
	.w8(32'hbae7e51d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819817),
	.w1(32'h398e5aad),
	.w2(32'hbb269b5d),
	.w3(32'h3bef41fe),
	.w4(32'hbbe8c804),
	.w5(32'hbb4ce3ce),
	.w6(32'hbb6300f9),
	.w7(32'hb9ea9ead),
	.w8(32'hbbda5718),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1e31),
	.w1(32'hbc54e80d),
	.w2(32'hbc55bfac),
	.w3(32'h393f6482),
	.w4(32'hbc5af31c),
	.w5(32'hbc281ff1),
	.w6(32'hbbf978bc),
	.w7(32'hbbb63c61),
	.w8(32'h3a515198),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5af004),
	.w1(32'hba16ade0),
	.w2(32'hb830ed66),
	.w3(32'hbb13c3ba),
	.w4(32'hbb060709),
	.w5(32'hbbb65cd9),
	.w6(32'h3a4f9a48),
	.w7(32'hbb83a788),
	.w8(32'h3b0661e3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a454d8),
	.w1(32'h3b393fc4),
	.w2(32'h3bd2b7c5),
	.w3(32'hbbc612b1),
	.w4(32'hb9f3ac18),
	.w5(32'hbb02f1e7),
	.w6(32'h3ba785a7),
	.w7(32'h3b325505),
	.w8(32'h3bcb5d29),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b373ebd),
	.w1(32'h3b843078),
	.w2(32'hbbd02494),
	.w3(32'h3a240123),
	.w4(32'hbb008362),
	.w5(32'hbbe7a900),
	.w6(32'h3b059136),
	.w7(32'hbc04ba69),
	.w8(32'h3aba0642),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89bf132),
	.w1(32'hbbcb6b28),
	.w2(32'hbb6f840e),
	.w3(32'hbb72bb0d),
	.w4(32'hbc131cdb),
	.w5(32'hbb188cd0),
	.w6(32'hbc3ee623),
	.w7(32'hbbc6c434),
	.w8(32'hbbf3c819),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06718),
	.w1(32'h39105c9e),
	.w2(32'hbb08c5aa),
	.w3(32'hbae3a9f2),
	.w4(32'hba218957),
	.w5(32'hbbf69a50),
	.w6(32'hbbb71f34),
	.w7(32'hbbf96571),
	.w8(32'hbb26f913),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7df581),
	.w1(32'h3b04ff5a),
	.w2(32'h3a42a938),
	.w3(32'h3bcccc92),
	.w4(32'hbb13a41f),
	.w5(32'h3b1400c9),
	.w6(32'h3a28b590),
	.w7(32'h3ab47bca),
	.w8(32'hbaa866e7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f2817),
	.w1(32'h3b745da1),
	.w2(32'hbb25a9d6),
	.w3(32'hbb7974f7),
	.w4(32'h3b118912),
	.w5(32'hba244a92),
	.w6(32'h3b08eb87),
	.w7(32'hba9b89d9),
	.w8(32'hbb96e638),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3ba12),
	.w1(32'hbaa182fc),
	.w2(32'hbb3f5be7),
	.w3(32'hbbcac3f2),
	.w4(32'h39cce8a8),
	.w5(32'h3ac00843),
	.w6(32'h3b490f0f),
	.w7(32'h3bac99f1),
	.w8(32'h3bf03595),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005c71),
	.w1(32'h3b512c43),
	.w2(32'h3b5ff871),
	.w3(32'hba2cde12),
	.w4(32'h3ae6bf9f),
	.w5(32'hbb3acef7),
	.w6(32'h3b2ed690),
	.w7(32'h3b37a1d9),
	.w8(32'h39c02bdc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b99d1),
	.w1(32'hbaab8a65),
	.w2(32'hb9bf8010),
	.w3(32'h3b5e2fbe),
	.w4(32'hbbca93ab),
	.w5(32'hb99cf4ce),
	.w6(32'hbae88f6b),
	.w7(32'hbb8170cb),
	.w8(32'hbabc6fdd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891448),
	.w1(32'h3b06fd94),
	.w2(32'h3bbd0392),
	.w3(32'hbae0c655),
	.w4(32'h39fc56c2),
	.w5(32'h3b388953),
	.w6(32'h3b63d94b),
	.w7(32'h3abe4494),
	.w8(32'hbae8f1cd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a1e0e),
	.w1(32'hbac65395),
	.w2(32'hbadfd533),
	.w3(32'h3bbfbf6c),
	.w4(32'hbb3f003a),
	.w5(32'h3a3a0ab6),
	.w6(32'hbb7caec0),
	.w7(32'hbb2dfd03),
	.w8(32'h3ab745eb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65fccb),
	.w1(32'hba1c88af),
	.w2(32'hbb37378d),
	.w3(32'h3b16b431),
	.w4(32'hb8b49c52),
	.w5(32'hba80eee0),
	.w6(32'hbb5570ea),
	.w7(32'hbbc65c82),
	.w8(32'hbb00b7a4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d80e),
	.w1(32'h3b7a2d27),
	.w2(32'h3c1f6ee3),
	.w3(32'h3bde8a77),
	.w4(32'hbb1d5b2f),
	.w5(32'hba102f66),
	.w6(32'h3a11cb37),
	.w7(32'h3b5c16c0),
	.w8(32'hbad0e43f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9439dcf),
	.w1(32'h39971d72),
	.w2(32'h3bbab4b6),
	.w3(32'hba584996),
	.w4(32'h3a355b04),
	.w5(32'hb9c727d9),
	.w6(32'hbb431ed5),
	.w7(32'h3bcb0c1a),
	.w8(32'h3bcfc4a3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f312b),
	.w1(32'h3ba6adba),
	.w2(32'h3b8ed1d3),
	.w3(32'h3a982f05),
	.w4(32'h39846d0c),
	.w5(32'h3b36448b),
	.w6(32'h3bfc4b87),
	.w7(32'h3c15a271),
	.w8(32'h3c046a2b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9bcbe),
	.w1(32'h3af83b61),
	.w2(32'h3a74e593),
	.w3(32'h3b0af9c6),
	.w4(32'h3c41e95c),
	.w5(32'h3c1dff9c),
	.w6(32'hbb79a808),
	.w7(32'hbbfea4ce),
	.w8(32'hbbe34768),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d81899),
	.w1(32'hbad998e9),
	.w2(32'hbb80ac9f),
	.w3(32'h3bb7642c),
	.w4(32'hbbc5c463),
	.w5(32'hbbdfb7de),
	.w6(32'h3bc4cd52),
	.w7(32'h3bb2d218),
	.w8(32'h3b9aa0aa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba73f1e),
	.w1(32'hbad0e5cf),
	.w2(32'h39b2541d),
	.w3(32'hbc068ad1),
	.w4(32'hba957c9e),
	.w5(32'hbb25d57d),
	.w6(32'h3a9dffb3),
	.w7(32'hba10a5f7),
	.w8(32'hbb907657),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf15db9),
	.w1(32'hbb3a087a),
	.w2(32'hbadcd55f),
	.w3(32'hba4864af),
	.w4(32'h3a2d0ede),
	.w5(32'hbb44f695),
	.w6(32'h3a194ceb),
	.w7(32'hbb51b02b),
	.w8(32'hbb388727),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6fcaf),
	.w1(32'hbb9667f9),
	.w2(32'hbb170183),
	.w3(32'hba286493),
	.w4(32'h3ba19fb3),
	.w5(32'h3a2bf36d),
	.w6(32'hb997a670),
	.w7(32'h3a7072bc),
	.w8(32'hbb2ffd08),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2777c8),
	.w1(32'hbae9f4f6),
	.w2(32'h3bfba68c),
	.w3(32'h3aeea4cb),
	.w4(32'hbaea4e44),
	.w5(32'h3be44fe6),
	.w6(32'hbc099884),
	.w7(32'hba900e88),
	.w8(32'h3909f5f6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08a60d),
	.w1(32'h3ca2c250),
	.w2(32'h3d14bc37),
	.w3(32'h3bfc1d68),
	.w4(32'h3c774797),
	.w5(32'h3cf10f5d),
	.w6(32'h3bfa7a08),
	.w7(32'h3ca80600),
	.w8(32'h3c653a5b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3a213),
	.w1(32'hbae3648d),
	.w2(32'hbacc8fc8),
	.w3(32'h3cae6b69),
	.w4(32'hbb3ce3cc),
	.w5(32'h3b64245d),
	.w6(32'hba826ed6),
	.w7(32'h3b894ce2),
	.w8(32'hba1efff7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8df1f),
	.w1(32'h3be603c3),
	.w2(32'h3b33b127),
	.w3(32'hbb70c2cd),
	.w4(32'h3bc4eaf0),
	.w5(32'h3ab4bce2),
	.w6(32'h3c3602b1),
	.w7(32'h3ba0247d),
	.w8(32'h3b87f7f8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba491b68),
	.w1(32'hbadbee4d),
	.w2(32'h3af16396),
	.w3(32'hbb5076dc),
	.w4(32'hb9e78e83),
	.w5(32'hbbd71fef),
	.w6(32'h3a07a970),
	.w7(32'hb9a03ebe),
	.w8(32'hbbb3307b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadd1ff),
	.w1(32'hb931d170),
	.w2(32'hbbc4d402),
	.w3(32'h3c285a1c),
	.w4(32'h3a0b7b7a),
	.w5(32'hbb8a2246),
	.w6(32'hbb7fec57),
	.w7(32'hbb7198ba),
	.w8(32'hbb351d4e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7c943),
	.w1(32'h38f513b8),
	.w2(32'hbacb04aa),
	.w3(32'hbad0043b),
	.w4(32'h3ac10fa8),
	.w5(32'hbba46f52),
	.w6(32'h3b861480),
	.w7(32'hbb4442ee),
	.w8(32'hba93d1dd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01f54c),
	.w1(32'hbb3a97aa),
	.w2(32'h3a1a74d7),
	.w3(32'hbb284311),
	.w4(32'h3a8eaa39),
	.w5(32'hbae9a2e3),
	.w6(32'hbaacddcb),
	.w7(32'h3a19cbe7),
	.w8(32'h3a8ea7de),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dfd5),
	.w1(32'h3bb0f314),
	.w2(32'hba075235),
	.w3(32'hbafe274f),
	.w4(32'h3b114d6a),
	.w5(32'h3ba96ed2),
	.w6(32'h3a6de459),
	.w7(32'h3b9fd60c),
	.w8(32'hbb05c922),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab149d9),
	.w1(32'h3bc2f6d2),
	.w2(32'h3b7b95a7),
	.w3(32'hba8f14c4),
	.w4(32'h3afbe35e),
	.w5(32'hbb8002c1),
	.w6(32'h3b7f308d),
	.w7(32'h3b658e29),
	.w8(32'hba83d9d3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e374ff),
	.w1(32'h3b6ea42d),
	.w2(32'h3c1e9b37),
	.w3(32'hbbbf60ff),
	.w4(32'h3bb99337),
	.w5(32'h3bccd36d),
	.w6(32'h3a81be07),
	.w7(32'h3b9a0867),
	.w8(32'h3b097dce),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dbd82),
	.w1(32'hbba67652),
	.w2(32'hbbc8bf51),
	.w3(32'h3b535127),
	.w4(32'hbc01e4c8),
	.w5(32'hbb31a0fc),
	.w6(32'h3bc23120),
	.w7(32'h3a963bb8),
	.w8(32'h3b680d28),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a162116),
	.w1(32'h393decd4),
	.w2(32'h3a2f676a),
	.w3(32'hbb0fcc76),
	.w4(32'hbabdc14a),
	.w5(32'h3a3b56ac),
	.w6(32'hbb24632c),
	.w7(32'h3a4338a5),
	.w8(32'hbbcb4b33),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865e50),
	.w1(32'h3c2c6f6a),
	.w2(32'h3c29d2c1),
	.w3(32'hba0b5471),
	.w4(32'h3c83ea3e),
	.w5(32'h3c8b75cc),
	.w6(32'h3c887172),
	.w7(32'h3c4bc860),
	.w8(32'h3c24bfa9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be85dbe),
	.w1(32'h3842bc98),
	.w2(32'hbaef96cb),
	.w3(32'h3c5f7eab),
	.w4(32'hb9c5792d),
	.w5(32'hbb1838f7),
	.w6(32'h3b891ca8),
	.w7(32'h3bf99897),
	.w8(32'h3bc7f0ea),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fe8a),
	.w1(32'h39e73431),
	.w2(32'hbb3c76bc),
	.w3(32'hba6c74e7),
	.w4(32'h3b9ff420),
	.w5(32'hbb06c25e),
	.w6(32'hbb31f54b),
	.w7(32'hbc38bc3e),
	.w8(32'hbbf0c660),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38706f),
	.w1(32'h3bb7ee17),
	.w2(32'h3b90efd0),
	.w3(32'h399f5363),
	.w4(32'h3c197f33),
	.w5(32'h3c1a45d4),
	.w6(32'h3be4e0f0),
	.w7(32'h3b9a4ae4),
	.w8(32'h3beb42b0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baac3fd),
	.w1(32'h3cf2a55c),
	.w2(32'h3d67befd),
	.w3(32'h3c0108b2),
	.w4(32'h3ca813e4),
	.w5(32'h3d2a8a96),
	.w6(32'h3c3fbc43),
	.w7(32'h3cf93084),
	.w8(32'h3ca6708e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d26e450),
	.w1(32'h3ba44938),
	.w2(32'h3aef2749),
	.w3(32'h3cf1b649),
	.w4(32'h3b84b2b8),
	.w5(32'h3a3cf78e),
	.w6(32'h3a11989e),
	.w7(32'hbbb4f989),
	.w8(32'h3b62c5a3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced8bc),
	.w1(32'hbb146097),
	.w2(32'hbbbdeb83),
	.w3(32'h3b770729),
	.w4(32'hba35f1a1),
	.w5(32'hbb966758),
	.w6(32'h3a90e2ab),
	.w7(32'hba0942f9),
	.w8(32'hbac7d7e2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6d119),
	.w1(32'hbbe1e7c0),
	.w2(32'hbc4dd4d5),
	.w3(32'hbbbe0995),
	.w4(32'hbc16a918),
	.w5(32'hbc5057b6),
	.w6(32'hbbe52fd6),
	.w7(32'hbc14d637),
	.w8(32'hbb0890cb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8e8de),
	.w1(32'h3b11b1ef),
	.w2(32'h3b026c76),
	.w3(32'hbc420534),
	.w4(32'h3b418a8e),
	.w5(32'h3b45a75e),
	.w6(32'h3a313732),
	.w7(32'h3c01f759),
	.w8(32'h3b59292f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba595f4),
	.w1(32'hbb73ddab),
	.w2(32'hbbb46da4),
	.w3(32'h3a0a0d01),
	.w4(32'hbc2bf962),
	.w5(32'hbc0b71a9),
	.w6(32'h3a62411d),
	.w7(32'h3b4eb934),
	.w8(32'h3c0ab542),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6323d3),
	.w1(32'h3ca31855),
	.w2(32'h3d1f2998),
	.w3(32'hbba04b15),
	.w4(32'h3c6e3cda),
	.w5(32'h3cf022f1),
	.w6(32'h3bf288fc),
	.w7(32'h3ca02088),
	.w8(32'h3c54e8f0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4c1c4),
	.w1(32'h3b459214),
	.w2(32'h3ac5a60b),
	.w3(32'h3caac332),
	.w4(32'hba2fa84b),
	.w5(32'hbb587907),
	.w6(32'h3b585681),
	.w7(32'h3bc65125),
	.w8(32'h3b7a46ca),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad6e56),
	.w1(32'hbbccab26),
	.w2(32'hbc08bf35),
	.w3(32'hbb87fc20),
	.w4(32'hbb91e2f0),
	.w5(32'hbbc2df8e),
	.w6(32'hbbdc755d),
	.w7(32'hbc2d0372),
	.w8(32'hbc115b7d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d57a5),
	.w1(32'h3b331e7e),
	.w2(32'h3a7e21a8),
	.w3(32'hbb8ec870),
	.w4(32'h3b59b40b),
	.w5(32'h3aefbb3f),
	.w6(32'h3aacd8ed),
	.w7(32'h3be63e36),
	.w8(32'hbadcd289),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2545b3),
	.w1(32'hbad543b4),
	.w2(32'hbb216425),
	.w3(32'h3b9d5d78),
	.w4(32'hbb4533a9),
	.w5(32'hba4fa028),
	.w6(32'hba53dc09),
	.w7(32'hba6aef7e),
	.w8(32'hbb59c3c2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6da35),
	.w1(32'hbb2bb872),
	.w2(32'h3b5ba7ad),
	.w3(32'hbb28a606),
	.w4(32'hb80fbcd8),
	.w5(32'h3b268463),
	.w6(32'h3bafb244),
	.w7(32'hb97a44c6),
	.w8(32'hbad4295a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cec4c),
	.w1(32'h3a17dc29),
	.w2(32'hbb8a3d38),
	.w3(32'h3b732934),
	.w4(32'hbab2cab3),
	.w5(32'hbb84ada9),
	.w6(32'hb921db9d),
	.w7(32'h3b53678a),
	.w8(32'hbaad696e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969bb16),
	.w1(32'h3c322022),
	.w2(32'h3d10c06f),
	.w3(32'hbae96f94),
	.w4(32'h3ae24ec1),
	.w5(32'h3cb1a1df),
	.w6(32'hbc06a93f),
	.w7(32'h3c09fd38),
	.w8(32'h3a58a969),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc05c0e),
	.w1(32'h3ad8a925),
	.w2(32'hbb8b8955),
	.w3(32'h3c362e47),
	.w4(32'h3a95c61d),
	.w5(32'hbb857e47),
	.w6(32'hba1c6341),
	.w7(32'hbba90dd0),
	.w8(32'hbbe4770e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaf7a7),
	.w1(32'hbb4852c3),
	.w2(32'hbb9ccb4e),
	.w3(32'hbb9880b2),
	.w4(32'hbb6fcf7e),
	.w5(32'h3b591ddf),
	.w6(32'hba1189d5),
	.w7(32'h3b6edf30),
	.w8(32'h3ad8d30b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1b837),
	.w1(32'hb9c8b286),
	.w2(32'h39dd7b5f),
	.w3(32'h3aba7e30),
	.w4(32'hbae8570a),
	.w5(32'h3c0792af),
	.w6(32'hba394064),
	.w7(32'hb6ff9d5d),
	.w8(32'h3a95162a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99346dc),
	.w1(32'h39ab7a7b),
	.w2(32'hbb9c8a5b),
	.w3(32'h3b2851c9),
	.w4(32'h3a8ff87e),
	.w5(32'hbafd4637),
	.w6(32'h3ac1f846),
	.w7(32'hb99b344f),
	.w8(32'h39b0acb7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1baf7),
	.w1(32'hbbca6bb1),
	.w2(32'hb95cd0e5),
	.w3(32'h3a3534dc),
	.w4(32'hbbafe437),
	.w5(32'h3b0c7b8f),
	.w6(32'hbb45f07e),
	.w7(32'h391cd993),
	.w8(32'h3be5ac7c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule