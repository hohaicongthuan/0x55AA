module layer_10_featuremap_0(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2496c1),
	.w1(32'hbb98451f),
	.w2(32'hbbec119d),
	.w3(32'hbbdbecd9),
	.w4(32'h3a98f310),
	.w5(32'h3ae6a0d1),
	.w6(32'hbc0777b5),
	.w7(32'h3a1dbe99),
	.w8(32'h3b7ab3f0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b8519),
	.w1(32'hbbc0f9ee),
	.w2(32'hbc073d4a),
	.w3(32'h3bf5b85f),
	.w4(32'h3bec7d34),
	.w5(32'hbc123922),
	.w6(32'h3c71463b),
	.w7(32'h3c33c010),
	.w8(32'hbb98696a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89736d),
	.w1(32'h3b0d8dd5),
	.w2(32'h3c0932f6),
	.w3(32'hba8e84d7),
	.w4(32'hbaa024fd),
	.w5(32'hbb0df89f),
	.w6(32'hbb328488),
	.w7(32'hbba92ec1),
	.w8(32'hb9a01786),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc37a0),
	.w1(32'h3bad2162),
	.w2(32'h3c46c935),
	.w3(32'hbacdedfc),
	.w4(32'h3afdefa0),
	.w5(32'h3c1c831c),
	.w6(32'hbbbc35e9),
	.w7(32'hbad92c23),
	.w8(32'hba1d438c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773e23),
	.w1(32'hbc6db2a4),
	.w2(32'h390aec6d),
	.w3(32'hbb80e893),
	.w4(32'h3a2f98ee),
	.w5(32'h3c1e94d9),
	.w6(32'hbba166c5),
	.w7(32'h3a951d4c),
	.w8(32'h3bfa79d2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04005b),
	.w1(32'h3ba7f90d),
	.w2(32'h3b7910b8),
	.w3(32'h3c6f8d20),
	.w4(32'h3c33d101),
	.w5(32'h3b79a95e),
	.w6(32'h3c066a6d),
	.w7(32'h3c4d821b),
	.w8(32'h3b5d9275),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c7f45),
	.w1(32'hbc83c1ae),
	.w2(32'hbae62e73),
	.w3(32'hbc19a417),
	.w4(32'hbcbcb1e9),
	.w5(32'hbcb5d484),
	.w6(32'hbb99b7d0),
	.w7(32'hbc98a986),
	.w8(32'hbcd8c7ec),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b94f6),
	.w1(32'hbc519174),
	.w2(32'h3beb9895),
	.w3(32'hbd3a452f),
	.w4(32'hbc955a59),
	.w5(32'hbc2f296b),
	.w6(32'hbd4f4c21),
	.w7(32'hbbd23965),
	.w8(32'hbbb74974),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e01c4),
	.w1(32'h3b413ebf),
	.w2(32'h3c24315f),
	.w3(32'hbc44ac7f),
	.w4(32'h3aecd80f),
	.w5(32'h3b9ef0fc),
	.w6(32'hbbd0d935),
	.w7(32'hbacdf427),
	.w8(32'h3b6b77b5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273a2f),
	.w1(32'h3b87b0cd),
	.w2(32'hb93295c8),
	.w3(32'hbc28531e),
	.w4(32'hbb0adacf),
	.w5(32'h3c3c8e36),
	.w6(32'hbc28519d),
	.w7(32'h3bd51f9c),
	.w8(32'h3c6b595f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37470fb0),
	.w1(32'hbbf29ae4),
	.w2(32'hbb436fc7),
	.w3(32'hbaa6b805),
	.w4(32'hbc350c67),
	.w5(32'h3b6ba303),
	.w6(32'hba159236),
	.w7(32'hbc012725),
	.w8(32'h3b3b3f3e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1471f9),
	.w1(32'hbb494163),
	.w2(32'h3c870f15),
	.w3(32'hbba4559d),
	.w4(32'h3bf06e32),
	.w5(32'h3c047b1b),
	.w6(32'hbc156475),
	.w7(32'hbc24fdf4),
	.w8(32'hba8d0edd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb31b8e),
	.w1(32'h3a752adc),
	.w2(32'hbbd9a159),
	.w3(32'hbccc04ef),
	.w4(32'hb79e7a80),
	.w5(32'h3c2b32b6),
	.w6(32'hbc564263),
	.w7(32'h3bffd7be),
	.w8(32'h3c856fb8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bba09),
	.w1(32'hbb746eeb),
	.w2(32'hbc89462a),
	.w3(32'hbb98f9b8),
	.w4(32'hb9ad8119),
	.w5(32'hbb205a35),
	.w6(32'hbb58342e),
	.w7(32'hba316ec2),
	.w8(32'h3c1fe30a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edb94d),
	.w1(32'h3c1a7aa1),
	.w2(32'hbb22a70e),
	.w3(32'hbb8240e6),
	.w4(32'hbbd26d57),
	.w5(32'h3b18915f),
	.w6(32'h3c0d5f55),
	.w7(32'hbbb91573),
	.w8(32'hbb8e7e54),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad958b),
	.w1(32'h3ccc564a),
	.w2(32'h3b099879),
	.w3(32'hbbb9655f),
	.w4(32'h3d146eaa),
	.w5(32'h3c8d6445),
	.w6(32'hbb231649),
	.w7(32'h3d29fed2),
	.w8(32'h3ca323a0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab29df3),
	.w1(32'hbbddf275),
	.w2(32'h3ab85435),
	.w3(32'h39ab5f57),
	.w4(32'hbc259d25),
	.w5(32'hbb37b77e),
	.w6(32'h3a9a13b8),
	.w7(32'hbbfca815),
	.w8(32'hbc3d30e4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd02c2a8),
	.w1(32'h3bd3e621),
	.w2(32'h3c2c02a6),
	.w3(32'hbc4a2a83),
	.w4(32'h3d0a89e1),
	.w5(32'h3c144863),
	.w6(32'hbc53caff),
	.w7(32'h3d21e620),
	.w8(32'h3c95aaeb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc827948),
	.w1(32'h3b0792d5),
	.w2(32'hbc79c97f),
	.w3(32'hbc43ad30),
	.w4(32'h3c39f5a1),
	.w5(32'hbc470580),
	.w6(32'hbc08377f),
	.w7(32'h3c0ca47e),
	.w8(32'h3acf70b5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60ee59),
	.w1(32'hbc61efb9),
	.w2(32'hb9e6df3a),
	.w3(32'hbc7680b7),
	.w4(32'hbbf6ae41),
	.w5(32'hb94384b5),
	.w6(32'hbc3df0db),
	.w7(32'hbbf53044),
	.w8(32'hba79f1ce),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab83a46),
	.w1(32'h3c2d015e),
	.w2(32'h3b1bb95d),
	.w3(32'h3c31953b),
	.w4(32'h3caedc2b),
	.w5(32'hbbaafd47),
	.w6(32'h3babccc4),
	.w7(32'h3c49fa17),
	.w8(32'hbb0067a0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79d58c),
	.w1(32'hbbd0aad9),
	.w2(32'hbc2667bf),
	.w3(32'h3a6ecbf1),
	.w4(32'hbbe2e672),
	.w5(32'hbc47fd64),
	.w6(32'h3b671662),
	.w7(32'hbb59bcc3),
	.w8(32'hbc2ce488),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19779d),
	.w1(32'hba4fd673),
	.w2(32'h3c81d041),
	.w3(32'hbd4bfdb8),
	.w4(32'h3bb96945),
	.w5(32'h3caa0488),
	.w6(32'hbce0a041),
	.w7(32'h3c097ed0),
	.w8(32'h3ccf8c6a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af3c9),
	.w1(32'h3bb871e1),
	.w2(32'hbb087532),
	.w3(32'hbbc46942),
	.w4(32'h3bba016a),
	.w5(32'h3a1afa93),
	.w6(32'hbb00c18c),
	.w7(32'h3c651dfb),
	.w8(32'h3b853045),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051d5f),
	.w1(32'h3af8002b),
	.w2(32'hbcb98bf0),
	.w3(32'h3bf16f73),
	.w4(32'h3b927eb6),
	.w5(32'hbce8a073),
	.w6(32'h3bd7b8a7),
	.w7(32'h3c098163),
	.w8(32'hbccdedda),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0282),
	.w1(32'hbb52c708),
	.w2(32'hbb17fe51),
	.w3(32'hbc0b9b9d),
	.w4(32'hbb5ee7f9),
	.w5(32'hbb340558),
	.w6(32'hbac173d8),
	.w7(32'h39be21c4),
	.w8(32'hba8b1c3c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736361),
	.w1(32'hbb35379c),
	.w2(32'h39a4314d),
	.w3(32'h3aa332fd),
	.w4(32'h3ae31a5d),
	.w5(32'h3981b884),
	.w6(32'h3b26d17f),
	.w7(32'hbb63bd61),
	.w8(32'h3968200f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd43107),
	.w1(32'h3c4ee242),
	.w2(32'hbc5183fe),
	.w3(32'hbc9690b2),
	.w4(32'h3c08502d),
	.w5(32'h3aea01a3),
	.w6(32'hbc09f975),
	.w7(32'h3d05f62d),
	.w8(32'h3c37360f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cd37a),
	.w1(32'h3a7a435b),
	.w2(32'hb9d5a74b),
	.w3(32'hbb3c2019),
	.w4(32'h3aa7b91e),
	.w5(32'h3aa08b16),
	.w6(32'hbba97362),
	.w7(32'h39ecf81b),
	.w8(32'h3a8199c3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e5b19),
	.w1(32'h3c920469),
	.w2(32'hbc69f668),
	.w3(32'hbb7f2fb0),
	.w4(32'h3c0c881c),
	.w5(32'hbc9cf076),
	.w6(32'h3bc9db91),
	.w7(32'h3ca83990),
	.w8(32'hbc85ca66),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76c0fb),
	.w1(32'h39a2900a),
	.w2(32'hb8c1ec35),
	.w3(32'h3a80bc28),
	.w4(32'h3a3e69ee),
	.w5(32'hb9f92e02),
	.w6(32'h39c9de2c),
	.w7(32'h391190ab),
	.w8(32'hba56cff1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ddc353),
	.w1(32'h37b14ed2),
	.w2(32'hb9f1c236),
	.w3(32'hba89ddd2),
	.w4(32'h39848e99),
	.w5(32'hb9b5a819),
	.w6(32'hba761b43),
	.w7(32'hb9959205),
	.w8(32'hba3395a6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a7670),
	.w1(32'hba86cad2),
	.w2(32'hb9e17722),
	.w3(32'hbb9a8840),
	.w4(32'h3b93b2af),
	.w5(32'h3b89fbac),
	.w6(32'hbb7982b3),
	.w7(32'h3bcbcb06),
	.w8(32'h3bd89e7f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb689215f),
	.w1(32'h3b2e73d8),
	.w2(32'hbbceab0b),
	.w3(32'hb8d173cb),
	.w4(32'h3b7464e3),
	.w5(32'hbbb05ae5),
	.w6(32'h3a8890bd),
	.w7(32'h3b7b94bb),
	.w8(32'hbb40139d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba935666),
	.w1(32'h393935da),
	.w2(32'h3b5d3628),
	.w3(32'hb9c68ea0),
	.w4(32'h3a7acdc3),
	.w5(32'h3b801180),
	.w6(32'hbb382dde),
	.w7(32'hba6edbeb),
	.w8(32'h3ae403e5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec72c9),
	.w1(32'hbc1745e0),
	.w2(32'hbb8fba31),
	.w3(32'hbbdbb90e),
	.w4(32'hbc14e139),
	.w5(32'hba9b8489),
	.w6(32'hbbaec7da),
	.w7(32'hbb4db67b),
	.w8(32'h3b65c65e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8f13f),
	.w1(32'hbce2831b),
	.w2(32'hbc6c3ec8),
	.w3(32'hbcd0fef1),
	.w4(32'hbb997e22),
	.w5(32'h3cca2d2f),
	.w6(32'hbbc41bc2),
	.w7(32'hbaf00928),
	.w8(32'hbbb319db),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814dc8),
	.w1(32'h3b83457a),
	.w2(32'hbcd47d9e),
	.w3(32'hbb03bd65),
	.w4(32'hbac9c5cc),
	.w5(32'hbcf61fe0),
	.w6(32'h3a500671),
	.w7(32'hb8b3cd05),
	.w8(32'hbd05b036),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2e14),
	.w1(32'h3c3c68bc),
	.w2(32'hbc83df05),
	.w3(32'hbbcd2504),
	.w4(32'h3a9efeb2),
	.w5(32'hbd0726ab),
	.w6(32'hbb908310),
	.w7(32'h3bbab0b5),
	.w8(32'hbd1e147e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089435),
	.w1(32'hbb391918),
	.w2(32'hbb375b90),
	.w3(32'hbb6c9d15),
	.w4(32'hbb8c2ced),
	.w5(32'hbb4383c5),
	.w6(32'hbb9b7598),
	.w7(32'hbba2171b),
	.w8(32'hbbc5c428),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f15ff),
	.w1(32'h37e6e6d3),
	.w2(32'hb9c4345b),
	.w3(32'h3a28d225),
	.w4(32'h397e4813),
	.w5(32'hba9b2603),
	.w6(32'h3a1ee567),
	.w7(32'h3a0653bb),
	.w8(32'hba14c5d9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0013a),
	.w1(32'hb6e866e4),
	.w2(32'h39d8d91d),
	.w3(32'hb9ad14a4),
	.w4(32'hba3b40fb),
	.w5(32'h38ae8a1d),
	.w6(32'h3a199b47),
	.w7(32'h39261a5c),
	.w8(32'h39422007),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb835a3d),
	.w1(32'h3b27d0a9),
	.w2(32'h3a4084ef),
	.w3(32'hbb4cb21f),
	.w4(32'h3a990723),
	.w5(32'hbaa9de79),
	.w6(32'hbab4cca0),
	.w7(32'h3ad5c7d2),
	.w8(32'hbad365df),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2fc88a),
	.w1(32'h3c5d6f07),
	.w2(32'h3c4a3e14),
	.w3(32'hbd2b495c),
	.w4(32'h3c561d46),
	.w5(32'h3ca7c13f),
	.w6(32'hbce3a8d0),
	.w7(32'h3c8f15ba),
	.w8(32'h3cf794b7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a268bcd),
	.w1(32'h3c1e52a8),
	.w2(32'hbbc73fd4),
	.w3(32'hba6babff),
	.w4(32'h3c388ffe),
	.w5(32'hbaf526e5),
	.w6(32'h3b9223f7),
	.w7(32'h3c7a30bc),
	.w8(32'hb9867b2b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c7e7),
	.w1(32'h3b82bcea),
	.w2(32'hba107380),
	.w3(32'hbb191b82),
	.w4(32'h3c7d2104),
	.w5(32'h3bcf1cf9),
	.w6(32'hb88b188b),
	.w7(32'h3c8231d6),
	.w8(32'h3c2cb081),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5ce36),
	.w1(32'h3c134dc6),
	.w2(32'h3a85cc68),
	.w3(32'hbc0d6824),
	.w4(32'h3be925de),
	.w5(32'h3b043ee3),
	.w6(32'hbb8c5d0d),
	.w7(32'h3c286bff),
	.w8(32'h3b7994f8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceb0341),
	.w1(32'hbc2dae2e),
	.w2(32'h3bca7ba8),
	.w3(32'hbcc878df),
	.w4(32'hba842482),
	.w5(32'h3c7c11b3),
	.w6(32'hbcb8240b),
	.w7(32'h3c502b54),
	.w8(32'h3d09f5f6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9910f),
	.w1(32'h39327c7d),
	.w2(32'h369b03b1),
	.w3(32'hb9ab63e7),
	.w4(32'h398a2045),
	.w5(32'h3a688896),
	.w6(32'hb906cf84),
	.w7(32'h399d0b79),
	.w8(32'hba01355a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b833f),
	.w1(32'h3a4a53ea),
	.w2(32'h3b05d777),
	.w3(32'h3a2c34d2),
	.w4(32'h3a1ef76c),
	.w5(32'h3abbfce9),
	.w6(32'h396cc1b4),
	.w7(32'h3969a40a),
	.w8(32'h3a398fd1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5f690),
	.w1(32'h3a24ad50),
	.w2(32'h3ae152cf),
	.w3(32'h3b23f571),
	.w4(32'h3a8e3818),
	.w5(32'h39cdd425),
	.w6(32'h3b105355),
	.w7(32'h3aabdebd),
	.w8(32'h3a1783be),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55745e),
	.w1(32'hbae2db1e),
	.w2(32'hbb755741),
	.w3(32'hbc586e84),
	.w4(32'h3b85abf7),
	.w5(32'h3993b2ba),
	.w6(32'hbb4a1d1b),
	.w7(32'h3bc2ea1d),
	.w8(32'h3aa1b689),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03ab0),
	.w1(32'hba0ceb5b),
	.w2(32'hba9052e6),
	.w3(32'hbb42a422),
	.w4(32'h3b40728c),
	.w5(32'h3a1532e1),
	.w6(32'hbb5e88c9),
	.w7(32'h3b632303),
	.w8(32'h3b7e5aa9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd144b26),
	.w1(32'h39a32da9),
	.w2(32'h3c0d5789),
	.w3(32'hbcb3f52d),
	.w4(32'h3c7ed561),
	.w5(32'h3c89bd8a),
	.w6(32'hbca9cebd),
	.w7(32'h3ca588ba),
	.w8(32'h3d00f290),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07105d),
	.w1(32'h3bc91aa5),
	.w2(32'h3be7d20c),
	.w3(32'hbbd5181a),
	.w4(32'h3bc5e38a),
	.w5(32'h3bd6c50d),
	.w6(32'hbab22f25),
	.w7(32'h3c216c96),
	.w8(32'h3c0ea04d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93452ee),
	.w1(32'hb973f796),
	.w2(32'h383baa3b),
	.w3(32'hb908bdea),
	.w4(32'hba447fb2),
	.w5(32'h3977b6b5),
	.w6(32'hb99908b1),
	.w7(32'hb9c141eb),
	.w8(32'h39728882),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a863091),
	.w1(32'h3a6fbaa5),
	.w2(32'hb940af8b),
	.w3(32'h3ad17541),
	.w4(32'h3a772167),
	.w5(32'hba11479b),
	.w6(32'h3aa6b0b1),
	.w7(32'h3a88271a),
	.w8(32'hba3bd297),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac401a3),
	.w1(32'h3a0ae680),
	.w2(32'hba3b5814),
	.w3(32'hba3d9cab),
	.w4(32'hba5867b3),
	.w5(32'hbadcf75e),
	.w6(32'hba24d523),
	.w7(32'hba8a200b),
	.w8(32'hbac22398),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91d19e),
	.w1(32'h3ac0b6db),
	.w2(32'hb9dcbe1a),
	.w3(32'h3a44ae9e),
	.w4(32'h3a891904),
	.w5(32'hba592980),
	.w6(32'hba92724b),
	.w7(32'hb99f124c),
	.w8(32'hbab31ecd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7b052),
	.w1(32'h38959c63),
	.w2(32'hb95e2b9b),
	.w3(32'hbac1cc92),
	.w4(32'h39ff8c15),
	.w5(32'hb9b3abeb),
	.w6(32'hba869f1d),
	.w7(32'h3a68bc8b),
	.w8(32'h39e24a03),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94cfe2),
	.w1(32'hb88e089e),
	.w2(32'h3b8a203d),
	.w3(32'hbc8277af),
	.w4(32'h3b87c48f),
	.w5(32'h3bf6a30a),
	.w6(32'hbc3ba704),
	.w7(32'h3bf54651),
	.w8(32'h3c39254b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6a244),
	.w1(32'h3c411f24),
	.w2(32'h3c70be5a),
	.w3(32'hbcd2ac5e),
	.w4(32'h3c870efd),
	.w5(32'h3c8cb666),
	.w6(32'hbc423813),
	.w7(32'h3cb81504),
	.w8(32'h3c90000d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca5055),
	.w1(32'hbaaacbfb),
	.w2(32'hb9db8634),
	.w3(32'hbab91d6f),
	.w4(32'hba95dadf),
	.w5(32'hba5d7a32),
	.w6(32'hba9b78c2),
	.w7(32'hba9411d2),
	.w8(32'hb9af6564),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983213c),
	.w1(32'hb9a85cf5),
	.w2(32'h390a0592),
	.w3(32'hba114441),
	.w4(32'hba3b96e1),
	.w5(32'h3900822c),
	.w6(32'hb9508457),
	.w7(32'hba0a1a02),
	.w8(32'hba124a95),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6c6ab),
	.w1(32'h3a1f52f2),
	.w2(32'hba193081),
	.w3(32'h3a53e7d6),
	.w4(32'h3a17039c),
	.w5(32'hba03423c),
	.w6(32'hb909eba2),
	.w7(32'hb96ccf46),
	.w8(32'hba0482b2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be4e3d),
	.w1(32'hb9fad6b0),
	.w2(32'hba57bb7d),
	.w3(32'hb9f60487),
	.w4(32'hba6eaeee),
	.w5(32'hba9c4e99),
	.w6(32'hba18a615),
	.w7(32'hba4e504d),
	.w8(32'hba872ab2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd355e29),
	.w1(32'h3c14c814),
	.w2(32'h3cbc3c1e),
	.w3(32'hbd22fd87),
	.w4(32'h3c1e4bf8),
	.w5(32'h3cf24445),
	.w6(32'hbd179a70),
	.w7(32'h3bfa6dce),
	.w8(32'h3cc39398),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7d414),
	.w1(32'hbb54a375),
	.w2(32'hba851e49),
	.w3(32'hbc9054d1),
	.w4(32'h3c89c9a9),
	.w5(32'h3bb44882),
	.w6(32'hbca7dba2),
	.w7(32'h3c42cdbe),
	.w8(32'h3c7abc6b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf6d25a),
	.w1(32'h3c28acff),
	.w2(32'h3bd7b4e4),
	.w3(32'hbcef656a),
	.w4(32'h3caae259),
	.w5(32'h3c63dff7),
	.w6(32'hbc98b095),
	.w7(32'h3cbfcbb7),
	.w8(32'h3c98f1a9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c2221),
	.w1(32'h3c36a281),
	.w2(32'hbd023315),
	.w3(32'h3a4d0e26),
	.w4(32'h3c24e627),
	.w5(32'hbccef7d8),
	.w6(32'h3b26a966),
	.w7(32'h3c50495c),
	.w8(32'hbcddd1e8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385bf9d4),
	.w1(32'hba827b9a),
	.w2(32'hb903921d),
	.w3(32'hb92385a1),
	.w4(32'hba21bd84),
	.w5(32'hb97a551d),
	.w6(32'hb9bdb64b),
	.w7(32'hba655e50),
	.w8(32'hb934e04b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9468c48),
	.w1(32'hb9abe30e),
	.w2(32'h39b3fa45),
	.w3(32'hb78d0f24),
	.w4(32'hba0adf73),
	.w5(32'h372c4bd5),
	.w6(32'h386b68aa),
	.w7(32'hb9ff98ef),
	.w8(32'h3994b9b7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39013ae4),
	.w1(32'hb997e482),
	.w2(32'h3a785e34),
	.w3(32'hb96fd813),
	.w4(32'hba33f59c),
	.w5(32'h3a6294a6),
	.w6(32'h371d1ae2),
	.w7(32'hb97c5af4),
	.w8(32'h3abe5644),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02040f),
	.w1(32'h3b365249),
	.w2(32'h3b6c04af),
	.w3(32'hbbba6e7d),
	.w4(32'h3b8a9e53),
	.w5(32'h3b92803e),
	.w6(32'hbb960eca),
	.w7(32'h3bb79149),
	.w8(32'h3be68d22),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa010e3),
	.w1(32'h39e3470b),
	.w2(32'hb827f5b7),
	.w3(32'h3ac98804),
	.w4(32'h3a320512),
	.w5(32'hb8d9e9d5),
	.w6(32'h3ac39fc8),
	.w7(32'h3a41f412),
	.w8(32'h38501a97),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b4f4b),
	.w1(32'hbbdebe91),
	.w2(32'h3be173fc),
	.w3(32'hbc8cec7d),
	.w4(32'hbc649a28),
	.w5(32'h3c0af602),
	.w6(32'hbc6b7bd5),
	.w7(32'hbb7189a7),
	.w8(32'h3be99e5a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda5765),
	.w1(32'hbca4e384),
	.w2(32'h3b1cf192),
	.w3(32'hbcb0d2e8),
	.w4(32'hbc298c2c),
	.w5(32'h3c6fe7c0),
	.w6(32'hbcd03336),
	.w7(32'hbc169d14),
	.w8(32'h3cc6fc9d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aaa3d),
	.w1(32'h3b4ac977),
	.w2(32'hbc5caa12),
	.w3(32'hbb02675e),
	.w4(32'h3b79ed24),
	.w5(32'hbc00b494),
	.w6(32'h3bd8fad2),
	.w7(32'h3c105e8f),
	.w8(32'hbbc77c4b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc424205),
	.w1(32'h3bb07f9b),
	.w2(32'h3a6f7cd4),
	.w3(32'hbc028185),
	.w4(32'h3c2faa83),
	.w5(32'h3b8c96bd),
	.w6(32'hbbe91d36),
	.w7(32'h3c429f97),
	.w8(32'h3c00f942),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3485c9),
	.w1(32'hbbf61dc2),
	.w2(32'h3b862295),
	.w3(32'hbbfe2431),
	.w4(32'hbbf0a3bb),
	.w5(32'h3bf765ca),
	.w6(32'hbc21bd1a),
	.w7(32'hbbe0beaa),
	.w8(32'h3b91d245),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa00fc),
	.w1(32'h3c10e410),
	.w2(32'h389ff965),
	.w3(32'hbb8f0334),
	.w4(32'h3c18b497),
	.w5(32'h3b518395),
	.w6(32'hb94a00df),
	.w7(32'h3c20321a),
	.w8(32'h3bce2441),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc362ba0),
	.w1(32'hbb41acef),
	.w2(32'hb9ad2136),
	.w3(32'hbc21ef52),
	.w4(32'hbb418cad),
	.w5(32'h3b1d1b3d),
	.w6(32'hbbdd2fd0),
	.w7(32'h3b7f8d73),
	.w8(32'h3c189db4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1aafb),
	.w1(32'h39d1437a),
	.w2(32'h38dcd0b0),
	.w3(32'h3a99f53c),
	.w4(32'h3a0f7556),
	.w5(32'h3a2b1d3e),
	.w6(32'h3984c999),
	.w7(32'hb538fb94),
	.w8(32'hb9a155cc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919b6ae),
	.w1(32'hb9757199),
	.w2(32'h39c10aa1),
	.w3(32'h3a038af2),
	.w4(32'h3a1f125b),
	.w5(32'h3a95877e),
	.w6(32'hb98b6988),
	.w7(32'hb8c7facc),
	.w8(32'h3a6085fc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389283fe),
	.w1(32'h391773ef),
	.w2(32'h399b3083),
	.w3(32'h39f5fc18),
	.w4(32'h39e409b4),
	.w5(32'hb9147c84),
	.w6(32'h3997891f),
	.w7(32'h397e8b94),
	.w8(32'hb95eb454),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec11ee),
	.w1(32'hbaf2f681),
	.w2(32'hba61f3af),
	.w3(32'h3a6a104b),
	.w4(32'hbb212b5a),
	.w5(32'hbb2123c5),
	.w6(32'h3a862a4b),
	.w7(32'hbb25f667),
	.w8(32'hbb3c5a0e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e02ac),
	.w1(32'h3bc6619e),
	.w2(32'hbbb8be7a),
	.w3(32'hbc00e85e),
	.w4(32'h3afadeb7),
	.w5(32'hbbd2de4d),
	.w6(32'hba988380),
	.w7(32'h3bdc164a),
	.w8(32'hbc193598),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4f78b),
	.w1(32'h38f58d2e),
	.w2(32'h3abfb94a),
	.w3(32'h3a37227a),
	.w4(32'h3a2e8dff),
	.w5(32'h3b010d45),
	.w6(32'hb9f1dabd),
	.w7(32'hb8d56acd),
	.w8(32'h3a90a462),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a35d8),
	.w1(32'hba84a353),
	.w2(32'hbbe76eb7),
	.w3(32'hb8e75c8d),
	.w4(32'h3c20b0d7),
	.w5(32'hbbb2df97),
	.w6(32'hb9b3c016),
	.w7(32'h3b1ce53a),
	.w8(32'hbb786089),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc944fd3),
	.w1(32'h39288d2e),
	.w2(32'h3bfef08c),
	.w3(32'hbc987ad4),
	.w4(32'h39dbbc02),
	.w5(32'h3c2bce35),
	.w6(32'hbc72d21c),
	.w7(32'h3bc400cf),
	.w8(32'h3c934f4f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c409c1f),
	.w1(32'h3bd36ef8),
	.w2(32'hbc445ef4),
	.w3(32'h39ab9050),
	.w4(32'hb92f16e4),
	.w5(32'hbc89766c),
	.w6(32'h3bdb8622),
	.w7(32'h3b7f75f6),
	.w8(32'hbc8fac4f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd160fb1),
	.w1(32'hbca8e94a),
	.w2(32'h3c66d828),
	.w3(32'hbd0bdd5f),
	.w4(32'hbc1ef2bc),
	.w5(32'h3cb29604),
	.w6(32'hbca8833d),
	.w7(32'hbc8d789e),
	.w8(32'h3ccffd77),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55f9d1),
	.w1(32'h3aa49278),
	.w2(32'hba98eedf),
	.w3(32'h3c1793a3),
	.w4(32'hbb124098),
	.w5(32'hbac04ba8),
	.w6(32'h3bb50de5),
	.w7(32'h39c92adc),
	.w8(32'hbbcc41cc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdfda46),
	.w1(32'h3c560924),
	.w2(32'h3c20cf2c),
	.w3(32'hbc8a296a),
	.w4(32'h3cc13882),
	.w5(32'h3c9a18ac),
	.w6(32'hbc9a6e8d),
	.w7(32'h3cbe12cd),
	.w8(32'h3cdc4b4a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952ae3),
	.w1(32'h3b2a08c3),
	.w2(32'hbaf91b93),
	.w3(32'hbbbac45b),
	.w4(32'h3c33ba19),
	.w5(32'h3c17926f),
	.w6(32'hbb039501),
	.w7(32'h3b905e42),
	.w8(32'h3b56fbb8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1611),
	.w1(32'h3b807fc7),
	.w2(32'hbc78ad8b),
	.w3(32'hbb8f8a86),
	.w4(32'hbb4224d8),
	.w5(32'hbcad5a84),
	.w6(32'hbab50c64),
	.w7(32'hb96ae6da),
	.w8(32'hbc8aafc9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a212653),
	.w1(32'hba24fff8),
	.w2(32'h3a71ffd8),
	.w3(32'h395f383b),
	.w4(32'h396b05ac),
	.w5(32'h3ad01798),
	.w6(32'h398d3af3),
	.w7(32'h3a701097),
	.w8(32'h3a8f19c9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb19359),
	.w1(32'h3ba17acd),
	.w2(32'h3be47b09),
	.w3(32'hbc585291),
	.w4(32'h3c813e65),
	.w5(32'h3c3e75b8),
	.w6(32'hbc71a839),
	.w7(32'h3c80a74f),
	.w8(32'h3c74f2e2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc19f7b),
	.w1(32'h3b9d0d25),
	.w2(32'h3c97050e),
	.w3(32'hbcc2b369),
	.w4(32'h3b323fc4),
	.w5(32'h3ca5a0f3),
	.w6(32'hbc62ba37),
	.w7(32'h3b58d820),
	.w8(32'h3b9815ec),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce505fc),
	.w1(32'hbce976b5),
	.w2(32'hbcbbb146),
	.w3(32'hbd19d6a5),
	.w4(32'hbc91b8e4),
	.w5(32'h3cbed9f5),
	.w6(32'hbbd124d9),
	.w7(32'hbb4d10d3),
	.w8(32'h3cb820cd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4feddb),
	.w1(32'hbbc5a563),
	.w2(32'hbbe14401),
	.w3(32'hbcb7510f),
	.w4(32'hbc318d4f),
	.w5(32'hbc49cf4b),
	.w6(32'hbc3710f9),
	.w7(32'hbc2d7c09),
	.w8(32'hbc849622),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8330e2),
	.w1(32'h3bbdd564),
	.w2(32'hbc962241),
	.w3(32'hb9f09359),
	.w4(32'h3bd528e7),
	.w5(32'hbc50e0ae),
	.w6(32'h3adda649),
	.w7(32'h3c449c37),
	.w8(32'hbc3a2ab3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcece265),
	.w1(32'hbcc75a5d),
	.w2(32'h3c8d2a9c),
	.w3(32'hbcc36d9f),
	.w4(32'hbc041699),
	.w5(32'h3d0ecdd6),
	.w6(32'hbbbf62fb),
	.w7(32'hbc3719b8),
	.w8(32'h3d1441ce),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d484d),
	.w1(32'hb9c9e30b),
	.w2(32'hba380066),
	.w3(32'hbac78837),
	.w4(32'hb9332f0e),
	.w5(32'hba7b4b88),
	.w6(32'hbb02a5fd),
	.w7(32'hba0b8e34),
	.w8(32'hba376ecf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d3278),
	.w1(32'hbc9b4a03),
	.w2(32'hbcd5af83),
	.w3(32'hbd27e581),
	.w4(32'hbb7f94fd),
	.w5(32'h3c06e195),
	.w6(32'hbb7515b6),
	.w7(32'h3c77b1c3),
	.w8(32'hbcc0d4d7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa02c04),
	.w1(32'hbbb3cef4),
	.w2(32'h3bc3f018),
	.w3(32'hbc249e49),
	.w4(32'hb99f8cd7),
	.w5(32'hb94bebc4),
	.w6(32'hbabbfdb9),
	.w7(32'h3b7a43eb),
	.w8(32'hbc012766),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88171fb),
	.w1(32'hba871f73),
	.w2(32'hba8b8ce2),
	.w3(32'hb89a22cb),
	.w4(32'hba61bfdb),
	.w5(32'hba42ef29),
	.w6(32'hb8cebba8),
	.w7(32'hba852a19),
	.w8(32'hbac02320),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1bb6e),
	.w1(32'h3aeb5549),
	.w2(32'hbb440ae6),
	.w3(32'hbb04d0bd),
	.w4(32'h3af79a57),
	.w5(32'h3b01a68a),
	.w6(32'hba95b6e6),
	.w7(32'hb9d88ef6),
	.w8(32'h3b5dc344),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69c71b),
	.w1(32'hbaca58e8),
	.w2(32'hbb708972),
	.w3(32'hbc4571f7),
	.w4(32'hba010e9a),
	.w5(32'hbb38569f),
	.w6(32'hbc3274bf),
	.w7(32'h3b5195a7),
	.w8(32'h3b846812),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f28fc),
	.w1(32'h3ba37c68),
	.w2(32'hbc13b254),
	.w3(32'hbb63e2ea),
	.w4(32'h3b1621ea),
	.w5(32'hbc16c9dd),
	.w6(32'h3af6960e),
	.w7(32'h3c057ec4),
	.w8(32'hbbb16856),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ab0eb),
	.w1(32'hbad8faa8),
	.w2(32'hbbd2b711),
	.w3(32'hbb9653cd),
	.w4(32'hba315265),
	.w5(32'hbc4805b5),
	.w6(32'hb70c9d8c),
	.w7(32'h3bff83e8),
	.w8(32'hbc4e3172),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eb393),
	.w1(32'h3b7e5c98),
	.w2(32'hbbde5e05),
	.w3(32'hba58a15e),
	.w4(32'h3ba5ce8c),
	.w5(32'hbb7869ef),
	.w6(32'h3b24a11b),
	.w7(32'h3b9b0ecc),
	.w8(32'hbbe01ee5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c168),
	.w1(32'h3bddb6e4),
	.w2(32'h38381ec0),
	.w3(32'hb9bca613),
	.w4(32'h3c737f1f),
	.w5(32'h3bbaf238),
	.w6(32'hbc483236),
	.w7(32'h3c1e15a8),
	.w8(32'h3c3b85ec),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6a96d),
	.w1(32'h3c54f67e),
	.w2(32'hbab33317),
	.w3(32'hbc101278),
	.w4(32'h3c8beea8),
	.w5(32'h3ca10220),
	.w6(32'hbb8dc0e6),
	.w7(32'h3c724911),
	.w8(32'h3c956814),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b1239),
	.w1(32'h3b8681bd),
	.w2(32'hba09deba),
	.w3(32'hba9a1e6d),
	.w4(32'h3b5dafeb),
	.w5(32'hba2a2033),
	.w6(32'hb8d07286),
	.w7(32'h3bd1d5de),
	.w8(32'h39dc8335),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914acc6),
	.w1(32'h39056f0f),
	.w2(32'hbaf0212f),
	.w3(32'hb9b40865),
	.w4(32'hb83d340e),
	.w5(32'hbae7763c),
	.w6(32'hb97fbe16),
	.w7(32'hb9a686d2),
	.w8(32'hbac0b150),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6ea7),
	.w1(32'h3ad4f83c),
	.w2(32'hba5ba831),
	.w3(32'hbaf506b3),
	.w4(32'hba02330a),
	.w5(32'hb9f8fc9b),
	.w6(32'hbb1927ac),
	.w7(32'hba02de94),
	.w8(32'hb95bbb4c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d8fd8),
	.w1(32'h3a23b95c),
	.w2(32'hb9f937d5),
	.w3(32'hb9b699ab),
	.w4(32'h399b5c38),
	.w5(32'hb7db7d75),
	.w6(32'h3903867f),
	.w7(32'h39febe94),
	.w8(32'hb9ffc8f5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08c1b8),
	.w1(32'hb8801642),
	.w2(32'hb8bb5079),
	.w3(32'hb9f8508a),
	.w4(32'h3939a52d),
	.w5(32'h398596b1),
	.w6(32'hba620ec9),
	.w7(32'h3a0ed596),
	.w8(32'h39a76938),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba953a40),
	.w1(32'h3bcc73e4),
	.w2(32'hbab06a9c),
	.w3(32'hbad86385),
	.w4(32'h3c02b4aa),
	.w5(32'hb9eaf8b1),
	.w6(32'h399f309f),
	.w7(32'h3c1b0e24),
	.w8(32'h3a85b033),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8b44),
	.w1(32'hbacb77d8),
	.w2(32'hbacf03c4),
	.w3(32'hba19f7b0),
	.w4(32'hb9cce5c5),
	.w5(32'hba4c9f07),
	.w6(32'hb9748065),
	.w7(32'h398f2cbb),
	.w8(32'hb9c73f40),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc544226),
	.w1(32'hbb963436),
	.w2(32'h3b436387),
	.w3(32'hbc4e3fcd),
	.w4(32'hbbc62c28),
	.w5(32'h3b842cdc),
	.w6(32'hbc152df2),
	.w7(32'h39b2f187),
	.w8(32'h3c39074d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95c33),
	.w1(32'h3a95c4d6),
	.w2(32'hbc9a8128),
	.w3(32'hbaa4e96b),
	.w4(32'hbaf3cc96),
	.w5(32'hbc9b895a),
	.w6(32'h3b3bfb52),
	.w7(32'h3a056bad),
	.w8(32'hbca601b6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5e52),
	.w1(32'h3a1b92fc),
	.w2(32'h39ee65ea),
	.w3(32'h3aba35bf),
	.w4(32'h3a957109),
	.w5(32'h39df2d31),
	.w6(32'h39badf59),
	.w7(32'hb7b1f569),
	.w8(32'h38631767),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba6491),
	.w1(32'hb91fa205),
	.w2(32'hb91e01e4),
	.w3(32'h39501ea5),
	.w4(32'h39019bbb),
	.w5(32'h398f27c3),
	.w6(32'hb9d27edb),
	.w7(32'hba15db83),
	.w8(32'hba2ffb2b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92185e),
	.w1(32'h3a5f954b),
	.w2(32'hb97e4cbd),
	.w3(32'h39499bb6),
	.w4(32'h3946f710),
	.w5(32'hb8f217aa),
	.w6(32'hb9bc5e98),
	.w7(32'h3a2a9ffe),
	.w8(32'hb9d27a50),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1942dd),
	.w1(32'hba8555fb),
	.w2(32'hba2b70dd),
	.w3(32'hbb123a65),
	.w4(32'hb9d76062),
	.w5(32'hba4008f8),
	.w6(32'hbb55173a),
	.w7(32'hbb0ee75d),
	.w8(32'hbae42765),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca44d1e),
	.w1(32'hbccb43ec),
	.w2(32'h3b27f1d3),
	.w3(32'hbc11e156),
	.w4(32'hbb3824f4),
	.w5(32'h3c465363),
	.w6(32'hbcb36fe6),
	.w7(32'hbb50b035),
	.w8(32'h3c32df11),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7984b),
	.w1(32'h3b0b5f68),
	.w2(32'h3b9030c8),
	.w3(32'hbc456894),
	.w4(32'h3c6c3637),
	.w5(32'h3c31757f),
	.w6(32'hbc613a7b),
	.w7(32'h3c8e10df),
	.w8(32'h3c820ab8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb151f34),
	.w1(32'hb9576659),
	.w2(32'h3b183096),
	.w3(32'hbb196f1e),
	.w4(32'hba478bda),
	.w5(32'h3b22498c),
	.w6(32'hbadba928),
	.w7(32'h3ae58598),
	.w8(32'h3b83e527),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd666),
	.w1(32'h39ae2466),
	.w2(32'h3a0f8278),
	.w3(32'hbba2ea49),
	.w4(32'h3b3b6156),
	.w5(32'h3a16dcb0),
	.w6(32'hbbb5f5c5),
	.w7(32'h3adcdd56),
	.w8(32'h3b2b9207),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d321cb),
	.w1(32'h3ae92ca7),
	.w2(32'hba64403f),
	.w3(32'hba02b2b9),
	.w4(32'h3aa36ff0),
	.w5(32'hbb0bd043),
	.w6(32'h3b09442f),
	.w7(32'h3b7b5e7d),
	.w8(32'hba45304a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16a4aa),
	.w1(32'h3b9156dc),
	.w2(32'h3b6bdc19),
	.w3(32'hbc0cafc6),
	.w4(32'h3bd430ad),
	.w5(32'h3bb79118),
	.w6(32'hbbd83f83),
	.w7(32'h3c17b004),
	.w8(32'h3c16aac0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbd0f9),
	.w1(32'h3c58a615),
	.w2(32'hbb86c33d),
	.w3(32'h3a5ce2ee),
	.w4(32'h3c951afb),
	.w5(32'h3b8de519),
	.w6(32'h3b83363f),
	.w7(32'h3c77d8df),
	.w8(32'h3bc43176),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b90d4),
	.w1(32'hbbe258cc),
	.w2(32'h3c1aa3c1),
	.w3(32'hbcbf9e9a),
	.w4(32'h3b8f6868),
	.w5(32'h3c4cd4d1),
	.w6(32'hbc91edaf),
	.w7(32'h3bdcea93),
	.w8(32'h3c6cec5c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a0741),
	.w1(32'h39c1a9b5),
	.w2(32'hbc176ee2),
	.w3(32'hbb984c6e),
	.w4(32'hbb0b1ed0),
	.w5(32'hbc21da69),
	.w6(32'hba5dfe9d),
	.w7(32'hb9a10c91),
	.w8(32'hbc3725be),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8333a2),
	.w1(32'hbb4a4fd2),
	.w2(32'h3ad4f071),
	.w3(32'hbc5a3d82),
	.w4(32'h3baa6715),
	.w5(32'h3c36bb45),
	.w6(32'hbc280aff),
	.w7(32'hba9c3f20),
	.w8(32'h3bafeec0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1241f),
	.w1(32'hbb9c355c),
	.w2(32'h3bac857b),
	.w3(32'hbc9dfe75),
	.w4(32'h3b8ee3a0),
	.w5(32'h3c1541d4),
	.w6(32'hbc30f320),
	.w7(32'h3bf72c59),
	.w8(32'h3ca66e51),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7bea),
	.w1(32'hbb067a83),
	.w2(32'hbbd13833),
	.w3(32'hba87945b),
	.w4(32'h3b5d06da),
	.w5(32'hbaa4f9df),
	.w6(32'hbba369bc),
	.w7(32'h3a1c9763),
	.w8(32'hbb065408),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64a88e),
	.w1(32'hbb06dc90),
	.w2(32'h3b3e715b),
	.w3(32'hbc1efcf8),
	.w4(32'h3b5d6a82),
	.w5(32'h3c0370f9),
	.w6(32'hbc11018c),
	.w7(32'h3b5740a1),
	.w8(32'h3c20ffb7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b93c58),
	.w1(32'h3ad426cd),
	.w2(32'hba8c5089),
	.w3(32'h3a56f675),
	.w4(32'h3b1b1a97),
	.w5(32'h39c8cde1),
	.w6(32'h3aa730f0),
	.w7(32'h3b448068),
	.w8(32'h390ffee2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c853a01),
	.w1(32'h3b9efad7),
	.w2(32'hbc4a54da),
	.w3(32'hbbd93e11),
	.w4(32'hbc2c9535),
	.w5(32'hbcd4b746),
	.w6(32'h3b21d1e2),
	.w7(32'h3b2ce7eb),
	.w8(32'hbce8372f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b55e8),
	.w1(32'h3b99a5af),
	.w2(32'h3bf0504a),
	.w3(32'hbb979874),
	.w4(32'h3bc02afb),
	.w5(32'h3bf0d750),
	.w6(32'hbb54012d),
	.w7(32'h3c079b38),
	.w8(32'h3bc870c6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a45221),
	.w1(32'h3a660f91),
	.w2(32'hba459877),
	.w3(32'h37b510b2),
	.w4(32'h3a201dd0),
	.w5(32'hba92b779),
	.w6(32'h388ffa2c),
	.w7(32'h397cce74),
	.w8(32'hba372510),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516b3d),
	.w1(32'hbaef76d4),
	.w2(32'hba096c9f),
	.w3(32'hba45a6aa),
	.w4(32'hbabac2a3),
	.w5(32'hba5709a4),
	.w6(32'hba41f840),
	.w7(32'hbad72f14),
	.w8(32'hba1c3a49),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb377cf2),
	.w1(32'hbb3a6e2c),
	.w2(32'hba5bc6c3),
	.w3(32'hbbbc645c),
	.w4(32'hba7536c1),
	.w5(32'hb9eb8a91),
	.w6(32'hbbcca64a),
	.w7(32'h3a567ac4),
	.w8(32'hbacc7ea0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f2e50),
	.w1(32'h3a08b417),
	.w2(32'hbc3753e0),
	.w3(32'hbac86b2b),
	.w4(32'hb9611b5d),
	.w5(32'hbbf51fea),
	.w6(32'h3ac0f63c),
	.w7(32'h3aba5adc),
	.w8(32'hbc6a0989),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12f7d2),
	.w1(32'h3ae52b66),
	.w2(32'hbba3e818),
	.w3(32'hbc53064d),
	.w4(32'h3b1616a8),
	.w5(32'hbadbbffc),
	.w6(32'hbbcb3bf2),
	.w7(32'h3be14480),
	.w8(32'h3b911671),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d8d7f),
	.w1(32'h388601e0),
	.w2(32'h3ad0b2f9),
	.w3(32'hb9f2ad66),
	.w4(32'hb9b772a9),
	.w5(32'h3ad9d80b),
	.w6(32'hba23b527),
	.w7(32'hb9ed0ee6),
	.w8(32'h3addfce2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7da019),
	.w1(32'h3b89d036),
	.w2(32'h3a178c8b),
	.w3(32'hbc44a22a),
	.w4(32'h3bda71b3),
	.w5(32'h3b9ee068),
	.w6(32'hbc2b00c6),
	.w7(32'h3c0cfc00),
	.w8(32'h3c29cff3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478301),
	.w1(32'h3abc978a),
	.w2(32'hbb33907b),
	.w3(32'hbaec0987),
	.w4(32'h3b5ca51c),
	.w5(32'h39cfb1a5),
	.w6(32'hba8973e2),
	.w7(32'h3b682723),
	.w8(32'h3a928363),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1e487),
	.w1(32'hbbd48261),
	.w2(32'h3bc9c253),
	.w3(32'hbc7966aa),
	.w4(32'hbc14a9bb),
	.w5(32'h3c2fcc37),
	.w6(32'hbc164479),
	.w7(32'hbbda0534),
	.w8(32'h3cb6d2f0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b89e),
	.w1(32'h3c57e756),
	.w2(32'hbc45973e),
	.w3(32'hbc0146b2),
	.w4(32'h3c330df8),
	.w5(32'hbbc9959a),
	.w6(32'h3b4602e5),
	.w7(32'h3cfae3cc),
	.w8(32'h3b3a5a46),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b7b7),
	.w1(32'h3a0cb75f),
	.w2(32'hbb16ec76),
	.w3(32'hb8a0f408),
	.w4(32'h3b0af541),
	.w5(32'hbb5a55f6),
	.w6(32'h3a0ffc11),
	.w7(32'h3b78a7a2),
	.w8(32'hbb8ed067),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ade05),
	.w1(32'h3a58e1f6),
	.w2(32'h3b4271b7),
	.w3(32'h3a494bb9),
	.w4(32'h3a882522),
	.w5(32'h3b8ebc60),
	.w6(32'h3a820a1f),
	.w7(32'h3a60f71a),
	.w8(32'h3ab1cf8d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6db5b),
	.w1(32'h3bff70de),
	.w2(32'h3cb568d0),
	.w3(32'hbad997e8),
	.w4(32'h3be5b5e4),
	.w5(32'h3cebdae8),
	.w6(32'hbb4fdb6a),
	.w7(32'h3bd37add),
	.w8(32'h3c2c94ff),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31db76),
	.w1(32'hba603980),
	.w2(32'h3c4dbb5d),
	.w3(32'hbcd05bf9),
	.w4(32'h3960eec4),
	.w5(32'h3bab07c1),
	.w6(32'hbcd3204a),
	.w7(32'h3b1e6353),
	.w8(32'h3b721b48),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e9831),
	.w1(32'h3c830962),
	.w2(32'hbbd85517),
	.w3(32'h3b72ab5e),
	.w4(32'h3b34d980),
	.w5(32'hbbda388c),
	.w6(32'h3bb4a307),
	.w7(32'h3c172f9d),
	.w8(32'hbbbc08a4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296d64),
	.w1(32'hbbdc9b5d),
	.w2(32'h39e7c6c0),
	.w3(32'h3af8d56e),
	.w4(32'hbbb89cd3),
	.w5(32'hbbb59cb6),
	.w6(32'hb9fd636a),
	.w7(32'hbbe2af36),
	.w8(32'h3b19a308),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61888),
	.w1(32'hbb60a9b5),
	.w2(32'h3ab4a63a),
	.w3(32'h3babf7ba),
	.w4(32'h3b661240),
	.w5(32'h3b054a29),
	.w6(32'h3c4278e5),
	.w7(32'hbb7efca3),
	.w8(32'hbbbcf369),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9d063),
	.w1(32'hbbb9bfb6),
	.w2(32'h3b2fa587),
	.w3(32'hbcbdc2c3),
	.w4(32'h3b947200),
	.w5(32'h3c3bc9bb),
	.w6(32'hbc318ee1),
	.w7(32'hbb33a411),
	.w8(32'h3c4510cf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb387fd3),
	.w1(32'hba8c224f),
	.w2(32'hbc60c921),
	.w3(32'hbb802709),
	.w4(32'h3b4df08f),
	.w5(32'h3c26fbda),
	.w6(32'hbb3973fe),
	.w7(32'h3b72ff17),
	.w8(32'h3c346c8f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c881701),
	.w1(32'hbbfdf868),
	.w2(32'h3b89ffe5),
	.w3(32'h3ce6fd0a),
	.w4(32'hbcb31f65),
	.w5(32'h3c0ce3db),
	.w6(32'h3c85d178),
	.w7(32'hbc9f0d0f),
	.w8(32'h3b83fc0a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bddb),
	.w1(32'hba3a078c),
	.w2(32'h3c1f55b3),
	.w3(32'hbbe17ffa),
	.w4(32'h3af920d3),
	.w5(32'h3b97b437),
	.w6(32'hbb9282d9),
	.w7(32'h3b842594),
	.w8(32'h3c7f6aba),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b887ab0),
	.w1(32'hbc4541ca),
	.w2(32'hbb7bb38f),
	.w3(32'h3a3870ed),
	.w4(32'hbc42fc0e),
	.w5(32'h3a504686),
	.w6(32'h3b9cb150),
	.w7(32'hbca325e1),
	.w8(32'hbb815594),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53d46f),
	.w1(32'hba65b7cb),
	.w2(32'h3c2c84ca),
	.w3(32'hbc57022e),
	.w4(32'h3c4912eb),
	.w5(32'h3c56e4df),
	.w6(32'hbbeb4e8a),
	.w7(32'h3c54fa23),
	.w8(32'h3c31aadd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096610),
	.w1(32'hbb9aba08),
	.w2(32'hbbeee297),
	.w3(32'h3ac3afba),
	.w4(32'hbc144967),
	.w5(32'h3a94ba30),
	.w6(32'h3bff6f5f),
	.w7(32'h3b9995ef),
	.w8(32'h3b411bee),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10d4ad),
	.w1(32'hbb0b9c03),
	.w2(32'hbbf3a988),
	.w3(32'h3c178e10),
	.w4(32'hbc24380b),
	.w5(32'hbb172272),
	.w6(32'h3bfc2c94),
	.w7(32'h38959079),
	.w8(32'h3ab56adf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca69d21),
	.w1(32'hbcad3972),
	.w2(32'h3cbd5ed1),
	.w3(32'hbc96f9b0),
	.w4(32'hbc9c39b3),
	.w5(32'h3c1dd489),
	.w6(32'hbc669694),
	.w7(32'hbbc2ec93),
	.w8(32'h3cca423c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b255d68),
	.w1(32'hb983958d),
	.w2(32'h3a226d51),
	.w3(32'hbaed331b),
	.w4(32'hbba83b93),
	.w5(32'h3aaf189b),
	.w6(32'h3b837d62),
	.w7(32'hbb933dc8),
	.w8(32'hbb158347),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fa3b6),
	.w1(32'h3c18af94),
	.w2(32'hbb60a58f),
	.w3(32'h3c224f38),
	.w4(32'hbb134084),
	.w5(32'hbb9e87f3),
	.w6(32'h3c330cce),
	.w7(32'h3b464a04),
	.w8(32'hbbe21637),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00396a),
	.w1(32'h3c0f8b07),
	.w2(32'h3b7e5452),
	.w3(32'hbc8244fc),
	.w4(32'h3be67127),
	.w5(32'h3c10320a),
	.w6(32'hbbb0f437),
	.w7(32'h3c45050e),
	.w8(32'h3b2e7a51),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a37f7),
	.w1(32'h3baf2fc0),
	.w2(32'h3b767dce),
	.w3(32'hbd44a612),
	.w4(32'h3ca476e6),
	.w5(32'h3c853ff0),
	.w6(32'hbd2ea19b),
	.w7(32'h3c868778),
	.w8(32'h3be991e7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dad2f),
	.w1(32'hbad7c207),
	.w2(32'hbbb64ee2),
	.w3(32'hbc3b4f3d),
	.w4(32'h3c0bdb93),
	.w5(32'h3b106adb),
	.w6(32'h3a27d7cc),
	.w7(32'h3c2b5049),
	.w8(32'hbbcffca0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce14c0c),
	.w1(32'hbc7c6c1b),
	.w2(32'hbc69a2b5),
	.w3(32'hbc6867d0),
	.w4(32'hb943ebcb),
	.w5(32'hbc70dba4),
	.w6(32'hbc1cdf22),
	.w7(32'h3b93ef94),
	.w8(32'hbb091319),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe83fab),
	.w1(32'h3a1a4d7e),
	.w2(32'h3b8bbb69),
	.w3(32'h3be09216),
	.w4(32'h3c676acd),
	.w5(32'h3bb868f0),
	.w6(32'h3b804c45),
	.w7(32'h3c6cdcc2),
	.w8(32'h3bcfb338),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1360f4),
	.w1(32'h3c41f3ae),
	.w2(32'hbc4403ea),
	.w3(32'hbc1495cc),
	.w4(32'h3c749f83),
	.w5(32'h3b06995d),
	.w6(32'hbb8a2161),
	.w7(32'h3ca7a241),
	.w8(32'h3c3c8125),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b64f5),
	.w1(32'h3af12753),
	.w2(32'hb9974fc8),
	.w3(32'hbc7a66c4),
	.w4(32'hbbf5a50d),
	.w5(32'hbc800baf),
	.w6(32'hbc27534a),
	.w7(32'hbb954497),
	.w8(32'hbc3300d1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8aea1c),
	.w1(32'hbc1bd5fc),
	.w2(32'hbc5bb7f1),
	.w3(32'hbc393cee),
	.w4(32'hbc19eb9c),
	.w5(32'hbc07c6d7),
	.w6(32'hbc2cb64a),
	.w7(32'hbc98b010),
	.w8(32'hbbe9592f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31183a),
	.w1(32'h3b5d91c2),
	.w2(32'hbbb7eef7),
	.w3(32'h3cf5b367),
	.w4(32'h3c0d665e),
	.w5(32'hbb152c18),
	.w6(32'h3c819265),
	.w7(32'hbc2f8082),
	.w8(32'h3b0d01d5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf23c3e),
	.w1(32'h39e14f0d),
	.w2(32'hbb009ff5),
	.w3(32'hbc99b563),
	.w4(32'h3b671e35),
	.w5(32'hbb6e7a91),
	.w6(32'hbc8ef966),
	.w7(32'h3c045919),
	.w8(32'h3c15a59b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d577c),
	.w1(32'h3c4c86c4),
	.w2(32'hbc1b01a2),
	.w3(32'h3c427f75),
	.w4(32'h3c2983af),
	.w5(32'hbc36f143),
	.w6(32'h3c8af7e1),
	.w7(32'h3befeb03),
	.w8(32'h3ab8e1da),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3596be),
	.w1(32'h3bd18fc2),
	.w2(32'hbc43e652),
	.w3(32'hbc371330),
	.w4(32'hb9d52112),
	.w5(32'hbc23e956),
	.w6(32'hba584626),
	.w7(32'h3b31af3c),
	.w8(32'hbb9551bc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc437382),
	.w1(32'hba692022),
	.w2(32'hbb5f2a25),
	.w3(32'hbbad8e83),
	.w4(32'hb9c84a29),
	.w5(32'h3babc531),
	.w6(32'hbbc43525),
	.w7(32'h3c0704b8),
	.w8(32'h3b92a260),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb171f1),
	.w1(32'h3b3d8d35),
	.w2(32'h3c116a7a),
	.w3(32'hbcc43c6e),
	.w4(32'h3c06317b),
	.w5(32'h3cc9ec72),
	.w6(32'hbcc1aa50),
	.w7(32'hbb13c086),
	.w8(32'h3c97917f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852e30),
	.w1(32'hbd0adc05),
	.w2(32'hbbbc7397),
	.w3(32'hbc35e396),
	.w4(32'hbd1914a0),
	.w5(32'h3b66af20),
	.w6(32'hbc7c76d6),
	.w7(32'hbc9e4244),
	.w8(32'h3b21a7f8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a741e89),
	.w1(32'h3b8dadd9),
	.w2(32'hbb29e221),
	.w3(32'hbbb9d11f),
	.w4(32'h3b17be11),
	.w5(32'h3c3fe08a),
	.w6(32'h3c00a7f7),
	.w7(32'h3c73bd08),
	.w8(32'h3c457347),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd41f3e5),
	.w1(32'hbc356426),
	.w2(32'hbc025592),
	.w3(32'hbd240b67),
	.w4(32'hbb2449ae),
	.w5(32'h3ac5ee42),
	.w6(32'hbcf90cb6),
	.w7(32'h3c23e083),
	.w8(32'h3cc0bbf5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9445),
	.w1(32'h3cbeb03d),
	.w2(32'hbbd53cb5),
	.w3(32'hbca8911e),
	.w4(32'h3c8cbde6),
	.w5(32'h3a6d4a7f),
	.w6(32'hbaf06c7c),
	.w7(32'h3cd6bb72),
	.w8(32'hb9875a7b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99f8c3),
	.w1(32'hbca87829),
	.w2(32'hbb4e05ac),
	.w3(32'hbc97e06b),
	.w4(32'hbca53d83),
	.w5(32'hbbc1a1e7),
	.w6(32'hbc92d812),
	.w7(32'hbba4be85),
	.w8(32'hbc1ec36d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dda67),
	.w1(32'h3c128bc8),
	.w2(32'h3cd26124),
	.w3(32'hbb6eca25),
	.w4(32'h3b77b9d6),
	.w5(32'h3cc289c6),
	.w6(32'h3a9ebfd9),
	.w7(32'h3b0c4885),
	.w8(32'h3c91bb4b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d7160),
	.w1(32'hbb9527a4),
	.w2(32'hbab56751),
	.w3(32'h3a9d7084),
	.w4(32'hbc491425),
	.w5(32'h3889329c),
	.w6(32'h3b9cbf6d),
	.w7(32'hbc05e050),
	.w8(32'hbb96572b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a0616),
	.w1(32'hba14d394),
	.w2(32'h3c7cdffa),
	.w3(32'hbb9a7167),
	.w4(32'h3ac8224e),
	.w5(32'h3c49d481),
	.w6(32'hbab7c53b),
	.w7(32'h3b398214),
	.w8(32'h3bcb4f07),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565a88),
	.w1(32'hbc6a4937),
	.w2(32'h3b729541),
	.w3(32'hbc2be396),
	.w4(32'hbcb695c5),
	.w5(32'h3b78553d),
	.w6(32'hbc83168b),
	.w7(32'hbc9b6c1a),
	.w8(32'hbbb8d887),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc884a03),
	.w1(32'hb9554546),
	.w2(32'h3c3493e5),
	.w3(32'hbc9c3026),
	.w4(32'h3bf87990),
	.w5(32'h3c8b2fc5),
	.w6(32'hbc7083a4),
	.w7(32'h3be46db8),
	.w8(32'h3bd352c1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e74dd),
	.w1(32'hbc0a58c0),
	.w2(32'hbcab5d16),
	.w3(32'h3bf85e88),
	.w4(32'hbc09438d),
	.w5(32'hbc7ebca4),
	.w6(32'h3bf9e2f9),
	.w7(32'h3bda9436),
	.w8(32'hbc51c8c8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe05e0),
	.w1(32'h3c0fa6c5),
	.w2(32'h3b0776b5),
	.w3(32'hbb943bd4),
	.w4(32'h3c28a190),
	.w5(32'h3b5bde96),
	.w6(32'hbc0ba8d2),
	.w7(32'h3bd75ac4),
	.w8(32'h3bedec21),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9afbbd),
	.w1(32'hbac5e373),
	.w2(32'hbcde9157),
	.w3(32'hbc7f6176),
	.w4(32'h3b2307b8),
	.w5(32'hbcd95342),
	.w6(32'hbc6527f5),
	.w7(32'h3b9acaab),
	.w8(32'hbc2005db),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd24469),
	.w1(32'h3c1e98d9),
	.w2(32'h3b7e2df9),
	.w3(32'h3c10cb24),
	.w4(32'h3c90bdd0),
	.w5(32'h3c4a0581),
	.w6(32'h3c6fac0e),
	.w7(32'h3c37de24),
	.w8(32'h3c5016fa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842dbd),
	.w1(32'hbc70c2aa),
	.w2(32'h3b52d094),
	.w3(32'h3a2a804f),
	.w4(32'hbcb9b28a),
	.w5(32'h3a4cd524),
	.w6(32'hbb6a6491),
	.w7(32'hbc89dff0),
	.w8(32'hbc117e19),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270a09),
	.w1(32'hbc15c6d5),
	.w2(32'hbcc3c6e7),
	.w3(32'hbc90bd2a),
	.w4(32'hbc3a8a7d),
	.w5(32'hbc62da30),
	.w6(32'hbc6f883e),
	.w7(32'hbba27eba),
	.w8(32'hbc12f607),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f7e9a),
	.w1(32'hba509873),
	.w2(32'hb9cf5b7d),
	.w3(32'hbbd8ba1c),
	.w4(32'hbab56ad4),
	.w5(32'hbb0911c5),
	.w6(32'hbc0515ec),
	.w7(32'h3ba802f6),
	.w8(32'h39ebfffc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc613ff4),
	.w1(32'hbaa4d055),
	.w2(32'hbaca2650),
	.w3(32'hbc74a8a1),
	.w4(32'hbacf5171),
	.w5(32'h3bdce0e4),
	.w6(32'hbc1aec68),
	.w7(32'h3b15e630),
	.w8(32'h3b62c7c6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed610a),
	.w1(32'h3b849c24),
	.w2(32'hbc0668eb),
	.w3(32'hbc288591),
	.w4(32'h3acf8a37),
	.w5(32'hbc95540c),
	.w6(32'hbbfcab45),
	.w7(32'hbaa8482e),
	.w8(32'hbc23163f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f3f76),
	.w1(32'h3b27f778),
	.w2(32'hbca0dc82),
	.w3(32'hbb491176),
	.w4(32'h3b0314ea),
	.w5(32'hbc0cf5eb),
	.w6(32'hb98309e1),
	.w7(32'h3bd2649d),
	.w8(32'hbc2c903f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e1bf0),
	.w1(32'hbc8279dc),
	.w2(32'hbc1ccc13),
	.w3(32'hbc597f35),
	.w4(32'hbbd70291),
	.w5(32'h393fda04),
	.w6(32'hbc24f3bd),
	.w7(32'hbbe7ce40),
	.w8(32'hbbb18611),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2081f6),
	.w1(32'hbb6f81e5),
	.w2(32'hbc24060d),
	.w3(32'h3af54c4b),
	.w4(32'hb9b3c7b8),
	.w5(32'hbb29eaac),
	.w6(32'h3b20bafc),
	.w7(32'h3bbfbcf0),
	.w8(32'hbbd5d1c3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3faab7),
	.w1(32'h3b75dc65),
	.w2(32'hbc8c34af),
	.w3(32'hbbf3cb28),
	.w4(32'h3c49c24f),
	.w5(32'hbc5d8c47),
	.w6(32'hbc7c0c1c),
	.w7(32'h3be6caa0),
	.w8(32'h3b569cc2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e2255),
	.w1(32'h3c22b785),
	.w2(32'h3b16f059),
	.w3(32'hbb951f3c),
	.w4(32'h3cb61c72),
	.w5(32'h3bfd5d38),
	.w6(32'h3b49ba24),
	.w7(32'h3c9dc4f5),
	.w8(32'h3b6fa333),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d6aa),
	.w1(32'hbb06de03),
	.w2(32'h3b46a916),
	.w3(32'h3b6558bb),
	.w4(32'hbab16f98),
	.w5(32'h3bbd8174),
	.w6(32'hbb6066f4),
	.w7(32'hbbc20654),
	.w8(32'h3bd53ea7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78158d),
	.w1(32'hbb4acd3b),
	.w2(32'hbc532a08),
	.w3(32'h3c922a98),
	.w4(32'hbc4f8267),
	.w5(32'hbc4d0ffe),
	.w6(32'h3c8ce04e),
	.w7(32'hbc6e7f4c),
	.w8(32'hbc82eb75),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd001a63),
	.w1(32'hbc9205ed),
	.w2(32'h3b2eef70),
	.w3(32'hbce31092),
	.w4(32'h3b66d961),
	.w5(32'h3beb49a7),
	.w6(32'hbcd94469),
	.w7(32'h3b476ab3),
	.w8(32'h3c5bdf40),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0300d6),
	.w1(32'hbbb570be),
	.w2(32'h3c86c03a),
	.w3(32'hbd0d748e),
	.w4(32'hba65f7e5),
	.w5(32'h3d05f2dd),
	.w6(32'hbca40588),
	.w7(32'h3beb6481),
	.w8(32'h3ccb30fd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba4c6b),
	.w1(32'hbc74e741),
	.w2(32'h3c67d119),
	.w3(32'hbcff32b7),
	.w4(32'hbc53129f),
	.w5(32'h3c9671d5),
	.w6(32'hbd09a07c),
	.w7(32'h3b72de15),
	.w8(32'h3cb21278),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63d342),
	.w1(32'hbcbca078),
	.w2(32'h3cbd4aef),
	.w3(32'hbcd47f25),
	.w4(32'hbd0b1351),
	.w5(32'h3c82aa47),
	.w6(32'hbcde46b3),
	.w7(32'hbd1c86cf),
	.w8(32'h3c3c47cd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ebeff),
	.w1(32'hbaec294d),
	.w2(32'hbbfea64b),
	.w3(32'hbb467e3e),
	.w4(32'hbb8ac393),
	.w5(32'hbb98d6bb),
	.w6(32'hbab9b77b),
	.w7(32'hbb8d4f11),
	.w8(32'hbb0bb2c7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972ac5),
	.w1(32'hbc24faf9),
	.w2(32'hbc2c1e79),
	.w3(32'hbab7dec0),
	.w4(32'hbc23bdc5),
	.w5(32'hbbad3665),
	.w6(32'hbce055ae),
	.w7(32'h3b5560da),
	.w8(32'h3b29fc48),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c3680),
	.w1(32'hbc815cd1),
	.w2(32'h3b031193),
	.w3(32'hbc09978b),
	.w4(32'hbbb92921),
	.w5(32'hbb901cd8),
	.w6(32'hbb206031),
	.w7(32'hbb76eec6),
	.w8(32'h3bcbd6ac),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03c24c),
	.w1(32'h3c68021e),
	.w2(32'hbad8a84b),
	.w3(32'hbcc2dffc),
	.w4(32'h3d14975d),
	.w5(32'h3c832857),
	.w6(32'hbc23964d),
	.w7(32'h3d06ba81),
	.w8(32'h3cdd8f7e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fb7e5),
	.w1(32'hbcb83ab4),
	.w2(32'h3c187b12),
	.w3(32'hbc5adf35),
	.w4(32'hbc9e9840),
	.w5(32'h3c82e1b0),
	.w6(32'hbc1c7ecb),
	.w7(32'hbc57ca08),
	.w8(32'h3ce645e1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f44b),
	.w1(32'h3bca9be7),
	.w2(32'hbba7b8d4),
	.w3(32'hbbab3c5d),
	.w4(32'hbb45932d),
	.w5(32'hbbd7fc7d),
	.w6(32'h3a616b87),
	.w7(32'h3b5e1671),
	.w8(32'hbbfdb107),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beff787),
	.w1(32'h3acb33a1),
	.w2(32'hbb56445d),
	.w3(32'h3b94ba87),
	.w4(32'hbb4fbbd9),
	.w5(32'hbc56c6e3),
	.w6(32'h3bfb0ece),
	.w7(32'h394775b3),
	.w8(32'hbc743ba9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfaaf6),
	.w1(32'hbba4b4ef),
	.w2(32'h3c469bc6),
	.w3(32'hbbd3dc09),
	.w4(32'hbaed5cba),
	.w5(32'h3bf43be8),
	.w6(32'hbbadaf4e),
	.w7(32'h3a131b78),
	.w8(32'hbba886c7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bb846),
	.w1(32'hba81e69e),
	.w2(32'hbc5fddc1),
	.w3(32'h3a9f3cdb),
	.w4(32'h3be4f644),
	.w5(32'hbc259b41),
	.w6(32'h3b4675c4),
	.w7(32'h3c4bb0eb),
	.w8(32'hbc0d775b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea5e33),
	.w1(32'h3b1b1058),
	.w2(32'h3b9e9bde),
	.w3(32'hbbe04b8f),
	.w4(32'h3c84b831),
	.w5(32'h3bd7e4cf),
	.w6(32'h37f24018),
	.w7(32'h3bea5129),
	.w8(32'hbaea67b8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8159c4),
	.w1(32'h3b91de35),
	.w2(32'hbba2013e),
	.w3(32'h3c84369e),
	.w4(32'h3bac30b9),
	.w5(32'h3babd4ad),
	.w6(32'h3c229020),
	.w7(32'h3c1b76ea),
	.w8(32'hbc116460),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9bed),
	.w1(32'hbc7372c0),
	.w2(32'hbc150d73),
	.w3(32'hbabbd3df),
	.w4(32'hbc0fed12),
	.w5(32'hbca8e97e),
	.w6(32'hbc61288a),
	.w7(32'hbc2757f1),
	.w8(32'hbc5db9c4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafc51b),
	.w1(32'h3b1c293e),
	.w2(32'h3b951ccd),
	.w3(32'hbc79f586),
	.w4(32'h3cf3779d),
	.w5(32'h3c281a05),
	.w6(32'hbb6f5e46),
	.w7(32'h3c9ee669),
	.w8(32'h3b6f4659),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c83971),
	.w1(32'h3bdc1cbf),
	.w2(32'hbbf1e6c5),
	.w3(32'hbb8b14a1),
	.w4(32'h3b455483),
	.w5(32'hbc6d49b4),
	.w6(32'hbaa60fe0),
	.w7(32'h3bce7c1f),
	.w8(32'h3b5f48f7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c6018),
	.w1(32'h3b3e8e55),
	.w2(32'h3c6b9fcc),
	.w3(32'hbabcca48),
	.w4(32'h3b0d2e41),
	.w5(32'h3c711c96),
	.w6(32'hbae54b9a),
	.w7(32'h39e01d7e),
	.w8(32'h3bed163f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf7fefd),
	.w1(32'hbd2ad0cc),
	.w2(32'hbc87774b),
	.w3(32'hbd149ed1),
	.w4(32'hbcf9e942),
	.w5(32'hbaf7842a),
	.w6(32'hbd3bcbbc),
	.w7(32'hbc998d32),
	.w8(32'h3cce3a20),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ce060),
	.w1(32'hbb3ead14),
	.w2(32'h3c63af41),
	.w3(32'h3b0926a0),
	.w4(32'h3c26a78f),
	.w5(32'h3ce99acf),
	.w6(32'h3c128ce2),
	.w7(32'h3c313cac),
	.w8(32'h3cc6d96b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc017b),
	.w1(32'h3c79c151),
	.w2(32'h3c02758c),
	.w3(32'h3c189197),
	.w4(32'h3cbfdee2),
	.w5(32'h3c63ebf3),
	.w6(32'h3c2d289c),
	.w7(32'h3c522dfe),
	.w8(32'h3c152669),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31a063),
	.w1(32'hbcafd28d),
	.w2(32'h3c4f1c83),
	.w3(32'hbc4bcb0d),
	.w4(32'hbccd83c7),
	.w5(32'h3cc07ed4),
	.w6(32'hbca6d1c2),
	.w7(32'hbca0fdd4),
	.w8(32'h3ccb7a84),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b275f65),
	.w1(32'hbbdc9229),
	.w2(32'hbc14d717),
	.w3(32'h3b314247),
	.w4(32'hbbb76bdf),
	.w5(32'hbb496e48),
	.w6(32'hbb65a343),
	.w7(32'hbbc118d8),
	.w8(32'hbb890af6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e0c69),
	.w1(32'h3c20de56),
	.w2(32'hbc160fef),
	.w3(32'h3ba9cf84),
	.w4(32'h3c70e65f),
	.w5(32'hbba8b3ae),
	.w6(32'h3bf66bc3),
	.w7(32'h3bfc45b3),
	.w8(32'hbb853478),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00886),
	.w1(32'hbac93e08),
	.w2(32'hbb800890),
	.w3(32'hbc352f9d),
	.w4(32'hbb978e47),
	.w5(32'hbbe94947),
	.w6(32'hbb410ab9),
	.w7(32'h3b91bad3),
	.w8(32'hb7e58eb4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e592c),
	.w1(32'hba0d4c9e),
	.w2(32'hba10cf3b),
	.w3(32'h3a886788),
	.w4(32'h3ba97b42),
	.w5(32'h3ad12206),
	.w6(32'hbb69f33a),
	.w7(32'hbb670e6f),
	.w8(32'hbab918c8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c50e),
	.w1(32'h3b8433a2),
	.w2(32'hbbc0713a),
	.w3(32'h3ad8991c),
	.w4(32'h3b76c00a),
	.w5(32'hba82c34d),
	.w6(32'h3bc6ea18),
	.w7(32'h3b5e7127),
	.w8(32'h3b132b77),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f3606),
	.w1(32'h3c2a21ff),
	.w2(32'h3a684962),
	.w3(32'h3c3220a3),
	.w4(32'h3c899265),
	.w5(32'h3b876f0f),
	.w6(32'hbb6d31ea),
	.w7(32'h3c438c41),
	.w8(32'h39cf4f9d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c1dff),
	.w1(32'hbb9dff3d),
	.w2(32'hbbc40d45),
	.w3(32'hbd0db5ed),
	.w4(32'h3c1a66fd),
	.w5(32'h3b11f6c0),
	.w6(32'hbce1a6fd),
	.w7(32'h3bba4ff8),
	.w8(32'h3c80b70a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd980eb),
	.w1(32'h3b6df4ed),
	.w2(32'h3c00a929),
	.w3(32'hbc6b3b1d),
	.w4(32'h3c1504a3),
	.w5(32'h3c72d639),
	.w6(32'hbc58c8b7),
	.w7(32'h3c1832c2),
	.w8(32'h3c7a45a5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a9fa),
	.w1(32'hbb8fd92b),
	.w2(32'hba1783bd),
	.w3(32'h3c57e686),
	.w4(32'hbc69aec4),
	.w5(32'hba864091),
	.w6(32'h3a61fb98),
	.w7(32'hbc914f38),
	.w8(32'h3bb4d7dd),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37fde5),
	.w1(32'hb970ee62),
	.w2(32'hbc0b15e4),
	.w3(32'hba968f31),
	.w4(32'hbb4c41c2),
	.w5(32'hbc3e408f),
	.w6(32'h3bf886ca),
	.w7(32'h3ab6f6b5),
	.w8(32'hbbbe67e3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a878bf3),
	.w1(32'h3a575a24),
	.w2(32'h3c034dd1),
	.w3(32'h3be90b8c),
	.w4(32'hb8997ca1),
	.w5(32'h3c032e08),
	.w6(32'h3b5cb964),
	.w7(32'hbc01f6ae),
	.w8(32'h3c5676cf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b6870),
	.w1(32'hbb426326),
	.w2(32'hbc2334be),
	.w3(32'hbbca9552),
	.w4(32'hbc534de4),
	.w5(32'h3bd0c432),
	.w6(32'h3bfa4cbd),
	.w7(32'hb9c4206d),
	.w8(32'h3a305220),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7ba92),
	.w1(32'h3c389259),
	.w2(32'h3c119284),
	.w3(32'hbba4dbc0),
	.w4(32'h3c58f857),
	.w5(32'h3be38797),
	.w6(32'hbaa542d9),
	.w7(32'h3c887289),
	.w8(32'h3c5a9c8d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac45d),
	.w1(32'h3c015ca1),
	.w2(32'hbbf54f5b),
	.w3(32'h3a2b1746),
	.w4(32'hba6c939f),
	.w5(32'hbb7eb6da),
	.w6(32'h3b272ba5),
	.w7(32'hbae1c9cc),
	.w8(32'hbb832018),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0b6d),
	.w1(32'h3b74c31b),
	.w2(32'h3b29ca0b),
	.w3(32'hbbe78ba6),
	.w4(32'h3a9056f1),
	.w5(32'h3af1cd3a),
	.w6(32'hbb898e5b),
	.w7(32'h3b67e282),
	.w8(32'h3a09b9ef),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b312),
	.w1(32'h3ade3554),
	.w2(32'hbbe14409),
	.w3(32'hbab7d041),
	.w4(32'h3ae690a7),
	.w5(32'hbb54899f),
	.w6(32'h3ab4a5c5),
	.w7(32'h3bd03d3e),
	.w8(32'h3b02a593),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0ce3),
	.w1(32'hbbbf28b5),
	.w2(32'h3cc0cf3d),
	.w3(32'h3b87bd0a),
	.w4(32'hbbdba957),
	.w5(32'h3d06e831),
	.w6(32'hb797df73),
	.w7(32'hbc249d1a),
	.w8(32'h3c94c24a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb19a82),
	.w1(32'hbbc12f4a),
	.w2(32'h3caa2fe6),
	.w3(32'h3cd5637a),
	.w4(32'hbcea4b77),
	.w5(32'h3c946aa4),
	.w6(32'h3a408768),
	.w7(32'hbd08f10f),
	.w8(32'h3c6edf42),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baa55b),
	.w1(32'hbc371a21),
	.w2(32'hbc9253a4),
	.w3(32'hbc2d3a19),
	.w4(32'hbc9dcfb7),
	.w5(32'hbb66dd93),
	.w6(32'hbc555e36),
	.w7(32'hbc42f425),
	.w8(32'h3b95c9fe),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd27cee3),
	.w1(32'h3cbcc127),
	.w2(32'h3b765ac9),
	.w3(32'hbcc72d87),
	.w4(32'h3d03eb17),
	.w5(32'h3caa8d4e),
	.w6(32'hbccc18ca),
	.w7(32'h3cdcb3eb),
	.w8(32'h3ce8a25e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0257b1),
	.w1(32'hbc97f1de),
	.w2(32'h3c0516e6),
	.w3(32'hbc2bf455),
	.w4(32'hbba98ef9),
	.w5(32'h3c11d868),
	.w6(32'hbc3b66de),
	.w7(32'hbb79e866),
	.w8(32'h3c036f78),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e01c),
	.w1(32'hbc3da70e),
	.w2(32'h3cbfb6e2),
	.w3(32'hbb4c8a9d),
	.w4(32'hbc077094),
	.w5(32'h3cb63cc3),
	.w6(32'hbc90529e),
	.w7(32'hbc633165),
	.w8(32'h3c574b22),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule