module layer_6_featuremap_125(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb41e8a),
	.w1(32'h3bbb8c54),
	.w2(32'h3c1e0313),
	.w3(32'h3b9fda2c),
	.w4(32'h3b69130f),
	.w5(32'h3c4e8646),
	.w6(32'h3b77e292),
	.w7(32'h3bd07bed),
	.w8(32'h3c880615),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a3ab3),
	.w1(32'h3bdc38c8),
	.w2(32'h3b1ab759),
	.w3(32'hb9f611a1),
	.w4(32'h39c77e5d),
	.w5(32'hbaa75af3),
	.w6(32'h3c3196ac),
	.w7(32'h3b18e33e),
	.w8(32'hbc27bf8d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4983db),
	.w1(32'h3c9a72eb),
	.w2(32'hbbe2b6e6),
	.w3(32'h3caa00b7),
	.w4(32'h3ca1f52d),
	.w5(32'hbc13fd71),
	.w6(32'h3d15b96a),
	.w7(32'h3c724f9d),
	.w8(32'hbba1dbb0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe17af9),
	.w1(32'h3c7c96e9),
	.w2(32'h3c74364d),
	.w3(32'h3c2abdb3),
	.w4(32'h3c415bd6),
	.w5(32'hba5a0ec4),
	.w6(32'h3c83fdb0),
	.w7(32'h3c6ae258),
	.w8(32'hbb90a271),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbcd2e),
	.w1(32'hbc990d51),
	.w2(32'hbbf086b3),
	.w3(32'hbc605607),
	.w4(32'hbc390fd1),
	.w5(32'h39e143f5),
	.w6(32'hbcfb162f),
	.w7(32'hbc2c077d),
	.w8(32'h3c526ea9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560943),
	.w1(32'hbc80a6ba),
	.w2(32'hbb20730c),
	.w3(32'hbc2b8684),
	.w4(32'hbb52b580),
	.w5(32'h3bc237aa),
	.w6(32'hbc88b2d1),
	.w7(32'hbb058054),
	.w8(32'h3c4bb972),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bfba5),
	.w1(32'h3c35c0cf),
	.w2(32'hbb5cfc3b),
	.w3(32'h3c1bf76a),
	.w4(32'h3b22d9bd),
	.w5(32'hbc87333e),
	.w6(32'h3c94a367),
	.w7(32'hbb3d6ebd),
	.w8(32'hbcef1e98),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccaf353),
	.w1(32'h3cacf668),
	.w2(32'h3bc0bb1b),
	.w3(32'h3c9f2d6b),
	.w4(32'hbb248f48),
	.w5(32'hbba9493a),
	.w6(32'h3cb710e0),
	.w7(32'h3ca5a8e6),
	.w8(32'hbcc33ca0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f7a0f),
	.w1(32'hbbe7cc3c),
	.w2(32'h3a1599e5),
	.w3(32'hbc11a4f9),
	.w4(32'h3c1daf1c),
	.w5(32'hbc0f6b7b),
	.w6(32'hbb85cec0),
	.w7(32'h3b1a91cf),
	.w8(32'hbbb1e96a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0b84c),
	.w1(32'hbb6c2c9e),
	.w2(32'h3c33f12c),
	.w3(32'hbc000893),
	.w4(32'h3b531043),
	.w5(32'h3c7b4c99),
	.w6(32'hbc122f4b),
	.w7(32'h3c054155),
	.w8(32'h3ca7b993),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21b3e3),
	.w1(32'hbc2ec16a),
	.w2(32'hbc02f53f),
	.w3(32'hbb897f3e),
	.w4(32'h3b1cbffe),
	.w5(32'hbca1f6cf),
	.w6(32'h3ad32b59),
	.w7(32'hbc09dc6a),
	.w8(32'hbcb72e95),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb466e8),
	.w1(32'hbc332908),
	.w2(32'h3b5be985),
	.w3(32'hbb2e33be),
	.w4(32'h39f70375),
	.w5(32'h3c9b8a28),
	.w6(32'hbc4bdc40),
	.w7(32'hbbe775c9),
	.w8(32'h3c56f0d3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92b625),
	.w1(32'hbb5c8451),
	.w2(32'h3c638329),
	.w3(32'hbb8bdd31),
	.w4(32'h3c71a434),
	.w5(32'hbb7738fa),
	.w6(32'hba429b64),
	.w7(32'h3c7aec17),
	.w8(32'hbc0d6a4f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d271f),
	.w1(32'h3cc30cce),
	.w2(32'h3c5df920),
	.w3(32'h3c5d3b8e),
	.w4(32'h3c87e149),
	.w5(32'h3bb2995b),
	.w6(32'h3cc3df9a),
	.w7(32'h3c9ad185),
	.w8(32'hbb05aa12),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3531),
	.w1(32'h3b79ebdc),
	.w2(32'hbb03c673),
	.w3(32'h3bfa4858),
	.w4(32'h3bc407c5),
	.w5(32'h39a2bdc4),
	.w6(32'h3c0b9c63),
	.w7(32'h3bc1f022),
	.w8(32'hbb3bb468),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b7beb),
	.w1(32'hbb82754e),
	.w2(32'hbb9c1e0b),
	.w3(32'hbb301507),
	.w4(32'hbb13658f),
	.w5(32'hbb29cadd),
	.w6(32'h3b1b51b0),
	.w7(32'hbb2fb7d0),
	.w8(32'hbbb0cc15),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c49f),
	.w1(32'h3c9f6c5a),
	.w2(32'h3bcc676f),
	.w3(32'h3cdcdfcf),
	.w4(32'h3c40f9f9),
	.w5(32'hbcda3dbb),
	.w6(32'h3d12aa49),
	.w7(32'h3c47d658),
	.w8(32'hbcf3f52f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c18eb),
	.w1(32'hbaf69e8a),
	.w2(32'h3b90b470),
	.w3(32'hbb84e030),
	.w4(32'hbae98e86),
	.w5(32'h3bf1562f),
	.w6(32'hbb52203d),
	.w7(32'h39e76f93),
	.w8(32'h3c19749f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4968a5),
	.w1(32'hba387a2f),
	.w2(32'h3ab9a7c5),
	.w3(32'h3b05fe61),
	.w4(32'h3b4e8109),
	.w5(32'h3ac9b47f),
	.w6(32'h3b142ed1),
	.w7(32'h3b25bce9),
	.w8(32'h3abdba6a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a421279),
	.w1(32'h3ca5f0f4),
	.w2(32'hbc5f423c),
	.w3(32'h3c17784b),
	.w4(32'hbc302362),
	.w5(32'hbc80127a),
	.w6(32'h3c4d4472),
	.w7(32'hbc872a50),
	.w8(32'hbc1cdb75),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd616e),
	.w1(32'h3bc72701),
	.w2(32'hbb30bc2c),
	.w3(32'h3bb53f6d),
	.w4(32'hbacec21b),
	.w5(32'hbbb67293),
	.w6(32'h3bead556),
	.w7(32'hbb48d453),
	.w8(32'hbc0d0e2e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58a704),
	.w1(32'h3c85e082),
	.w2(32'hbc02c01e),
	.w3(32'h3c97834e),
	.w4(32'hbc3d1b66),
	.w5(32'hbce1aa1f),
	.w6(32'h3cdb53b4),
	.w7(32'h3a44279e),
	.w8(32'hbcc88476),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b79d6),
	.w1(32'h3c9a529a),
	.w2(32'h3d86184c),
	.w3(32'hbc767db8),
	.w4(32'h3ca87f7c),
	.w5(32'h3bd9b5b4),
	.w6(32'h3bc20175),
	.w7(32'h3d7a7874),
	.w8(32'h3d0bd924),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfdd3c0),
	.w1(32'hbb8ba325),
	.w2(32'hbc886af6),
	.w3(32'hbca28571),
	.w4(32'hbc7c87c6),
	.w5(32'hbd33cc71),
	.w6(32'h3bb21726),
	.w7(32'hbc25cfd1),
	.w8(32'hbd18c6b7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce78503),
	.w1(32'h3b98394c),
	.w2(32'h3c6db84c),
	.w3(32'h3cb38391),
	.w4(32'h3c1f5c8d),
	.w5(32'hbcb5f5de),
	.w6(32'h3c8ec399),
	.w7(32'h3c30f78f),
	.w8(32'hbb6953b0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc382ece),
	.w1(32'hbae1e33f),
	.w2(32'hb9ff6e10),
	.w3(32'h3c881e3d),
	.w4(32'hba81acc4),
	.w5(32'hbc438ae8),
	.w6(32'h3c86d160),
	.w7(32'h3b65089b),
	.w8(32'hbc64e1e2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1bd8),
	.w1(32'hbbcf5140),
	.w2(32'hbc0204ea),
	.w3(32'h3c2906c0),
	.w4(32'h3bcdc116),
	.w5(32'hbc3710a9),
	.w6(32'h3b30fcc0),
	.w7(32'hbba8406c),
	.w8(32'hbc2f614c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84e7f8),
	.w1(32'hb9fc3c82),
	.w2(32'hbc2666dd),
	.w3(32'h3bd110ad),
	.w4(32'hba597da4),
	.w5(32'hbc6f126b),
	.w6(32'h3c2ba4e5),
	.w7(32'hbb8fef95),
	.w8(32'hbcae4729),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ea3c7),
	.w1(32'h3b8d6d75),
	.w2(32'hbb70f26e),
	.w3(32'h3b651ad4),
	.w4(32'hb9079cc4),
	.w5(32'hbba4d308),
	.w6(32'h3b9603f3),
	.w7(32'hbb3c1744),
	.w8(32'hbc27f113),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd3342),
	.w1(32'hbb60aed9),
	.w2(32'h3cbffa49),
	.w3(32'hbb905998),
	.w4(32'hbc904c6d),
	.w5(32'h3c873faa),
	.w6(32'h3c43842b),
	.w7(32'hbac2711f),
	.w8(32'hbc97efc4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25da17),
	.w1(32'hbccf9aa3),
	.w2(32'hbd2d4b17),
	.w3(32'h3c698abc),
	.w4(32'h3cf57df1),
	.w5(32'h3c19c92c),
	.w6(32'h3bb93797),
	.w7(32'h394c56f5),
	.w8(32'hbbc6de83),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc726466),
	.w1(32'hbcdec9ca),
	.w2(32'hbc031751),
	.w3(32'hbce45b74),
	.w4(32'hbc858441),
	.w5(32'hba77a1cf),
	.w6(32'hbd1a1b21),
	.w7(32'hbccba2c8),
	.w8(32'h3c0268b0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c7b5a),
	.w1(32'h3c2f959e),
	.w2(32'hbc87a6b9),
	.w3(32'h3c3c64d6),
	.w4(32'hbc55c3e0),
	.w5(32'hbcbc3ea9),
	.w6(32'h3cff4a6d),
	.w7(32'hbc3e25fa),
	.w8(32'hbd089914),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca23365),
	.w1(32'h3c42ac48),
	.w2(32'h3c3ca489),
	.w3(32'h3abba59c),
	.w4(32'hbaa59787),
	.w5(32'hbb2a66d4),
	.w6(32'h3c02f3aa),
	.w7(32'h3b227b26),
	.w8(32'hbbc5dbba),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3898a5),
	.w1(32'hbbae4797),
	.w2(32'h3bf4c19a),
	.w3(32'hbbab17e5),
	.w4(32'h3a2c66ee),
	.w5(32'h3c092657),
	.w6(32'hbc00e934),
	.w7(32'h3bc43b6d),
	.w8(32'h3c79422b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfb82),
	.w1(32'hb7e38992),
	.w2(32'h3bcc3908),
	.w3(32'h3ad92988),
	.w4(32'hbb078f81),
	.w5(32'hbbb106c9),
	.w6(32'h3b80f6c5),
	.w7(32'h3b02e34c),
	.w8(32'hbc788631),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c045365),
	.w1(32'hbc1db63b),
	.w2(32'hbc1126d0),
	.w3(32'h3abd8ff1),
	.w4(32'hbb05e822),
	.w5(32'h39884173),
	.w6(32'hbc24160e),
	.w7(32'hbb8f0ea0),
	.w8(32'h3bb84f3c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a68389),
	.w1(32'h3bd5213f),
	.w2(32'h3b7576cd),
	.w3(32'h3c00d30c),
	.w4(32'h3a1e709b),
	.w5(32'hbaf5ccf3),
	.w6(32'h3c1a6963),
	.w7(32'h3b60dddb),
	.w8(32'hbb89befc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc63897),
	.w1(32'h3c80a811),
	.w2(32'h3c259d54),
	.w3(32'h3c6f3740),
	.w4(32'h3c9c3b32),
	.w5(32'h3c59b6a1),
	.w6(32'h3c97a763),
	.w7(32'h3c7f912d),
	.w8(32'h3cb75d93),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d168d59),
	.w1(32'hbc791752),
	.w2(32'hbcca74d2),
	.w3(32'h3c5eca45),
	.w4(32'h3bb745c6),
	.w5(32'hbc3f59d3),
	.w6(32'h3c51df13),
	.w7(32'hbcd9e85e),
	.w8(32'hbc0c99f7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba41350),
	.w1(32'hbc20ac7f),
	.w2(32'hbcabcbca),
	.w3(32'hbbf7e3da),
	.w4(32'hbc4584db),
	.w5(32'hbab35d39),
	.w6(32'hbb043211),
	.w7(32'hbc8c7785),
	.w8(32'hbb759a5c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e4fee),
	.w1(32'h3c3f3fc6),
	.w2(32'h3bd79cce),
	.w3(32'h3c0764c1),
	.w4(32'h3bb19f7b),
	.w5(32'hbbb956b0),
	.w6(32'h3c7f7d8a),
	.w7(32'h3bc6f9b0),
	.w8(32'hbc4fdaf7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfebc0e),
	.w1(32'h3be0ae46),
	.w2(32'h3c1b85e7),
	.w3(32'h3b06531f),
	.w4(32'hbb6b7a36),
	.w5(32'hbac28df3),
	.w6(32'h3a020956),
	.w7(32'h3b8a8d58),
	.w8(32'h3bfcdcbb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae094a7),
	.w1(32'h3b44fad1),
	.w2(32'h3c20aaca),
	.w3(32'h3c1dff99),
	.w4(32'h3b17815a),
	.w5(32'hbacf2869),
	.w6(32'h3c7fd3bf),
	.w7(32'hbb952ab1),
	.w8(32'hbcdefcd2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b122d63),
	.w1(32'h3aa9de48),
	.w2(32'hbc352d35),
	.w3(32'h3b6ec757),
	.w4(32'hba866062),
	.w5(32'hbc140d5c),
	.w6(32'h3bfc53d0),
	.w7(32'hbb118a0d),
	.w8(32'hbbc18712),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205ef7),
	.w1(32'h3b8a802b),
	.w2(32'h39ffd9cc),
	.w3(32'h3c541b90),
	.w4(32'h3bb00858),
	.w5(32'hbcad4631),
	.w6(32'h3c537d3e),
	.w7(32'h3aa806c9),
	.w8(32'hbbe19c2c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a1675),
	.w1(32'h3c9eaaa3),
	.w2(32'h3cb35a12),
	.w3(32'h3b87e58e),
	.w4(32'h3c76767d),
	.w5(32'h3c8a1191),
	.w6(32'h3c6a784f),
	.w7(32'h3cfaf9fe),
	.w8(32'hbac1a56b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dc449),
	.w1(32'h3d15ad6a),
	.w2(32'hbbf3dc9a),
	.w3(32'h3ce00719),
	.w4(32'hbbc67442),
	.w5(32'hbcd416ea),
	.w6(32'h3d31c932),
	.w7(32'hbc6876cd),
	.w8(32'hbd1799c1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd062880),
	.w1(32'hbba960fb),
	.w2(32'h3b663be6),
	.w3(32'hbc088289),
	.w4(32'hbb5875b5),
	.w5(32'h3b8d226e),
	.w6(32'hbb6e1684),
	.w7(32'h3ae5d5ac),
	.w8(32'h3b8907d1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6ce14),
	.w1(32'hbbeaf6d4),
	.w2(32'h3b18e486),
	.w3(32'hbc96c212),
	.w4(32'hbb3a1570),
	.w5(32'h3b04ed8a),
	.w6(32'hba273915),
	.w7(32'h3b93850f),
	.w8(32'hba8ef8d5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ed706),
	.w1(32'h3c48ace6),
	.w2(32'h3c9ee4d1),
	.w3(32'h3c21e71b),
	.w4(32'h3c889ee6),
	.w5(32'hbbf371cd),
	.w6(32'h3cb3aaac),
	.w7(32'h3cc6cb6c),
	.w8(32'hbc31e52d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17ceca),
	.w1(32'h3c58553e),
	.w2(32'h3bd6d930),
	.w3(32'h3c6a8acc),
	.w4(32'h3c1f1d0c),
	.w5(32'hbb9fc47e),
	.w6(32'h3cc18454),
	.w7(32'h3c70764e),
	.w8(32'hbbd06366),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18f64e),
	.w1(32'h3c8901d1),
	.w2(32'hbb962e91),
	.w3(32'h3ca40184),
	.w4(32'h3c55167b),
	.w5(32'hbc8ae443),
	.w6(32'h3d112723),
	.w7(32'h3c5db7b3),
	.w8(32'hbc8ddbd4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd2682),
	.w1(32'h3c07238f),
	.w2(32'hb9f207bc),
	.w3(32'hbafbbc9c),
	.w4(32'hb9718df0),
	.w5(32'hbc0993ad),
	.w6(32'h3c4026c2),
	.w7(32'h3b97448e),
	.w8(32'hbc905319),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3708d),
	.w1(32'h3bc08248),
	.w2(32'h3c384e9e),
	.w3(32'h3b229bf1),
	.w4(32'h3c1d2aaf),
	.w5(32'h39f98beb),
	.w6(32'h3c6240e4),
	.w7(32'h3c86a2c5),
	.w8(32'hbb9a4d9f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2572c7),
	.w1(32'h3b0bf98b),
	.w2(32'h3c18dd43),
	.w3(32'h3b26851a),
	.w4(32'h3aff2a8e),
	.w5(32'h3b5941c1),
	.w6(32'h3b80e2ac),
	.w7(32'h3ac82e40),
	.w8(32'hbb905d89),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6550c5),
	.w1(32'hbb8cebe6),
	.w2(32'hbb59b7ed),
	.w3(32'hbbce7cd7),
	.w4(32'hbb97c703),
	.w5(32'hbb66834b),
	.w6(32'hbbbcdedb),
	.w7(32'hbb7f0e99),
	.w8(32'hbb489e67),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3d0f0),
	.w1(32'h3b62c8b8),
	.w2(32'h3b41c44e),
	.w3(32'h3b748342),
	.w4(32'h3b44b8db),
	.w5(32'h3b3ed210),
	.w6(32'h3b8eeabd),
	.w7(32'h3b57df54),
	.w8(32'h3b237e30),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca4ff),
	.w1(32'h3b0bff13),
	.w2(32'h3afab802),
	.w3(32'h3b297a04),
	.w4(32'h3b3d83e3),
	.w5(32'h3b37771b),
	.w6(32'h3b1abb26),
	.w7(32'h3b124e2c),
	.w8(32'h3aeec0c1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f7576),
	.w1(32'h3c0319d2),
	.w2(32'h3be3c8a5),
	.w3(32'h3c58205f),
	.w4(32'h3c3133e9),
	.w5(32'hbb1f2107),
	.w6(32'h3c7bb118),
	.w7(32'h3c386dfc),
	.w8(32'h3b6b99e8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34e7ed),
	.w1(32'h3bf01b80),
	.w2(32'h3bc94e15),
	.w3(32'h3c378561),
	.w4(32'h3c101084),
	.w5(32'h3b8fa318),
	.w6(32'h3c18fb96),
	.w7(32'h3bd731fe),
	.w8(32'h3b89e9e6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1ee8b),
	.w1(32'h3a9b0619),
	.w2(32'h3bb0a92f),
	.w3(32'h3bb12793),
	.w4(32'h3ba426ab),
	.w5(32'hbb2a78e1),
	.w6(32'h3c2fb499),
	.w7(32'h3bf05c65),
	.w8(32'hbb049d46),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc796cdb),
	.w1(32'hbbe471bd),
	.w2(32'hb9a7ccea),
	.w3(32'hbbe1d472),
	.w4(32'hbc0fd167),
	.w5(32'h3aa04753),
	.w6(32'hbbdd281a),
	.w7(32'hbb2d4ea2),
	.w8(32'hbc3c30e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d358),
	.w1(32'h3baccb77),
	.w2(32'h3ade48bc),
	.w3(32'h3bfcb8d3),
	.w4(32'h3bf28475),
	.w5(32'h3b929575),
	.w6(32'h3be4b030),
	.w7(32'h3bc52292),
	.w8(32'h3b46b6bc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule