module layer_8_featuremap_83(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b624212),
	.w1(32'hba30d38c),
	.w2(32'h3ba2d756),
	.w3(32'h3aa53f28),
	.w4(32'h3b899c5b),
	.w5(32'h3adde6ea),
	.w6(32'h3b2f2741),
	.w7(32'h3a1f4f2a),
	.w8(32'hba20bca9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacbf96),
	.w1(32'h3977bba5),
	.w2(32'h3a284dc6),
	.w3(32'hba34616c),
	.w4(32'h3a8cf018),
	.w5(32'hbabaa22f),
	.w6(32'h39aa714b),
	.w7(32'hb9d487b0),
	.w8(32'h3a11bd6b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec56e6),
	.w1(32'hbb20b673),
	.w2(32'h3aa79e14),
	.w3(32'hb9cbb1ae),
	.w4(32'hb9d66c57),
	.w5(32'hb8b7b77a),
	.w6(32'hb88fba2e),
	.w7(32'h39dabb68),
	.w8(32'hbb7c9d8c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab924b5),
	.w1(32'hbc1ba2e3),
	.w2(32'h3b947099),
	.w3(32'h3b12b9d9),
	.w4(32'hbbcb256d),
	.w5(32'hbbecf427),
	.w6(32'h3be5a751),
	.w7(32'h3b0ea05e),
	.w8(32'hbb119bd4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba742a3f),
	.w1(32'hbbb550c6),
	.w2(32'hbab10432),
	.w3(32'h3a8ab6ac),
	.w4(32'hba59d037),
	.w5(32'hbac4f970),
	.w6(32'hbb45d830),
	.w7(32'hbb01a352),
	.w8(32'hbb6485fa),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbd54c),
	.w1(32'hbb6a21b3),
	.w2(32'h3c3a80b7),
	.w3(32'h3bc2a6a0),
	.w4(32'h3b49467f),
	.w5(32'h3acfd680),
	.w6(32'hbaddf03a),
	.w7(32'h3c0b8341),
	.w8(32'h3b14c402),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa33fb),
	.w1(32'h3afe65b7),
	.w2(32'h3b1d310b),
	.w3(32'hb813d744),
	.w4(32'h3ac09a59),
	.w5(32'h3a844f82),
	.w6(32'h39e1f098),
	.w7(32'hbac0118f),
	.w8(32'hbb564a99),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8621e),
	.w1(32'hbbe3f8c1),
	.w2(32'hbb1083b4),
	.w3(32'h39e07e61),
	.w4(32'h3aacc853),
	.w5(32'hba7deacf),
	.w6(32'hbb813936),
	.w7(32'hbb185bda),
	.w8(32'h38198cf7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841006),
	.w1(32'h3a24ecb9),
	.w2(32'h38a59c60),
	.w3(32'hba4da7d3),
	.w4(32'h389cba3b),
	.w5(32'hbacfd9ca),
	.w6(32'hbac071fb),
	.w7(32'hbb9ee987),
	.w8(32'hbc82298f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d780),
	.w1(32'h3c1a6d5a),
	.w2(32'hbc9e774e),
	.w3(32'hb95d7ab8),
	.w4(32'h3af8aa82),
	.w5(32'hbbac6e51),
	.w6(32'hbc8d3550),
	.w7(32'hbc7b9bc5),
	.w8(32'hbbc3e551),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ab68),
	.w1(32'hbb9e5b11),
	.w2(32'hbba1257f),
	.w3(32'hbc1e4f15),
	.w4(32'hbaa109e2),
	.w5(32'hbb859e82),
	.w6(32'hbb998964),
	.w7(32'hbc18d8d6),
	.w8(32'h3affbb46),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89512a),
	.w1(32'h38e9e160),
	.w2(32'h3b565b47),
	.w3(32'h3939c765),
	.w4(32'h3ac61a31),
	.w5(32'h395aa0e7),
	.w6(32'h3b0b4239),
	.w7(32'h3af251f9),
	.w8(32'h37c34514),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9030d3),
	.w1(32'h39d6d3c3),
	.w2(32'h3aa07862),
	.w3(32'hbb02b35d),
	.w4(32'hb9dc6717),
	.w5(32'hba3b4b1c),
	.w6(32'hb9c1a539),
	.w7(32'hbb12c144),
	.w8(32'hbb418ec3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02981b),
	.w1(32'hbb87574f),
	.w2(32'h3c67d3ca),
	.w3(32'h3bfd0146),
	.w4(32'h3b75d752),
	.w5(32'h3b4562c9),
	.w6(32'hbacd2b26),
	.w7(32'h3c2e8304),
	.w8(32'hbad015e3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069f5f),
	.w1(32'hbb251168),
	.w2(32'h3b7c86ef),
	.w3(32'h3b7d8638),
	.w4(32'h39f1ad3c),
	.w5(32'h397e6140),
	.w6(32'hbac09391),
	.w7(32'h3bc43274),
	.w8(32'hbb03fa11),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bce63),
	.w1(32'h3af8f338),
	.w2(32'h3a2f5626),
	.w3(32'hbb1381ef),
	.w4(32'hbab626f2),
	.w5(32'h3a223be5),
	.w6(32'hba60ad56),
	.w7(32'hbaf69353),
	.w8(32'h3b7bf633),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee5fb),
	.w1(32'hbc9e1fa3),
	.w2(32'hbb1a7a0e),
	.w3(32'h3c01079c),
	.w4(32'h3cf9b452),
	.w5(32'h3b606f41),
	.w6(32'h3c63de77),
	.w7(32'h3b8f0c0c),
	.w8(32'hbaf5c7b5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7861bf),
	.w1(32'hb90dc111),
	.w2(32'h3b3d4813),
	.w3(32'hbaae5de2),
	.w4(32'h3b4041ab),
	.w5(32'hba0147a9),
	.w6(32'hba6b8bbd),
	.w7(32'hbb7a54ed),
	.w8(32'hbc3505a3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8902),
	.w1(32'hbc17769c),
	.w2(32'hbadd2717),
	.w3(32'hbb80d468),
	.w4(32'hbaaf766a),
	.w5(32'hbb8850af),
	.w6(32'hbbda9782),
	.w7(32'hbbdb5418),
	.w8(32'hbc220329),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf69e5d),
	.w1(32'h3caaea49),
	.w2(32'hbbb1fbe7),
	.w3(32'h3affcd43),
	.w4(32'hbb68fd6b),
	.w5(32'hb9127918),
	.w6(32'h3b9b517d),
	.w7(32'hbbd509f1),
	.w8(32'hbae814f8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724138),
	.w1(32'hba8182ab),
	.w2(32'hba2622e7),
	.w3(32'hbb837395),
	.w4(32'hbaef4142),
	.w5(32'h3b3d78eb),
	.w6(32'hba81da34),
	.w7(32'h3b086a81),
	.w8(32'h3b0256f3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec4720),
	.w1(32'hbbb553bb),
	.w2(32'h3a593b69),
	.w3(32'h3b8baef1),
	.w4(32'h3af62acd),
	.w5(32'h3ad68d6b),
	.w6(32'hbaca1c16),
	.w7(32'h3aa81abe),
	.w8(32'h3c4ecc61),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b371536),
	.w1(32'h3ab5ae4e),
	.w2(32'h3b17ce77),
	.w3(32'h3b7a09fb),
	.w4(32'hb8b96510),
	.w5(32'h3c1a1cb6),
	.w6(32'h3b73de52),
	.w7(32'h3b5ee927),
	.w8(32'hbab32cff),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24aaf),
	.w1(32'hbb6a4a5f),
	.w2(32'h3ba8f928),
	.w3(32'h3c01dbab),
	.w4(32'h3c0fca56),
	.w5(32'h39650748),
	.w6(32'h3b118ac2),
	.w7(32'hbaa32256),
	.w8(32'hbca35f43),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3962e7),
	.w1(32'h3bff59b1),
	.w2(32'h3c0e4392),
	.w3(32'hbc52b183),
	.w4(32'h3b78a8a3),
	.w5(32'h3b8ed0ac),
	.w6(32'h3a003eef),
	.w7(32'hbaa27ec3),
	.w8(32'h3c40a804),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3745e0),
	.w1(32'h3ab7d36a),
	.w2(32'h3b0d3ffd),
	.w3(32'h3b7b6735),
	.w4(32'h38820ad4),
	.w5(32'h3c125afd),
	.w6(32'h3b71bff7),
	.w7(32'h3b59caa8),
	.w8(32'h3c22d0d3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22956e),
	.w1(32'h3aa6ddf2),
	.w2(32'h3af6c264),
	.w3(32'h3b5af5f0),
	.w4(32'h390e2b9b),
	.w5(32'h3bfd0e4b),
	.w6(32'h3b52a558),
	.w7(32'h3b41a1af),
	.w8(32'hbb976cd0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4619a6),
	.w1(32'hbc26c78a),
	.w2(32'hbbd1b0dd),
	.w3(32'hbc3af52b),
	.w4(32'hbc6ae531),
	.w5(32'hbc0d3b40),
	.w6(32'hbbfd22ba),
	.w7(32'hbb4654d1),
	.w8(32'hbbdb4191),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f09b),
	.w1(32'h3c35631a),
	.w2(32'hbbc02fd5),
	.w3(32'h3b9a60d2),
	.w4(32'h3b9365a9),
	.w5(32'h39a7fd72),
	.w6(32'h3b81e117),
	.w7(32'hbc00e6fc),
	.w8(32'h397eb095),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a761be5),
	.w1(32'hbae27d4a),
	.w2(32'h3ad9ecee),
	.w3(32'hb9bbdbf2),
	.w4(32'hb984f0a1),
	.w5(32'hb9815b7f),
	.w6(32'h3a1bcad2),
	.w7(32'h3ab9c886),
	.w8(32'hbc707c5e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b86e6),
	.w1(32'h3b08c6bc),
	.w2(32'h3af0a06d),
	.w3(32'hbc874021),
	.w4(32'hbbd6524a),
	.w5(32'hbc411016),
	.w6(32'hbc5a0215),
	.w7(32'hbb91dee3),
	.w8(32'hbb78bd21),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2032cf),
	.w1(32'hbb906be7),
	.w2(32'h3b5fe98f),
	.w3(32'hbc02a3e6),
	.w4(32'hb945480d),
	.w5(32'h3bbb10a6),
	.w6(32'h3ab6f8c3),
	.w7(32'h3b64d8ab),
	.w8(32'h3c30401a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b5cd7),
	.w1(32'h3c2307b2),
	.w2(32'h3c1c53cd),
	.w3(32'hbb42672c),
	.w4(32'h3c270d0c),
	.w5(32'hbbbab922),
	.w6(32'h3c97b026),
	.w7(32'h3c9a3031),
	.w8(32'hbc1ecd3a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc968944),
	.w1(32'hbc1b854a),
	.w2(32'hbd073256),
	.w3(32'hbcdb13b3),
	.w4(32'hbd5a7b48),
	.w5(32'hbcd19e7f),
	.w6(32'h3c561b29),
	.w7(32'hbc2250aa),
	.w8(32'hbb2bad78),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be583b7),
	.w1(32'hbb6b23b9),
	.w2(32'h3c4aca24),
	.w3(32'h3bdd59ab),
	.w4(32'h3b59d78c),
	.w5(32'h3b2cfd67),
	.w6(32'hbab2d7e1),
	.w7(32'h3c1944fe),
	.w8(32'hbb8237d7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17bbc3),
	.w1(32'hbab1cbe0),
	.w2(32'h3acb373b),
	.w3(32'h3afedd76),
	.w4(32'h3b5f21ba),
	.w5(32'hbb62aeaa),
	.w6(32'h355af51d),
	.w7(32'hbb56b5af),
	.w8(32'h3bd2ff60),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcca70a),
	.w1(32'h3b501a63),
	.w2(32'hba3622d4),
	.w3(32'h3bdb6260),
	.w4(32'h3b367de2),
	.w5(32'hbbc127a0),
	.w6(32'h3ba036bb),
	.w7(32'hbc0d307f),
	.w8(32'h3a10f743),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add2593),
	.w1(32'hbbc15e69),
	.w2(32'h3b42550f),
	.w3(32'h3a3a67d4),
	.w4(32'hb99f9542),
	.w5(32'h3aa556c8),
	.w6(32'hba082a97),
	.w7(32'h3b1b0119),
	.w8(32'hbabb30d8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b997a16),
	.w1(32'hbb5a76eb),
	.w2(32'h3b9b5d5f),
	.w3(32'h3c4dd71e),
	.w4(32'h3a99c4e8),
	.w5(32'h3a6d9a09),
	.w6(32'hbadd4a61),
	.w7(32'h3c3f9549),
	.w8(32'hbbce5e63),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36851e),
	.w1(32'hbba46b1a),
	.w2(32'hbb50dc5e),
	.w3(32'hbc2b532e),
	.w4(32'hbc0ec85d),
	.w5(32'hbbb4307f),
	.w6(32'hbb9be449),
	.w7(32'hbb1d4e76),
	.w8(32'h3b96db25),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a061988),
	.w1(32'h39c3361c),
	.w2(32'h3982d14d),
	.w3(32'h3a760a57),
	.w4(32'hb9aa46b9),
	.w5(32'h3b505586),
	.w6(32'h3a88b3c3),
	.w7(32'h3a382038),
	.w8(32'hb9c69173),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a116d2d),
	.w1(32'h3b79be69),
	.w2(32'h3a503376),
	.w3(32'hbaa35a00),
	.w4(32'h3a880059),
	.w5(32'h3a91587a),
	.w6(32'h3aa24f33),
	.w7(32'hbacdb3d6),
	.w8(32'hbb35a6d2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebf91c),
	.w1(32'hbb139281),
	.w2(32'h3ba9f375),
	.w3(32'hbb9ef4d3),
	.w4(32'h3b2bc7ea),
	.w5(32'h3bae020c),
	.w6(32'h3b113dcb),
	.w7(32'h3baa9a94),
	.w8(32'hbab5e454),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a760e14),
	.w1(32'h3bb153c9),
	.w2(32'h3b26f4f7),
	.w3(32'hba7d3202),
	.w4(32'h3b1c966b),
	.w5(32'h3abd9ce5),
	.w6(32'h3b2c1330),
	.w7(32'h3a2f30e9),
	.w8(32'hbb99b284),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e6b9),
	.w1(32'h3a1dbb26),
	.w2(32'hbabb92a8),
	.w3(32'hbb04d2f4),
	.w4(32'hb9c4f6c2),
	.w5(32'hba6c6cd0),
	.w6(32'hbb37e6fe),
	.w7(32'hbb661c3b),
	.w8(32'h39721796),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75563),
	.w1(32'h3a940454),
	.w2(32'h39da1456),
	.w3(32'h3b660b5c),
	.w4(32'hba363c3e),
	.w5(32'h3a1ce88e),
	.w6(32'h3a720f3b),
	.w7(32'h3b5a1dd0),
	.w8(32'hbc2ac6bb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb444a54),
	.w1(32'h3b5e9931),
	.w2(32'h3af8608b),
	.w3(32'h3b38b635),
	.w4(32'h3b4d9199),
	.w5(32'hbb674c7f),
	.w6(32'hbc07fcdb),
	.w7(32'hbb33ecfd),
	.w8(32'h3ba5b7ad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4363ee),
	.w1(32'h3b076e6d),
	.w2(32'h3b5c0999),
	.w3(32'h3b3c0c72),
	.w4(32'h3b1eb707),
	.w5(32'h3be12131),
	.w6(32'h3b2d8f29),
	.w7(32'h3b80df05),
	.w8(32'hbab42ca4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd981b5),
	.w1(32'hbc222939),
	.w2(32'hbb1c52aa),
	.w3(32'hbb74477b),
	.w4(32'hbbaf7a6b),
	.w5(32'h3972e7ea),
	.w6(32'hbb5976fc),
	.w7(32'h3a958f0d),
	.w8(32'hbb9fccaa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18ad00),
	.w1(32'hb8bc9105),
	.w2(32'hbac270af),
	.w3(32'hbb1d70af),
	.w4(32'hbae8b33a),
	.w5(32'hba88a31c),
	.w6(32'hbb4c14ed),
	.w7(32'hbb2ada47),
	.w8(32'h3a794b0e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bde7b),
	.w1(32'h3b698d3e),
	.w2(32'h3af7d98e),
	.w3(32'h3b03f666),
	.w4(32'h3b142113),
	.w5(32'h3a90e0b2),
	.w6(32'h3ade8355),
	.w7(32'h3a85bada),
	.w8(32'h3b344c2e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc454b8),
	.w1(32'h3c0749f7),
	.w2(32'h3b882e75),
	.w3(32'h3b7ea28c),
	.w4(32'h3ba6097f),
	.w5(32'h3b296879),
	.w6(32'h3b8eb5a4),
	.w7(32'h3ad3be49),
	.w8(32'h3c0ac8aa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b8d01),
	.w1(32'hbc055d8b),
	.w2(32'hbb0a5598),
	.w3(32'h3c1cd773),
	.w4(32'h3a99a6d6),
	.w5(32'hb9fba5bf),
	.w6(32'hbb220d5b),
	.w7(32'hbb441628),
	.w8(32'hbacc22d5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4916b9),
	.w1(32'hbb33e5c6),
	.w2(32'hbb159218),
	.w3(32'hbb232672),
	.w4(32'hbb63a071),
	.w5(32'hbb3fe617),
	.w6(32'hbb1fdce9),
	.w7(32'hbaed713f),
	.w8(32'hbaf07d40),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6dbde),
	.w1(32'h3b1554ea),
	.w2(32'h3ac99186),
	.w3(32'hbb1bdd76),
	.w4(32'h3c0af207),
	.w5(32'h3b3205fd),
	.w6(32'h3b8cb86b),
	.w7(32'h3b6a3dde),
	.w8(32'hbac9b832),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b683020),
	.w1(32'hbaab2a15),
	.w2(32'hbb9a77be),
	.w3(32'h3a7594a3),
	.w4(32'hba166857),
	.w5(32'hbac52fab),
	.w6(32'hbb3ea8f5),
	.w7(32'h3965316b),
	.w8(32'hbc1ba44e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6b6f4),
	.w1(32'h39f98372),
	.w2(32'hbafd075c),
	.w3(32'hbb29a44a),
	.w4(32'hbb44c843),
	.w5(32'hbbbc656b),
	.w6(32'h3954d24d),
	.w7(32'h3aeb53ee),
	.w8(32'h3b331b1a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8443b0),
	.w1(32'h3bcaa6aa),
	.w2(32'h3a55e67b),
	.w3(32'hbc750ba2),
	.w4(32'h3b19e607),
	.w5(32'h3b462c53),
	.w6(32'hba3dfcab),
	.w7(32'hbbef598c),
	.w8(32'h3903ca9c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd11c),
	.w1(32'h3a141ccc),
	.w2(32'h3b430c11),
	.w3(32'h3aac8744),
	.w4(32'h3ae2c441),
	.w5(32'h3b88ca60),
	.w6(32'h3a2c1d09),
	.w7(32'h3af30b5e),
	.w8(32'hbbade62b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1f98b),
	.w1(32'hbbbf3e07),
	.w2(32'hbb681274),
	.w3(32'hbbe996a0),
	.w4(32'hbbcff810),
	.w5(32'hbb3e8923),
	.w6(32'hbb9c213b),
	.w7(32'hbb838245),
	.w8(32'hbc095c37),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14eed7),
	.w1(32'hbbae607e),
	.w2(32'hbb9f7b02),
	.w3(32'h3b77f666),
	.w4(32'h3b8a6abb),
	.w5(32'hba8c7b06),
	.w6(32'hbb945d2c),
	.w7(32'h39498f35),
	.w8(32'h3a44f18c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183682),
	.w1(32'h3b1ad930),
	.w2(32'h3b93ee32),
	.w3(32'h3bca29d4),
	.w4(32'h3b63d263),
	.w5(32'h3be050a9),
	.w6(32'h3ab040ed),
	.w7(32'h3b9e4189),
	.w8(32'hb9f1a917),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55853),
	.w1(32'h3957bb6c),
	.w2(32'h3b2f5845),
	.w3(32'h3b143afb),
	.w4(32'hb8922ad9),
	.w5(32'h3b2f4797),
	.w6(32'hb9ef80af),
	.w7(32'h3b6791f2),
	.w8(32'h3bf0bf13),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70c62f),
	.w1(32'h3af37798),
	.w2(32'h3becbd7b),
	.w3(32'hbc09ca5e),
	.w4(32'hba4c2c12),
	.w5(32'h3b9a35b9),
	.w6(32'h3b84e938),
	.w7(32'h3b4f3a1d),
	.w8(32'hbaf29819),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdd03a),
	.w1(32'h3b20f19e),
	.w2(32'h3ad7d26c),
	.w3(32'hba290d0f),
	.w4(32'h3aa26240),
	.w5(32'h3ab1f627),
	.w6(32'h3ae54a8a),
	.w7(32'h3a7011c7),
	.w8(32'h39a9763d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dc2b5),
	.w1(32'h3bb410d1),
	.w2(32'h3b0f40a9),
	.w3(32'h3a1a61f5),
	.w4(32'h3b30d735),
	.w5(32'h3a97f1a3),
	.w6(32'h3b3c4719),
	.w7(32'h39ac780d),
	.w8(32'h393b1bc2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1cc15),
	.w1(32'h3b22c6bc),
	.w2(32'h3a630054),
	.w3(32'h3a88d5cd),
	.w4(32'h3acadc4c),
	.w5(32'h3a04c0fa),
	.w6(32'h3aa2d5af),
	.w7(32'h38f09a45),
	.w8(32'hbb74d270),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94ddb8),
	.w1(32'h3ab43cb8),
	.w2(32'h3b2b8cf5),
	.w3(32'h39b11699),
	.w4(32'h3a9d98da),
	.w5(32'h3b5c78d9),
	.w6(32'hbb3332f4),
	.w7(32'hbb310f46),
	.w8(32'hbb828268),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf09cb3),
	.w1(32'hb943121c),
	.w2(32'hbacfc395),
	.w3(32'hbb1bfcfb),
	.w4(32'hbada71c0),
	.w5(32'hbaa66c7a),
	.w6(32'hbb3d2ae3),
	.w7(32'hbb4aa119),
	.w8(32'h3a84991e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122650),
	.w1(32'h3c472b97),
	.w2(32'h3c02bd89),
	.w3(32'h3bd4bd27),
	.w4(32'h3c1574a9),
	.w5(32'h3bed488e),
	.w6(32'h3b85175e),
	.w7(32'h3b07c537),
	.w8(32'hba47915c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4da963),
	.w1(32'h3b825147),
	.w2(32'h3a9a712e),
	.w3(32'hba581998),
	.w4(32'h3ac42961),
	.w5(32'h3a41053b),
	.w6(32'h3aaa10c0),
	.w7(32'hbab35e1d),
	.w8(32'hbb943eb7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca2e7),
	.w1(32'hbac0b770),
	.w2(32'hbb3004fb),
	.w3(32'hbb659394),
	.w4(32'hbb1e9a01),
	.w5(32'hbaad63c2),
	.w6(32'hbb62f613),
	.w7(32'hbb81f49e),
	.w8(32'hb96c57f7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67030f),
	.w1(32'h3bf57249),
	.w2(32'h3b070a5e),
	.w3(32'h3a132d1e),
	.w4(32'h3b5f9406),
	.w5(32'h39f147e2),
	.w6(32'h3b457902),
	.w7(32'hba89be02),
	.w8(32'hbbaf0d61),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac94dd),
	.w1(32'h3b91e373),
	.w2(32'hbb565d87),
	.w3(32'h3b9a3dd6),
	.w4(32'h3bae8787),
	.w5(32'h3adf24b7),
	.w6(32'hbc22237a),
	.w7(32'hbc4405d6),
	.w8(32'hbaab613a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949a4db),
	.w1(32'h3a46ef54),
	.w2(32'hba8aa6a9),
	.w3(32'hba5caba2),
	.w4(32'hba8430b9),
	.w5(32'hba9ad939),
	.w6(32'hbac27841),
	.w7(32'hbb2a756f),
	.w8(32'hb89126e9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa17f22),
	.w1(32'h3b87a914),
	.w2(32'h3af87afb),
	.w3(32'h389e1c43),
	.w4(32'h3b00cdd2),
	.w5(32'h3ab2eaef),
	.w6(32'h3b1404d1),
	.w7(32'h3a023f78),
	.w8(32'hb90a28f1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a822b49),
	.w1(32'h3b437cad),
	.w2(32'h39f2260d),
	.w3(32'h399608ce),
	.w4(32'h3a94682b),
	.w5(32'h3a024350),
	.w6(32'h3a75c889),
	.w7(32'hbaa17b2d),
	.w8(32'h3a8acde7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21b3fb),
	.w1(32'h3c5aebc0),
	.w2(32'h3c178baf),
	.w3(32'h3bf337d2),
	.w4(32'h3c289998),
	.w5(32'h3c10deb0),
	.w6(32'h3b91c171),
	.w7(32'h3b2ece18),
	.w8(32'hba0fd8e5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1a9d0),
	.w1(32'h3be4d609),
	.w2(32'h3b386eac),
	.w3(32'h3b38b8e4),
	.w4(32'h3b87c2f4),
	.w5(32'h3b0e32b3),
	.w6(32'h3a658904),
	.w7(32'hb9e665ca),
	.w8(32'hbaca1cec),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a658),
	.w1(32'h3b0359a2),
	.w2(32'h39af86d5),
	.w3(32'hbad09e1c),
	.w4(32'hb92c877e),
	.w5(32'h39d8d4c3),
	.w6(32'h3ac76bb3),
	.w7(32'hb9fbc084),
	.w8(32'hbbc00436),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba020339),
	.w1(32'h3a1becef),
	.w2(32'hbb0f67e9),
	.w3(32'h3c0f0aab),
	.w4(32'h3bff7f8b),
	.w5(32'h3c0a6257),
	.w6(32'hbb1fd51f),
	.w7(32'hbbc9e5ea),
	.w8(32'h397c4e6b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cf9a9),
	.w1(32'h3ad95efc),
	.w2(32'h3aed00dd),
	.w3(32'h3ad36ef7),
	.w4(32'h3a8f87c5),
	.w5(32'h3ad9a8af),
	.w6(32'h3ac7216c),
	.w7(32'h3b1c8a5f),
	.w8(32'hbbc97d2a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d5ad),
	.w1(32'h38fe21fd),
	.w2(32'hbaaf0740),
	.w3(32'hbaa63f9d),
	.w4(32'hb9c9c8e2),
	.w5(32'hb98278f8),
	.w6(32'hbabe26a8),
	.w7(32'hba7ede42),
	.w8(32'h3b3a0cd1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4a8a1),
	.w1(32'h3b2e5d44),
	.w2(32'h3b5061f3),
	.w3(32'h3b7b963e),
	.w4(32'hbac05ff6),
	.w5(32'h3a9abe76),
	.w6(32'h3c06062c),
	.w7(32'h3c07c3d4),
	.w8(32'hbafd24e5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb235763),
	.w1(32'hbb32c677),
	.w2(32'hbb0ed8fb),
	.w3(32'hbb1d2cde),
	.w4(32'hbb4ee301),
	.w5(32'hbb3c7073),
	.w6(32'hbb1c0e66),
	.w7(32'hbb0cdca6),
	.w8(32'hbb956260),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7448c),
	.w1(32'hb883b280),
	.w2(32'hbac4b7a9),
	.w3(32'hbb0ef02c),
	.w4(32'hba9cc94e),
	.w5(32'hba29c4b7),
	.w6(32'hbb6578d5),
	.w7(32'hbb5afee8),
	.w8(32'hbadd7a84),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc90b),
	.w1(32'hbc5718c9),
	.w2(32'hbb4f3ea6),
	.w3(32'hbba13a5c),
	.w4(32'hbbe89f37),
	.w5(32'h39a5cb11),
	.w6(32'hbb90a340),
	.w7(32'h3ac21ac0),
	.w8(32'h39dfaffa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab3896),
	.w1(32'h3a2fa90d),
	.w2(32'h3a6b9d4d),
	.w3(32'h3a0ea4dc),
	.w4(32'hb9e2db4e),
	.w5(32'h3abb3139),
	.w6(32'h3b053e73),
	.w7(32'h3a93814c),
	.w8(32'hbb5ff7d8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad4a3),
	.w1(32'hbc0973be),
	.w2(32'hbb727c6b),
	.w3(32'hbbc1c875),
	.w4(32'hbc110d73),
	.w5(32'hbbdb1760),
	.w6(32'hbb63c831),
	.w7(32'hbb75b351),
	.w8(32'hbad4e8bd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067f23),
	.w1(32'hbc48d3b5),
	.w2(32'hbb3fa5ac),
	.w3(32'hbb96f845),
	.w4(32'hbbd8d502),
	.w5(32'h39ad0b36),
	.w6(32'hbb8703ca),
	.w7(32'h3ab8bdd2),
	.w8(32'hbaaf6196),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe572df),
	.w1(32'hbc2b73fb),
	.w2(32'hbb2897af),
	.w3(32'hbb81641a),
	.w4(32'hbbbb2855),
	.w5(32'h396f1a18),
	.w6(32'hbb663c32),
	.w7(32'h3a9e28f7),
	.w8(32'hbb1dabaa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f22e9),
	.w1(32'hbb3620df),
	.w2(32'hbb8b7902),
	.w3(32'hbb68f05a),
	.w4(32'hbb8cfecd),
	.w5(32'hbba525fc),
	.w6(32'hbb4895af),
	.w7(32'hbb83e20a),
	.w8(32'hbbbe5248),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1413f1),
	.w1(32'hbbc72631),
	.w2(32'hbb965872),
	.w3(32'hbbfcf3d8),
	.w4(32'hbb68f037),
	.w5(32'hbaa1d4f2),
	.w6(32'h387222a3),
	.w7(32'hbba8e51f),
	.w8(32'h3a476a8e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5a0b4),
	.w1(32'h3b2efcf0),
	.w2(32'h3abb5672),
	.w3(32'h3aae62aa),
	.w4(32'h3add7f25),
	.w5(32'h3a6ca3bb),
	.w6(32'h3aa93417),
	.w7(32'h3a375ac6),
	.w8(32'hb9e1c973),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06e1c5),
	.w1(32'hbaf4e5ff),
	.w2(32'hbaefd3c8),
	.w3(32'hbba170b7),
	.w4(32'hbbb9e6e5),
	.w5(32'hbbc8f03a),
	.w6(32'hbb0a6b2d),
	.w7(32'hb90aa99d),
	.w8(32'hbb20aa87),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2815e),
	.w1(32'hbbdc85cc),
	.w2(32'hbb932ffc),
	.w3(32'hbbc4b2af),
	.w4(32'hbbe8dab6),
	.w5(32'hbbbc6e80),
	.w6(32'hbb896932),
	.w7(32'hbb557a7b),
	.w8(32'h3b7626d1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947adb),
	.w1(32'h3b373594),
	.w2(32'h3b20512f),
	.w3(32'h3b7034c4),
	.w4(32'h3b31da47),
	.w5(32'h3b8071dd),
	.w6(32'h3b80ad41),
	.w7(32'h3bb9b244),
	.w8(32'h3b3505e7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd60cd),
	.w1(32'hbb2d213d),
	.w2(32'hbb8cc43c),
	.w3(32'hbc3bc4c6),
	.w4(32'hbc427f9c),
	.w5(32'hbc20c7be),
	.w6(32'h3b5f4a5d),
	.w7(32'h3b57a3fc),
	.w8(32'h3a74462a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100cac),
	.w1(32'h3c419ed0),
	.w2(32'h3c05d348),
	.w3(32'h3bdb3b65),
	.w4(32'h3c1664f2),
	.w5(32'h3c011c07),
	.w6(32'h3b83ee15),
	.w7(32'h3b218402),
	.w8(32'hbb378691),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9591fcd),
	.w1(32'h3b39a93a),
	.w2(32'h3a54e469),
	.w3(32'hbaa3d5cc),
	.w4(32'h3a153c4a),
	.w5(32'h3a324547),
	.w6(32'h3b2d9cda),
	.w7(32'h3a136d03),
	.w8(32'hbb371ca1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfe618),
	.w1(32'hbb9ae07e),
	.w2(32'hbb62163b),
	.w3(32'hbbb7ed93),
	.w4(32'hbbd2d86e),
	.w5(32'hbb6c631b),
	.w6(32'hbb3cd268),
	.w7(32'hbac2ac11),
	.w8(32'h3a602b84),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a352d),
	.w1(32'h3b766402),
	.w2(32'h3aeb6f5d),
	.w3(32'h3b1e38ae),
	.w4(32'h3b2ec529),
	.w5(32'h3aa3f37e),
	.w6(32'h3aebc6f8),
	.w7(32'h3a860254),
	.w8(32'hbac4b4c4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c088c7d),
	.w1(32'h3c4528e5),
	.w2(32'h3b5d2bea),
	.w3(32'h3b818db2),
	.w4(32'h3bc14f5f),
	.w5(32'h3af572cd),
	.w6(32'h3914c48b),
	.w7(32'hbadace28),
	.w8(32'hbb3ad0bf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb606eed),
	.w1(32'hbb838905),
	.w2(32'hbb959596),
	.w3(32'hbb94abbe),
	.w4(32'hbbae9f89),
	.w5(32'hbbad543e),
	.w6(32'hbb79c1ef),
	.w7(32'hbb93a23e),
	.w8(32'hba212ed9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee549),
	.w1(32'hbba593f0),
	.w2(32'hbab371df),
	.w3(32'hbb009e37),
	.w4(32'hbb383c9f),
	.w5(32'hb8e9758e),
	.w6(32'hbadea114),
	.w7(32'h39fe9e74),
	.w8(32'h380187ed),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8c4a0),
	.w1(32'hb893ead8),
	.w2(32'hb75ef70f),
	.w3(32'hb8eb7f5f),
	.w4(32'hb89fc58d),
	.w5(32'hb85c8514),
	.w6(32'hb88892db),
	.w7(32'hb8a96398),
	.w8(32'hb881d4d6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a53cac),
	.w1(32'h37a3aae9),
	.w2(32'h3808370e),
	.w3(32'hb798cb05),
	.w4(32'hb7638942),
	.w5(32'h38133ab3),
	.w6(32'hb76edac5),
	.w7(32'hb76c402b),
	.w8(32'h37931b3b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d3424e),
	.w1(32'h37d0ed22),
	.w2(32'h376fc473),
	.w3(32'h37aa68b1),
	.w4(32'h372104da),
	.w5(32'h37acdc6a),
	.w6(32'h37a7c007),
	.w7(32'h37cf23af),
	.w8(32'h380e49da),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b235e6),
	.w1(32'h3803d46f),
	.w2(32'h382fbc3e),
	.w3(32'h37c199f2),
	.w4(32'h3824cc25),
	.w5(32'h383ae759),
	.w6(32'h37da68c2),
	.w7(32'h386ff491),
	.w8(32'h386f25ed),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7025ff2),
	.w1(32'h36993c00),
	.w2(32'h37db1230),
	.w3(32'hb80618f9),
	.w4(32'hb84e8178),
	.w5(32'hb458bf59),
	.w6(32'hb7539ae9),
	.w7(32'hb7b4cf31),
	.w8(32'h367be583),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84bb598),
	.w1(32'hb6cf82f8),
	.w2(32'hb863590f),
	.w3(32'hb8217de3),
	.w4(32'hb849b835),
	.w5(32'hb85e3229),
	.w6(32'hb793e7c3),
	.w7(32'hb7bb5cde),
	.w8(32'hb89f705f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7937e3c),
	.w1(32'hb80eb4c6),
	.w2(32'hb8353785),
	.w3(32'hb7eda7aa),
	.w4(32'hb81afc38),
	.w5(32'hb82f4e35),
	.w6(32'h350d179b),
	.w7(32'h3685581c),
	.w8(32'h36954d9a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70b6dbf),
	.w1(32'h36897a17),
	.w2(32'h37cfea3d),
	.w3(32'h369434e5),
	.w4(32'h3806e6a1),
	.w5(32'h383563af),
	.w6(32'h37bcf54d),
	.w7(32'h389d021f),
	.w8(32'h38a06fb1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5913e8d),
	.w1(32'h3664da5e),
	.w2(32'h365aefa0),
	.w3(32'hb556b7e5),
	.w4(32'h36929118),
	.w5(32'h36574b69),
	.w6(32'hb5c52046),
	.w7(32'h33d8957d),
	.w8(32'h369cd6ef),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c90947),
	.w1(32'hb713876e),
	.w2(32'hb7d4c971),
	.w3(32'hb76b8a3c),
	.w4(32'hb7118ce3),
	.w5(32'hb75ee447),
	.w6(32'hb7a37343),
	.w7(32'hb7c805ca),
	.w8(32'hb70520e0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ecb478),
	.w1(32'hb832699d),
	.w2(32'hb818d5c9),
	.w3(32'hb828ce67),
	.w4(32'hb879981e),
	.w5(32'hb80af179),
	.w6(32'hb718ad39),
	.w7(32'hb82eb83b),
	.w8(32'hb7de932c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77a84b4),
	.w1(32'hb7c02493),
	.w2(32'hb74c9fe4),
	.w3(32'hb701c175),
	.w4(32'hb798b9b5),
	.w5(32'hb73071f8),
	.w6(32'h36d178f0),
	.w7(32'h38018fea),
	.w8(32'h3750ea7e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e04b01),
	.w1(32'hb8a18b57),
	.w2(32'hb8986fd6),
	.w3(32'hb90e1e9b),
	.w4(32'hb8e47444),
	.w5(32'hb8beae98),
	.w6(32'hb8b9db24),
	.w7(32'hb89809d8),
	.w8(32'hb8927781),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb704de71),
	.w1(32'h371ac837),
	.w2(32'hb65f74af),
	.w3(32'hb70eff58),
	.w4(32'h37070e3d),
	.w5(32'hb5fb5232),
	.w6(32'h370a8f5e),
	.w7(32'hb65e6762),
	.w8(32'hb368ef7b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb706c238),
	.w1(32'hb730fec2),
	.w2(32'hb7620f6a),
	.w3(32'hb78ebedd),
	.w4(32'hb7b056b6),
	.w5(32'hb788563a),
	.w6(32'hb77886dd),
	.w7(32'hb7634deb),
	.w8(32'hb716e881),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b6407c),
	.w1(32'hb84307db),
	.w2(32'hb7bbc993),
	.w3(32'hb804854d),
	.w4(32'hb8299514),
	.w5(32'hb7587996),
	.w6(32'hb807aeb3),
	.w7(32'hb85a5264),
	.w8(32'hb8968c1d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69d9dc1),
	.w1(32'h372b4346),
	.w2(32'h3702b13d),
	.w3(32'hb6a055aa),
	.w4(32'hb6ef143b),
	.w5(32'h370e135a),
	.w6(32'h3738afd9),
	.w7(32'h3386432a),
	.w8(32'hb66b65ea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3774304a),
	.w1(32'h36f8ebc3),
	.w2(32'h369f433e),
	.w3(32'h376a97cb),
	.w4(32'h36dc7006),
	.w5(32'h369cbd20),
	.w6(32'h37b505a1),
	.w7(32'h35e3802a),
	.w8(32'hb60842f0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82dccd9),
	.w1(32'hb83acd75),
	.w2(32'hb7d536be),
	.w3(32'hb819537a),
	.w4(32'hb7e62bb2),
	.w5(32'hb785fca8),
	.w6(32'hb749b6a5),
	.w7(32'hb6ae505e),
	.w8(32'h36b4845c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37849fa3),
	.w1(32'h36648762),
	.w2(32'hb65151ad),
	.w3(32'h370f77bc),
	.w4(32'hb6a77f34),
	.w5(32'hb71a78f7),
	.w6(32'h375f0df9),
	.w7(32'hb42ea95b),
	.w8(32'hb7395f52),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5634d),
	.w1(32'h3618f8b1),
	.w2(32'hb7e16265),
	.w3(32'hb7954a23),
	.w4(32'hb7b312c9),
	.w5(32'hb871654b),
	.w6(32'hb7d4063b),
	.w7(32'hb7fc2c16),
	.w8(32'hb7dc4125),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acf096),
	.w1(32'hb8789123),
	.w2(32'hb86dac5f),
	.w3(32'hb8a2a5b9),
	.w4(32'hb89eede5),
	.w5(32'hb86200e1),
	.w6(32'hb882843a),
	.w7(32'hb8957a33),
	.w8(32'hb87d5b54),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869af40),
	.w1(32'hb8125a65),
	.w2(32'hb6a59eaf),
	.w3(32'hb8784100),
	.w4(32'hb87466ee),
	.w5(32'hb850eaca),
	.w6(32'hb7a53a45),
	.w7(32'hb8354256),
	.w8(32'hb7ca8cf0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule