module layer_6_featuremap_11(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a841),
	.w1(32'hbb10f096),
	.w2(32'hb9baf5ee),
	.w3(32'h3b82e5a3),
	.w4(32'h3b26e578),
	.w5(32'h3be606c2),
	.w6(32'hbbeb68e7),
	.w7(32'hbc0ec6f6),
	.w8(32'hbc40ab54),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891717),
	.w1(32'hbbb6b0e7),
	.w2(32'hbab4c869),
	.w3(32'h3c204798),
	.w4(32'hbc089a6c),
	.w5(32'hbb431dd1),
	.w6(32'hbbcf5d2b),
	.w7(32'hbba30699),
	.w8(32'hbb8fa201),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92a4b9),
	.w1(32'h3c7ab5c9),
	.w2(32'hbade36db),
	.w3(32'hbb6980d1),
	.w4(32'h3c009d41),
	.w5(32'h3b99f99c),
	.w6(32'hbb2ce1fc),
	.w7(32'hbc3b37f5),
	.w8(32'hbc53442a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe58e6a),
	.w1(32'hb9bf8eed),
	.w2(32'h3ba4b456),
	.w3(32'hbac53ba0),
	.w4(32'h3b9081ee),
	.w5(32'h3b45ba33),
	.w6(32'h3c1d457d),
	.w7(32'h3b94bb56),
	.w8(32'h3c415fad),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefcaa1),
	.w1(32'h3cc5d86e),
	.w2(32'h3d63d632),
	.w3(32'h3be9beb6),
	.w4(32'h3cb91ff7),
	.w5(32'h3d3efb87),
	.w6(32'h3c543258),
	.w7(32'h3d0d2a93),
	.w8(32'h3d187470),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5fc72e),
	.w1(32'hba9487da),
	.w2(32'hbbae50d7),
	.w3(32'h3d31e93a),
	.w4(32'h3b7ff26c),
	.w5(32'hb918f485),
	.w6(32'h3b6e3d8c),
	.w7(32'hbb033846),
	.w8(32'h3bbff9d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8697b),
	.w1(32'hb9c94649),
	.w2(32'h3a1d8a15),
	.w3(32'h3b3a6fbb),
	.w4(32'hbad5a6f6),
	.w5(32'hba1bc80a),
	.w6(32'hbb2da193),
	.w7(32'hbaf461bc),
	.w8(32'hbb818b6b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d2f3),
	.w1(32'h3ba2801c),
	.w2(32'h3b2af708),
	.w3(32'hbb3a9087),
	.w4(32'hbae96e6d),
	.w5(32'hbbcac107),
	.w6(32'hbbe73a68),
	.w7(32'hbc1c5593),
	.w8(32'hbc0141f5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb3648),
	.w1(32'h3c4132a7),
	.w2(32'h3c366a96),
	.w3(32'hbc246acf),
	.w4(32'h3c2eee63),
	.w5(32'h3c09546c),
	.w6(32'h3bd21bb6),
	.w7(32'h3b50cd11),
	.w8(32'h3a1fbb43),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fd6c6),
	.w1(32'hba221d0b),
	.w2(32'h392b1313),
	.w3(32'h39bb33ac),
	.w4(32'h394a9384),
	.w5(32'h3a689119),
	.w6(32'hba8f3e38),
	.w7(32'h3ab5e1ac),
	.w8(32'h3b1ccbbe),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61619b),
	.w1(32'h3c9b2ceb),
	.w2(32'h3c67bdf6),
	.w3(32'h3c044759),
	.w4(32'h3c97774a),
	.w5(32'h3c9cd04b),
	.w6(32'h3c103576),
	.w7(32'h3bc21487),
	.w8(32'h3c109659),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91054b),
	.w1(32'h3b13307e),
	.w2(32'h3bbaa553),
	.w3(32'hbacbb1b8),
	.w4(32'hbafecc24),
	.w5(32'h3c674be2),
	.w6(32'h3bb2de14),
	.w7(32'hbbab3177),
	.w8(32'hbbeea410),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a1c22),
	.w1(32'hba891d8e),
	.w2(32'h3c0810af),
	.w3(32'h3c08e72b),
	.w4(32'h3b31c1bb),
	.w5(32'h3c0724b4),
	.w6(32'h3934a968),
	.w7(32'h3b8a1cbd),
	.w8(32'h3b2e87a2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0feaa),
	.w1(32'h3cac7e75),
	.w2(32'h3c590941),
	.w3(32'h3b997566),
	.w4(32'h3c2eb692),
	.w5(32'h3be6fe23),
	.w6(32'h3c41010c),
	.w7(32'h3c0896e5),
	.w8(32'h3c39a12a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea27b3),
	.w1(32'hbc086d44),
	.w2(32'hbc0537d2),
	.w3(32'hbb5698f9),
	.w4(32'h3b63db82),
	.w5(32'h3b18027b),
	.w6(32'hbbef9d1f),
	.w7(32'hbb7243b3),
	.w8(32'h3c172b6b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f99ac),
	.w1(32'h3b88c793),
	.w2(32'hbb16209d),
	.w3(32'h3c01a9fa),
	.w4(32'h3b463226),
	.w5(32'hbb1c84e9),
	.w6(32'h3c57a1d4),
	.w7(32'h3c2e52e6),
	.w8(32'h3c4ef534),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16af1a),
	.w1(32'h3c08d325),
	.w2(32'hbb5f31b2),
	.w3(32'h3b32efd1),
	.w4(32'h3cb48c89),
	.w5(32'h3cbd1fd6),
	.w6(32'hbb63aef8),
	.w7(32'h3c47291c),
	.w8(32'h3c462b65),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed413d),
	.w1(32'h3c71c6ba),
	.w2(32'h3a472daf),
	.w3(32'h3b959eb1),
	.w4(32'h3c4abb73),
	.w5(32'hba885822),
	.w6(32'h3c3f70ef),
	.w7(32'h38e8db96),
	.w8(32'hbc8c4217),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4273f),
	.w1(32'h3c244f00),
	.w2(32'h3c62908b),
	.w3(32'hbcb24b26),
	.w4(32'h3bddc7a3),
	.w5(32'h3be4956b),
	.w6(32'h3b2e8ebb),
	.w7(32'h3bb0c0cc),
	.w8(32'h3b261dd7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c7646),
	.w1(32'h3a4f8cdd),
	.w2(32'h3aa68f8f),
	.w3(32'h3c10b642),
	.w4(32'hbb356106),
	.w5(32'h3b3aa451),
	.w6(32'h3a161b30),
	.w7(32'hba3c4997),
	.w8(32'hbb9e5e92),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7faa),
	.w1(32'hbb42ae6b),
	.w2(32'hbbbadb52),
	.w3(32'hbacf2b87),
	.w4(32'h3b5a4f83),
	.w5(32'hbb2acb81),
	.w6(32'hbaa325d5),
	.w7(32'hbb923287),
	.w8(32'hbb1259fb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf37f6),
	.w1(32'h3d056e18),
	.w2(32'h3d5262d7),
	.w3(32'hbba12ed3),
	.w4(32'h3cf33d9c),
	.w5(32'h3d30d848),
	.w6(32'h3c6c7fba),
	.w7(32'h3cd029a6),
	.w8(32'h3cf28285),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03b96e),
	.w1(32'hbb3ebfcb),
	.w2(32'hbb5b6f4b),
	.w3(32'h3ccddeb5),
	.w4(32'hbba3b535),
	.w5(32'hbb697f4f),
	.w6(32'hbb207bee),
	.w7(32'hbc2cf753),
	.w8(32'hbc8bcae3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756ebd),
	.w1(32'h3cc211c4),
	.w2(32'h3c08ca93),
	.w3(32'hbb98afd1),
	.w4(32'h3c8eb5f7),
	.w5(32'h3d05fe87),
	.w6(32'h3c8b68dc),
	.w7(32'h3beaeae7),
	.w8(32'h3c8acaab),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c841b9c),
	.w1(32'h3b74f4d9),
	.w2(32'hba4c3f13),
	.w3(32'h3ca22141),
	.w4(32'h3c68f2bc),
	.w5(32'h3b256d20),
	.w6(32'hbbf0ea45),
	.w7(32'hbbc034c5),
	.w8(32'h3afb4434),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a075570),
	.w1(32'h3a89f32f),
	.w2(32'hbb5eda32),
	.w3(32'h3c1d5358),
	.w4(32'h3badfbaf),
	.w5(32'h3bdd3e4d),
	.w6(32'h3afa22e5),
	.w7(32'hbb21fa64),
	.w8(32'h3b8a4602),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3617fe),
	.w1(32'h3b4ee95b),
	.w2(32'hbba7735b),
	.w3(32'h3c1a6be0),
	.w4(32'h3b69ef2b),
	.w5(32'h3bc7ef6e),
	.w6(32'h3c26843c),
	.w7(32'hbb0bbf84),
	.w8(32'hbb5c4acb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c7f9),
	.w1(32'h398fb4e5),
	.w2(32'hbc28afe9),
	.w3(32'h3bacd164),
	.w4(32'h3c11b722),
	.w5(32'h3a0f3c7f),
	.w6(32'h3ac0bf63),
	.w7(32'hbc15492d),
	.w8(32'h3b1ef1af),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b49fa),
	.w1(32'h3b0829c8),
	.w2(32'hb9f5f824),
	.w3(32'h3b2b8942),
	.w4(32'h3b9daca8),
	.w5(32'h3b867dad),
	.w6(32'hbb9a6039),
	.w7(32'hbafe9dc4),
	.w8(32'h3c010c81),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36d9a4),
	.w1(32'h3a67e4b1),
	.w2(32'hbc402fdd),
	.w3(32'h3d8e9ae3),
	.w4(32'hbc88c706),
	.w5(32'hbd77bc96),
	.w6(32'hbc2efeb0),
	.w7(32'hbcb5573d),
	.w8(32'hbc065966),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1478a9),
	.w1(32'h3b7e3956),
	.w2(32'hbc117543),
	.w3(32'hbc1fd146),
	.w4(32'h3c2ec4f5),
	.w5(32'hbc9ae404),
	.w6(32'h3cb694d2),
	.w7(32'h3c0df6d6),
	.w8(32'h3b0ea728),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb418ec),
	.w1(32'hbb6c5f05),
	.w2(32'h3ce2254d),
	.w3(32'h3c48523d),
	.w4(32'hbb72864a),
	.w5(32'hbc22c398),
	.w6(32'hbb64fad3),
	.w7(32'hba991cd4),
	.w8(32'h3c3f5c60),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451787),
	.w1(32'hba075efc),
	.w2(32'hbbe98b79),
	.w3(32'h3c1c60de),
	.w4(32'hbc35a27e),
	.w5(32'h3bbba9db),
	.w6(32'h3cb867c9),
	.w7(32'hbb90c6f0),
	.w8(32'hbc09b8f4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0ad05),
	.w1(32'h3d256e8c),
	.w2(32'h3aa03179),
	.w3(32'h3b4447c9),
	.w4(32'hb8ac6a92),
	.w5(32'h38fb9d3a),
	.w6(32'hbc1b42dd),
	.w7(32'hbc10b1d9),
	.w8(32'hbbb50608),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8e515),
	.w1(32'hbc3662f6),
	.w2(32'hbc9f93b6),
	.w3(32'h3ad8c36b),
	.w4(32'hbc74d268),
	.w5(32'hbcce9a60),
	.w6(32'hbc8cf3df),
	.w7(32'hbcfc0c16),
	.w8(32'hbc5ba223),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb43abf),
	.w1(32'h3c9873e5),
	.w2(32'hbca4bffd),
	.w3(32'hb9b4daf7),
	.w4(32'h3b2968c6),
	.w5(32'hbcc1d4b4),
	.w6(32'hbc0d1619),
	.w7(32'hbc54bafd),
	.w8(32'h3bc5f618),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cbeb3),
	.w1(32'h3c38c90c),
	.w2(32'hbaf479f5),
	.w3(32'h3b3f12f8),
	.w4(32'h3bf57a15),
	.w5(32'h3a6b99b1),
	.w6(32'h3c2d8846),
	.w7(32'h3bef4877),
	.w8(32'hb9dc0928),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64fa02),
	.w1(32'hba13938e),
	.w2(32'hbc480ba0),
	.w3(32'h3ae90f83),
	.w4(32'hb902d6a2),
	.w5(32'hbcfc3f06),
	.w6(32'hbb8fbf84),
	.w7(32'hbbff11ce),
	.w8(32'h3c8ba752),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885ecf),
	.w1(32'hbb84ddac),
	.w2(32'h39bdffac),
	.w3(32'h3c69789f),
	.w4(32'h3a4931aa),
	.w5(32'h3b72c068),
	.w6(32'hba4db3e1),
	.w7(32'h3b2566f9),
	.w8(32'h3aac5154),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d014346),
	.w1(32'hbbfeff88),
	.w2(32'h3c1214f7),
	.w3(32'hba9fec23),
	.w4(32'h3bc52147),
	.w5(32'h3d0a8b52),
	.w6(32'hbc4f44af),
	.w7(32'h3b3f8d3f),
	.w8(32'h3b85c368),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cbe5d),
	.w1(32'hbc1cd092),
	.w2(32'hbc3e8b4d),
	.w3(32'h3c122bb8),
	.w4(32'hbbff6e94),
	.w5(32'h3adfffe2),
	.w6(32'hbcb14ffc),
	.w7(32'hbb65db9a),
	.w8(32'hbb41148f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a739c),
	.w1(32'hbba439be),
	.w2(32'hbb4a0095),
	.w3(32'h3b8f709f),
	.w4(32'hbaa4c581),
	.w5(32'hbadb0e4c),
	.w6(32'hba2f2e7c),
	.w7(32'h3b936944),
	.w8(32'h3b3f5a0b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908ad3),
	.w1(32'hba84d6b5),
	.w2(32'hbc7b49d0),
	.w3(32'h39635ef1),
	.w4(32'h3adf1d77),
	.w5(32'hbb0e2eef),
	.w6(32'h3c0c0016),
	.w7(32'hbb14945b),
	.w8(32'h399ec751),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2fa39b),
	.w1(32'hbc39932e),
	.w2(32'hbd25fcd2),
	.w3(32'h3d8c4a67),
	.w4(32'hbbc24319),
	.w5(32'hbdbd670f),
	.w6(32'hbcdefa71),
	.w7(32'h3c55535c),
	.w8(32'h3c4367ac),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6b71a),
	.w1(32'h39d648fc),
	.w2(32'h3cd65f11),
	.w3(32'h3b7269eb),
	.w4(32'hbc53e543),
	.w5(32'hbc29ab06),
	.w6(32'hbcd34a65),
	.w7(32'hbc651a9a),
	.w8(32'h3b8e7773),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b44c),
	.w1(32'hbcef52c5),
	.w2(32'h3c46491e),
	.w3(32'hbc8fca6b),
	.w4(32'hbb41c424),
	.w5(32'h3b66df33),
	.w6(32'hbc8b9995),
	.w7(32'hbaf9d9d7),
	.w8(32'h3bd342d2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca82408),
	.w1(32'hbbd1e9c0),
	.w2(32'h3b907c6e),
	.w3(32'hbc277fa2),
	.w4(32'h3b3c5b81),
	.w5(32'h3c1297ee),
	.w6(32'h3bbd1f03),
	.w7(32'hbcdaa3da),
	.w8(32'hbc3668d7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43730c),
	.w1(32'h3a5ab9bc),
	.w2(32'hbc2fda4a),
	.w3(32'h3cf25814),
	.w4(32'h3bfb1fbc),
	.w5(32'h3c4f4de5),
	.w6(32'h3cb196ea),
	.w7(32'h3c7940b6),
	.w8(32'h3bd1d96a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7abba),
	.w1(32'h3c7e7aa2),
	.w2(32'h3d589f41),
	.w3(32'h3ccdb0d7),
	.w4(32'h3ba3f7e3),
	.w5(32'hbbe81302),
	.w6(32'h3b8ecadf),
	.w7(32'hbc6e6d13),
	.w8(32'hbba00b2e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801d6e),
	.w1(32'h3c3680ba),
	.w2(32'hbd7b1d83),
	.w3(32'hbbb5771e),
	.w4(32'h3b554a26),
	.w5(32'h3c9c63af),
	.w6(32'hb9cd0b64),
	.w7(32'h3bc8f18f),
	.w8(32'h3ca94852),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc337434),
	.w1(32'h3919014a),
	.w2(32'hba289d4f),
	.w3(32'h3cbd3910),
	.w4(32'h3bc5901f),
	.w5(32'h3bf07b0f),
	.w6(32'h3afb71d3),
	.w7(32'h3c1a3467),
	.w8(32'h3b9e392c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494d76),
	.w1(32'h3b46b785),
	.w2(32'h3b641128),
	.w3(32'h3bac8ed1),
	.w4(32'h3c298c26),
	.w5(32'hbc6563c0),
	.w6(32'h3b8102f4),
	.w7(32'hbc84f39a),
	.w8(32'hbb787af0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d208327),
	.w1(32'hbbc3e912),
	.w2(32'h3ad812a6),
	.w3(32'hbcbaa68f),
	.w4(32'h3be34df9),
	.w5(32'h3cd05bb2),
	.w6(32'h3a1aa4e9),
	.w7(32'h3bd3afb4),
	.w8(32'h3b69e3a5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ba28),
	.w1(32'h3bc41fb2),
	.w2(32'hbbff38e9),
	.w3(32'h3ac2b3da),
	.w4(32'h3c021b6f),
	.w5(32'h3ab28555),
	.w6(32'hb9c9b0ab),
	.w7(32'hbb149abf),
	.w8(32'hbc23570d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80d4b8),
	.w1(32'hbba7b099),
	.w2(32'hbbccf9ba),
	.w3(32'hbc27c629),
	.w4(32'hbb94913d),
	.w5(32'hbbfc1ad9),
	.w6(32'hbbce4b8f),
	.w7(32'hbc18177b),
	.w8(32'hbc0deeec),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a18957),
	.w1(32'hbcf727a7),
	.w2(32'h3b9cd6b7),
	.w3(32'h3c9a0e39),
	.w4(32'hbc683291),
	.w5(32'hbc6b56e0),
	.w6(32'hbc10604f),
	.w7(32'h3b668c1c),
	.w8(32'hb91440ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdff87e),
	.w1(32'h3cb7438a),
	.w2(32'h3b0f8cbc),
	.w3(32'h3ac41988),
	.w4(32'h3c145a59),
	.w5(32'hbcb33f97),
	.w6(32'hbb49007b),
	.w7(32'hbc4f9d72),
	.w8(32'h3cc0594c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9547ad),
	.w1(32'hb7f3e5b5),
	.w2(32'h3c0313cb),
	.w3(32'hbcac7547),
	.w4(32'h3c1d829c),
	.w5(32'h3c881246),
	.w6(32'hbc12df0a),
	.w7(32'h3c1ad9bf),
	.w8(32'h3c9453dd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35f080),
	.w1(32'hbc9630b0),
	.w2(32'h3d3fd1ae),
	.w3(32'h3c922803),
	.w4(32'hbcb7c802),
	.w5(32'hbc0045fd),
	.w6(32'hbcaa4e9c),
	.w7(32'hbc9c0f75),
	.w8(32'hbcc264d1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c702749),
	.w1(32'hbb786a03),
	.w2(32'hbc85eba7),
	.w3(32'hbcf2c748),
	.w4(32'h3a99b056),
	.w5(32'hbcac87aa),
	.w6(32'hbbae6a75),
	.w7(32'hbcf87b5a),
	.w8(32'h3ae310d3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccba86c),
	.w1(32'hbc8d0dd7),
	.w2(32'h3c24e0a5),
	.w3(32'h3bb14b96),
	.w4(32'hbbf3b8a1),
	.w5(32'h3c9e2489),
	.w6(32'h3ac8a575),
	.w7(32'h3cae16ca),
	.w8(32'h3b3eef9b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1b290),
	.w1(32'hbc0d8530),
	.w2(32'hbc4a5daf),
	.w3(32'h3ccb025f),
	.w4(32'hbbc37db4),
	.w5(32'hbc52439d),
	.w6(32'hbc904d89),
	.w7(32'hbb004630),
	.w8(32'hbbbbbf2d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8dc47),
	.w1(32'h3c828d2a),
	.w2(32'h3d137f41),
	.w3(32'h3c90dbc3),
	.w4(32'hbcbda423),
	.w5(32'hbbeac6e6),
	.w6(32'hba318368),
	.w7(32'hbb109b31),
	.w8(32'hbb61bb24),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c5a5b),
	.w1(32'hbaf79684),
	.w2(32'hbd2c3e5b),
	.w3(32'hbc2f5439),
	.w4(32'hbca798dc),
	.w5(32'hbc9a2eec),
	.w6(32'h3d2088e4),
	.w7(32'h3cc281c7),
	.w8(32'h3d48791d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule