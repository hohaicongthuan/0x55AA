module layer_10_featuremap_247(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b8f2a),
	.w1(32'hbaa043de),
	.w2(32'hba82bfe6),
	.w3(32'hba7062ba),
	.w4(32'hb9e1d5d5),
	.w5(32'h3a27f868),
	.w6(32'h3a56d725),
	.w7(32'hba4e8a0e),
	.w8(32'h39c1610f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9849310),
	.w1(32'hba0d484d),
	.w2(32'h3a53047b),
	.w3(32'h3a859586),
	.w4(32'h38216820),
	.w5(32'hba37a385),
	.w6(32'h3ad41ea9),
	.w7(32'hb8a53b78),
	.w8(32'h3903841a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba062b7d),
	.w1(32'hba0d9e28),
	.w2(32'h3ab14162),
	.w3(32'h3a80f7d2),
	.w4(32'h3acd3ccd),
	.w5(32'h3a1c7191),
	.w6(32'h3aa79c64),
	.w7(32'h3a6da489),
	.w8(32'h3a295720),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed17cc),
	.w1(32'h3942620c),
	.w2(32'h3a17c24d),
	.w3(32'h390b6d2c),
	.w4(32'h386f3007),
	.w5(32'hb9d9e95e),
	.w6(32'hb97331cf),
	.w7(32'h39664708),
	.w8(32'h389119ec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecbc50),
	.w1(32'hba7febc3),
	.w2(32'h399932d6),
	.w3(32'hbb5e67a5),
	.w4(32'hbb23ea99),
	.w5(32'h3a44dda3),
	.w6(32'hbb3c85ac),
	.w7(32'hbb3967e4),
	.w8(32'h3a8a80a8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2a16b),
	.w1(32'h3a9b62e3),
	.w2(32'h3ac01f11),
	.w3(32'h39b77a50),
	.w4(32'h39bd0795),
	.w5(32'h3a2db8b9),
	.w6(32'hb85ed95c),
	.w7(32'h3a2ad983),
	.w8(32'h38801425),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4c96f),
	.w1(32'h3a6c4de4),
	.w2(32'h3aa47a83),
	.w3(32'h391935c6),
	.w4(32'h39662407),
	.w5(32'hbac6ab72),
	.w6(32'hb9d5cb9b),
	.w7(32'h3a81d50a),
	.w8(32'hba5a5af6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8318f40),
	.w1(32'h3a33fb56),
	.w2(32'h3705c3a8),
	.w3(32'hba550ddc),
	.w4(32'h39fbe637),
	.w5(32'h3616a9b1),
	.w6(32'hbabe5b10),
	.w7(32'h3a318a77),
	.w8(32'hb907ce28),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882c51),
	.w1(32'hba7fd280),
	.w2(32'hb8ca3910),
	.w3(32'hbb34dfd9),
	.w4(32'hbab240bf),
	.w5(32'h3a8d862e),
	.w6(32'hbb1f1b19),
	.w7(32'hba31b36a),
	.w8(32'h3ad2ca4a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca1f8e),
	.w1(32'hbabf5c25),
	.w2(32'h3b0e4c06),
	.w3(32'hbb186fec),
	.w4(32'hbb0dd994),
	.w5(32'h3b1c685e),
	.w6(32'hbafb12e2),
	.w7(32'hba3d6b14),
	.w8(32'h3af30a0e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaae5fd),
	.w1(32'h3a7ebe88),
	.w2(32'h3ace003a),
	.w3(32'h394e544c),
	.w4(32'h398c3591),
	.w5(32'h3ab8a374),
	.w6(32'hb9d6da29),
	.w7(32'h3a4f71ce),
	.w8(32'h39c77d60),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3d604),
	.w1(32'h3b3a4e10),
	.w2(32'h3bd52b4d),
	.w3(32'h3ae84dd9),
	.w4(32'h3b39ad30),
	.w5(32'h3b79d6b0),
	.w6(32'h3a926cb5),
	.w7(32'h3b5a22aa),
	.w8(32'h3b1ffa3f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a7573),
	.w1(32'hbb367bf0),
	.w2(32'h3b370898),
	.w3(32'hbb871466),
	.w4(32'hba9c9332),
	.w5(32'h3b50f736),
	.w6(32'hbb7d41a2),
	.w7(32'hba5bb1b1),
	.w8(32'h3b5621dc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa53fed),
	.w1(32'hbb26b7c8),
	.w2(32'hbb5bc8ab),
	.w3(32'hbb1878cf),
	.w4(32'hbb70f999),
	.w5(32'hbadf9193),
	.w6(32'hb9867a3f),
	.w7(32'hbb6fdac7),
	.w8(32'hb9dc8b3a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a3f3),
	.w1(32'h3a90aef3),
	.w2(32'h3b31aa78),
	.w3(32'hb87dfe58),
	.w4(32'h3a2b244a),
	.w5(32'h3968ddbe),
	.w6(32'h39e38e6f),
	.w7(32'h3ac5e395),
	.w8(32'h3a351ded),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac22524),
	.w1(32'hbb3bab45),
	.w2(32'h3a01b5fa),
	.w3(32'hbb03f40c),
	.w4(32'hbb2bfc53),
	.w5(32'hba1100a4),
	.w6(32'hb97478c0),
	.w7(32'h3a12cdb8),
	.w8(32'hba46602b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3778d5e1),
	.w1(32'hb96e3312),
	.w2(32'h398e5dc4),
	.w3(32'hba692dd5),
	.w4(32'hb8bf85ec),
	.w5(32'h39e75372),
	.w6(32'hb9a173a5),
	.w7(32'h3a0f543b),
	.w8(32'h3a0df23f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11ee5),
	.w1(32'hbae2d3a2),
	.w2(32'h3ab75c2d),
	.w3(32'hbb1f06c9),
	.w4(32'hb9867b0e),
	.w5(32'h3b28edf3),
	.w6(32'h39665e1c),
	.w7(32'h3b293bf6),
	.w8(32'h3927a36f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1678),
	.w1(32'hbafc3838),
	.w2(32'h3a2673ad),
	.w3(32'hbb6ec381),
	.w4(32'hbadc7776),
	.w5(32'h39945cd0),
	.w6(32'hbb184f2f),
	.w7(32'h3a8c5e24),
	.w8(32'h3a155469),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7ca62),
	.w1(32'h39943591),
	.w2(32'h3aa0d2b3),
	.w3(32'hb8ff68d3),
	.w4(32'hba9a8e58),
	.w5(32'hbaca32ff),
	.w6(32'h3a411a64),
	.w7(32'h3a565d90),
	.w8(32'hb98304d8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e03a13),
	.w1(32'h37eea570),
	.w2(32'h3a83b577),
	.w3(32'h394c659d),
	.w4(32'hb91a17b8),
	.w5(32'hba5113bd),
	.w6(32'h3a2a8799),
	.w7(32'h3a9dce84),
	.w8(32'hb997555e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4458b),
	.w1(32'hba04028a),
	.w2(32'h37546f0a),
	.w3(32'hba917e8b),
	.w4(32'hbad4e809),
	.w5(32'h3b0864a8),
	.w6(32'hbac7bc63),
	.w7(32'hba9c48fe),
	.w8(32'h3a8de97e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d1bde),
	.w1(32'h3ac040bc),
	.w2(32'h3ba8f2d4),
	.w3(32'hba11d850),
	.w4(32'h3aad04ee),
	.w5(32'h3b9f9a5f),
	.w6(32'h3acf06d6),
	.w7(32'h3b3c58db),
	.w8(32'h3bccf36e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab74b1e),
	.w1(32'hbb82a120),
	.w2(32'h3a17d703),
	.w3(32'hbacb190f),
	.w4(32'hbb378c4d),
	.w5(32'h3a89ef2c),
	.w6(32'hbb047d9f),
	.w7(32'hbb099b2b),
	.w8(32'h3b099119),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeff382),
	.w1(32'hbab28493),
	.w2(32'h3af95f2f),
	.w3(32'h39dbda0e),
	.w4(32'h3ab34875),
	.w5(32'h3a99f077),
	.w6(32'h3ad49efb),
	.w7(32'hb900e3f1),
	.w8(32'h3ab5f9f5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928e8bb),
	.w1(32'h3ac8e027),
	.w2(32'h3aae7085),
	.w3(32'h3a862c38),
	.w4(32'h39b43dc9),
	.w5(32'h3987d801),
	.w6(32'h3ab86233),
	.w7(32'h3ae9f548),
	.w8(32'h39d32ca8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba166faf),
	.w1(32'hba19be32),
	.w2(32'hba18b057),
	.w3(32'h39be94a4),
	.w4(32'hb7055ea8),
	.w5(32'hbac8e855),
	.w6(32'hb9cf9d57),
	.w7(32'hb7f5fdd7),
	.w8(32'hb9dfd6cf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba153c4c),
	.w1(32'hb96f6a0b),
	.w2(32'h3a134882),
	.w3(32'hba518a76),
	.w4(32'h39d18662),
	.w5(32'h3ad150a8),
	.w6(32'hba26d260),
	.w7(32'hb9e544d4),
	.w8(32'h3a9ad9e3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6b7ee),
	.w1(32'h3aff882b),
	.w2(32'h3b46dba2),
	.w3(32'hb9085ff5),
	.w4(32'h3a2378bd),
	.w5(32'h3b899ec6),
	.w6(32'hb8fe2e1d),
	.w7(32'hb9ccd940),
	.w8(32'h3b47db55),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc7ad),
	.w1(32'hbb78904a),
	.w2(32'h3a318539),
	.w3(32'hba72abf6),
	.w4(32'hba94afe3),
	.w5(32'h3afe8955),
	.w6(32'hbab89779),
	.w7(32'hb9e5e37b),
	.w8(32'h3adffd97),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf4fee),
	.w1(32'h3a2ba04c),
	.w2(32'hb9967954),
	.w3(32'h3b1717dc),
	.w4(32'h39fc7324),
	.w5(32'hbab31c66),
	.w6(32'h3a6dc8eb),
	.w7(32'hb9665cdf),
	.w8(32'hba76c9e3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80d1998),
	.w1(32'h39a1e547),
	.w2(32'hba7b833b),
	.w3(32'hbb033154),
	.w4(32'hbabc5205),
	.w5(32'h3b4c4246),
	.w6(32'h3982d8ed),
	.w7(32'hba112035),
	.w8(32'h3a90eda3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba936372),
	.w1(32'hba92cc49),
	.w2(32'h3b07a603),
	.w3(32'h3ac2477a),
	.w4(32'h3a137ecb),
	.w5(32'h3a06be7a),
	.w6(32'h3a8db584),
	.w7(32'h3985738f),
	.w8(32'hba66859d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11c712),
	.w1(32'h3acb1770),
	.w2(32'h3b35d899),
	.w3(32'h3a133ec3),
	.w4(32'h3af7c9b7),
	.w5(32'hb934dd8f),
	.w6(32'h3a20f7ae),
	.w7(32'h3a967054),
	.w8(32'hba0df498),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6766f),
	.w1(32'hbab25cfa),
	.w2(32'hb96c5ae3),
	.w3(32'hba1987c1),
	.w4(32'hba5d7b26),
	.w5(32'h3abc2d2f),
	.w6(32'h39e56448),
	.w7(32'h3a2db5d8),
	.w8(32'h3ad18a5e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115c68),
	.w1(32'hb9199771),
	.w2(32'h39a1717a),
	.w3(32'h3b020da7),
	.w4(32'h3b00c740),
	.w5(32'h3aa88eb0),
	.w6(32'h3abd9ce8),
	.w7(32'hba2e1819),
	.w8(32'h3a23b445),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f10d1b),
	.w1(32'hba39cbfc),
	.w2(32'h3922358e),
	.w3(32'h38c68c7e),
	.w4(32'hb8bb7bad),
	.w5(32'hb95336d2),
	.w6(32'hb98f42e9),
	.w7(32'hba1f4e8c),
	.w8(32'h3a8577ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35f23),
	.w1(32'h3b92b999),
	.w2(32'h3bda3b24),
	.w3(32'h3b2b0558),
	.w4(32'h3a8a17ea),
	.w5(32'h3bc2a93e),
	.w6(32'h3a883018),
	.w7(32'hb9fa77fb),
	.w8(32'h3b7a8064),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31819b),
	.w1(32'h3bbf778f),
	.w2(32'h3c2241e4),
	.w3(32'h3ba71350),
	.w4(32'h3bcea820),
	.w5(32'h3bd2c0c9),
	.w6(32'h3b90f166),
	.w7(32'h3a69cb68),
	.w8(32'h3be7c3bd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4324b),
	.w1(32'hbb26ea6e),
	.w2(32'hbb95d106),
	.w3(32'hbb47cb24),
	.w4(32'hbb990f5a),
	.w5(32'hbabbf5b9),
	.w6(32'hbb436c5a),
	.w7(32'hbb6e2644),
	.w8(32'hbb18d17c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba012fbb),
	.w1(32'h3a6affc2),
	.w2(32'h3a483dcb),
	.w3(32'hbaa5e580),
	.w4(32'h3a86101c),
	.w5(32'hba63c909),
	.w6(32'h3a814dce),
	.w7(32'h3aa3a157),
	.w8(32'hb978c575),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c096a),
	.w1(32'h3a88a279),
	.w2(32'h3a9325e8),
	.w3(32'h389aa4ea),
	.w4(32'h380e9854),
	.w5(32'h3a977473),
	.w6(32'hb9f9165a),
	.w7(32'h3a453432),
	.w8(32'h3aa417b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65cc3b),
	.w1(32'h39847d19),
	.w2(32'h3b0dcd19),
	.w3(32'h39fe1cbd),
	.w4(32'hb9c71e69),
	.w5(32'h3b190e7e),
	.w6(32'h39b8880b),
	.w7(32'h39a0f162),
	.w8(32'h3aff00de),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b5921),
	.w1(32'hbb0a87ef),
	.w2(32'h3aaf7790),
	.w3(32'hbb94750e),
	.w4(32'hbb134788),
	.w5(32'hbb0122c4),
	.w6(32'hbb4d15f1),
	.w7(32'hbab7ee53),
	.w8(32'hba98e42c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907fef),
	.w1(32'hbb69ef77),
	.w2(32'hb9be876d),
	.w3(32'hbb36ee6d),
	.w4(32'hbb89bc0e),
	.w5(32'h3a385f0f),
	.w6(32'hbb99ea95),
	.w7(32'hbb55a4e7),
	.w8(32'h3a1ef1ef),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1ba7),
	.w1(32'hbb74a470),
	.w2(32'h39c5d0f4),
	.w3(32'hbb3127de),
	.w4(32'hbb14d6fc),
	.w5(32'h3ada491c),
	.w6(32'hbb5622b8),
	.w7(32'hbaa4d1b6),
	.w8(32'h39978c11),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995f71),
	.w1(32'hbaccc0cc),
	.w2(32'h3a199be5),
	.w3(32'hb86b2ef6),
	.w4(32'hba5e3f86),
	.w5(32'hb9afa3be),
	.w6(32'hbaf4967b),
	.w7(32'hbad3da1e),
	.w8(32'hbaa4791e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e643b),
	.w1(32'hbb61752a),
	.w2(32'h3a689270),
	.w3(32'hbbbd03a0),
	.w4(32'hbaf8926c),
	.w5(32'h3a094abf),
	.w6(32'hbba55902),
	.w7(32'h3a4f636d),
	.w8(32'hba792718),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74d66),
	.w1(32'hbaf15df5),
	.w2(32'hba19f08b),
	.w3(32'hb9cde543),
	.w4(32'h39ae7ff4),
	.w5(32'hba553d8a),
	.w6(32'hba6c23c0),
	.w7(32'hb981ad7a),
	.w8(32'hba2d029e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba939dd9),
	.w1(32'hb94d984e),
	.w2(32'h3a02f053),
	.w3(32'hba3eec98),
	.w4(32'hbac1f9b0),
	.w5(32'hb9257e3c),
	.w6(32'hba0c790e),
	.w7(32'hb85c3323),
	.w8(32'hb926a248),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab938a7),
	.w1(32'hb955b6e2),
	.w2(32'h3ae8f12f),
	.w3(32'hb9cc3da4),
	.w4(32'h3a599e30),
	.w5(32'h39dc0a94),
	.w6(32'hb9e9f3d0),
	.w7(32'h3adbc25b),
	.w8(32'hba90127c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385886b3),
	.w1(32'hb9da439a),
	.w2(32'h3ada782d),
	.w3(32'hba7d7f6e),
	.w4(32'h3a30a3ac),
	.w5(32'hb9a6d67b),
	.w6(32'hbb02072f),
	.w7(32'hba46670a),
	.w8(32'h39d7363b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67ccaa),
	.w1(32'h39b0c51a),
	.w2(32'h38d45a66),
	.w3(32'hbad90409),
	.w4(32'h381ed59b),
	.w5(32'hb98dfac3),
	.w6(32'h3a3d172c),
	.w7(32'h3a87da93),
	.w8(32'hb9270ea4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33defb),
	.w1(32'hb9d3c844),
	.w2(32'h3a27b88a),
	.w3(32'hba2fb3e0),
	.w4(32'h390de445),
	.w5(32'hb9cbd640),
	.w6(32'h3a06ee44),
	.w7(32'h3b34d2bd),
	.w8(32'hba9245f1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42e14),
	.w1(32'h3abc249e),
	.w2(32'h3b08ffaa),
	.w3(32'h3a98d2e0),
	.w4(32'h3a881f24),
	.w5(32'h39388b06),
	.w6(32'h3aa4fa6a),
	.w7(32'h3b1f80ec),
	.w8(32'h3a2c2182),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd296e),
	.w1(32'h39ff7b88),
	.w2(32'h3a3c4a13),
	.w3(32'h39ca49e8),
	.w4(32'h39c84cba),
	.w5(32'hba2c1264),
	.w6(32'h3aba5695),
	.w7(32'h3ae225a7),
	.w8(32'hb9272f63),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39234f8e),
	.w1(32'hba2ed84c),
	.w2(32'hba8443bf),
	.w3(32'hba88691c),
	.w4(32'hba503f4e),
	.w5(32'hb8a93c36),
	.w6(32'hb887c1c7),
	.w7(32'hba3743e6),
	.w8(32'h3aa61b9a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfd408),
	.w1(32'h3ac2ab76),
	.w2(32'h3a9a8b11),
	.w3(32'h3ac57d74),
	.w4(32'h3a492465),
	.w5(32'hba0745a0),
	.w6(32'h3ae3c894),
	.w7(32'h3ace191b),
	.w8(32'hba269f83),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e4058),
	.w1(32'hb9b48040),
	.w2(32'h3a9a3789),
	.w3(32'hb93c54f1),
	.w4(32'hb986ec67),
	.w5(32'h397a2e53),
	.w6(32'hba19723b),
	.w7(32'h3a0f4192),
	.w8(32'h3a2cea7e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cf6b5),
	.w1(32'hba86278b),
	.w2(32'hbb11877d),
	.w3(32'hbb02a83d),
	.w4(32'hbb29b22e),
	.w5(32'h3a03241d),
	.w6(32'hbb6da3fb),
	.w7(32'hbb593dff),
	.w8(32'hb9cf4f3a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1682f7),
	.w1(32'hbb106f64),
	.w2(32'hb98fb358),
	.w3(32'hbae8532b),
	.w4(32'hbab6fdbd),
	.w5(32'hba1eaede),
	.w6(32'hbaf61e23),
	.w7(32'hbb0dd9d8),
	.w8(32'hba0bd42c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a361b76),
	.w1(32'h3a83cf4b),
	.w2(32'h3a9c9b61),
	.w3(32'hba4d580e),
	.w4(32'h39e609b1),
	.w5(32'hba1b8d55),
	.w6(32'h3825c2d5),
	.w7(32'h3a83ffef),
	.w8(32'hba16b0ad),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3db0a5),
	.w1(32'hba836647),
	.w2(32'hba06dc1f),
	.w3(32'hb94e1511),
	.w4(32'h3a471fca),
	.w5(32'h39013650),
	.w6(32'h3ab542d4),
	.w7(32'h3abceb37),
	.w8(32'hb9b0d47c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c78a0d),
	.w1(32'h3a5d8d7f),
	.w2(32'h39db7213),
	.w3(32'h39d1092a),
	.w4(32'h39de1549),
	.w5(32'hb9b16bfb),
	.w6(32'h3ab4abed),
	.w7(32'h391b78c9),
	.w8(32'h388fa568),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a39d2),
	.w1(32'hb9b7efc6),
	.w2(32'hb9072af9),
	.w3(32'h3954e07b),
	.w4(32'hbac90ead),
	.w5(32'hbaca0669),
	.w6(32'h39d52ada),
	.w7(32'h3a161df0),
	.w8(32'hbae7d5e6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3ee52),
	.w1(32'h3ac19e5d),
	.w2(32'h3ab6ecaa),
	.w3(32'hba4cd2a9),
	.w4(32'h3a7ea86e),
	.w5(32'hba6a07be),
	.w6(32'h3a35fc0f),
	.w7(32'h3a987320),
	.w8(32'hbaa25dd6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e1289),
	.w1(32'hbaf8a640),
	.w2(32'hbafe427b),
	.w3(32'hba928398),
	.w4(32'hbae1ddf4),
	.w5(32'hbb077480),
	.w6(32'hbad00924),
	.w7(32'hba322f22),
	.w8(32'hbb2d6962),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5468f),
	.w1(32'hbaa03a12),
	.w2(32'h3b09b696),
	.w3(32'hbb4115e7),
	.w4(32'hba200f86),
	.w5(32'h3b303ac9),
	.w6(32'hbb1e5e4b),
	.w7(32'hba2e8beb),
	.w8(32'h3b5d829b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab77573),
	.w1(32'hba3ca979),
	.w2(32'h3b784b4f),
	.w3(32'h3b29e97b),
	.w4(32'h39b1c8d7),
	.w5(32'h3aff6d0e),
	.w6(32'hb91d232e),
	.w7(32'hb8eb127d),
	.w8(32'hb88f1088),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875b51),
	.w1(32'hbb3eb93a),
	.w2(32'h3af1651e),
	.w3(32'hbb1395a4),
	.w4(32'hba49fe13),
	.w5(32'h3b708e82),
	.w6(32'hbb756140),
	.w7(32'hbaddceb4),
	.w8(32'h3b4c755e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ef39),
	.w1(32'h3a814ce9),
	.w2(32'h3946fd09),
	.w3(32'h39ebb060),
	.w4(32'h39851eee),
	.w5(32'hb936815a),
	.w6(32'h3aa8bdf9),
	.w7(32'h3a2a4f5e),
	.w8(32'h3b023fb0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b614640),
	.w1(32'hba28f234),
	.w2(32'hbb148179),
	.w3(32'h3b1dfe77),
	.w4(32'h3a8613b6),
	.w5(32'hb8f67ed8),
	.w6(32'h3b13b81b),
	.w7(32'hbb2146b5),
	.w8(32'hb9f3cc59),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9475ee2),
	.w1(32'hba84dfbf),
	.w2(32'hbb02fdcc),
	.w3(32'h3afdf209),
	.w4(32'h3b8207fa),
	.w5(32'h3a07ab0b),
	.w6(32'h3a63f925),
	.w7(32'hba0fed46),
	.w8(32'h39a410d6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38182b1f),
	.w1(32'h3a2a7573),
	.w2(32'h3a87c99b),
	.w3(32'h38f11abc),
	.w4(32'h3aab7093),
	.w5(32'h3a07d822),
	.w6(32'h39e222f5),
	.w7(32'h39a7cef7),
	.w8(32'hb8e447d9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f78502),
	.w1(32'h3a8cda0c),
	.w2(32'h39f0bca3),
	.w3(32'hba8e0536),
	.w4(32'hba6e9872),
	.w5(32'h39c65110),
	.w6(32'h3984ec8e),
	.w7(32'h3a8dd4b0),
	.w8(32'h3a1f05db),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab514ea),
	.w1(32'h39a2ec6e),
	.w2(32'h3a1eebe1),
	.w3(32'h3a42a67f),
	.w4(32'h3b412ace),
	.w5(32'h3a66c873),
	.w6(32'h3aac49e0),
	.w7(32'h3b0d3209),
	.w8(32'hbaa77d08),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d85f),
	.w1(32'hbabf60ce),
	.w2(32'hba519687),
	.w3(32'hbb1794e5),
	.w4(32'hba81c78e),
	.w5(32'h3a98258b),
	.w6(32'hb9d026ae),
	.w7(32'hba842400),
	.w8(32'h39e897eb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883c9d3),
	.w1(32'hb865f976),
	.w2(32'h3b524fc6),
	.w3(32'hbab8dcf8),
	.w4(32'h3a2ba65a),
	.w5(32'h3ad3520c),
	.w6(32'hbb83f189),
	.w7(32'hb946be1f),
	.w8(32'h3ac0c242),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b70fb9),
	.w1(32'hb9dc7c15),
	.w2(32'hba91f2a6),
	.w3(32'hbb1a5ce8),
	.w4(32'hba10f6ee),
	.w5(32'hba938e93),
	.w6(32'hbacf4490),
	.w7(32'hb95ef549),
	.w8(32'hba9ff48f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a30ee),
	.w1(32'hba962f4d),
	.w2(32'h393b47c5),
	.w3(32'hbad277ed),
	.w4(32'hba98ff0c),
	.w5(32'h39d6883f),
	.w6(32'hbacf5892),
	.w7(32'hba9ea579),
	.w8(32'h3a739afe),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a322720),
	.w1(32'h3aa26b0b),
	.w2(32'h39bfcca9),
	.w3(32'h3ac71a23),
	.w4(32'h3abfd6c3),
	.w5(32'h3aef2d66),
	.w6(32'h3a84998c),
	.w7(32'h38f67507),
	.w8(32'h3a99371b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d9776),
	.w1(32'hba42f86b),
	.w2(32'h3a59d92f),
	.w3(32'hb9bbbe41),
	.w4(32'h3a61254f),
	.w5(32'h39a44965),
	.w6(32'hb990bc1f),
	.w7(32'h3a13fa35),
	.w8(32'h3aba1bd0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5d5ee),
	.w1(32'hb9f66140),
	.w2(32'h3a12238b),
	.w3(32'h3b01d2fe),
	.w4(32'h3a78a00c),
	.w5(32'h3a9fbc6a),
	.w6(32'h3af285fa),
	.w7(32'hba06cc1f),
	.w8(32'h3a398329),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac259a0),
	.w1(32'h3900f5c2),
	.w2(32'h395eeade),
	.w3(32'hb9e8273c),
	.w4(32'hba96b474),
	.w5(32'hb8f13845),
	.w6(32'hbab43d15),
	.w7(32'h3a80044e),
	.w8(32'h381b61df),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6c410),
	.w1(32'h3a9836a1),
	.w2(32'h3a1efa74),
	.w3(32'hb8341e93),
	.w4(32'hb6c5bf97),
	.w5(32'hba2d7eb0),
	.w6(32'h3ae775ab),
	.w7(32'h39ac0f07),
	.w8(32'h3912bbb4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8efc2c0),
	.w1(32'h3a4d46b5),
	.w2(32'h3a851237),
	.w3(32'hb91d2d0e),
	.w4(32'h3a18d66b),
	.w5(32'h38120290),
	.w6(32'hb9e67fd1),
	.w7(32'h3986a7d5),
	.w8(32'h3a94441f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c69b50),
	.w1(32'h3b0c5a6d),
	.w2(32'h3b36855a),
	.w3(32'h3b8093fa),
	.w4(32'h3ab72db2),
	.w5(32'h3a9800dc),
	.w6(32'h3b569f51),
	.w7(32'h3a34ef6c),
	.w8(32'hb9db75a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa489c1),
	.w1(32'h3a922577),
	.w2(32'h3b286d43),
	.w3(32'h3a30f289),
	.w4(32'hb9e060f0),
	.w5(32'h3a5a7991),
	.w6(32'h3aa6a0e3),
	.w7(32'h3a20de8a),
	.w8(32'h392fd737),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60b014),
	.w1(32'hbaad9d5b),
	.w2(32'hb89dd15d),
	.w3(32'hbb020258),
	.w4(32'hbb3b6da3),
	.w5(32'hbb25f2b8),
	.w6(32'hbb070034),
	.w7(32'hba009111),
	.w8(32'hbb4c4330),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332d68),
	.w1(32'hbb82c28b),
	.w2(32'h397c2244),
	.w3(32'hbab39f41),
	.w4(32'h3a1c4a3b),
	.w5(32'h3b009eac),
	.w6(32'hba0b543e),
	.w7(32'h3a9fd05a),
	.w8(32'h39916c0c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f01bc),
	.w1(32'h3a6175bd),
	.w2(32'h3b2d88ee),
	.w3(32'h371ff718),
	.w4(32'h3901c991),
	.w5(32'h3b18587d),
	.w6(32'hb9d7d9ed),
	.w7(32'hb9ab9581),
	.w8(32'h399fa5e4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91baf94),
	.w1(32'hbb2006ac),
	.w2(32'h3a88a167),
	.w3(32'hb9f55f3d),
	.w4(32'hbadf5120),
	.w5(32'h3aac2754),
	.w6(32'hba15eaaf),
	.w7(32'hb9d3602a),
	.w8(32'h39c85e44),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c910b),
	.w1(32'hba615b07),
	.w2(32'h3a82f800),
	.w3(32'hb9e45bca),
	.w4(32'hbaf0d00f),
	.w5(32'hb984c02a),
	.w6(32'hb9b09a12),
	.w7(32'hba7db0da),
	.w8(32'hb8eb8df4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3814f95e),
	.w1(32'hb9b122b1),
	.w2(32'hb9d2aaa4),
	.w3(32'h3aa937fa),
	.w4(32'hba5e7fc5),
	.w5(32'hbb7900ee),
	.w6(32'h3a368583),
	.w7(32'hbad268e8),
	.w8(32'hbb18b71e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f6da),
	.w1(32'h3a0ff210),
	.w2(32'hba8f594c),
	.w3(32'h3a7fc748),
	.w4(32'hbae6e69e),
	.w5(32'hbad133ba),
	.w6(32'h3b070f7d),
	.w7(32'hba5a968a),
	.w8(32'hbb1ad440),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef8bed),
	.w1(32'h3a6944bb),
	.w2(32'h3a8c1218),
	.w3(32'hb896468d),
	.w4(32'hbaab77b8),
	.w5(32'hba65db0c),
	.w6(32'h3a452d92),
	.w7(32'h3af929ef),
	.w8(32'h378b2e77),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e701e),
	.w1(32'h398c93ee),
	.w2(32'hba8ec2f0),
	.w3(32'hbac4a9b8),
	.w4(32'hba19caa3),
	.w5(32'h3a994eaa),
	.w6(32'hbacb2f50),
	.w7(32'hba5aaf6e),
	.w8(32'hb8bc0ef5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161d38),
	.w1(32'hbb217262),
	.w2(32'h39bc83a1),
	.w3(32'hbb1f5c9b),
	.w4(32'hbadd0a1c),
	.w5(32'hba9f37a3),
	.w6(32'hb9ed01a4),
	.w7(32'h39b12473),
	.w8(32'hbaab4d49),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f7d0),
	.w1(32'hba8487f6),
	.w2(32'h3b167dae),
	.w3(32'hba1fa74a),
	.w4(32'h39158570),
	.w5(32'hbb6dd088),
	.w6(32'hba17dcf6),
	.w7(32'h3a5c0ac3),
	.w8(32'hbb83df09),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb481f2),
	.w1(32'hbba1260c),
	.w2(32'hbb1c7fda),
	.w3(32'hbbb833e7),
	.w4(32'hbb1408d9),
	.w5(32'h3b144f3f),
	.w6(32'hbb496951),
	.w7(32'hba957e69),
	.w8(32'h3b27bd86),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd6cda),
	.w1(32'h3badbe53),
	.w2(32'h3bd243cc),
	.w3(32'h3b273a5e),
	.w4(32'h3b113f78),
	.w5(32'h3b7f5422),
	.w6(32'h3a35ae4d),
	.w7(32'h39a5d8b6),
	.w8(32'h3b77391b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd391c),
	.w1(32'hba44382f),
	.w2(32'h3ad68433),
	.w3(32'hbb48da7c),
	.w4(32'hbb4732e5),
	.w5(32'hba304c7c),
	.w6(32'hba9f70c5),
	.w7(32'h3a4ab615),
	.w8(32'hb9c947a4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f984a),
	.w1(32'h39ada88a),
	.w2(32'h3a6de275),
	.w3(32'hb9c9f4f0),
	.w4(32'hbaf415c9),
	.w5(32'h39956045),
	.w6(32'hb9f1805a),
	.w7(32'hba1b9750),
	.w8(32'hbab1a645),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0939e),
	.w1(32'h38b85a99),
	.w2(32'hba134cb1),
	.w3(32'h38ed6a8f),
	.w4(32'hb9c0b932),
	.w5(32'h3a02b66b),
	.w6(32'hba1ec380),
	.w7(32'hba8f9f95),
	.w8(32'h3a8fcd4b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88ac3d),
	.w1(32'h3ad3632c),
	.w2(32'h3ab5ef19),
	.w3(32'h375a81f5),
	.w4(32'h3ab88af5),
	.w5(32'h3b1037ee),
	.w6(32'h3a8cf1b3),
	.w7(32'h3b16ab83),
	.w8(32'h3ab5625b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afdb2d),
	.w1(32'h3a2b6b92),
	.w2(32'h3a96488d),
	.w3(32'h3a6b0d7e),
	.w4(32'h3b30ef39),
	.w5(32'hba3b5bae),
	.w6(32'hba707575),
	.w7(32'h3909d922),
	.w8(32'hbadf2709),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95e685),
	.w1(32'hbbc98ab3),
	.w2(32'hbba729bb),
	.w3(32'hbb49bcb2),
	.w4(32'hbb22897e),
	.w5(32'h3a42b0bf),
	.w6(32'hbb99f43e),
	.w7(32'hbb83ee18),
	.w8(32'h39dae9c6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a276c),
	.w1(32'h3aab62ce),
	.w2(32'h39c703fb),
	.w3(32'h3ab08c20),
	.w4(32'h3a22273e),
	.w5(32'hbb6bb3d7),
	.w6(32'h3a3ecf97),
	.w7(32'h39d9e917),
	.w8(32'hbb30d678),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba672ec),
	.w1(32'hbba69922),
	.w2(32'h3aca5aeb),
	.w3(32'hbbcd1421),
	.w4(32'hba97285c),
	.w5(32'h3a012c3e),
	.w6(32'hbb9dad7f),
	.w7(32'h3a9acb59),
	.w8(32'h3a39d2bc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9898c5),
	.w1(32'hbafc4ba5),
	.w2(32'hb98db6e2),
	.w3(32'hbab29ae9),
	.w4(32'hbac0f607),
	.w5(32'h3a09e155),
	.w6(32'hba42693b),
	.w7(32'hb9f87d5a),
	.w8(32'h3a585aaa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f4695),
	.w1(32'h3a933604),
	.w2(32'h3b28e4a5),
	.w3(32'hb9e085f8),
	.w4(32'h3a494b94),
	.w5(32'h3b07c4b3),
	.w6(32'h3a6c4c28),
	.w7(32'h3b1e25b4),
	.w8(32'h3b0a06e4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a554ad3),
	.w1(32'h3a48236b),
	.w2(32'h3ad3a84a),
	.w3(32'h39de57b6),
	.w4(32'hba00f32f),
	.w5(32'h3ac656a9),
	.w6(32'h39f196eb),
	.w7(32'h389c37ca),
	.w8(32'h3a5c4fe3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7891d0),
	.w1(32'h3a5c56d9),
	.w2(32'h3ac193ed),
	.w3(32'h3a758a65),
	.w4(32'h3a052238),
	.w5(32'h3ae8255c),
	.w6(32'h38c8b11e),
	.w7(32'h37b004f8),
	.w8(32'h3aca2f54),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf91f2),
	.w1(32'hba21370a),
	.w2(32'h39cc7418),
	.w3(32'hbae9c684),
	.w4(32'hbacc3ca8),
	.w5(32'hbaa27dd2),
	.w6(32'hba9509b6),
	.w7(32'hba2271f8),
	.w8(32'hbb351c0f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ceda3),
	.w1(32'hbb771224),
	.w2(32'hba568b56),
	.w3(32'hba72d3ab),
	.w4(32'hb947a3d7),
	.w5(32'h39c91a7b),
	.w6(32'hbb2c153d),
	.w7(32'hb9feb8a8),
	.w8(32'h3a78bf0c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387025de),
	.w1(32'h39152599),
	.w2(32'h399dae84),
	.w3(32'hba586b68),
	.w4(32'hba69c4db),
	.w5(32'h395446fd),
	.w6(32'h372d47ef),
	.w7(32'h396ec1e2),
	.w8(32'h398401c2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1bf10),
	.w1(32'h3818f57e),
	.w2(32'hba0a23b8),
	.w3(32'h38dc20fa),
	.w4(32'hb9577dc9),
	.w5(32'hbb518974),
	.w6(32'h397f892a),
	.w7(32'hba37e86c),
	.w8(32'hbaf9e981),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf59b73),
	.w1(32'hbb0857db),
	.w2(32'hbb34d946),
	.w3(32'hbb957322),
	.w4(32'hbb9260f1),
	.w5(32'hbb1f71e5),
	.w6(32'hbb469995),
	.w7(32'hbb55767f),
	.w8(32'hbab251ec),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc817f),
	.w1(32'hba96e208),
	.w2(32'hba6984cb),
	.w3(32'hba9b0c97),
	.w4(32'hb9fba665),
	.w5(32'hbb89edd5),
	.w6(32'hb9b7d1d4),
	.w7(32'h3910e54a),
	.w8(32'hbba4a0d2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f61bc),
	.w1(32'hbbcf7747),
	.w2(32'hbae7b703),
	.w3(32'hbbedd66a),
	.w4(32'hbb8db13f),
	.w5(32'h3b016c75),
	.w6(32'hbc06e46c),
	.w7(32'hbbb33588),
	.w8(32'h3a4f6156),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941ff9a),
	.w1(32'hbab0bfae),
	.w2(32'hbaa0fed3),
	.w3(32'hb6c4bff5),
	.w4(32'hba43092d),
	.w5(32'h39de2b3c),
	.w6(32'hba42f71d),
	.w7(32'hbb020310),
	.w8(32'h396dc57c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bac14),
	.w1(32'h392da799),
	.w2(32'h3a712109),
	.w3(32'hb89038b1),
	.w4(32'hb92988b2),
	.w5(32'h3aa094c8),
	.w6(32'hba3c5e40),
	.w7(32'h3a4b8ef7),
	.w8(32'h3a155686),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bacae5),
	.w1(32'h39891300),
	.w2(32'h39c7e859),
	.w3(32'hb9841f80),
	.w4(32'hb7b4bddf),
	.w5(32'h3acb694e),
	.w6(32'hba08c34d),
	.w7(32'hb98350dc),
	.w8(32'h3a7cdbc2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a020e69),
	.w1(32'h395b3e90),
	.w2(32'h394096ff),
	.w3(32'h39c4685d),
	.w4(32'h39c4064d),
	.w5(32'h39c3f03b),
	.w6(32'h38972066),
	.w7(32'h3980e11a),
	.w8(32'h3a87013e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c7e1e),
	.w1(32'h39db9122),
	.w2(32'h37082f6d),
	.w3(32'h3863a46a),
	.w4(32'h37a03263),
	.w5(32'hb933c90f),
	.w6(32'hb9995ba6),
	.w7(32'h378fa834),
	.w8(32'h39abfc16),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a654d23),
	.w1(32'h3a88a091),
	.w2(32'h39a5dadc),
	.w3(32'h380ac5fb),
	.w4(32'hb9eee70b),
	.w5(32'h3af6a1fe),
	.w6(32'h390bc5ed),
	.w7(32'hb956df9f),
	.w8(32'h3a8fd4ee),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872112),
	.w1(32'h3acdd0bd),
	.w2(32'h3ad5985e),
	.w3(32'h3b009425),
	.w4(32'h3a3c9969),
	.w5(32'hba8e71a1),
	.w6(32'h3a979f95),
	.w7(32'h3a1d89da),
	.w8(32'hbb0ab24f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07446c),
	.w1(32'hbb5f5131),
	.w2(32'hba8e81b7),
	.w3(32'hbb1da484),
	.w4(32'hba28645d),
	.w5(32'h3b0e6dc3),
	.w6(32'hbb7fee3c),
	.w7(32'hbaec630f),
	.w8(32'h3b050513),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f2c17),
	.w1(32'hba71d494),
	.w2(32'hbb0b2179),
	.w3(32'hbab52f3d),
	.w4(32'hbb3b0899),
	.w5(32'hba96b230),
	.w6(32'h3a1d599f),
	.w7(32'hba86968c),
	.w8(32'hb96de0f0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f709),
	.w1(32'h3ad9ea59),
	.w2(32'h3a83d920),
	.w3(32'h3abb7e5b),
	.w4(32'h3aa3db4f),
	.w5(32'hb9b57720),
	.w6(32'h3ae0a0af),
	.w7(32'h3ae60e82),
	.w8(32'hba71e68d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d9540),
	.w1(32'hbabbfd31),
	.w2(32'hba654e57),
	.w3(32'hba1a35f2),
	.w4(32'hba83f57d),
	.w5(32'h36d63bfc),
	.w6(32'hbafac753),
	.w7(32'hbababc76),
	.w8(32'h3a0712de),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5f035),
	.w1(32'h3ac344ee),
	.w2(32'h3ad7284a),
	.w3(32'h3719e1b2),
	.w4(32'h38eb36c3),
	.w5(32'hbb1bdc6a),
	.w6(32'h3aa62e5e),
	.w7(32'h3a8184f3),
	.w8(32'hbb21accb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39827e),
	.w1(32'hbb73e64e),
	.w2(32'hbb2502b9),
	.w3(32'hbb410407),
	.w4(32'hbb415919),
	.w5(32'hb8a56541),
	.w6(32'hbb39d631),
	.w7(32'hbb56a5cc),
	.w8(32'h39380f79),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b77c),
	.w1(32'hba4c0900),
	.w2(32'hbad2cc16),
	.w3(32'hba17a440),
	.w4(32'hbaaca474),
	.w5(32'hbab20c46),
	.w6(32'hbab5eb04),
	.w7(32'hbadeb9a5),
	.w8(32'hbb13decd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c04d),
	.w1(32'hbb3026e5),
	.w2(32'hbab91ebf),
	.w3(32'hbaf5a806),
	.w4(32'hbade1114),
	.w5(32'h3a3e384f),
	.w6(32'hbb180d04),
	.w7(32'hbaaeb3b1),
	.w8(32'h3a0179f9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e3b31),
	.w1(32'hbad79cae),
	.w2(32'hbacda0f6),
	.w3(32'hba4c0a1a),
	.w4(32'hba2d03e3),
	.w5(32'hb9105bd6),
	.w6(32'hba692eba),
	.w7(32'hbae8d23a),
	.w8(32'hba1595ec),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b58e),
	.w1(32'hb90c60bc),
	.w2(32'hb94a07af),
	.w3(32'hbac0ada2),
	.w4(32'hbb3d3f52),
	.w5(32'h3a811e95),
	.w6(32'h381ba3c0),
	.w7(32'hbb01fc5b),
	.w8(32'h3a367ab4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e80e9a),
	.w1(32'hb93f5aed),
	.w2(32'hb9a029aa),
	.w3(32'h39625abc),
	.w4(32'hba7272fc),
	.w5(32'hba81de56),
	.w6(32'h3a97b96a),
	.w7(32'h380b191d),
	.w8(32'hba661100),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24c30c),
	.w1(32'hba727a1d),
	.w2(32'hbad09dbb),
	.w3(32'hb9e0387f),
	.w4(32'hba86422f),
	.w5(32'h39bdf28e),
	.w6(32'hb8fc3e86),
	.w7(32'hba18e773),
	.w8(32'hba3844df),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ef812),
	.w1(32'hbafa9d53),
	.w2(32'hb965e77e),
	.w3(32'hb884040d),
	.w4(32'hba3fb5d9),
	.w5(32'h3a96915c),
	.w6(32'hbad520a9),
	.w7(32'hbadc8661),
	.w8(32'h39166436),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03c7c6),
	.w1(32'hba942e4d),
	.w2(32'h3a86f4c1),
	.w3(32'h3a360ffb),
	.w4(32'h3ac1b6ec),
	.w5(32'h399d9e00),
	.w6(32'hba4b4519),
	.w7(32'h3762b0b5),
	.w8(32'h3a998cf6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982994f),
	.w1(32'h3a7b4d0f),
	.w2(32'h3b125b25),
	.w3(32'hb9d73062),
	.w4(32'h394d246e),
	.w5(32'h3a7c4639),
	.w6(32'h3a447705),
	.w7(32'h3a8b682c),
	.w8(32'hba268321),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a69a94),
	.w1(32'hba243121),
	.w2(32'hbafabb11),
	.w3(32'h3a800d90),
	.w4(32'hba48940b),
	.w5(32'hba4c6164),
	.w6(32'h3ab02877),
	.w7(32'hba1d80a6),
	.w8(32'h396ede41),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af29668),
	.w1(32'h3b129eea),
	.w2(32'h3acd2fef),
	.w3(32'h3ad96eaa),
	.w4(32'h3a456a84),
	.w5(32'h3a71fd2d),
	.w6(32'h3b0030e8),
	.w7(32'h3ace4087),
	.w8(32'h3acba5ab),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17b49),
	.w1(32'h3af6386a),
	.w2(32'h3a89ccaf),
	.w3(32'h3ab49bb9),
	.w4(32'h3a82d706),
	.w5(32'hba1005ce),
	.w6(32'h3ae6da32),
	.w7(32'h3aad66b4),
	.w8(32'hba86fe94),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae718),
	.w1(32'hba90be5e),
	.w2(32'hba3b2ace),
	.w3(32'hba0e56eb),
	.w4(32'h3906e446),
	.w5(32'hba9e47db),
	.w6(32'hbaa1e1fa),
	.w7(32'hba1c011b),
	.w8(32'hba3d28e3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913671),
	.w1(32'hbac54bb3),
	.w2(32'hbaf26424),
	.w3(32'hbad9ddd2),
	.w4(32'hbb279fda),
	.w5(32'hb9eae622),
	.w6(32'hba0157c5),
	.w7(32'hba80efc2),
	.w8(32'hba8491ff),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28d22),
	.w1(32'h3a0af99f),
	.w2(32'h3b6249fa),
	.w3(32'hbadaa96e),
	.w4(32'h3a7004cb),
	.w5(32'h3b92547c),
	.w6(32'hbabb88d5),
	.w7(32'h3ac72857),
	.w8(32'h3b647d09),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae0b45),
	.w1(32'h3ac95449),
	.w2(32'h3aac6b75),
	.w3(32'h3a50e304),
	.w4(32'h3968d50b),
	.w5(32'h3a7ff2f6),
	.w6(32'h3a4dfd30),
	.w7(32'h3a3d81f8),
	.w8(32'h3a8dc905),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2e8da),
	.w1(32'hb7fba333),
	.w2(32'h3ac9ea8e),
	.w3(32'hba214e93),
	.w4(32'hb9fbcb3e),
	.w5(32'hba4c2607),
	.w6(32'h3a3d6cc5),
	.w7(32'h3a065d4e),
	.w8(32'hba90bced),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace9c47),
	.w1(32'hbae46839),
	.w2(32'hb9243de1),
	.w3(32'hbade019b),
	.w4(32'hbb01f272),
	.w5(32'h3a3fd93b),
	.w6(32'hbac73caa),
	.w7(32'hb955f3bb),
	.w8(32'h3a9e1d3d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbbf70),
	.w1(32'hb87c1613),
	.w2(32'h3a316544),
	.w3(32'hba364219),
	.w4(32'hb9b1cc3e),
	.w5(32'h3a78f4ae),
	.w6(32'hbb02cbc8),
	.w7(32'hba824ada),
	.w8(32'h3a0244d7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de8126),
	.w1(32'h3a56b8b2),
	.w2(32'h3aec188f),
	.w3(32'hb9a2e2aa),
	.w4(32'hba1f065a),
	.w5(32'h3ad8b4b6),
	.w6(32'h3941b0eb),
	.w7(32'h39d34b6a),
	.w8(32'h3a52efcf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2db6a9),
	.w1(32'h3a65b401),
	.w2(32'hba1e4013),
	.w3(32'h3ad15247),
	.w4(32'h3a72891e),
	.w5(32'hbb0c1058),
	.w6(32'h3a57a21b),
	.w7(32'h397fb41a),
	.w8(32'hba29fab6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b26995),
	.w1(32'hba1bbb83),
	.w2(32'h3ad15846),
	.w3(32'hba88d006),
	.w4(32'h3ac01afa),
	.w5(32'h3a896571),
	.w6(32'hb91004ec),
	.w7(32'h3b097cc8),
	.w8(32'h3a826f00),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d4bed),
	.w1(32'hb9c88df6),
	.w2(32'h38fc5ba5),
	.w3(32'hba6f675c),
	.w4(32'hbad61e29),
	.w5(32'h3abb7778),
	.w6(32'hbab07ad3),
	.w7(32'hbb23d76e),
	.w8(32'h3ac370d6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b467e38),
	.w1(32'h3a7ae2d8),
	.w2(32'hbb26e6c0),
	.w3(32'h3b20324a),
	.w4(32'hbafcf547),
	.w5(32'hba94a340),
	.w6(32'h3b8ee338),
	.w7(32'hbabb369a),
	.w8(32'hbb63283f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dc878),
	.w1(32'h3aeb1d27),
	.w2(32'h3b6445f5),
	.w3(32'h3ab3fa59),
	.w4(32'h3afd03db),
	.w5(32'h3b178f04),
	.w6(32'h3a41b227),
	.w7(32'h3a8bf302),
	.w8(32'h3b020f70),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16b8fe),
	.w1(32'h3a1da84e),
	.w2(32'h3a6f1fdf),
	.w3(32'hb9da92d1),
	.w4(32'hb97bf446),
	.w5(32'h393b9f47),
	.w6(32'hbaca47df),
	.w7(32'h3920b1f7),
	.w8(32'hba889385),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9dfea),
	.w1(32'h375161e8),
	.w2(32'hba22bb2b),
	.w3(32'h3a0f4d27),
	.w4(32'hb855fcc4),
	.w5(32'hba425f70),
	.w6(32'hbadfb675),
	.w7(32'hbad55b4d),
	.w8(32'hbac77e94),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14d46f),
	.w1(32'hbaafb076),
	.w2(32'h3aa1ab87),
	.w3(32'hbb5b8a2d),
	.w4(32'hbb128dc2),
	.w5(32'hba9d92af),
	.w6(32'hbb83cd89),
	.w7(32'hba440cfd),
	.w8(32'hbab1526d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06ddc6),
	.w1(32'hbac512e9),
	.w2(32'hbaa25f6b),
	.w3(32'hbabae9c0),
	.w4(32'hba5093dc),
	.w5(32'hb9b0fa0e),
	.w6(32'hbacd2ef7),
	.w7(32'hba88572f),
	.w8(32'hb8f32a5c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ad887),
	.w1(32'hb94fbaed),
	.w2(32'h3a951343),
	.w3(32'hb9e13b77),
	.w4(32'hba4872ef),
	.w5(32'hbad0eb7e),
	.w6(32'hb89a62ed),
	.w7(32'h393a59d6),
	.w8(32'hbabe553a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb063a87),
	.w1(32'hbac937e8),
	.w2(32'hb9f6a28e),
	.w3(32'hbadf521c),
	.w4(32'hba8f6455),
	.w5(32'hba6eda42),
	.w6(32'hbb19b71f),
	.w7(32'hba02fb0a),
	.w8(32'hbb12bf0c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962aae4),
	.w1(32'h3a1e2165),
	.w2(32'h3b4d8f00),
	.w3(32'hbb0b2e8a),
	.w4(32'hbb0a6b97),
	.w5(32'h3b94d916),
	.w6(32'hbba5d11e),
	.w7(32'hbb838b39),
	.w8(32'h3b9b85a4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc657f),
	.w1(32'hb9f21744),
	.w2(32'h39817f1e),
	.w3(32'hba497445),
	.w4(32'hb8b6ceae),
	.w5(32'hb88aebdd),
	.w6(32'hb8968b13),
	.w7(32'h3a86a2b1),
	.w8(32'h39e70121),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2be1d4),
	.w1(32'hb78cb49a),
	.w2(32'hba24fd43),
	.w3(32'h389dcffb),
	.w4(32'h38628953),
	.w5(32'hb9c59886),
	.w6(32'hba094cfa),
	.w7(32'hb9b284ed),
	.w8(32'h3801a0b1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae784eb),
	.w1(32'h3ab8fee0),
	.w2(32'h3965ac32),
	.w3(32'hb95641cd),
	.w4(32'hbb15a43a),
	.w5(32'hbb233685),
	.w6(32'h3acb0969),
	.w7(32'hb95ffd8d),
	.w8(32'hbb2dccec),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b88b8),
	.w1(32'hbaf1fae7),
	.w2(32'h3a8648c5),
	.w3(32'hbae26ce5),
	.w4(32'hbb0bb357),
	.w5(32'hb947cbf9),
	.w6(32'hba951ab2),
	.w7(32'hba72a02b),
	.w8(32'hbb260a15),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b33970),
	.w1(32'h3909028b),
	.w2(32'h3b0637f3),
	.w3(32'hb995fbae),
	.w4(32'h3a82951e),
	.w5(32'h3ad006c6),
	.w6(32'hbb239d9b),
	.w7(32'hbaa988e7),
	.w8(32'h3a8f4e48),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e57c),
	.w1(32'hbb149858),
	.w2(32'hba227c93),
	.w3(32'hbb28322e),
	.w4(32'hbb30cdd0),
	.w5(32'hba8d5fa9),
	.w6(32'hbb00ac81),
	.w7(32'hbabcf535),
	.w8(32'h3ab4a9e4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba255123),
	.w1(32'hb8ed2eb5),
	.w2(32'hba013047),
	.w3(32'h3966f972),
	.w4(32'h38fa09fc),
	.w5(32'hba5c3693),
	.w6(32'h3ae6b82d),
	.w7(32'h3b0d79ac),
	.w8(32'hbade5112),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb422c77),
	.w1(32'hbb61951e),
	.w2(32'hba04b158),
	.w3(32'hbb9b73c6),
	.w4(32'hbb7968cd),
	.w5(32'h3b470fd6),
	.w6(32'hbb65df00),
	.w7(32'hbb634370),
	.w8(32'h39803a48),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1cb68),
	.w1(32'h39ea151e),
	.w2(32'h3a8e25c1),
	.w3(32'h3a8918d1),
	.w4(32'h3987836c),
	.w5(32'h3a29b878),
	.w6(32'hb9ec89a7),
	.w7(32'hba919157),
	.w8(32'h3a03eb1b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f4718),
	.w1(32'hbb6c98b8),
	.w2(32'hbabfb611),
	.w3(32'hbb39be3c),
	.w4(32'hbb139079),
	.w5(32'h3b446899),
	.w6(32'hbb004137),
	.w7(32'hba91c6d6),
	.w8(32'h3b26ce2f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1788),
	.w1(32'h3b472e85),
	.w2(32'h3b201b91),
	.w3(32'h3b54e973),
	.w4(32'h3b0acd98),
	.w5(32'h3b16068f),
	.w6(32'h3b6809e6),
	.w7(32'h3b14da18),
	.w8(32'h3a9f2e09),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae431e1),
	.w1(32'h39ebd640),
	.w2(32'h392acf36),
	.w3(32'h3acdb975),
	.w4(32'h3a839a02),
	.w5(32'hba723cf7),
	.w6(32'h3a2b364f),
	.w7(32'h394964a4),
	.w8(32'hbafb5f6c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b097),
	.w1(32'h3b224359),
	.w2(32'h3b0fbff7),
	.w3(32'h3b07fcc0),
	.w4(32'h3af8da19),
	.w5(32'hbb298e29),
	.w6(32'h3b01e177),
	.w7(32'h3adcce9e),
	.w8(32'hbb0c397d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61b810),
	.w1(32'hbb85bfab),
	.w2(32'hbac196fe),
	.w3(32'hbb6bf960),
	.w4(32'hbb286b8e),
	.w5(32'hbb056eff),
	.w6(32'hbb5371bd),
	.w7(32'hbaf47235),
	.w8(32'hbabb5b08),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4f11),
	.w1(32'hbb198278),
	.w2(32'hbb1a013f),
	.w3(32'hbb10f397),
	.w4(32'hbad60048),
	.w5(32'h3a3d2e5f),
	.w6(32'hbacc3944),
	.w7(32'hbaae125b),
	.w8(32'h3a8a25dc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95beef),
	.w1(32'hba215169),
	.w2(32'hb9277ff4),
	.w3(32'hb9deadbf),
	.w4(32'h39a91e06),
	.w5(32'h3b303656),
	.w6(32'hbad76011),
	.w7(32'hba8cea89),
	.w8(32'h3ab44df8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac83a73),
	.w1(32'hba0f31e0),
	.w2(32'h3a58325e),
	.w3(32'hba5e1075),
	.w4(32'h38a52d0e),
	.w5(32'h389c77f5),
	.w6(32'hbb0c5b80),
	.w7(32'hb956ab5f),
	.w8(32'h3a0af88a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eddb71),
	.w1(32'h397a90f6),
	.w2(32'h385d49a6),
	.w3(32'h3a39263a),
	.w4(32'h3a145951),
	.w5(32'h38c37824),
	.w6(32'h39a29f0d),
	.w7(32'h3a76736e),
	.w8(32'h39fe474d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19f92d),
	.w1(32'h3a3ab3fd),
	.w2(32'h3a5185e1),
	.w3(32'h39f5f390),
	.w4(32'h39e6ac3e),
	.w5(32'h3b16855e),
	.w6(32'h3a26d39b),
	.w7(32'h39bbc64a),
	.w8(32'h3b007c58),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33ac10),
	.w1(32'h3ad6a794),
	.w2(32'h3b8898c3),
	.w3(32'h3ac68598),
	.w4(32'h3ae1983a),
	.w5(32'h3b23b8b5),
	.w6(32'h3a128a22),
	.w7(32'h3aaf17ce),
	.w8(32'h3b1464fc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37a0e2),
	.w1(32'h398f269b),
	.w2(32'h391bcd2a),
	.w3(32'hb9381d5c),
	.w4(32'hb938592e),
	.w5(32'h3a8722fa),
	.w6(32'hb9d17138),
	.w7(32'h3921d753),
	.w8(32'h3a3d0e34),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8035b0),
	.w1(32'h3a3f9c7d),
	.w2(32'h3a3fbf4e),
	.w3(32'h39ea99fd),
	.w4(32'h3a273a5f),
	.w5(32'h3a0e6e0b),
	.w6(32'h395d06f3),
	.w7(32'h37ba4043),
	.w8(32'hb9d5f16e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb49f),
	.w1(32'hbc0bd7c3),
	.w2(32'hb9a440aa),
	.w3(32'hbc17980f),
	.w4(32'hbbdd0dc5),
	.w5(32'h3b642cfb),
	.w6(32'hbc29495c),
	.w7(32'hbbb6a2c2),
	.w8(32'h3a1045a9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b3313d),
	.w1(32'hb8447dc9),
	.w2(32'hbafca170),
	.w3(32'h3b1c9ba5),
	.w4(32'hbb0787ae),
	.w5(32'hbb4b2096),
	.w6(32'h3ae7395b),
	.w7(32'hbb74e08c),
	.w8(32'hbbc23543),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7b67c),
	.w1(32'h3b11e2fd),
	.w2(32'h3aa1f809),
	.w3(32'h3ae60223),
	.w4(32'h3a903480),
	.w5(32'h398d2683),
	.w6(32'h3aafec10),
	.w7(32'h3a4cb053),
	.w8(32'h398ffe8b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393085b1),
	.w1(32'h3824911b),
	.w2(32'hba80cca4),
	.w3(32'h3a547da7),
	.w4(32'h399c2d50),
	.w5(32'hba90a849),
	.w6(32'h395ebb73),
	.w7(32'hba040aab),
	.w8(32'hba893648),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e7232),
	.w1(32'hbac557d3),
	.w2(32'hba2cb3e9),
	.w3(32'hbaafb83a),
	.w4(32'hbaa5ec97),
	.w5(32'hb9ca08f8),
	.w6(32'hbaca0aaa),
	.w7(32'hba2d5669),
	.w8(32'hb88777aa),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ff7a8),
	.w1(32'h398b3036),
	.w2(32'h3a38bffb),
	.w3(32'hb6307275),
	.w4(32'h39b171c9),
	.w5(32'h3a084099),
	.w6(32'h355cc16e),
	.w7(32'h3a04e36c),
	.w8(32'h3b03cc01),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0fa36),
	.w1(32'h3a9ae1e5),
	.w2(32'hb93f6db8),
	.w3(32'h3ad5d750),
	.w4(32'h39fcc246),
	.w5(32'hb38024ed),
	.w6(32'h3aff4b2d),
	.w7(32'h3aa9d35f),
	.w8(32'hb9fed041),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f5f3),
	.w1(32'h3965c216),
	.w2(32'hba3e7d42),
	.w3(32'h3b17757a),
	.w4(32'h3a68ef48),
	.w5(32'hbb37d145),
	.w6(32'h3a8b7f16),
	.w7(32'h3ac85e34),
	.w8(32'hbb55869d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba001f2),
	.w1(32'hbbabe733),
	.w2(32'hb8ff97dc),
	.w3(32'hbb8b000c),
	.w4(32'hbb018f92),
	.w5(32'h3a4a2776),
	.w6(32'hbb3081e7),
	.w7(32'h3984ae2c),
	.w8(32'h39f9dac5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918f3a5),
	.w1(32'h38548635),
	.w2(32'h3ac512a8),
	.w3(32'hba261cd8),
	.w4(32'h3a1361de),
	.w5(32'hbabe98d4),
	.w6(32'hb9a70178),
	.w7(32'h3b02e880),
	.w8(32'hba3b183e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903b64),
	.w1(32'hbb68ad3d),
	.w2(32'h3afdc738),
	.w3(32'hbb466f3d),
	.w4(32'hba2bc636),
	.w5(32'h3afe8ab3),
	.w6(32'hbb6b5cfd),
	.w7(32'hba2246dc),
	.w8(32'h3aa0d58c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba112e66),
	.w1(32'h3a9c395b),
	.w2(32'h3aa6058f),
	.w3(32'hbaf5b17e),
	.w4(32'h39eeddd1),
	.w5(32'h3b4fdc15),
	.w6(32'hbaa157f1),
	.w7(32'h39b28232),
	.w8(32'h3b82e639),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affa710),
	.w1(32'h3af61ba4),
	.w2(32'h3a6a7e97),
	.w3(32'h3add96af),
	.w4(32'h3abbda9b),
	.w5(32'h3a987512),
	.w6(32'h3ab1f11d),
	.w7(32'h3a7bf3a8),
	.w8(32'h3a048408),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb8ad2),
	.w1(32'hb929cdc9),
	.w2(32'h39378349),
	.w3(32'h3a990c7c),
	.w4(32'h3a8e9dfc),
	.w5(32'h3910e3de),
	.w6(32'hb9432f70),
	.w7(32'h3a10440c),
	.w8(32'h393038ae),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03c4d3),
	.w1(32'h3a54502c),
	.w2(32'hb8902841),
	.w3(32'h3a19f43c),
	.w4(32'h3a8aae45),
	.w5(32'h39976f2c),
	.w6(32'hba784b72),
	.w7(32'hba3b4bbb),
	.w8(32'h3a05016b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393cdbc1),
	.w1(32'h3a8680eb),
	.w2(32'h3b103355),
	.w3(32'h3a7a8555),
	.w4(32'h3a850894),
	.w5(32'h3b6aa389),
	.w6(32'h3a204e06),
	.w7(32'h3adc7777),
	.w8(32'h3b385a0d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a27b4),
	.w1(32'h3a416bea),
	.w2(32'hb994b0ef),
	.w3(32'h3b9e6ff9),
	.w4(32'h3ac19b61),
	.w5(32'hbb3bc5b6),
	.w6(32'h3b4ce6b9),
	.w7(32'hba3189b1),
	.w8(32'hbaf89b0e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fc79c),
	.w1(32'hba922922),
	.w2(32'h392bc624),
	.w3(32'hba2ee5c7),
	.w4(32'hbac1e93f),
	.w5(32'hbaff7425),
	.w6(32'hb996a808),
	.w7(32'hb97588b6),
	.w8(32'hbac906a9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcb0e0),
	.w1(32'h3974498a),
	.w2(32'h3a3fe723),
	.w3(32'hba50b3c1),
	.w4(32'hb845f62f),
	.w5(32'h3b3e5739),
	.w6(32'h395b4133),
	.w7(32'h38beed7c),
	.w8(32'h3b2aa037),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cd8ab),
	.w1(32'hba33e301),
	.w2(32'h3a8e5c0e),
	.w3(32'hba874f0f),
	.w4(32'hba06de3c),
	.w5(32'h3a2c5c57),
	.w6(32'h39bf727e),
	.w7(32'h3a2bf680),
	.w8(32'h3a96e972),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba596cbf),
	.w1(32'hba898626),
	.w2(32'hba34eb69),
	.w3(32'hb9658d6a),
	.w4(32'hbaa42e2f),
	.w5(32'h3b863bc9),
	.w6(32'hb949800a),
	.w7(32'hba028329),
	.w8(32'h3b5f364d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831d63),
	.w1(32'h3b9d20d4),
	.w2(32'h3c0dfc1c),
	.w3(32'h3b36a5d8),
	.w4(32'h3bc54594),
	.w5(32'h3befd3c1),
	.w6(32'h3a42b739),
	.w7(32'h3b59c91e),
	.w8(32'h3b910b04),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2930b),
	.w1(32'h3a5d5639),
	.w2(32'h3aeaa951),
	.w3(32'h3a830f4a),
	.w4(32'h3ad137d7),
	.w5(32'hba3be2af),
	.w6(32'hba4ba04e),
	.w7(32'h3a04fb9d),
	.w8(32'hba29baa2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72d92d),
	.w1(32'h3770c37f),
	.w2(32'h3a8d6eab),
	.w3(32'hb9b62767),
	.w4(32'hb5eef51e),
	.w5(32'hbb3a1b2c),
	.w6(32'hba04538b),
	.w7(32'h3a6cfcef),
	.w8(32'hba96f833),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa5aa4),
	.w1(32'hba24ef5a),
	.w2(32'h3aff87d9),
	.w3(32'hbb117ae7),
	.w4(32'hbaca48b8),
	.w5(32'h3affda50),
	.w6(32'hbaa3008f),
	.w7(32'hb80ce786),
	.w8(32'h3ada1ec0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca161),
	.w1(32'hba8fd633),
	.w2(32'h3b112be6),
	.w3(32'hba88698d),
	.w4(32'hbaa3200c),
	.w5(32'h3b0ce155),
	.w6(32'hbaaab080),
	.w7(32'hb9826fe5),
	.w8(32'h3adcabe3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02ce9d),
	.w1(32'h39b7824c),
	.w2(32'h39fd9bbc),
	.w3(32'hb8bdf600),
	.w4(32'hba20104c),
	.w5(32'h3aa4b66a),
	.w6(32'h39457799),
	.w7(32'hba0d8d61),
	.w8(32'h3a56e1c7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5f30d),
	.w1(32'h39995802),
	.w2(32'h3a8fb2a5),
	.w3(32'h39f08e7f),
	.w4(32'h3aec359e),
	.w5(32'hba1e3820),
	.w6(32'hb986b464),
	.w7(32'h3a9f81ef),
	.w8(32'hb971e9bd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f36e0),
	.w1(32'h3a17a7bb),
	.w2(32'hb937b8fb),
	.w3(32'hb9755890),
	.w4(32'hba0a401b),
	.w5(32'hb93210ff),
	.w6(32'h38c0d052),
	.w7(32'hb943515d),
	.w8(32'hb80d351a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4ddaf),
	.w1(32'hb9c17a1f),
	.w2(32'hba7b85d9),
	.w3(32'hb97d319e),
	.w4(32'hba352e6e),
	.w5(32'h3a9f7da6),
	.w6(32'hb932662d),
	.w7(32'hba306de1),
	.w8(32'h3a1f8c7b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606844),
	.w1(32'h3a3622e2),
	.w2(32'h3b06e790),
	.w3(32'h3a2472ee),
	.w4(32'h3a980897),
	.w5(32'h3ae13885),
	.w6(32'hb98095c4),
	.w7(32'h3a9ea2a0),
	.w8(32'h3b00bca4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2af258),
	.w1(32'hbae1ebe6),
	.w2(32'h39ea7b61),
	.w3(32'hbaf17679),
	.w4(32'hbad97ab1),
	.w5(32'h37fe9682),
	.w6(32'hba927f97),
	.w7(32'hba0ce884),
	.w8(32'h3a0049f0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6dd2),
	.w1(32'hb9fecd96),
	.w2(32'hb9c086e2),
	.w3(32'hbb22b4bf),
	.w4(32'hbb26e823),
	.w5(32'h3ab9cf2a),
	.w6(32'hbb2a32cb),
	.w7(32'hbab5e0af),
	.w8(32'h3a26a1e2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdd26b),
	.w1(32'h3afd28f3),
	.w2(32'h3b2a1ab7),
	.w3(32'h3af4adee),
	.w4(32'h3b3fbb03),
	.w5(32'hbb065e64),
	.w6(32'h3aef2c02),
	.w7(32'h3b149ad1),
	.w8(32'hbabd9698),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163254),
	.w1(32'hbaf158e0),
	.w2(32'h3ab77e0f),
	.w3(32'hbb455554),
	.w4(32'hbaafd252),
	.w5(32'h3bcbcf7c),
	.w6(32'hbb694ffe),
	.w7(32'hbb005f76),
	.w8(32'h3bb5d3b4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420a48),
	.w1(32'h3b2dc74c),
	.w2(32'h3b2f2b7e),
	.w3(32'h3b0ee75a),
	.w4(32'h3b1873e0),
	.w5(32'h3a41c242),
	.w6(32'h3b3e268d),
	.w7(32'h3b481024),
	.w8(32'h39221035),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e44ff),
	.w1(32'hbaadd098),
	.w2(32'hba610c55),
	.w3(32'h3a8fa66f),
	.w4(32'h3ad89f55),
	.w5(32'h3aff5825),
	.w6(32'hb9cb2f28),
	.w7(32'h39ad157e),
	.w8(32'h3b2065c7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab872),
	.w1(32'h3b060e05),
	.w2(32'h3acc3e2c),
	.w3(32'h3ac87257),
	.w4(32'h3a077baa),
	.w5(32'h3ae072c4),
	.w6(32'h3b103312),
	.w7(32'h3aa831bf),
	.w8(32'h3b106419),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab36137),
	.w1(32'h3a53ca0d),
	.w2(32'h39f71db0),
	.w3(32'h3a69f692),
	.w4(32'h3a312227),
	.w5(32'h3b5160c8),
	.w6(32'h39aba35c),
	.w7(32'h3a31c33f),
	.w8(32'h3ae14b62),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39a2a3),
	.w1(32'hbb62328f),
	.w2(32'hbb0a82b6),
	.w3(32'hbb4f76d9),
	.w4(32'hba18a045),
	.w5(32'hbb3ad7cb),
	.w6(32'hbbbe4a44),
	.w7(32'hbb4959fa),
	.w8(32'hbb2f9643),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6363a2),
	.w1(32'hbb30d497),
	.w2(32'h3a133858),
	.w3(32'h3ae38602),
	.w4(32'hbbb50043),
	.w5(32'h3b4668c0),
	.w6(32'h3b17586b),
	.w7(32'hba7060d4),
	.w8(32'h3aeaf778),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba62e1d),
	.w1(32'h3b9dd3a3),
	.w2(32'h3b944df9),
	.w3(32'hbad272d6),
	.w4(32'h3ab024ca),
	.w5(32'h392f239e),
	.w6(32'hbbdc8329),
	.w7(32'hbb4d8078),
	.w8(32'hb9624045),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb372469),
	.w1(32'hbbf2f56f),
	.w2(32'hbbbed643),
	.w3(32'h3b7a9ead),
	.w4(32'h37ae51c1),
	.w5(32'hbac3de91),
	.w6(32'hbb6556b5),
	.w7(32'hbbb35993),
	.w8(32'hba4801a6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f1fd39),
	.w1(32'hbad28afa),
	.w2(32'hb95a93e1),
	.w3(32'hbb8397de),
	.w4(32'h37ece624),
	.w5(32'hbaa928e6),
	.w6(32'hbb9e5e5e),
	.w7(32'h3ac267e6),
	.w8(32'h3b1468da),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba57e),
	.w1(32'hbb079986),
	.w2(32'hbab68516),
	.w3(32'hbb279a9e),
	.w4(32'hbb33d2cf),
	.w5(32'hbb749eab),
	.w6(32'hbb21bc6e),
	.w7(32'hba80228e),
	.w8(32'hbb352ed6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c9ab9),
	.w1(32'hbaa0e148),
	.w2(32'h3bdb0a08),
	.w3(32'h3a0308ce),
	.w4(32'h3b42e8fd),
	.w5(32'hbaf2141a),
	.w6(32'hbb4244f8),
	.w7(32'h3ba9c539),
	.w8(32'hbae5ce1f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb653b81),
	.w1(32'hbae65548),
	.w2(32'h3a605d72),
	.w3(32'h3998da46),
	.w4(32'hba3b32d0),
	.w5(32'hbb430966),
	.w6(32'h3b11d397),
	.w7(32'h3b1c4b50),
	.w8(32'hbad066be),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a153c64),
	.w1(32'hbb46893d),
	.w2(32'hbac71ab6),
	.w3(32'hbbf7599b),
	.w4(32'hbb33d03d),
	.w5(32'hbad9cde7),
	.w6(32'hba779a31),
	.w7(32'hbafedf0f),
	.w8(32'hbb3ba22e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcf0ec),
	.w1(32'h3b6221e0),
	.w2(32'h380e5285),
	.w3(32'h3ae56e79),
	.w4(32'hbb0b5bc7),
	.w5(32'h3c0e6cc1),
	.w6(32'h3b7c9ca3),
	.w7(32'h3a3f0cb7),
	.w8(32'h3bcbc1d5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be37ef2),
	.w1(32'hbaa4a879),
	.w2(32'hbb036515),
	.w3(32'hbaabe007),
	.w4(32'hba501444),
	.w5(32'h3a6bc0a9),
	.w6(32'hbb662ca4),
	.w7(32'hbb016676),
	.w8(32'h3b70e1f8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5efd48),
	.w1(32'h3af04f92),
	.w2(32'hbb38382b),
	.w3(32'h3aa38b8a),
	.w4(32'h3a69a84b),
	.w5(32'hbb9c6bbc),
	.w6(32'h3b0f4338),
	.w7(32'hbafc2919),
	.w8(32'hbb35fa38),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2c89),
	.w1(32'h3b03d69c),
	.w2(32'h3a5f5bd4),
	.w3(32'hbb9e8994),
	.w4(32'h3a8d4ef8),
	.w5(32'hbaf6b3a1),
	.w6(32'h3aa26a2e),
	.w7(32'h3aa684c3),
	.w8(32'hbb87ff6a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ec95),
	.w1(32'hbb578dba),
	.w2(32'h393ad7be),
	.w3(32'hbb27b510),
	.w4(32'hbbb20b30),
	.w5(32'h37bc5ed9),
	.w6(32'hbaebebf1),
	.w7(32'hbbad6cbe),
	.w8(32'hb8d25654),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c29cd),
	.w1(32'hba6eb440),
	.w2(32'h3a6d9acf),
	.w3(32'hbbe74606),
	.w4(32'hba17b746),
	.w5(32'hbb1bdacc),
	.w6(32'hbb9a053f),
	.w7(32'h3b8c51b5),
	.w8(32'hba3b7f92),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab68d0f),
	.w1(32'h3b83465a),
	.w2(32'h3b499166),
	.w3(32'hbbdc0650),
	.w4(32'hbb83f545),
	.w5(32'hbad3b206),
	.w6(32'hbb9531a3),
	.w7(32'hbb10457a),
	.w8(32'hbbb21d40),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ad35),
	.w1(32'h3c1de2e8),
	.w2(32'h3b15d780),
	.w3(32'h3b986d83),
	.w4(32'hbbc66478),
	.w5(32'hb98ef1c1),
	.w6(32'h3c1908bd),
	.w7(32'hbbd8408a),
	.w8(32'hba15a2d9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f64fc),
	.w1(32'hbb964b86),
	.w2(32'hbb004283),
	.w3(32'hba88bfff),
	.w4(32'hbbbf42f5),
	.w5(32'h3c3fd96f),
	.w6(32'hba9c97fb),
	.w7(32'hbbca25a3),
	.w8(32'h3bf35a90),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2aa82),
	.w1(32'h39f8d023),
	.w2(32'hba220f54),
	.w3(32'h3b59c92c),
	.w4(32'h3b89b176),
	.w5(32'h3b463a6c),
	.w6(32'hbb62e478),
	.w7(32'hbadf274e),
	.w8(32'h3c0c1b8b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce920b),
	.w1(32'hbbec72e9),
	.w2(32'h3bfbef58),
	.w3(32'h3b8c487d),
	.w4(32'h3b71f60a),
	.w5(32'h3b41d807),
	.w6(32'h3bf2f61e),
	.w7(32'h3bdc3846),
	.w8(32'h3b26c1dd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5d258),
	.w1(32'h3b7129fe),
	.w2(32'h3bb041cd),
	.w3(32'h3ae90883),
	.w4(32'h3b9837f1),
	.w5(32'h373984ad),
	.w6(32'hbb0a53e9),
	.w7(32'h3b17146b),
	.w8(32'hbbba9aac),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e1b4),
	.w1(32'hbb40827c),
	.w2(32'h3a424877),
	.w3(32'hbbaaa056),
	.w4(32'h3b0ccf09),
	.w5(32'hba1518eb),
	.w6(32'hbc196e71),
	.w7(32'h3ae0289a),
	.w8(32'hb9351286),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75e79c),
	.w1(32'hbb7bdb36),
	.w2(32'hbb4bd138),
	.w3(32'hbad229de),
	.w4(32'hbb8b3276),
	.w5(32'hbb99f231),
	.w6(32'h38bac324),
	.w7(32'hbb73b490),
	.w8(32'hbb24b47a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac56c01),
	.w1(32'hba2727cb),
	.w2(32'h3abe19d3),
	.w3(32'hbba7312b),
	.w4(32'hbafa7ce7),
	.w5(32'hbb892930),
	.w6(32'hbb89c114),
	.w7(32'h3b14786d),
	.w8(32'hbb6bd4ea),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbe380),
	.w1(32'hbb03df5c),
	.w2(32'hbbb1c4e9),
	.w3(32'hbb4f003e),
	.w4(32'hbb414d5f),
	.w5(32'hbb0c7468),
	.w6(32'h3bbc6213),
	.w7(32'h3b2b20e1),
	.w8(32'hbb4f28e8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bdb9d),
	.w1(32'h38b5ebcb),
	.w2(32'hbbf90306),
	.w3(32'hbaea401b),
	.w4(32'hbb6c7824),
	.w5(32'hbba7957c),
	.w6(32'hbb8c30a5),
	.w7(32'hbb8efbab),
	.w8(32'h3a1f0aa9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94a337),
	.w1(32'h3a0b9fa3),
	.w2(32'hbbbbd556),
	.w3(32'hbb05ef17),
	.w4(32'h39157a75),
	.w5(32'h3a1c3b3a),
	.w6(32'h3bcce5fc),
	.w7(32'hba0ba7da),
	.w8(32'hba23305f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad25b62),
	.w1(32'hbaa9c3c3),
	.w2(32'hbb7ae874),
	.w3(32'h3b2186e7),
	.w4(32'h3ac1004c),
	.w5(32'h3b927377),
	.w6(32'h3ad288d8),
	.w7(32'hbb43c22f),
	.w8(32'hbb268ea4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b5cf),
	.w1(32'hbaa43bdc),
	.w2(32'hbb1b9e8e),
	.w3(32'h3b170c84),
	.w4(32'hbb0fcaf0),
	.w5(32'h3b51869f),
	.w6(32'hbbd0beab),
	.w7(32'hbbdc7133),
	.w8(32'h3b4e37d7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e771),
	.w1(32'h3c3e0d4d),
	.w2(32'h3b86e45d),
	.w3(32'h3ba07ddc),
	.w4(32'hba2333a6),
	.w5(32'h3b11a923),
	.w6(32'h3bf6e607),
	.w7(32'hb9758a42),
	.w8(32'h3b5141bc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule