module layer_6_featuremap_126(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c535),
	.w1(32'hbb6a680a),
	.w2(32'hbb2961de),
	.w3(32'hbb7b57c4),
	.w4(32'hbb71c582),
	.w5(32'hbb331e5f),
	.w6(32'hbb7231b6),
	.w7(32'hbb79a315),
	.w8(32'hbb1d843a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa655e4),
	.w1(32'hb8926104),
	.w2(32'hb9a8e8a6),
	.w3(32'h39f43be3),
	.w4(32'h3a2f637e),
	.w5(32'h3a11428b),
	.w6(32'h3a9e6162),
	.w7(32'h3a857abf),
	.w8(32'h3961c89e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654417),
	.w1(32'hbb06a5a8),
	.w2(32'hbb6202cc),
	.w3(32'hbb17df88),
	.w4(32'h3b080447),
	.w5(32'h3b1a03e1),
	.w6(32'hbbcafead),
	.w7(32'hbb109356),
	.w8(32'hbaeac96c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad87de),
	.w1(32'hbb4df204),
	.w2(32'hbbc06116),
	.w3(32'hb8cc2f8a),
	.w4(32'hbaf072c2),
	.w5(32'hbb9aaa7a),
	.w6(32'h38eb1556),
	.w7(32'hbb0d739b),
	.w8(32'hbb5bfbe1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a23b1d),
	.w1(32'h3ac4a01b),
	.w2(32'hb777f9d6),
	.w3(32'h3ab1e75c),
	.w4(32'h399e0f41),
	.w5(32'h393f48d8),
	.w6(32'h3a6aa0f8),
	.w7(32'h3ad4be6d),
	.w8(32'hba5b70b8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874b622),
	.w1(32'hbb228473),
	.w2(32'hba90aeb7),
	.w3(32'hbb8c532f),
	.w4(32'hbb53a158),
	.w5(32'hbb092594),
	.w6(32'hbb6fef14),
	.w7(32'hbb1efe54),
	.w8(32'hba7b06cc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bcd74),
	.w1(32'h3c0c76d0),
	.w2(32'h3bf1435a),
	.w3(32'h3c16d503),
	.w4(32'h3c326105),
	.w5(32'h3c1a5afa),
	.w6(32'h3becda6b),
	.w7(32'h3c035ffa),
	.w8(32'h3bd41362),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada3c08),
	.w1(32'h3b43ec6e),
	.w2(32'h3b8371c1),
	.w3(32'h3b7f5475),
	.w4(32'h3b540df1),
	.w5(32'h3b77b457),
	.w6(32'h3b05e367),
	.w7(32'h3b9115c4),
	.w8(32'h3b21cbd4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14bf93),
	.w1(32'h3ab2bfbb),
	.w2(32'hbb0c2131),
	.w3(32'hb8da77d4),
	.w4(32'h3b16c95a),
	.w5(32'h3af3fa3d),
	.w6(32'h39c39836),
	.w7(32'h3b0a6203),
	.w8(32'hba156db2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23b66),
	.w1(32'h3a66ffd6),
	.w2(32'h3b4b1501),
	.w3(32'h38ee5606),
	.w4(32'h3a278517),
	.w5(32'h3acff4fe),
	.w6(32'h38e79548),
	.w7(32'h3acd65a1),
	.w8(32'h3b340005),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1f0e2),
	.w1(32'hbaa67757),
	.w2(32'hbb6b2da0),
	.w3(32'hb92f9242),
	.w4(32'hba622e76),
	.w5(32'h3accf512),
	.w6(32'hba7c6e62),
	.w7(32'hba68a0f5),
	.w8(32'h3a452e1c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fa4b4),
	.w1(32'h3928e31f),
	.w2(32'h3a1cb452),
	.w3(32'h38163b29),
	.w4(32'h3a1b0dac),
	.w5(32'h3ad3cd77),
	.w6(32'hba3f240a),
	.w7(32'hb94fcd96),
	.w8(32'h3ac841c2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038acd),
	.w1(32'h3a9b524a),
	.w2(32'h3ab8664d),
	.w3(32'h3a9e1802),
	.w4(32'h3ae1c8f8),
	.w5(32'h3a53f034),
	.w6(32'h3aef1ad3),
	.w7(32'h3b07b7ba),
	.w8(32'h3a532ab5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeed9a),
	.w1(32'h3ba4e4bb),
	.w2(32'h3b073b5a),
	.w3(32'h3b69d7d8),
	.w4(32'h3c092330),
	.w5(32'h3c23f87d),
	.w6(32'h3ba09437),
	.w7(32'h3bd7a45b),
	.w8(32'h3c02ee5b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade5b94),
	.w1(32'hba9378bc),
	.w2(32'hba99186f),
	.w3(32'hb9dc0484),
	.w4(32'hbaa8e69a),
	.w5(32'hba521b9b),
	.w6(32'hba579504),
	.w7(32'hba6c913c),
	.w8(32'h3948c616),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c3809),
	.w1(32'hbafbbe6a),
	.w2(32'hbb211f26),
	.w3(32'hbaadf1d8),
	.w4(32'hbabfaab0),
	.w5(32'hbaa9d413),
	.w6(32'hbaa692e9),
	.w7(32'hba316fc5),
	.w8(32'hba5c0749),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191877),
	.w1(32'hbaae12c9),
	.w2(32'hbb905e05),
	.w3(32'hbae4a9e3),
	.w4(32'h3c069252),
	.w5(32'h3c1691a7),
	.w6(32'hba0c68ef),
	.w7(32'h3c674905),
	.w8(32'h3c780dad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997e3ba),
	.w1(32'hb9b7c95e),
	.w2(32'h3975a38b),
	.w3(32'hbaae3e6f),
	.w4(32'hba855c2a),
	.w5(32'hb915bc3f),
	.w6(32'hbaaa273b),
	.w7(32'hba53a9bb),
	.w8(32'h392b0cb4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ac92),
	.w1(32'h3acba057),
	.w2(32'h3ab50f6f),
	.w3(32'h3b64d1a1),
	.w4(32'h3b0a2b08),
	.w5(32'h3a8be314),
	.w6(32'h3b3266b1),
	.w7(32'h3ae46748),
	.w8(32'h3aafd2ce),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84fbfef),
	.w1(32'hb9b4bb50),
	.w2(32'h3a30f8a0),
	.w3(32'h3a11e2af),
	.w4(32'h3a466c76),
	.w5(32'h3b1f3f21),
	.w6(32'h398be7cc),
	.w7(32'h3b12e7c2),
	.w8(32'h3b2c1d01),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38529385),
	.w1(32'hb9ae329b),
	.w2(32'hbae5ffdc),
	.w3(32'h385dc446),
	.w4(32'h399bd759),
	.w5(32'hba9b06b8),
	.w6(32'hb9251435),
	.w7(32'hb899cf05),
	.w8(32'hbaabc860),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87afde),
	.w1(32'hba6c5125),
	.w2(32'hbb8f5001),
	.w3(32'hba6ce8fd),
	.w4(32'h3a125b21),
	.w5(32'h3a82ce1c),
	.w6(32'hbb2ff19a),
	.w7(32'hba7c6fcf),
	.w8(32'hb8fee856),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc9cd6),
	.w1(32'h3a520436),
	.w2(32'h3b84ea0c),
	.w3(32'hbac8e115),
	.w4(32'h3aab5248),
	.w5(32'h3a0dfacf),
	.w6(32'h396138e5),
	.w7(32'h3b18eb1a),
	.w8(32'h3b2b803d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b120dea),
	.w1(32'h39fa12fa),
	.w2(32'hbb11b9cb),
	.w3(32'hbba6b472),
	.w4(32'hbb5bdf0a),
	.w5(32'h3a9d5d9c),
	.w6(32'hbb23a4c4),
	.w7(32'hba617ed7),
	.w8(32'h3ad90386),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974eb1),
	.w1(32'hba76aeb7),
	.w2(32'hbb8752ca),
	.w3(32'h3a9f63e1),
	.w4(32'h3b6b90e8),
	.w5(32'h3a2fd100),
	.w6(32'hbb4b32d7),
	.w7(32'h38a25bb9),
	.w8(32'h3b8b77d8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2e17f),
	.w1(32'h3b02450b),
	.w2(32'hb6ee4ad0),
	.w3(32'h3ab42cc6),
	.w4(32'hba6d59a4),
	.w5(32'hbb38ed9c),
	.w6(32'hba44ce22),
	.w7(32'hb9fadf63),
	.w8(32'h3b1187d2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc906d),
	.w1(32'h3b29a28e),
	.w2(32'hba8961cf),
	.w3(32'hb9816366),
	.w4(32'h3b219ce0),
	.w5(32'h3b6a849a),
	.w6(32'h39b9e0b2),
	.w7(32'hbb0de0f7),
	.w8(32'hb9610d1a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ae334),
	.w1(32'h3b242aa4),
	.w2(32'h3acdb4fe),
	.w3(32'h3b86e435),
	.w4(32'h3b8d1b75),
	.w5(32'h3aff1cda),
	.w6(32'h3b51000f),
	.w7(32'h3b1bebeb),
	.w8(32'h3972aa95),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8511c4),
	.w1(32'h398fdc9d),
	.w2(32'hb7d69ebb),
	.w3(32'h3a1c27be),
	.w4(32'h398b3cec),
	.w5(32'h39e3b34b),
	.w6(32'h398b7c86),
	.w7(32'hb8d31001),
	.w8(32'h395c94b3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc177b3),
	.w1(32'hbb8da4e9),
	.w2(32'hbb02f8a2),
	.w3(32'h3bcacda1),
	.w4(32'hbb8c9b5a),
	.w5(32'hbc3f0415),
	.w6(32'h3c307f18),
	.w7(32'hbc056f1a),
	.w8(32'hbb109c8e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa047a0),
	.w1(32'hbae4da12),
	.w2(32'hbb628524),
	.w3(32'hb92ab215),
	.w4(32'hba341955),
	.w5(32'hb9a6619e),
	.w6(32'hbaf06229),
	.w7(32'hbb6874f4),
	.w8(32'hbb479a55),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb585c),
	.w1(32'hbafe7403),
	.w2(32'hbb2876b1),
	.w3(32'hbb838f9d),
	.w4(32'hbb6cb0e1),
	.w5(32'hbb14b580),
	.w6(32'hbb766168),
	.w7(32'hbb383312),
	.w8(32'hba0c0841),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0667ed),
	.w1(32'hba70b389),
	.w2(32'hbb4c1be1),
	.w3(32'hba1c4489),
	.w4(32'hbacefac3),
	.w5(32'hba843454),
	.w6(32'hba835a86),
	.w7(32'hbb187810),
	.w8(32'hbb0553fb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35b367),
	.w1(32'h3aae3d6a),
	.w2(32'h3aadd306),
	.w3(32'h38438bba),
	.w4(32'h3aa0634e),
	.w5(32'h3a37a25b),
	.w6(32'h3b0c3708),
	.w7(32'h3aa2b58f),
	.w8(32'h3b09cf10),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fffc4),
	.w1(32'hbaf2650b),
	.w2(32'hba279b75),
	.w3(32'hbb63c37c),
	.w4(32'hbb1dfd68),
	.w5(32'hbac7239d),
	.w6(32'hbb32eb08),
	.w7(32'hbacb86c3),
	.w8(32'hb9a36ba1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e56b08),
	.w1(32'hba9a3d0b),
	.w2(32'hbb0874b1),
	.w3(32'hba05bd13),
	.w4(32'hb817c68d),
	.w5(32'hbacf4518),
	.w6(32'hb846089e),
	.w7(32'h3ab1ae29),
	.w8(32'h3a8e126c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2777ce),
	.w1(32'h3a255fa4),
	.w2(32'h3a841935),
	.w3(32'h39afec99),
	.w4(32'h38f92e83),
	.w5(32'h3a244f72),
	.w6(32'hba1309ed),
	.w7(32'hba23cafc),
	.w8(32'h3a12749f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16a640),
	.w1(32'h3b5acbee),
	.w2(32'h3b15d859),
	.w3(32'h3ba0a86b),
	.w4(32'h3bb712a6),
	.w5(32'h3b6b62ce),
	.w6(32'h3b95c1ae),
	.w7(32'h3bc7e690),
	.w8(32'h3bc5930f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6a907),
	.w1(32'h3a80e2d5),
	.w2(32'h3a7561fa),
	.w3(32'h3b27b119),
	.w4(32'h3b31753b),
	.w5(32'h37dbd668),
	.w6(32'h3afde6eb),
	.w7(32'h3897aed6),
	.w8(32'hbab86c6c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36444),
	.w1(32'h38e56111),
	.w2(32'hbc4a7566),
	.w3(32'h3b305f37),
	.w4(32'h3c0e4794),
	.w5(32'h3c101cf5),
	.w6(32'hba4dac1a),
	.w7(32'h3aef1010),
	.w8(32'h3a63c153),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b7bca),
	.w1(32'hb9ca941f),
	.w2(32'hb947f7e3),
	.w3(32'h3b84a953),
	.w4(32'h3b5a6417),
	.w5(32'h3ba80d08),
	.w6(32'h3aa230cc),
	.w7(32'h3b3c3c08),
	.w8(32'h3bbe97d8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe599),
	.w1(32'h3b0bb4ec),
	.w2(32'h3a8fc5a1),
	.w3(32'h3b8f3264),
	.w4(32'h3b6a75b8),
	.w5(32'h3b00d93e),
	.w6(32'h3b80cc3c),
	.w7(32'h3b63790b),
	.w8(32'h3b2070f7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a44c14),
	.w1(32'hba0f1b77),
	.w2(32'hb97b2410),
	.w3(32'hbaac2a3f),
	.w4(32'hbaaacc7d),
	.w5(32'hba4faed0),
	.w6(32'hbaacc023),
	.w7(32'hba7efeab),
	.w8(32'hb8d827b8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5bdde),
	.w1(32'hbbc86ddd),
	.w2(32'hbb7d9063),
	.w3(32'h3ac812d8),
	.w4(32'hbb30ac49),
	.w5(32'hbc6bac9f),
	.w6(32'h3a412f03),
	.w7(32'hbb3f96d3),
	.w8(32'hbb46c453),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4f84),
	.w1(32'h3b7cd847),
	.w2(32'hba5f87a2),
	.w3(32'h3a0a15ae),
	.w4(32'h3b9a118c),
	.w5(32'h3bb03b3d),
	.w6(32'hbaa2c720),
	.w7(32'h3adc3553),
	.w8(32'h3b3f7b99),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975ae54),
	.w1(32'hbb87ca7e),
	.w2(32'hbb7979ab),
	.w3(32'hbb4d646b),
	.w4(32'hbb0279bd),
	.w5(32'hbb53779e),
	.w6(32'hbac647f3),
	.w7(32'hbb23c869),
	.w8(32'hbb003522),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031ae0),
	.w1(32'h3a333c01),
	.w2(32'hb991384c),
	.w3(32'h3a6dd848),
	.w4(32'h3a31a737),
	.w5(32'h3a5a5a9f),
	.w6(32'h3ad899ab),
	.w7(32'h3a9df729),
	.w8(32'hba03dafe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc957b1),
	.w1(32'hbb23d01f),
	.w2(32'hba354d76),
	.w3(32'hba933c1f),
	.w4(32'h3a28c02c),
	.w5(32'h3a587b67),
	.w6(32'h3ac5394b),
	.w7(32'h3b30f4c4),
	.w8(32'h3b14af80),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d8c28),
	.w1(32'hbabc619b),
	.w2(32'hbabfcb6e),
	.w3(32'h3b0d42f8),
	.w4(32'h3aa467aa),
	.w5(32'h3aba01cb),
	.w6(32'h3aba86eb),
	.w7(32'h3ae6c69f),
	.w8(32'h3aec859a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab4cf),
	.w1(32'hbba7821f),
	.w2(32'hbbae9f85),
	.w3(32'hbbb34eee),
	.w4(32'hbb131bf9),
	.w5(32'hbb242611),
	.w6(32'hbba4ac6a),
	.w7(32'hbb800674),
	.w8(32'hbb19cab2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc7a4),
	.w1(32'h3a06d6c2),
	.w2(32'hbae24a2e),
	.w3(32'h3a2d9409),
	.w4(32'h3b179bd4),
	.w5(32'h39e1024e),
	.w6(32'h383a28c3),
	.w7(32'h3afb12f7),
	.w8(32'h3adab033),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fe00b),
	.w1(32'hbaf01043),
	.w2(32'h394193d9),
	.w3(32'h3aaed261),
	.w4(32'h3a888038),
	.w5(32'h3b026ebd),
	.w6(32'h3ac986c7),
	.w7(32'h3b248a62),
	.w8(32'h3b2f43ae),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2589ea),
	.w1(32'h3bc0b852),
	.w2(32'h3b10c9fa),
	.w3(32'h3b8c00ec),
	.w4(32'h3c343715),
	.w5(32'h3c25aa10),
	.w6(32'h3b9bf417),
	.w7(32'h3c1d5ddf),
	.w8(32'h3be488be),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398be31f),
	.w1(32'h3b9e3413),
	.w2(32'h3b86b913),
	.w3(32'h3c13f5fb),
	.w4(32'h3c21e311),
	.w5(32'h3c29c5f8),
	.w6(32'h3c194b40),
	.w7(32'h3c0f2fb3),
	.w8(32'h3be20f20),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522441),
	.w1(32'h3ba80f64),
	.w2(32'h3bd933b1),
	.w3(32'h3bdd48c5),
	.w4(32'h3c093107),
	.w5(32'h3c085d29),
	.w6(32'h3bc96a53),
	.w7(32'h3bd80291),
	.w8(32'h3bd2dddd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98a76d),
	.w1(32'hbd0160c8),
	.w2(32'hbc332358),
	.w3(32'hba2f94b5),
	.w4(32'hbc358610),
	.w5(32'hbc6e0f6e),
	.w6(32'hbbc3cd63),
	.w7(32'hbca897e1),
	.w8(32'h3a4f7cd8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be25ad9),
	.w1(32'h3b96b5f9),
	.w2(32'h3b651086),
	.w3(32'hbb2e6073),
	.w4(32'h3b0f93fb),
	.w5(32'h3bb261d9),
	.w6(32'hb8f58ea5),
	.w7(32'h3bae1f7f),
	.w8(32'h3b5c7bf5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ed1c2),
	.w1(32'h3ba5c579),
	.w2(32'hbb880b03),
	.w3(32'h3c82dc97),
	.w4(32'h3af3ae93),
	.w5(32'h3c319a9f),
	.w6(32'h3c4bd2cc),
	.w7(32'hbc5dd72c),
	.w8(32'h3ccdc1c6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda1690),
	.w1(32'hbb29df25),
	.w2(32'hbbde0109),
	.w3(32'h3adfe69a),
	.w4(32'hbabe495a),
	.w5(32'hbb69526e),
	.w6(32'h3a6d32d7),
	.w7(32'hbb34b0a1),
	.w8(32'hbb999bdd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f9701),
	.w1(32'hbb94b479),
	.w2(32'h3cacd4ed),
	.w3(32'hbd3e54f2),
	.w4(32'h3bbe6bcd),
	.w5(32'h3d400754),
	.w6(32'hbd262a41),
	.w7(32'h3d1e3d0f),
	.w8(32'h3d75e769),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94336e),
	.w1(32'h3b0efe99),
	.w2(32'hbc68690f),
	.w3(32'h3c2402d8),
	.w4(32'hbb51e61c),
	.w5(32'hbc3b2722),
	.w6(32'h3c4d9f54),
	.w7(32'hbc1cc6e0),
	.w8(32'hbc3ece95),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc440ab0),
	.w1(32'hbc35df25),
	.w2(32'hbd1b5bac),
	.w3(32'h3bfc066f),
	.w4(32'hbd24923e),
	.w5(32'hbcc6f8f7),
	.w6(32'hbb9c5f3a),
	.w7(32'hbd43ac4a),
	.w8(32'h39b1ee45),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ecd0),
	.w1(32'hbcf43017),
	.w2(32'h3b41f131),
	.w3(32'hbca503ba),
	.w4(32'h3bb0caf3),
	.w5(32'hbc10d908),
	.w6(32'hbc76476a),
	.w7(32'h3b8cb73d),
	.w8(32'hbcf7c36e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9400be),
	.w1(32'h3ba06430),
	.w2(32'hbb8e69fb),
	.w3(32'h3c9f7f4b),
	.w4(32'h3bd5d3ea),
	.w5(32'hbb26423a),
	.w6(32'h3c8c0f00),
	.w7(32'hbb34be00),
	.w8(32'hbab58f39),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule