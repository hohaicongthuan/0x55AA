module layer_6_featuremap_117(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cdf99),
	.w1(32'h39201779),
	.w2(32'hba811dfd),
	.w3(32'hba206341),
	.w4(32'hba6e2fe4),
	.w5(32'hbb175a49),
	.w6(32'hbab43888),
	.w7(32'hb99ec5cd),
	.w8(32'hba05bcd4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba659e32),
	.w1(32'hbb1118d6),
	.w2(32'hbaf9f1f4),
	.w3(32'hb9540164),
	.w4(32'hb97913e2),
	.w5(32'hb98851b0),
	.w6(32'h3a0c7f2c),
	.w7(32'h3a61866a),
	.w8(32'h3a90c4ae),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d5dcf),
	.w1(32'hbc6ab31b),
	.w2(32'hba297f16),
	.w3(32'h3c00aed8),
	.w4(32'hba73bca7),
	.w5(32'hbc278101),
	.w6(32'h3ae55691),
	.w7(32'h3b782bc6),
	.w8(32'h3b978cfc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2b66),
	.w1(32'hbb440e30),
	.w2(32'hbb6332c8),
	.w3(32'hba025de8),
	.w4(32'hbab1eba6),
	.w5(32'hba447c3b),
	.w6(32'h39c8254c),
	.w7(32'hba6af959),
	.w8(32'hbaf3fca4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaaf42),
	.w1(32'h3a68c2a2),
	.w2(32'h3ac05360),
	.w3(32'h3b190595),
	.w4(32'hb9486a37),
	.w5(32'hbab583f4),
	.w6(32'h3b74cf64),
	.w7(32'h3ae722e2),
	.w8(32'h3b3039b5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3860b6f1),
	.w1(32'h3a8742a2),
	.w2(32'h39c6165b),
	.w3(32'hbb3eef93),
	.w4(32'hbb719c3f),
	.w5(32'hbb926519),
	.w6(32'hba70b2b5),
	.w7(32'hbaaa4d22),
	.w8(32'hbb1da13d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38351c),
	.w1(32'hbaa5f5a4),
	.w2(32'h3914ee9f),
	.w3(32'h3b796531),
	.w4(32'h3bae31ba),
	.w5(32'h3bce5c16),
	.w6(32'h3ab33bea),
	.w7(32'h3b3e8ebb),
	.w8(32'h3b90ae91),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03cfe3),
	.w1(32'h3b31ec0a),
	.w2(32'h3b56e999),
	.w3(32'h3b3542ab),
	.w4(32'h3a7df2a2),
	.w5(32'h38f66368),
	.w6(32'h3a5244b5),
	.w7(32'h3b0dc0dd),
	.w8(32'h399e615e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4130ac),
	.w1(32'hbaeb3579),
	.w2(32'h3b67678d),
	.w3(32'h3bb9b7d3),
	.w4(32'hb94596f4),
	.w5(32'hbb0e63f3),
	.w6(32'hb8100a84),
	.w7(32'h3b9e61fa),
	.w8(32'hb9ea7fb9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e157),
	.w1(32'hb93168de),
	.w2(32'hba2600e8),
	.w3(32'hbb0757ee),
	.w4(32'hbb993c98),
	.w5(32'hbba41d72),
	.w6(32'h3ad13af8),
	.w7(32'hbaaeeaac),
	.w8(32'hbb7c89db),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa581a),
	.w1(32'hbb5ed168),
	.w2(32'hbb37809f),
	.w3(32'h3bdf3c5d),
	.w4(32'h3ab5c7d6),
	.w5(32'hbb3038a8),
	.w6(32'hba601ceb),
	.w7(32'hb990cb0e),
	.w8(32'h3ac68451),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8a9b),
	.w1(32'hb925ffd4),
	.w2(32'h385141bb),
	.w3(32'h39bc0ff1),
	.w4(32'h37e00019),
	.w5(32'h39a6b4d6),
	.w6(32'hba890e33),
	.w7(32'hba700664),
	.w8(32'hb8c5d30b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028ad7),
	.w1(32'hba1ec9bc),
	.w2(32'h3a0fc477),
	.w3(32'hb673061a),
	.w4(32'h3ac985f1),
	.w5(32'h3a85b059),
	.w6(32'hb9972580),
	.w7(32'h3a9dc708),
	.w8(32'h3a931d9a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b91e2),
	.w1(32'h3a39de5e),
	.w2(32'h3c175335),
	.w3(32'h3c50c6d5),
	.w4(32'h3bd5be04),
	.w5(32'hbb05d2d5),
	.w6(32'h3b758b1d),
	.w7(32'h3bf5c5a3),
	.w8(32'h3c167c2d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228b1b),
	.w1(32'hbabc54dd),
	.w2(32'hbb13bcdb),
	.w3(32'h3a314e51),
	.w4(32'hbaa69b4b),
	.w5(32'hbb01f482),
	.w6(32'h3b01f040),
	.w7(32'hba564b57),
	.w8(32'hbb369a41),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9abd96),
	.w1(32'hbb3497a2),
	.w2(32'hba9c2a2d),
	.w3(32'hbb858cea),
	.w4(32'hbb8ace8f),
	.w5(32'hbb76d014),
	.w6(32'hbb1f2e9c),
	.w7(32'hbb263a96),
	.w8(32'hbb4da3a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f6a9d),
	.w1(32'hbc4cb82a),
	.w2(32'hbb81797b),
	.w3(32'hbbd1fd70),
	.w4(32'hbc8da90b),
	.w5(32'hbc8056b2),
	.w6(32'hbb8d4c47),
	.w7(32'hbc3deef3),
	.w8(32'hbc74669e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9053379),
	.w1(32'h3a8e1aa4),
	.w2(32'h3a92abaa),
	.w3(32'hb9c0fa2f),
	.w4(32'hba67c8b4),
	.w5(32'hba79c7ba),
	.w6(32'hb92c903e),
	.w7(32'hb96b45c0),
	.w8(32'hb9d7b4f3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac828a9),
	.w1(32'hba34eb5e),
	.w2(32'hba17b21e),
	.w3(32'h3985b9d4),
	.w4(32'hba12ed31),
	.w5(32'h3a01c454),
	.w6(32'h3af48af7),
	.w7(32'h3a56f2cd),
	.w8(32'hb9927485),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0f25),
	.w1(32'hbaec1526),
	.w2(32'hbab9feeb),
	.w3(32'h398f2458),
	.w4(32'hbb3f4ed4),
	.w5(32'hbabee0d1),
	.w6(32'h3a3914e8),
	.w7(32'hba399416),
	.w8(32'hba7132f9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82ada21),
	.w1(32'hbacab232),
	.w2(32'hbaee105e),
	.w3(32'hb98f865b),
	.w4(32'hb8df6e74),
	.w5(32'h38018707),
	.w6(32'hb9ee76da),
	.w7(32'hba06f43a),
	.w8(32'hb9965102),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc688fb0),
	.w1(32'hbbe95089),
	.w2(32'h3b039493),
	.w3(32'h3abcb8bf),
	.w4(32'hbbd92b8b),
	.w5(32'hbc0eb94f),
	.w6(32'hbb5c5c40),
	.w7(32'hb9999d93),
	.w8(32'hba7ff41c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18704c),
	.w1(32'h3958e9ec),
	.w2(32'hba358156),
	.w3(32'hba8a65e4),
	.w4(32'hbaeb3ee5),
	.w5(32'hbb1c3196),
	.w6(32'hb65e10c9),
	.w7(32'hba22b41d),
	.w8(32'hba3591a8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7152fb),
	.w1(32'hbc0563e1),
	.w2(32'h3bc7cedb),
	.w3(32'h3b1366e6),
	.w4(32'h3badc7fe),
	.w5(32'hbbe1f698),
	.w6(32'hbc16aabf),
	.w7(32'h3b2c23d7),
	.w8(32'h3c3de9fb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd15c6),
	.w1(32'hbcb95a06),
	.w2(32'hbc344a38),
	.w3(32'hbc82537b),
	.w4(32'hbcb37f02),
	.w5(32'hbc63085b),
	.w6(32'hbc24983d),
	.w7(32'hbc158be0),
	.w8(32'hbc7a3b6b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7fd0),
	.w1(32'hba9143d8),
	.w2(32'h39a69638),
	.w3(32'hbad0de56),
	.w4(32'hbb8251e1),
	.w5(32'h3a727e01),
	.w6(32'h3bcc17b2),
	.w7(32'hb9ac1712),
	.w8(32'hbac5d46f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7c0b6),
	.w1(32'hbbc6a90d),
	.w2(32'hba21b9ea),
	.w3(32'h3b5829b6),
	.w4(32'h38b1fc10),
	.w5(32'hbbd88b86),
	.w6(32'hbbe98fad),
	.w7(32'hbb024b68),
	.w8(32'h3b557263),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb702d30),
	.w1(32'hb7c9e32e),
	.w2(32'h3aa52a17),
	.w3(32'h3b8bac4d),
	.w4(32'h3b15f3f5),
	.w5(32'h3b3d6238),
	.w6(32'h3b02208c),
	.w7(32'h3b7274b7),
	.w8(32'h3aaf1d31),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac992d5),
	.w1(32'hba137fee),
	.w2(32'hb9d2a378),
	.w3(32'h3a7eb540),
	.w4(32'h3a004213),
	.w5(32'h3a0919ef),
	.w6(32'hb9e52fdc),
	.w7(32'hb9e8831c),
	.w8(32'hb8fac31b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb872ec),
	.w1(32'h3c86cf0e),
	.w2(32'hbcbaebb1),
	.w3(32'hbcc7adef),
	.w4(32'h3c9149bb),
	.w5(32'h3d589d17),
	.w6(32'h3c5cd15a),
	.w7(32'hbbb4732c),
	.w8(32'h3cdcaf2d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b9911),
	.w1(32'hbac5175e),
	.w2(32'hbb92231a),
	.w3(32'h3a6361d2),
	.w4(32'hba7704be),
	.w5(32'hbb1ee615),
	.w6(32'hbab3ae7d),
	.w7(32'hbb98e593),
	.w8(32'hbbcf8e8a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ff36),
	.w1(32'hbbe07222),
	.w2(32'hbbc9860e),
	.w3(32'hbc2ee7a5),
	.w4(32'hbc13d13f),
	.w5(32'hbc052624),
	.w6(32'hbc08e0e4),
	.w7(32'hbc031f0a),
	.w8(32'hbbdc43b0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ea210),
	.w1(32'hb96f3ba3),
	.w2(32'hbaa38cd3),
	.w3(32'hbadeb4da),
	.w4(32'hbafc0e88),
	.w5(32'hbb5009e5),
	.w6(32'hba6abe21),
	.w7(32'h39d76d25),
	.w8(32'hbab23cac),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47d0bd),
	.w1(32'h3a5bb785),
	.w2(32'hbb6fba21),
	.w3(32'hbb2ed624),
	.w4(32'hbb035213),
	.w5(32'hba00577e),
	.w6(32'hba0a848d),
	.w7(32'hbb12c0f8),
	.w8(32'hbacd20e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946590),
	.w1(32'h3998c5a0),
	.w2(32'hb9821688),
	.w3(32'hbb3163f9),
	.w4(32'hbb503c5f),
	.w5(32'hbb5a8f55),
	.w6(32'hba912d7f),
	.w7(32'hbad58808),
	.w8(32'hbadf444b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97d669),
	.w1(32'h3b2f55d1),
	.w2(32'hba17ec78),
	.w3(32'hbb66704f),
	.w4(32'hbb4ab561),
	.w5(32'h3c169b40),
	.w6(32'h3ad5aca6),
	.w7(32'hbbe5c1ea),
	.w8(32'hb718b01e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89275e),
	.w1(32'hb98eb6a0),
	.w2(32'h37dff6a1),
	.w3(32'hba76524d),
	.w4(32'hba697e64),
	.w5(32'hba8195ad),
	.w6(32'hb99d9904),
	.w7(32'hba84308f),
	.w8(32'hba618678),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a1a40),
	.w1(32'hbabbfe35),
	.w2(32'hbba13830),
	.w3(32'hbbf4d1ed),
	.w4(32'hbbde1bd9),
	.w5(32'h3aeb256d),
	.w6(32'h3888070b),
	.w7(32'hbbe9a2b1),
	.w8(32'hbbada9c1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bc9ab),
	.w1(32'h3a89079b),
	.w2(32'h3ad73271),
	.w3(32'h3af4f086),
	.w4(32'h3b38bcf0),
	.w5(32'h398ea638),
	.w6(32'h3ad4f541),
	.w7(32'h39dcfa59),
	.w8(32'h3a2afe4c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99ff5e),
	.w1(32'hbc16427f),
	.w2(32'h3c1e4c80),
	.w3(32'h3c5a44f4),
	.w4(32'hbb15c277),
	.w5(32'hbc333c96),
	.w6(32'hbc600b46),
	.w7(32'h39896272),
	.w8(32'h3b21d9fb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae070af),
	.w1(32'hbb9a1e08),
	.w2(32'hbbc817d9),
	.w3(32'h3a373a40),
	.w4(32'hbb69175f),
	.w5(32'hbbaeb86a),
	.w6(32'h3bce3509),
	.w7(32'h3a06361c),
	.w8(32'hbb9cb023),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d855e),
	.w1(32'hbb4264ad),
	.w2(32'hbb648151),
	.w3(32'hbbe7292a),
	.w4(32'hbb75e3f3),
	.w5(32'h3b10edc0),
	.w6(32'hbb2d48fb),
	.w7(32'hbbf66817),
	.w8(32'hbb5740e2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ff99a),
	.w1(32'h3af9eb26),
	.w2(32'h3ac923cc),
	.w3(32'h39fbebd6),
	.w4(32'hba0134d2),
	.w5(32'hb943c0bc),
	.w6(32'h3abfe894),
	.w7(32'h3a9506a4),
	.w8(32'h3a6b7270),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce986c3),
	.w1(32'h3be17ef9),
	.w2(32'hbcfa0c1a),
	.w3(32'hbcd40859),
	.w4(32'hbc773b36),
	.w5(32'h3d03f25e),
	.w6(32'h3cedbbe7),
	.w7(32'hbc7d8210),
	.w8(32'h38a5c5b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5292d8),
	.w1(32'hbbf944f9),
	.w2(32'h3bcbf56f),
	.w3(32'h3c1b2a71),
	.w4(32'h3aac07d2),
	.w5(32'hbb8fac51),
	.w6(32'h3adba84e),
	.w7(32'h3bcfa8be),
	.w8(32'h3bd3854e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a252faf),
	.w1(32'hb9e9e4cf),
	.w2(32'h3ab0130a),
	.w3(32'h3b2909fc),
	.w4(32'h3a0b3521),
	.w5(32'hbb253d54),
	.w6(32'h3b6e5d4c),
	.w7(32'h3ad2af61),
	.w8(32'hb9b86c3c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f5e62),
	.w1(32'hbb11684e),
	.w2(32'hbb0bd790),
	.w3(32'h3a2b88b8),
	.w4(32'h39f61891),
	.w5(32'h3baefe22),
	.w6(32'h3a9ac4b8),
	.w7(32'h3aa0561a),
	.w8(32'h3b8b7a3f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc314959),
	.w1(32'hbc417276),
	.w2(32'hbc4adaac),
	.w3(32'hbc9be597),
	.w4(32'hbc92ac08),
	.w5(32'hbbf24273),
	.w6(32'hbc3fa93b),
	.w7(32'hbc9dba23),
	.w8(32'hbbd91c61),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bfc22),
	.w1(32'h3af74d5f),
	.w2(32'h3a7e9a3d),
	.w3(32'h3a1d2010),
	.w4(32'h3a1ec05c),
	.w5(32'hba51e3c2),
	.w6(32'hb92a402e),
	.w7(32'h38095994),
	.w8(32'hb9a81476),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a1e4),
	.w1(32'h3b979015),
	.w2(32'h3b3665c1),
	.w3(32'h3bf8527f),
	.w4(32'h3b881768),
	.w5(32'h3ad61a45),
	.w6(32'h3baefcf4),
	.w7(32'h3b25c4e8),
	.w8(32'h3b66a03f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967f38),
	.w1(32'hbb8e1750),
	.w2(32'hbb90dafa),
	.w3(32'hbafb4255),
	.w4(32'hbb3d91c7),
	.w5(32'hbacd5d29),
	.w6(32'h3893693c),
	.w7(32'hba466daa),
	.w8(32'hba7c1030),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9420f),
	.w1(32'hbb487b32),
	.w2(32'hbb99e4e6),
	.w3(32'h3abd58a5),
	.w4(32'hbb833ed1),
	.w5(32'hbb98d090),
	.w6(32'h3be3ce8e),
	.w7(32'hba1fca40),
	.w8(32'hbbdb5394),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d2c4b),
	.w1(32'hbbf67115),
	.w2(32'h3c0a2e47),
	.w3(32'h3c572eb1),
	.w4(32'h3bb7597b),
	.w5(32'h3b298e13),
	.w6(32'h3bb423c3),
	.w7(32'h3c5ab616),
	.w8(32'h3c4a859f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4a0d),
	.w1(32'h3b57cc79),
	.w2(32'h3b00e1f8),
	.w3(32'h3bcbb369),
	.w4(32'h3c002dbe),
	.w5(32'h3c0e05ff),
	.w6(32'h3bbb1131),
	.w7(32'h3bdcaad1),
	.w8(32'h3c06134e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b664429),
	.w1(32'h3ad07401),
	.w2(32'h39be27ed),
	.w3(32'h3b402359),
	.w4(32'h3b545795),
	.w5(32'h3b525fe1),
	.w6(32'h3b5120f9),
	.w7(32'h3b381e21),
	.w8(32'h3b936391),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1dfe),
	.w1(32'hbb24a943),
	.w2(32'hb99aab69),
	.w3(32'hbc6c5483),
	.w4(32'hbc062713),
	.w5(32'hbc1c5ba4),
	.w6(32'hbbf23f45),
	.w7(32'hbca7441a),
	.w8(32'hbc87f8f8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b039cd3),
	.w1(32'h3be7cec4),
	.w2(32'h3c8ecdad),
	.w3(32'h3cac345e),
	.w4(32'h3d0574a4),
	.w5(32'h3cd29e6d),
	.w6(32'h3cb101f8),
	.w7(32'h3d0d5044),
	.w8(32'h3cdbc3d8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a7e2c),
	.w1(32'hbb71d5ea),
	.w2(32'h3b9e80ba),
	.w3(32'hbc08c4d1),
	.w4(32'hba79c472),
	.w5(32'hb91c7d8d),
	.w6(32'hbc07247e),
	.w7(32'h3ba21771),
	.w8(32'hbb8776cd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe85c7),
	.w1(32'hbb78b59c),
	.w2(32'hbc20b2a8),
	.w3(32'hbbac6c78),
	.w4(32'hbc20cc32),
	.w5(32'hbc149675),
	.w6(32'hbbe5a3bc),
	.w7(32'hbc567e99),
	.w8(32'hbc2b5fba),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83530f),
	.w1(32'hbc09d265),
	.w2(32'h3b65b9e5),
	.w3(32'h3d1e7b52),
	.w4(32'h3c78542a),
	.w5(32'hbbd56cdc),
	.w6(32'h3c847e93),
	.w7(32'h3ca2b566),
	.w8(32'h3bfde0c9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9299d92),
	.w1(32'hbb81794f),
	.w2(32'hbb82ed82),
	.w3(32'hba52b005),
	.w4(32'hbbb3a983),
	.w5(32'hbbb9455e),
	.w6(32'hbbc6d9da),
	.w7(32'hbc198637),
	.w8(32'hbc21c8fd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8573),
	.w1(32'hbc1d4e81),
	.w2(32'hbb9690e7),
	.w3(32'hbc7c09a5),
	.w4(32'hbc97f644),
	.w5(32'hbb83fd59),
	.w6(32'hbadd0e8c),
	.w7(32'hbb8f59ad),
	.w8(32'hbaabcb64),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2853d4),
	.w1(32'h3c58cc11),
	.w2(32'hbd1cea63),
	.w3(32'h3c89b800),
	.w4(32'h3d03cdda),
	.w5(32'h3cf34d3f),
	.w6(32'hbc9dbdb3),
	.w7(32'hbce2d220),
	.w8(32'h3bd1ef88),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cde83),
	.w1(32'hbb47a5a0),
	.w2(32'hbd1312bf),
	.w3(32'hbd0c7d3d),
	.w4(32'hbd845cc7),
	.w5(32'hbd6eb6cb),
	.w6(32'hbd167847),
	.w7(32'hbd9a73a8),
	.w8(32'hbd8e77af),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule