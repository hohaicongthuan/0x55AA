module layer_10_featuremap_274(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaaba9),
	.w1(32'hbb696010),
	.w2(32'hbc2b1d8b),
	.w3(32'hbbe3ab12),
	.w4(32'hbc1eff02),
	.w5(32'h3be1a1a3),
	.w6(32'hbbbf22b7),
	.w7(32'hbc25990c),
	.w8(32'h3bda3fe8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21ec82),
	.w1(32'h3a3e209e),
	.w2(32'hbae5998c),
	.w3(32'h3bf1cf4f),
	.w4(32'h3b2938d1),
	.w5(32'hbc0d6c81),
	.w6(32'h3ae9f98b),
	.w7(32'h39fff41a),
	.w8(32'hbabf2109),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223c50),
	.w1(32'h3a25ad20),
	.w2(32'h3aca9e39),
	.w3(32'h3b4cc999),
	.w4(32'h3a6c10c3),
	.w5(32'hb8d618dd),
	.w6(32'h3bb898ac),
	.w7(32'h39f610ec),
	.w8(32'hbbb25f5e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23eb1d),
	.w1(32'h3a5dc7ec),
	.w2(32'h3bbbbf28),
	.w3(32'h3b57a7b2),
	.w4(32'h3bda7be2),
	.w5(32'h3b59916a),
	.w6(32'hba588ae5),
	.w7(32'h3c0a1f33),
	.w8(32'h3bd09892),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecde91),
	.w1(32'h3a103680),
	.w2(32'h394751c1),
	.w3(32'hba6ea080),
	.w4(32'h3a852155),
	.w5(32'hbb9c0d06),
	.w6(32'hbb44072d),
	.w7(32'hba721950),
	.w8(32'hbbfc3b47),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb601f6),
	.w1(32'h3a2dd52e),
	.w2(32'h3aef56d6),
	.w3(32'h39c4f995),
	.w4(32'h3b49bb8e),
	.w5(32'hbbb58e25),
	.w6(32'h3ab559ec),
	.w7(32'h3be29ce5),
	.w8(32'hbc20a316),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49245f),
	.w1(32'hbb6336ba),
	.w2(32'h3b8b4c35),
	.w3(32'hbacb83ae),
	.w4(32'h3b96f30b),
	.w5(32'hbab46ce5),
	.w6(32'h3ad87705),
	.w7(32'h3bfeaa72),
	.w8(32'hbbd7a4ee),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906bd3),
	.w1(32'h3b40b977),
	.w2(32'hb8132977),
	.w3(32'hba9feef1),
	.w4(32'h3abfa8b3),
	.w5(32'h3b46c7e2),
	.w6(32'h3a0927be),
	.w7(32'h3abf60bd),
	.w8(32'hb913c356),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07a848),
	.w1(32'h3a06ed0a),
	.w2(32'hbaede040),
	.w3(32'hba0d6fe8),
	.w4(32'hbb934bf4),
	.w5(32'hbb5da262),
	.w6(32'h3934ae68),
	.w7(32'hbb0a1446),
	.w8(32'hbc0f3dc6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcec2ec),
	.w1(32'h3a4654e1),
	.w2(32'h3b58f813),
	.w3(32'h3ab25b8a),
	.w4(32'h3b9a4f80),
	.w5(32'hbb32f11c),
	.w6(32'hba3afc5f),
	.w7(32'h3bfdb8b4),
	.w8(32'hbbebf203),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048960),
	.w1(32'h3a1a2857),
	.w2(32'h3b0c534f),
	.w3(32'h3b28e3e4),
	.w4(32'h3b6db5e3),
	.w5(32'hbbed6c8d),
	.w6(32'hba791753),
	.w7(32'h3b542158),
	.w8(32'hbb401fb4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60dfe1),
	.w1(32'hbb580450),
	.w2(32'h3b1aef42),
	.w3(32'h3907a37b),
	.w4(32'h3b27720f),
	.w5(32'h3b1101f2),
	.w6(32'h3bc0bee8),
	.w7(32'h3b4dc9d7),
	.w8(32'h3b2874bc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af295cc),
	.w1(32'hbb152fe9),
	.w2(32'hbbbcb4a3),
	.w3(32'hbb9b4caa),
	.w4(32'hbbfdf054),
	.w5(32'h3b51501a),
	.w6(32'hbb880f4f),
	.w7(32'hbc182bd3),
	.w8(32'h3ba78ee6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42cbc7),
	.w1(32'hb83a070e),
	.w2(32'h3b3941de),
	.w3(32'hba5a7bca),
	.w4(32'h3ae5fb75),
	.w5(32'hbb9135c1),
	.w6(32'hb999e705),
	.w7(32'h3b08fb7d),
	.w8(32'hbbbbc10e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54df5f),
	.w1(32'h3bbbc1d5),
	.w2(32'h3b6081a3),
	.w3(32'hbb5b38d9),
	.w4(32'hbb5877d9),
	.w5(32'h3a03bc2f),
	.w6(32'h3b129df5),
	.w7(32'h3b4b7303),
	.w8(32'hb865ca54),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03ef96),
	.w1(32'hbb3f34f9),
	.w2(32'h3908f2dc),
	.w3(32'hb9b7efd5),
	.w4(32'h3958ff59),
	.w5(32'hbb29df6b),
	.w6(32'hbbcaa8ba),
	.w7(32'hbaa877ff),
	.w8(32'hbb14e5eb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e885),
	.w1(32'h3add4675),
	.w2(32'h3b8ad8d4),
	.w3(32'h3bfb12b9),
	.w4(32'h3c03a896),
	.w5(32'hbb08139d),
	.w6(32'h3c2ed36e),
	.w7(32'h3c34d320),
	.w8(32'hbb442b6d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1deb),
	.w1(32'h399d45ce),
	.w2(32'h39bfa96e),
	.w3(32'hbb2fdcc8),
	.w4(32'hba1f395c),
	.w5(32'h396d2b36),
	.w6(32'h3a8195c1),
	.w7(32'hbae4266a),
	.w8(32'h3bd52786),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f97d),
	.w1(32'h3bd6f483),
	.w2(32'h3bb10dec),
	.w3(32'h3b248fee),
	.w4(32'h3ab94877),
	.w5(32'h3b93b6e0),
	.w6(32'h3b89875f),
	.w7(32'h3bb42c10),
	.w8(32'h3b069b54),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2929),
	.w1(32'hb9366092),
	.w2(32'hbae3ab0d),
	.w3(32'hb9216c8f),
	.w4(32'h3b966a73),
	.w5(32'h3abea690),
	.w6(32'h39ac8098),
	.w7(32'h3b006b38),
	.w8(32'h3b95cd4f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedca45),
	.w1(32'h39d9ea31),
	.w2(32'hbb87ac33),
	.w3(32'hb9ae3145),
	.w4(32'hbaadfdbf),
	.w5(32'hbb3f5dfd),
	.w6(32'hbb0ac427),
	.w7(32'hbb19570d),
	.w8(32'hbb7b806a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd84a5),
	.w1(32'h3bb09dd7),
	.w2(32'h3c3394c2),
	.w3(32'h3ba7e355),
	.w4(32'h3c1cf130),
	.w5(32'h393db97f),
	.w6(32'h3c0ff785),
	.w7(32'h3c4bcdd3),
	.w8(32'hba1246c7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f6f8),
	.w1(32'hbb020452),
	.w2(32'hbb5744a7),
	.w3(32'h3b6b1c79),
	.w4(32'h3a7df118),
	.w5(32'hb97081dc),
	.w6(32'h3b9dc830),
	.w7(32'hba3827d7),
	.w8(32'hba57f51d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6716f),
	.w1(32'h3a292a64),
	.w2(32'h3a27fd8e),
	.w3(32'hbbd84f5c),
	.w4(32'hbab155ab),
	.w5(32'hba5c5d5a),
	.w6(32'hbc00d2e1),
	.w7(32'hbb0d0439),
	.w8(32'h3b915c25),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0085),
	.w1(32'h39df34d8),
	.w2(32'h39013b0e),
	.w3(32'h3a95fc39),
	.w4(32'hbad80a45),
	.w5(32'hbba398e4),
	.w6(32'h39cc39b3),
	.w7(32'h3af0308e),
	.w8(32'hbbb1e078),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad5fc),
	.w1(32'h3c05c31e),
	.w2(32'h3c20cdcb),
	.w3(32'h3b7d2a30),
	.w4(32'h3be9dd15),
	.w5(32'hbbb4f35a),
	.w6(32'h3c0c38b6),
	.w7(32'h3c4692d4),
	.w8(32'hbc22c272),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62848),
	.w1(32'hba2dfc11),
	.w2(32'h3b09f222),
	.w3(32'h3b8720d8),
	.w4(32'h3bf63823),
	.w5(32'h39a7b340),
	.w6(32'h3b063c04),
	.w7(32'h3c024923),
	.w8(32'h3a67c68b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a95259),
	.w1(32'h3b42a255),
	.w2(32'hbbd2e484),
	.w3(32'hbb25c870),
	.w4(32'hbc19b401),
	.w5(32'hba8573f3),
	.w6(32'h3b388269),
	.w7(32'hbb9b5f33),
	.w8(32'hba4153b8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d5e0a),
	.w1(32'h3a162ef8),
	.w2(32'h3b85c39f),
	.w3(32'hbaeab96c),
	.w4(32'hbb118fc0),
	.w5(32'h3a089ac2),
	.w6(32'hbaa5e2cf),
	.w7(32'h3b431535),
	.w8(32'h3b073a07),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3657f0ac),
	.w1(32'hbb1461b5),
	.w2(32'hbb9a4853),
	.w3(32'hbb6a93ab),
	.w4(32'hbb3fe744),
	.w5(32'hbbe27534),
	.w6(32'hbb489dd4),
	.w7(32'hbbde8805),
	.w8(32'hbaa7200e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5137),
	.w1(32'h3c0679aa),
	.w2(32'h3c236f88),
	.w3(32'hbc0a9a26),
	.w4(32'hbb015ba2),
	.w5(32'hbaa51b67),
	.w6(32'hbb667ad5),
	.w7(32'h3c14aa8f),
	.w8(32'h3b88bb5e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbafd10),
	.w1(32'hbbeb6c06),
	.w2(32'hb9fd843e),
	.w3(32'h3b8c662c),
	.w4(32'h3bed7f1d),
	.w5(32'hbb4f9b46),
	.w6(32'h3b768a4f),
	.w7(32'h3b9e8307),
	.w8(32'h38fe40fe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb48fd),
	.w1(32'hbb60c987),
	.w2(32'h3bc41d90),
	.w3(32'hbb9a5db5),
	.w4(32'hbb8c7d29),
	.w5(32'hbc06cb5d),
	.w6(32'hbb916ecd),
	.w7(32'h3b99848a),
	.w8(32'hbc1ad4bb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd8476),
	.w1(32'hbb875a85),
	.w2(32'hba9e1a9b),
	.w3(32'hbb993cdc),
	.w4(32'hbaa88445),
	.w5(32'h3a861be9),
	.w6(32'hbba3202f),
	.w7(32'hba53c0c2),
	.w8(32'hbb2db10f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cb736),
	.w1(32'h3b816f97),
	.w2(32'h3b52a673),
	.w3(32'h3b0b97f9),
	.w4(32'hba6d0f74),
	.w5(32'h3af86db7),
	.w6(32'h3bafb6cb),
	.w7(32'h3b22776d),
	.w8(32'h39baa905),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7af41),
	.w1(32'h3adb6095),
	.w2(32'hba8b1bc1),
	.w3(32'hb9377afa),
	.w4(32'hbb1a5bce),
	.w5(32'hbb48a1ed),
	.w6(32'h3ad02018),
	.w7(32'h3a5086ea),
	.w8(32'hba903e5c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70ad5),
	.w1(32'h3b78842f),
	.w2(32'h3bfe4b4e),
	.w3(32'hbb4c654e),
	.w4(32'h3b8d25e0),
	.w5(32'hbb371c2f),
	.w6(32'hbb33b742),
	.w7(32'h3ba496d7),
	.w8(32'hbabe4bc7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d394d),
	.w1(32'hbb337d0a),
	.w2(32'hba664993),
	.w3(32'h3ae2836b),
	.w4(32'h3b89a3b1),
	.w5(32'h3bcca2f8),
	.w6(32'hbabe9d6d),
	.w7(32'h3bc9c2dc),
	.w8(32'h3b93f05c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f16a),
	.w1(32'hbb157ebd),
	.w2(32'hbb002f90),
	.w3(32'hba2b6933),
	.w4(32'hbb97494f),
	.w5(32'h3b094e6c),
	.w6(32'hbbb856fa),
	.w7(32'hbbe4dcb3),
	.w8(32'hbac78f45),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489281),
	.w1(32'h3aef1571),
	.w2(32'h3c30d14c),
	.w3(32'h3b2b7aa8),
	.w4(32'h3c476191),
	.w5(32'h3bcb335d),
	.w6(32'h390046d1),
	.w7(32'h3c25b6de),
	.w8(32'h3bbf822a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1274be),
	.w1(32'h3b15288f),
	.w2(32'h3a1befa5),
	.w3(32'hbab4290f),
	.w4(32'hbb45469b),
	.w5(32'hbc2ea4dc),
	.w6(32'h3b801e1e),
	.w7(32'hbabcde2b),
	.w8(32'hbc8c2e73),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f088d),
	.w1(32'h3bafcceb),
	.w2(32'h3c6a15cb),
	.w3(32'h3c0be0c5),
	.w4(32'h3c773e44),
	.w5(32'h3c088481),
	.w6(32'h3c40d565),
	.w7(32'h3c9f796b),
	.w8(32'h3c238fab),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf51922),
	.w1(32'h3b7e9bec),
	.w2(32'h3b24471d),
	.w3(32'h3b884405),
	.w4(32'hb9d96d01),
	.w5(32'hbc2d86b4),
	.w6(32'hbaa8bfd1),
	.w7(32'hbbbf8d2f),
	.w8(32'hbc445466),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5f2e),
	.w1(32'h3b5e9877),
	.w2(32'h3bb1d594),
	.w3(32'h3b80db3d),
	.w4(32'h387dda21),
	.w5(32'hbc1b2657),
	.w6(32'h3a2e94f1),
	.w7(32'h3bf0788e),
	.w8(32'hbc65819d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d2051),
	.w1(32'hbaf88045),
	.w2(32'h3ba6aafa),
	.w3(32'hbb9f2389),
	.w4(32'h3a17d503),
	.w5(32'hbb933260),
	.w6(32'hbb312b21),
	.w7(32'h3b9d0a25),
	.w8(32'h3b7c0b78),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7ed1),
	.w1(32'h3c866258),
	.w2(32'h3c07404f),
	.w3(32'h3c0c47f6),
	.w4(32'h3c135351),
	.w5(32'hbc066135),
	.w6(32'h3c894f60),
	.w7(32'h3c714f9e),
	.w8(32'hbc2142ba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc164752),
	.w1(32'h3aaa8bb9),
	.w2(32'h3b87bb20),
	.w3(32'h3abe33cd),
	.w4(32'h3b6f784b),
	.w5(32'h3c085914),
	.w6(32'h3a1b6f1f),
	.w7(32'h3b9a5213),
	.w8(32'h3c23f9fe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c262fb9),
	.w1(32'h3ba932ca),
	.w2(32'h3b84aad8),
	.w3(32'h3bd0ab4f),
	.w4(32'h39762b9b),
	.w5(32'hbad031d2),
	.w6(32'h3c148cce),
	.w7(32'h3ab7b616),
	.w8(32'hb90ece8a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d55a5d),
	.w1(32'hbb1113bd),
	.w2(32'hbb71f6c6),
	.w3(32'hbb97f7d4),
	.w4(32'hbc03498e),
	.w5(32'hbbd9093b),
	.w6(32'hbb6f1203),
	.w7(32'hbbda0321),
	.w8(32'hbc0a3400),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe14b91),
	.w1(32'h3a25a906),
	.w2(32'h3c294b0e),
	.w3(32'h3b063265),
	.w4(32'h3c0d4996),
	.w5(32'h3b9fed73),
	.w6(32'h3c0ce0bf),
	.w7(32'h3c4120f6),
	.w8(32'h3b46d465),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951fe5),
	.w1(32'hbb1bd4ac),
	.w2(32'h3a8afadd),
	.w3(32'hbb70e610),
	.w4(32'hbb3550c3),
	.w5(32'h3b8b8540),
	.w6(32'hbb3b055b),
	.w7(32'hbb204030),
	.w8(32'h3b063014),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2138e),
	.w1(32'hbab19b80),
	.w2(32'h39fd9410),
	.w3(32'h3c0b40f4),
	.w4(32'h3b8a77b4),
	.w5(32'hba488574),
	.w6(32'h3aada663),
	.w7(32'h3b32329f),
	.w8(32'hbbad065b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ebad8),
	.w1(32'h39864ea2),
	.w2(32'hba8216cc),
	.w3(32'hbb056f3b),
	.w4(32'hbb80d80a),
	.w5(32'h394ff72c),
	.w6(32'hbacb2eea),
	.w7(32'hbba97e5b),
	.w8(32'hbb9094a4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdb70c),
	.w1(32'hb9803b3d),
	.w2(32'h3bd321c3),
	.w3(32'hbb3c8cc7),
	.w4(32'h3ab732dc),
	.w5(32'h3b5930c5),
	.w6(32'h3ae2dc23),
	.w7(32'hba4bcd27),
	.w8(32'h39903f3e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb316fd2),
	.w1(32'hbb2c24ba),
	.w2(32'hbb56bc85),
	.w3(32'hba89a1ef),
	.w4(32'h3b6190b8),
	.w5(32'hb7f5016a),
	.w6(32'hbb230912),
	.w7(32'h3a7c71e5),
	.w8(32'h3a9abf11),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94445b),
	.w1(32'hbba774f6),
	.w2(32'hba26554c),
	.w3(32'h3a1a3c0c),
	.w4(32'hbb582e23),
	.w5(32'h3bc7c472),
	.w6(32'h3ab6e721),
	.w7(32'h3b5f51b0),
	.w8(32'h3ba150d6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67a507),
	.w1(32'h3aebb186),
	.w2(32'hbb2f9f23),
	.w3(32'hbaab0cb1),
	.w4(32'hbbebaed1),
	.w5(32'h3a3a89ca),
	.w6(32'h3b2cd9d9),
	.w7(32'hbb7c136e),
	.w8(32'hbb8949bd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87abfe0),
	.w1(32'hbc4e6248),
	.w2(32'h3b09296a),
	.w3(32'hbc537d73),
	.w4(32'hb9cbd0fc),
	.w5(32'hbbf6b7a1),
	.w6(32'hbc9c03fb),
	.w7(32'hbaff6786),
	.w8(32'hbc49050e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27e6cd),
	.w1(32'hb9eb98a5),
	.w2(32'h3c01fcb9),
	.w3(32'h3a43d1ec),
	.w4(32'h3be7310e),
	.w5(32'hbc51cb98),
	.w6(32'h3bbaf69a),
	.w7(32'h3c12291c),
	.w8(32'hbb9c9262),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e00e),
	.w1(32'hbbc869f2),
	.w2(32'h3b600f86),
	.w3(32'h3aabd029),
	.w4(32'h3b8b65b2),
	.w5(32'hbab124e6),
	.w6(32'hbb787f9d),
	.w7(32'h3bea3199),
	.w8(32'h39cf8fb1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca161),
	.w1(32'h3ad617c9),
	.w2(32'hba070fd8),
	.w3(32'hbb8e7eac),
	.w4(32'hbbeb9454),
	.w5(32'hbb9297cb),
	.w6(32'hba47dd40),
	.w7(32'hbbbfcf54),
	.w8(32'hbc0eb1bc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ceb2),
	.w1(32'h3b1d938f),
	.w2(32'h3be14680),
	.w3(32'h3b71785a),
	.w4(32'h3ae1dd58),
	.w5(32'h3a81d3f9),
	.w6(32'h3c04b5e5),
	.w7(32'h3c2d2a72),
	.w8(32'h3aaf4645),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c45f),
	.w1(32'hba4dc365),
	.w2(32'hb9cff778),
	.w3(32'h380334ce),
	.w4(32'h3a86bfbc),
	.w5(32'h3b839f72),
	.w6(32'hba0a3873),
	.w7(32'hba7d6124),
	.w8(32'h3b56f0c3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42da03),
	.w1(32'h3a62bb50),
	.w2(32'hbb60561f),
	.w3(32'h39eed567),
	.w4(32'hbbbb880f),
	.w5(32'h3b2a1365),
	.w6(32'h3b2eb47b),
	.w7(32'hbb949e07),
	.w8(32'h3aa56f07),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a5e02),
	.w1(32'h3ab34277),
	.w2(32'hbae4962e),
	.w3(32'hbb0f7e89),
	.w4(32'hbbb250e0),
	.w5(32'hbab2c148),
	.w6(32'hb89c7062),
	.w7(32'hbb5d86e9),
	.w8(32'hba37bfa5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc05fb),
	.w1(32'hbba0068f),
	.w2(32'hba8c668c),
	.w3(32'h3af2568a),
	.w4(32'h3bc75ca5),
	.w5(32'h3a25099a),
	.w6(32'hbb054c6b),
	.w7(32'h3ac67e69),
	.w8(32'h3a5444ea),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f3e26),
	.w1(32'h3c3b4e26),
	.w2(32'hba766b4a),
	.w3(32'h3b3e78b6),
	.w4(32'h3ab873ae),
	.w5(32'h3b735773),
	.w6(32'h3c1efd9a),
	.w7(32'h3ade37dc),
	.w8(32'h3c18a30e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb83f7),
	.w1(32'h3af107f2),
	.w2(32'h3b277f99),
	.w3(32'hb999674b),
	.w4(32'hbb36bc69),
	.w5(32'h3b867057),
	.w6(32'hbb591162),
	.w7(32'hbb09d3ca),
	.w8(32'hb9c950c4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27da69),
	.w1(32'hbb24f7ba),
	.w2(32'hb8bd929c),
	.w3(32'hbbb75dd6),
	.w4(32'h3a73269e),
	.w5(32'hbbf96651),
	.w6(32'hbbc4641c),
	.w7(32'hb9d7b36b),
	.w8(32'hbc29ad45),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8070c),
	.w1(32'h3a122948),
	.w2(32'h3b9488a6),
	.w3(32'h3a8e47d9),
	.w4(32'h3b74fb49),
	.w5(32'hba154ec4),
	.w6(32'h3b8afe19),
	.w7(32'h3c044811),
	.w8(32'hba557c15),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45124),
	.w1(32'h3b92a41f),
	.w2(32'h3bba336b),
	.w3(32'h3b14365c),
	.w4(32'h3b9b46c1),
	.w5(32'h3c35547b),
	.w6(32'h3a936b52),
	.w7(32'h3c022555),
	.w8(32'h3c295925),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93fa4a),
	.w1(32'h3ad59b37),
	.w2(32'hbadef037),
	.w3(32'hbab13481),
	.w4(32'hbb67769d),
	.w5(32'h3c00a913),
	.w6(32'hbb949310),
	.w7(32'hbb18d2f5),
	.w8(32'h3bb41705),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853147),
	.w1(32'hbbffe57e),
	.w2(32'hbc00f3f1),
	.w3(32'hb8d08301),
	.w4(32'hbc022457),
	.w5(32'h3aad4018),
	.w6(32'hbbb0b3b0),
	.w7(32'hbbe3bad8),
	.w8(32'hb9414dee),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078db5),
	.w1(32'hbb1240ac),
	.w2(32'hbabb48c8),
	.w3(32'h3a9ed6c5),
	.w4(32'hba081b68),
	.w5(32'hba2babc7),
	.w6(32'hba27d3bc),
	.w7(32'hba1e0131),
	.w8(32'hbb1ce372),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b23d6),
	.w1(32'h3b4b8834),
	.w2(32'hbb04ece7),
	.w3(32'h3b8d8d2a),
	.w4(32'h3ada4e42),
	.w5(32'h3b7e3ee4),
	.w6(32'h3b2d0d4e),
	.w7(32'h3a3b1f32),
	.w8(32'h3c1ca81e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075f58),
	.w1(32'h3ac261d2),
	.w2(32'hbbc4db1a),
	.w3(32'hbb935c36),
	.w4(32'hbc3f136c),
	.w5(32'hba62094f),
	.w6(32'hbaf64fae),
	.w7(32'hbc39b5a7),
	.w8(32'h3b28763b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ed5e),
	.w1(32'hba8d5a40),
	.w2(32'hbb3d3b51),
	.w3(32'h3a0320bd),
	.w4(32'hba662d96),
	.w5(32'hbb2471fa),
	.w6(32'h3abed82e),
	.w7(32'h398a2989),
	.w8(32'hbbd0b152),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2573),
	.w1(32'hbb8f572d),
	.w2(32'h3a1832ba),
	.w3(32'hbb92a941),
	.w4(32'hba8b8ae6),
	.w5(32'h3b675604),
	.w6(32'hbb4427c2),
	.w7(32'h3b327c23),
	.w8(32'h3be09e37),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ce436),
	.w1(32'h3b44bc0d),
	.w2(32'h3a800a48),
	.w3(32'hbaf501ed),
	.w4(32'hbae079bd),
	.w5(32'h3a861362),
	.w6(32'hbb2eaac5),
	.w7(32'hb713a4e9),
	.w8(32'h3ad30c96),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e6fc8),
	.w1(32'h3b9ae142),
	.w2(32'h38846791),
	.w3(32'h396ed2ae),
	.w4(32'hbb8df554),
	.w5(32'h3bb7abbf),
	.w6(32'h3bf367a1),
	.w7(32'h3b437fe2),
	.w8(32'h3b9a0a46),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55305c),
	.w1(32'h3bc10bc3),
	.w2(32'hba44209e),
	.w3(32'hbb047d62),
	.w4(32'hbab021e0),
	.w5(32'h380cc4fd),
	.w6(32'hbb66452b),
	.w7(32'hbbb1a2ce),
	.w8(32'h3ad2c5d2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53ec55),
	.w1(32'hbaad8315),
	.w2(32'hbace3910),
	.w3(32'hba6b163f),
	.w4(32'hbb1e6fdd),
	.w5(32'h3ac30967),
	.w6(32'h3ad9a5df),
	.w7(32'hbaa15874),
	.w8(32'h39c23679),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26242),
	.w1(32'hbba21fa1),
	.w2(32'hbb51963d),
	.w3(32'h3784facb),
	.w4(32'hba405b48),
	.w5(32'h3a752b30),
	.w6(32'hbad85ef9),
	.w7(32'hbb9c1e76),
	.w8(32'hb8905c79),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f70aa),
	.w1(32'hba943755),
	.w2(32'hbb1a77ba),
	.w3(32'h3b0c677a),
	.w4(32'h3bd10414),
	.w5(32'h3b04c6eb),
	.w6(32'hbbaa4335),
	.w7(32'hba2c7c7f),
	.w8(32'h3aeb8bd1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4314fb),
	.w1(32'hbb95ee43),
	.w2(32'hbb7fa1b1),
	.w3(32'h3b32050e),
	.w4(32'h3a4fc68e),
	.w5(32'hbba207d4),
	.w6(32'h3a97e78b),
	.w7(32'hbaa41ed9),
	.w8(32'hbbc8ae6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa5ac2),
	.w1(32'h3c15aa0f),
	.w2(32'h3c11fc43),
	.w3(32'h3baf0c07),
	.w4(32'h3aaa7420),
	.w5(32'hbbacaf43),
	.w6(32'h3bca935d),
	.w7(32'h3c14c6b5),
	.w8(32'hbc727517),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf89b6),
	.w1(32'hbb014fb5),
	.w2(32'h3c2614bc),
	.w3(32'hbb141c49),
	.w4(32'h3bec07ed),
	.w5(32'h3a814185),
	.w6(32'hba622b69),
	.w7(32'h3c1505c7),
	.w8(32'h3ae01bbb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f03a),
	.w1(32'hbb8bcf62),
	.w2(32'hbac8b22d),
	.w3(32'h3b27879a),
	.w4(32'h3b89b1af),
	.w5(32'hbbbe2497),
	.w6(32'hb9f76582),
	.w7(32'h3a6676db),
	.w8(32'hbbf121cc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf6f61),
	.w1(32'h38823219),
	.w2(32'h3b8d0783),
	.w3(32'h3a87a872),
	.w4(32'h3b6e7922),
	.w5(32'h3ba9cae7),
	.w6(32'h3bb139fa),
	.w7(32'h3bf98190),
	.w8(32'h3ba58364),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13c70e),
	.w1(32'h3adf7007),
	.w2(32'hba4d4527),
	.w3(32'hbb849136),
	.w4(32'hbaade064),
	.w5(32'h3b96878a),
	.w6(32'hbb506657),
	.w7(32'hbb11fcea),
	.w8(32'h3b41114f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b882d52),
	.w1(32'h3a89c983),
	.w2(32'h3ae7ca78),
	.w3(32'h3b6f9d5e),
	.w4(32'h381a9304),
	.w5(32'h37d5b86f),
	.w6(32'h3ba404df),
	.w7(32'h3af9dab2),
	.w8(32'hbaaa3f7d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e1d97),
	.w1(32'hbbe31370),
	.w2(32'h3ae75d42),
	.w3(32'hbb3b7518),
	.w4(32'h3ba41865),
	.w5(32'hbafec948),
	.w6(32'hbbefe557),
	.w7(32'hb8e4f82a),
	.w8(32'hbbbe28e8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeee9c7),
	.w1(32'hbae7b7ff),
	.w2(32'h3b94d5ff),
	.w3(32'h3b719812),
	.w4(32'h3b21f624),
	.w5(32'hbb9005e5),
	.w6(32'h3c07ee33),
	.w7(32'h3c3207ac),
	.w8(32'hbb753bc9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32f6a7),
	.w1(32'hb72261da),
	.w2(32'hbadae3ff),
	.w3(32'hbb018870),
	.w4(32'hbaa37d0f),
	.w5(32'h3a48f3c7),
	.w6(32'hbb49209d),
	.w7(32'h3a5878e1),
	.w8(32'hbaa5e969),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ecfae),
	.w1(32'hbb9e8c96),
	.w2(32'hbb9920c1),
	.w3(32'hbaf74e48),
	.w4(32'hbaad27a0),
	.w5(32'hbbf77316),
	.w6(32'hbb9b78f1),
	.w7(32'hbb214541),
	.w8(32'hb9cc5516),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3bf5b),
	.w1(32'h3ba733c6),
	.w2(32'h3ac492ac),
	.w3(32'h3bcdcc55),
	.w4(32'h3c695eaa),
	.w5(32'h3c1b4026),
	.w6(32'h39e156ae),
	.w7(32'h3b3165c5),
	.w8(32'h3c2b83d8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ec530),
	.w1(32'h3a5d2e9f),
	.w2(32'hba4f970c),
	.w3(32'h3b5c1103),
	.w4(32'h3b0eb48a),
	.w5(32'h3bc47fe5),
	.w6(32'hbb163ca9),
	.w7(32'hbb260692),
	.w8(32'h3b6ac99b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2603b9),
	.w1(32'hbaa60e96),
	.w2(32'h3bc7f944),
	.w3(32'hbaba3958),
	.w4(32'hba51736c),
	.w5(32'hba7e89cf),
	.w6(32'hbb4612a2),
	.w7(32'h3b6a1908),
	.w8(32'hba135e6e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d45a68),
	.w1(32'hba0d96c6),
	.w2(32'h3b59aac8),
	.w3(32'hbab8c4d0),
	.w4(32'h3af55506),
	.w5(32'h3a9a8a83),
	.w6(32'h3a606957),
	.w7(32'h3b4958bb),
	.w8(32'h3a1294b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66b8e5),
	.w1(32'h39178732),
	.w2(32'h3a14514a),
	.w3(32'h3ae93277),
	.w4(32'h39fefeb0),
	.w5(32'h3b000d0a),
	.w6(32'h3a96d206),
	.w7(32'h39a08c33),
	.w8(32'h3a11a92b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeee52),
	.w1(32'hbb423894),
	.w2(32'hbb6eb48a),
	.w3(32'hbaee4a55),
	.w4(32'hbb2701b4),
	.w5(32'hbaefbbbf),
	.w6(32'hbab225be),
	.w7(32'hbb1f2fd1),
	.w8(32'hbb424350),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac719d3),
	.w1(32'h3a1021bf),
	.w2(32'h3b156ee9),
	.w3(32'h3a55d47c),
	.w4(32'h3a84cfd1),
	.w5(32'hba9d5ff1),
	.w6(32'hb82736cf),
	.w7(32'hb7b503a8),
	.w8(32'h3ae09e19),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14ec06),
	.w1(32'h3b54e05e),
	.w2(32'h3b55f2bb),
	.w3(32'h39d6ee05),
	.w4(32'hba318f76),
	.w5(32'h3b1bc068),
	.w6(32'h3b4d1a1c),
	.w7(32'hb6f0dec1),
	.w8(32'h3af3f9d7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f549),
	.w1(32'hbb249bcd),
	.w2(32'hbb64cd15),
	.w3(32'h3a7b8235),
	.w4(32'hbacb6627),
	.w5(32'hb9580f0d),
	.w6(32'h3991c33b),
	.w7(32'hba98b5aa),
	.w8(32'h3a417923),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f3081),
	.w1(32'h3a5e16af),
	.w2(32'h3b5b27e1),
	.w3(32'h3a4026cf),
	.w4(32'h3b339be7),
	.w5(32'h3a0e27c5),
	.w6(32'h3b7b3028),
	.w7(32'h3ba2b886),
	.w8(32'hb94e857f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988c014),
	.w1(32'h3a92acdc),
	.w2(32'h39eac9bc),
	.w3(32'h3925d26d),
	.w4(32'h39ba79ab),
	.w5(32'hba239163),
	.w6(32'h3a370454),
	.w7(32'h37802611),
	.w8(32'hbaae5c81),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc4d68),
	.w1(32'hbb863b8a),
	.w2(32'hba4ae19d),
	.w3(32'hba99fbfa),
	.w4(32'h3970231e),
	.w5(32'h3a4eaeb6),
	.w6(32'hbb47d5c2),
	.w7(32'hbb4ca3af),
	.w8(32'hba2d6bbf),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbfb34),
	.w1(32'h3aa81703),
	.w2(32'h3a9b1d2f),
	.w3(32'h3aa9cc3a),
	.w4(32'h3977f4a9),
	.w5(32'h388882e0),
	.w6(32'h3a1a7842),
	.w7(32'h39625635),
	.w8(32'h3a9230be),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c1544),
	.w1(32'h3b2d199e),
	.w2(32'h3c0536c8),
	.w3(32'hb9f07739),
	.w4(32'h3bad48fe),
	.w5(32'h3b1608d8),
	.w6(32'h3ae53407),
	.w7(32'h3be18b49),
	.w8(32'h3a8b7532),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e38f0),
	.w1(32'hb9a8b327),
	.w2(32'hba4e3686),
	.w3(32'h3a19f054),
	.w4(32'h3926dd0b),
	.w5(32'hb93c80f1),
	.w6(32'hba831b59),
	.w7(32'hbabdd75e),
	.w8(32'hb923d180),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905e496),
	.w1(32'hba09cfa7),
	.w2(32'hba579c76),
	.w3(32'hb9f6f525),
	.w4(32'hb98fe016),
	.w5(32'hbb011e7a),
	.w6(32'hba7cdfc6),
	.w7(32'hba38bbe4),
	.w8(32'hba6d0bd0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3f5f),
	.w1(32'h3a7780ad),
	.w2(32'h3b71d3fc),
	.w3(32'hbb7ed118),
	.w4(32'hbb8a4c31),
	.w5(32'h3997815a),
	.w6(32'hbbacc7d5),
	.w7(32'hbaa3885e),
	.w8(32'hba0c64e3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23e358),
	.w1(32'h38190c16),
	.w2(32'h3a96da4a),
	.w3(32'hba4579e0),
	.w4(32'h3996b96d),
	.w5(32'hbbb4929b),
	.w6(32'hb9fa99dc),
	.w7(32'h382ab438),
	.w8(32'hbb90e81d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba859150),
	.w1(32'hba770193),
	.w2(32'h3b0f92d7),
	.w3(32'hbb99cb03),
	.w4(32'hbb53ea3e),
	.w5(32'h39ef564c),
	.w6(32'hba93a0de),
	.w7(32'hba3e9755),
	.w8(32'hbb3f3485),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a081b),
	.w1(32'hba348330),
	.w2(32'hbaa81ef5),
	.w3(32'h37a53a71),
	.w4(32'hb9bf4df1),
	.w5(32'hba925b7e),
	.w6(32'hba2a01f0),
	.w7(32'hba3cfacb),
	.w8(32'h3a5e8047),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c2413),
	.w1(32'h3ba2a9c4),
	.w2(32'h3bd252f1),
	.w3(32'hba870137),
	.w4(32'hba948f40),
	.w5(32'h39a37a99),
	.w6(32'hb963ef6b),
	.w7(32'h3a76913f),
	.w8(32'h38248202),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e36be),
	.w1(32'hb9cb2bf6),
	.w2(32'hba5d3c8f),
	.w3(32'h3a42b3b2),
	.w4(32'h3a436bcc),
	.w5(32'h3871bf8f),
	.w6(32'hb90b1f35),
	.w7(32'hb9ca56fa),
	.w8(32'hbab86238),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6f7f5),
	.w1(32'hbae9a1d7),
	.w2(32'hbaeac63e),
	.w3(32'hbb0daa79),
	.w4(32'hba3c9dc6),
	.w5(32'hbaa4b45b),
	.w6(32'hbafe4475),
	.w7(32'hba9c18a6),
	.w8(32'hbaeabcff),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0636e1),
	.w1(32'hba0abef8),
	.w2(32'h3aa086f2),
	.w3(32'hbaf5a4bc),
	.w4(32'hba9c85ae),
	.w5(32'hba1d23fd),
	.w6(32'hba7608a9),
	.w7(32'hb81610de),
	.w8(32'h3a1e60ed),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b2eae),
	.w1(32'h3b0e0886),
	.w2(32'h3b897d5d),
	.w3(32'hbade806d),
	.w4(32'h3a663a5b),
	.w5(32'h3b050a10),
	.w6(32'h3aae084d),
	.w7(32'h3b25f441),
	.w8(32'h3b90373c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810a08),
	.w1(32'h3b8eaa56),
	.w2(32'h3bbdc1a4),
	.w3(32'h3aad52f6),
	.w4(32'h3b84bdc7),
	.w5(32'h3add209c),
	.w6(32'h3a9d791e),
	.w7(32'h3bc5985f),
	.w8(32'h3a8a0f08),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74130c),
	.w1(32'h3a7b5b7c),
	.w2(32'h3a75b171),
	.w3(32'h3add0955),
	.w4(32'h3a3aec96),
	.w5(32'h3a053e29),
	.w6(32'h3abaf6c2),
	.w7(32'h38953b8f),
	.w8(32'hbaa14e2c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057cf7),
	.w1(32'hbb0fba67),
	.w2(32'hbaa82935),
	.w3(32'h39b7f201),
	.w4(32'h3a24711e),
	.w5(32'h39c9ef53),
	.w6(32'hbac0e7c5),
	.w7(32'hbb10d5e7),
	.w8(32'h39ecae08),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf86d3),
	.w1(32'h3ab13337),
	.w2(32'h38bdddfb),
	.w3(32'hba34431a),
	.w4(32'hba7d3c17),
	.w5(32'h3aad820b),
	.w6(32'h38fafa6f),
	.w7(32'hbab5b6a1),
	.w8(32'h39275d38),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d81be6),
	.w1(32'hbab0075c),
	.w2(32'hba8dc98d),
	.w3(32'h3910bdbd),
	.w4(32'hba30c8f9),
	.w5(32'hbabf1f0f),
	.w6(32'h39cac711),
	.w7(32'h387d20e7),
	.w8(32'hbae3824e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba822d76),
	.w1(32'hba82b94d),
	.w2(32'h3b2ba183),
	.w3(32'h3a7732dd),
	.w4(32'h3b381e35),
	.w5(32'h3a1d9ca8),
	.w6(32'h3af3c059),
	.w7(32'h3bd10682),
	.w8(32'hb8ed3591),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0ff9d),
	.w1(32'hb9c28fa5),
	.w2(32'h382ec001),
	.w3(32'h39133f2a),
	.w4(32'h3a10e47d),
	.w5(32'hbb794d3d),
	.w6(32'hb9597024),
	.w7(32'hba2e8d1a),
	.w8(32'hbb9f7557),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca23f),
	.w1(32'hba99c271),
	.w2(32'h3a29dde6),
	.w3(32'hbb452d6d),
	.w4(32'hbaac0e63),
	.w5(32'h3adca788),
	.w6(32'hbb26cbb8),
	.w7(32'h3aa13272),
	.w8(32'h3a9d60ae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58aaa0),
	.w1(32'h3a96e92c),
	.w2(32'h3a991137),
	.w3(32'h398b8ec6),
	.w4(32'h3a531859),
	.w5(32'h39fa3499),
	.w6(32'hbac92c9b),
	.w7(32'hba5a28cf),
	.w8(32'hb79d72a0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e4734),
	.w1(32'h3a5caa5e),
	.w2(32'h3a67553e),
	.w3(32'h3a440d01),
	.w4(32'h38fe2538),
	.w5(32'h3a0a7fbf),
	.w6(32'h3a56f90c),
	.w7(32'hb947adf4),
	.w8(32'h3a8e60db),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af69d61),
	.w1(32'hbb58604e),
	.w2(32'hbb51ee6e),
	.w3(32'h3a714af6),
	.w4(32'h3a2a4548),
	.w5(32'h388f9b86),
	.w6(32'hb99affc2),
	.w7(32'hbb3fd512),
	.w8(32'h3a07a522),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138020),
	.w1(32'h386cfad0),
	.w2(32'hb7b2f24b),
	.w3(32'h39ef10de),
	.w4(32'h3a5330e0),
	.w5(32'hba68d98c),
	.w6(32'h3aebea79),
	.w7(32'h3a2507f4),
	.w8(32'hbad68624),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021c6c),
	.w1(32'h3a3a1963),
	.w2(32'h3af2af2c),
	.w3(32'h3994432e),
	.w4(32'hb96ff6ee),
	.w5(32'hba68d4e7),
	.w6(32'h3a1a1053),
	.w7(32'h3af1c22e),
	.w8(32'hba7d0bdb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01dcaa),
	.w1(32'h3a36aed2),
	.w2(32'h3a4e7a60),
	.w3(32'hba9806e8),
	.w4(32'hba0db648),
	.w5(32'h3a43cb95),
	.w6(32'hb8fdde4a),
	.w7(32'hb8e7e6b3),
	.w8(32'h3991e788),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6edf9),
	.w1(32'h3a9b0cac),
	.w2(32'h3acb2d38),
	.w3(32'h3a33e19c),
	.w4(32'h3a7fc44c),
	.w5(32'hb8ba577a),
	.w6(32'h3addf4f5),
	.w7(32'h3a77af95),
	.w8(32'h39296668),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9021a0),
	.w1(32'h3902f88c),
	.w2(32'h38138039),
	.w3(32'h3a10573b),
	.w4(32'h3adbfd18),
	.w5(32'hba484f4a),
	.w6(32'hb9a1b9e1),
	.w7(32'h3a868a63),
	.w8(32'hba27105d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acc65d),
	.w1(32'h3a77d0fc),
	.w2(32'h3a937353),
	.w3(32'hbab898d5),
	.w4(32'hba348943),
	.w5(32'hb7146695),
	.w6(32'hba2a4707),
	.w7(32'hb7616c9f),
	.w8(32'hb9dfaa73),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8d409),
	.w1(32'h3983db58),
	.w2(32'h39de519f),
	.w3(32'hba3c0a81),
	.w4(32'hba168669),
	.w5(32'hbb084f4b),
	.w6(32'h3617e1ef),
	.w7(32'hba67bacf),
	.w8(32'hbae8e38d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac76463),
	.w1(32'hba170acd),
	.w2(32'hb9a543c8),
	.w3(32'hbb104c5d),
	.w4(32'hbb02c7e8),
	.w5(32'hba51f783),
	.w6(32'h39450e53),
	.w7(32'hba6cbe5c),
	.w8(32'hba5f2e5e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba192b2f),
	.w1(32'h3a7db32c),
	.w2(32'h3b36b6f1),
	.w3(32'hbb1cad0d),
	.w4(32'hb8143091),
	.w5(32'h3b1011c2),
	.w6(32'hb96f8f33),
	.w7(32'h3a596fbe),
	.w8(32'h3b03ab8a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6be9d),
	.w1(32'h39ec21fd),
	.w2(32'h3a2e4069),
	.w3(32'h3af16f1d),
	.w4(32'h3aecb6c5),
	.w5(32'hbb0c0d9a),
	.w6(32'h3a3b77e1),
	.w7(32'h3a42869f),
	.w8(32'hbb2ba57a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade5d35),
	.w1(32'hbb828ba7),
	.w2(32'hbb21afae),
	.w3(32'hbb66758f),
	.w4(32'hbb986e0a),
	.w5(32'hba2a0720),
	.w6(32'hbb8a9986),
	.w7(32'hbb2a8916),
	.w8(32'hba621a54),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0e63a),
	.w1(32'hb9796bfa),
	.w2(32'hb999fc46),
	.w3(32'hba12cb84),
	.w4(32'hb9d21a41),
	.w5(32'hba4acc06),
	.w6(32'h38e342da),
	.w7(32'hb9f7c2c6),
	.w8(32'hba9e01de),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f23f5),
	.w1(32'hbacd2527),
	.w2(32'hbac90fab),
	.w3(32'hba432f59),
	.w4(32'hba719de2),
	.w5(32'h3a159dea),
	.w6(32'hb9e68ca6),
	.w7(32'hba8905d0),
	.w8(32'hb8e0e471),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e2987),
	.w1(32'h3ad9cb81),
	.w2(32'h3b54c41d),
	.w3(32'h3a5c7502),
	.w4(32'h3b15c548),
	.w5(32'h39cc25bc),
	.w6(32'h3aa9be26),
	.w7(32'h3b14d8ef),
	.w8(32'h39ffa03b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906ef12),
	.w1(32'hb9e67e17),
	.w2(32'hb9148353),
	.w3(32'h38c74661),
	.w4(32'hb8d41541),
	.w5(32'h3a4f00f1),
	.w6(32'h39798a77),
	.w7(32'h37de58e9),
	.w8(32'h3a79e67d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383be751),
	.w1(32'h3983fbd3),
	.w2(32'h3937cdba),
	.w3(32'h3a828ee5),
	.w4(32'h3a88bf32),
	.w5(32'hbb18aaa9),
	.w6(32'h3ab2c6ee),
	.w7(32'h399b6196),
	.w8(32'hbb0b270e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fa6de),
	.w1(32'h3b7bef8c),
	.w2(32'h3bf98537),
	.w3(32'hba61f264),
	.w4(32'h3a771008),
	.w5(32'h3a81c254),
	.w6(32'h3b134f1d),
	.w7(32'h3bdaf0a4),
	.w8(32'h3a1b98c4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923d072),
	.w1(32'h3a629f20),
	.w2(32'hba22bd48),
	.w3(32'h3a79b5cf),
	.w4(32'h3a590b8c),
	.w5(32'h3983ce79),
	.w6(32'h3ac44135),
	.w7(32'h3985cb6c),
	.w8(32'h3a53e41d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9266d1),
	.w1(32'h3a995343),
	.w2(32'h39c3f093),
	.w3(32'h39c0c31e),
	.w4(32'h39c4bd61),
	.w5(32'hbbd2128a),
	.w6(32'h3a562070),
	.w7(32'h38c21ad2),
	.w8(32'hbb674664),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28d488),
	.w1(32'hbae790e7),
	.w2(32'hbad94940),
	.w3(32'hbb8eda09),
	.w4(32'hbbd5bbc2),
	.w5(32'hb944cde5),
	.w6(32'hba579084),
	.w7(32'hbbd937bf),
	.w8(32'h38252c97),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8849e73),
	.w1(32'h3a785f26),
	.w2(32'h3a0a6a20),
	.w3(32'hb7c1ef4d),
	.w4(32'hb8d00049),
	.w5(32'h3ac7376d),
	.w6(32'hb99e53df),
	.w7(32'hba7abc4c),
	.w8(32'h3b12ce73),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1319e),
	.w1(32'h3c1b7c3a),
	.w2(32'h3c025b62),
	.w3(32'h3951db50),
	.w4(32'h3a9b6bdf),
	.w5(32'hba154f88),
	.w6(32'h3b7490d9),
	.w7(32'h3b6e9345),
	.w8(32'hbaa011aa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25218),
	.w1(32'hbae8a2c9),
	.w2(32'hbaca0b3d),
	.w3(32'hba3fc74f),
	.w4(32'h39dc1e6d),
	.w5(32'h3b23a956),
	.w6(32'hbab8c47d),
	.w7(32'hba26e200),
	.w8(32'h3b3acb2d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b297a73),
	.w1(32'h3b1737ef),
	.w2(32'h3b8e76c1),
	.w3(32'h3aa7e09b),
	.w4(32'h3b87c2f8),
	.w5(32'h3b1d767d),
	.w6(32'h3b1a4e40),
	.w7(32'h3b994886),
	.w8(32'h3aba1fdf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5843),
	.w1(32'hb9b5bf89),
	.w2(32'hba2c07b6),
	.w3(32'hbab6c8f1),
	.w4(32'hba8ada0f),
	.w5(32'hba279f2d),
	.w6(32'hbb2adace),
	.w7(32'hbb19a512),
	.w8(32'hbabf0246),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe2b1),
	.w1(32'h3a9755f4),
	.w2(32'h3a731eb5),
	.w3(32'hbb157d5f),
	.w4(32'hbb2b27b5),
	.w5(32'h3a8d2d4b),
	.w6(32'hb85982a5),
	.w7(32'h3a7c9145),
	.w8(32'h3a55454d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39769c05),
	.w1(32'h394ea5ab),
	.w2(32'h3ab26293),
	.w3(32'h38b57e68),
	.w4(32'hb92d1a37),
	.w5(32'hba5854a3),
	.w6(32'hb917bf7b),
	.w7(32'hb9d44438),
	.w8(32'hba31ccd2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ae17a),
	.w1(32'hbb45554b),
	.w2(32'hbb677739),
	.w3(32'hbb2eff6c),
	.w4(32'hbafc2d47),
	.w5(32'h3b53a292),
	.w6(32'hbac683d3),
	.w7(32'hb8a78c3e),
	.w8(32'h3a4df4f3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec5c7),
	.w1(32'hba940df9),
	.w2(32'hbb008448),
	.w3(32'h3b4c84b6),
	.w4(32'h3b172cfc),
	.w5(32'hbb649001),
	.w6(32'h39fee735),
	.w7(32'hb9c7a87f),
	.w8(32'hbb33492e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c177),
	.w1(32'h3955ff5d),
	.w2(32'h3939e0e8),
	.w3(32'hbb768e72),
	.w4(32'hbb1d97e2),
	.w5(32'h396f0ae2),
	.w6(32'hba84c663),
	.w7(32'hb86a7581),
	.w8(32'hb98da5b4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a12917),
	.w1(32'hba1cc165),
	.w2(32'h3a345b55),
	.w3(32'hba5c493d),
	.w4(32'h3a21dfee),
	.w5(32'hbaea07a2),
	.w6(32'hb9e2bcf1),
	.w7(32'h3aa4a69d),
	.w8(32'hbb7022fa),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7759ed),
	.w1(32'h3bde39a6),
	.w2(32'h3b38fcb6),
	.w3(32'hbb2e53a3),
	.w4(32'hbac01221),
	.w5(32'hba5999cd),
	.w6(32'hbb052b77),
	.w7(32'hbb24cb9a),
	.w8(32'h3a89cbb7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62ca39),
	.w1(32'h3b583b36),
	.w2(32'h3b2303ea),
	.w3(32'h3a824e01),
	.w4(32'h3af923b8),
	.w5(32'hbb321ce0),
	.w6(32'h3b5cc65d),
	.w7(32'h3af936f8),
	.w8(32'hbb20e281),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134697),
	.w1(32'hbaf82056),
	.w2(32'hbb12a9b3),
	.w3(32'hbb56db17),
	.w4(32'hbb796021),
	.w5(32'h39f865d0),
	.w6(32'hbac8b8ce),
	.w7(32'hbb126fbe),
	.w8(32'h3a25fa0f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa79e8f),
	.w1(32'h39ae6a06),
	.w2(32'h3aad1560),
	.w3(32'hba4c0067),
	.w4(32'hb8794a15),
	.w5(32'hb9d1df47),
	.w6(32'h39b21869),
	.w7(32'h3a27555c),
	.w8(32'hb89635d2),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6d461),
	.w1(32'h38486869),
	.w2(32'hba42aa2d),
	.w3(32'hba690312),
	.w4(32'hba46f9ed),
	.w5(32'hbacde8f4),
	.w6(32'hba5906d9),
	.w7(32'hbab3122f),
	.w8(32'hbb04d427),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5047f),
	.w1(32'hb9a5a484),
	.w2(32'hbade988c),
	.w3(32'hbab6b0c9),
	.w4(32'hbb84ece3),
	.w5(32'hba450b18),
	.w6(32'hba6f76d5),
	.w7(32'hbb22c8d0),
	.w8(32'hba394b63),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea4e00),
	.w1(32'h39a5877e),
	.w2(32'h3a7e62de),
	.w3(32'hbac0c93c),
	.w4(32'hbb513b41),
	.w5(32'h39aaba14),
	.w6(32'hba8d578e),
	.w7(32'hbb260bd1),
	.w8(32'hbaabced4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33d744),
	.w1(32'hbaa6a052),
	.w2(32'hba2312c6),
	.w3(32'h3953d383),
	.w4(32'h3a5cd605),
	.w5(32'h3b2cf756),
	.w6(32'hba346a12),
	.w7(32'hb9f81ec0),
	.w8(32'h3a49ac17),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae5d2f),
	.w1(32'hb76c8403),
	.w2(32'hb896d17e),
	.w3(32'h3b03e8c0),
	.w4(32'h3aed3029),
	.w5(32'h3a243ee9),
	.w6(32'h3a5f36b8),
	.w7(32'h3a69fe79),
	.w8(32'hbb09b24b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd0fa),
	.w1(32'h3b2b375b),
	.w2(32'h3b422647),
	.w3(32'hb9ccb905),
	.w4(32'h3a23f3e5),
	.w5(32'h3b6346cd),
	.w6(32'h3a57eb7d),
	.w7(32'h3aaf7901),
	.w8(32'h3b157c7e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9213fd7),
	.w1(32'h3a63bbcf),
	.w2(32'hba67464a),
	.w3(32'h3b4e93ff),
	.w4(32'h3aa46a5b),
	.w5(32'h3b82f214),
	.w6(32'h3b4f448b),
	.w7(32'h3a8ed8c9),
	.w8(32'h3afb46a0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad015d1),
	.w1(32'hba411762),
	.w2(32'hb9e5e9de),
	.w3(32'h3b07fd04),
	.w4(32'h3b4b1463),
	.w5(32'h3b03128e),
	.w6(32'hb9b937ac),
	.w7(32'h3a9c2278),
	.w8(32'h3b3428a3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab92fa3),
	.w1(32'h3ad7ff3e),
	.w2(32'h3b638fff),
	.w3(32'hb8b052ce),
	.w4(32'h3abfcb79),
	.w5(32'hba2190ab),
	.w6(32'h3a9aebde),
	.w7(32'h3b4ace1e),
	.w8(32'h38eb0a17),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbfed5),
	.w1(32'h3aab9b61),
	.w2(32'h3a325fd6),
	.w3(32'hb969c963),
	.w4(32'hb8f68abc),
	.w5(32'h3a87b041),
	.w6(32'hb9e5c57e),
	.w7(32'hba1e2a95),
	.w8(32'h3a99850b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0809a),
	.w1(32'h3ac9638f),
	.w2(32'h3a782384),
	.w3(32'h39c48d59),
	.w4(32'h3a536fc8),
	.w5(32'h3a86f14b),
	.w6(32'h3a33fb33),
	.w7(32'h3a0a3ba9),
	.w8(32'h3a050dfc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9f78),
	.w1(32'h39ab5446),
	.w2(32'hb9faab27),
	.w3(32'h3a948767),
	.w4(32'h3a9f032b),
	.w5(32'hba25b4e5),
	.w6(32'h3a4bfd47),
	.w7(32'hb7b20609),
	.w8(32'h3b0f0a66),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6c0e),
	.w1(32'h3b877ea2),
	.w2(32'h3b850935),
	.w3(32'hbace074e),
	.w4(32'hb9e34081),
	.w5(32'hb9eeb41a),
	.w6(32'hbacc57a8),
	.w7(32'h3b17fcbb),
	.w8(32'hbab8283d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af65a9),
	.w1(32'hb81d28d8),
	.w2(32'h3a707d54),
	.w3(32'hb9fbe445),
	.w4(32'hba318c1f),
	.w5(32'h3b4e8fbf),
	.w6(32'hb9906a78),
	.w7(32'h396ac2f8),
	.w8(32'h3b870bb2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0987ce),
	.w1(32'hbb066144),
	.w2(32'hbaada8a9),
	.w3(32'h3b5e00df),
	.w4(32'h3b3e0e91),
	.w5(32'hbaa95bcb),
	.w6(32'h3aa9d711),
	.w7(32'h3ab65573),
	.w8(32'hbb111831),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad58c27),
	.w1(32'hb9fd2dfc),
	.w2(32'hba1b9860),
	.w3(32'hbaa5ba39),
	.w4(32'hba90531d),
	.w5(32'hba544add),
	.w6(32'hbaa9504c),
	.w7(32'hbaf34a3a),
	.w8(32'hbb36a742),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3af94d),
	.w1(32'h3ac3cad4),
	.w2(32'h3b8e2e07),
	.w3(32'hb94b9be7),
	.w4(32'h3b0d50ba),
	.w5(32'hbaa72400),
	.w6(32'h3a106c42),
	.w7(32'h3b94e105),
	.w8(32'hbb32973a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54aef9),
	.w1(32'h3b100e94),
	.w2(32'h38fb21ff),
	.w3(32'hbad81c18),
	.w4(32'hbb21d66f),
	.w5(32'h3aec0573),
	.w6(32'hb88da955),
	.w7(32'hba9e61f7),
	.w8(32'h3a4fcd3b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af81839),
	.w1(32'h3ba08568),
	.w2(32'h3b6725f6),
	.w3(32'h3b18d31a),
	.w4(32'h3a02da47),
	.w5(32'h3aab4edd),
	.w6(32'h3b0479bb),
	.w7(32'h3a9ce996),
	.w8(32'h3a935c2b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8368d2),
	.w1(32'h3a9a9f84),
	.w2(32'h3a8b4503),
	.w3(32'h3ac34c72),
	.w4(32'hba2fbbbc),
	.w5(32'h3a8e58ad),
	.w6(32'h3ac78850),
	.w7(32'hb995c450),
	.w8(32'h39c0461d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42c09c),
	.w1(32'hb8e4a0aa),
	.w2(32'hb9febeaf),
	.w3(32'hb817dc5d),
	.w4(32'h3a051946),
	.w5(32'hbac16ec1),
	.w6(32'hb9466d6e),
	.w7(32'hba1a8b18),
	.w8(32'h38f09b70),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0a207),
	.w1(32'hba19eea7),
	.w2(32'hbb12625a),
	.w3(32'hb9716eb4),
	.w4(32'hb8fc0440),
	.w5(32'hba996acd),
	.w6(32'hb9c89c7c),
	.w7(32'hb961d286),
	.w8(32'hba7409e6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99ea55),
	.w1(32'h3a4633d6),
	.w2(32'hb9f4b42b),
	.w3(32'hbaeae17b),
	.w4(32'hbaa9a7fe),
	.w5(32'h38905203),
	.w6(32'hba8df9a4),
	.w7(32'hbaad3b34),
	.w8(32'hb9a1bcc6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b5a8),
	.w1(32'hbaf81b91),
	.w2(32'hba85aa79),
	.w3(32'h3a4c4a24),
	.w4(32'h3aeb470d),
	.w5(32'h395c4c02),
	.w6(32'hb9eccb20),
	.w7(32'hba54628a),
	.w8(32'hbb518cc6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad30424),
	.w1(32'h3aac97c1),
	.w2(32'hb81195ac),
	.w3(32'h39872d26),
	.w4(32'h3ac3237d),
	.w5(32'hbb395b31),
	.w6(32'hbb875c7b),
	.w7(32'hbb50549a),
	.w8(32'hbb0b33da),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b21fd),
	.w1(32'h3b86a5d4),
	.w2(32'h3b271b1b),
	.w3(32'hbb5f6107),
	.w4(32'hbb9d7019),
	.w5(32'hbb002730),
	.w6(32'hba513c00),
	.w7(32'hbb4ed485),
	.w8(32'hbb831fd3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb447159),
	.w1(32'hbab10ef5),
	.w2(32'h3a955f72),
	.w3(32'hbb1cd3fa),
	.w4(32'hba3cebb3),
	.w5(32'h3ae65ec6),
	.w6(32'hbb5ce893),
	.w7(32'hba9a5cbc),
	.w8(32'h390f3f95),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae91209),
	.w1(32'h3ac57a75),
	.w2(32'h3b48dcbc),
	.w3(32'h3a2ecb47),
	.w4(32'h3adb89ff),
	.w5(32'h3a18d233),
	.w6(32'h3a928544),
	.w7(32'h3b19966a),
	.w8(32'h3a11f25b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a566e13),
	.w1(32'h3922051c),
	.w2(32'h3a2203db),
	.w3(32'h3a4b6967),
	.w4(32'h3affc0ed),
	.w5(32'hbb79b02b),
	.w6(32'hb9a6286b),
	.w7(32'h3a4184ce),
	.w8(32'hbb1cbe66),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba529866),
	.w1(32'hba3a046d),
	.w2(32'h3b1046b2),
	.w3(32'hbb3abf1d),
	.w4(32'h383e7ec9),
	.w5(32'hbb7a6d90),
	.w6(32'hba9441b7),
	.w7(32'h3a607c09),
	.w8(32'hbb950446),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa8f5),
	.w1(32'hbb35d80c),
	.w2(32'h3b990c72),
	.w3(32'hbba22199),
	.w4(32'h3a15298c),
	.w5(32'hb99e348e),
	.w6(32'hbb8ec904),
	.w7(32'h3b224bd6),
	.w8(32'hbb4845d7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c461),
	.w1(32'hbb08ef9e),
	.w2(32'h3994906f),
	.w3(32'h387a33d5),
	.w4(32'h3ab9bf4e),
	.w5(32'h39125514),
	.w6(32'hba959a5b),
	.w7(32'h3a4893b0),
	.w8(32'hba008852),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878fb7a),
	.w1(32'hb800185f),
	.w2(32'hba4721b4),
	.w3(32'hb952d705),
	.w4(32'h39e809a3),
	.w5(32'h3aceac73),
	.w6(32'h3a80805e),
	.w7(32'h398f6ba0),
	.w8(32'h3b01133d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96037e),
	.w1(32'h3a9ebd4a),
	.w2(32'h3a18d431),
	.w3(32'h3af9b355),
	.w4(32'h3b07fccb),
	.w5(32'hb818ab12),
	.w6(32'h3a27eb12),
	.w7(32'h3a1ea573),
	.w8(32'hb88b1201),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4a63e),
	.w1(32'h39f3a3b2),
	.w2(32'h3a111968),
	.w3(32'h395027ca),
	.w4(32'h3a9d4b9a),
	.w5(32'hba1e115a),
	.w6(32'hba6a40fd),
	.w7(32'hba9f67a8),
	.w8(32'hb9d8f77a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82ad074),
	.w1(32'h3a8aac59),
	.w2(32'h3a67820a),
	.w3(32'hbacc99d4),
	.w4(32'hbae4d8fb),
	.w5(32'hb9d9e40d),
	.w6(32'h37e8d4de),
	.w7(32'h3987f468),
	.w8(32'hb9c12e77),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae8bbb),
	.w1(32'hb7f52301),
	.w2(32'h3a18e5c0),
	.w3(32'hba38f913),
	.w4(32'h3993754f),
	.w5(32'h3939afe9),
	.w6(32'h393f0c5c),
	.w7(32'hb8d1a2be),
	.w8(32'h3a532349),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f9462),
	.w1(32'h3a199f75),
	.w2(32'hb9a411c0),
	.w3(32'h3917d9d1),
	.w4(32'hba52a06d),
	.w5(32'hba51230d),
	.w6(32'h3a44c95c),
	.w7(32'h38352390),
	.w8(32'h3af07900),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4029b),
	.w1(32'h3b17e1fe),
	.w2(32'h3b179da5),
	.w3(32'hb9ac0397),
	.w4(32'hbb053d72),
	.w5(32'h3abcd8a6),
	.w6(32'h3b464d34),
	.w7(32'hba45538d),
	.w8(32'hba5f4a24),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab31457),
	.w1(32'hbb0b0f17),
	.w2(32'hbaff72ae),
	.w3(32'h3a856b68),
	.w4(32'hb8a8915b),
	.w5(32'hb9a90aab),
	.w6(32'h39d11f09),
	.w7(32'hb9f65a5e),
	.w8(32'h3aea7d9f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5f8b),
	.w1(32'h3aabaf81),
	.w2(32'h3a8391b3),
	.w3(32'h3a0a2c42),
	.w4(32'hb930069b),
	.w5(32'hb9ae46e4),
	.w6(32'h3afdcfdb),
	.w7(32'h3ad5a081),
	.w8(32'hb9aea24d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa86174),
	.w1(32'h3a9a30a5),
	.w2(32'h3a69da36),
	.w3(32'hba4908d1),
	.w4(32'h3958e3fe),
	.w5(32'h36bdaad8),
	.w6(32'hba85dda6),
	.w7(32'hba5eee5f),
	.w8(32'h3a44119d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbf690),
	.w1(32'h3b1d3caf),
	.w2(32'h3a0e55da),
	.w3(32'h3aed876d),
	.w4(32'h3aba8601),
	.w5(32'h39652842),
	.w6(32'h3af9e447),
	.w7(32'h3b0ee748),
	.w8(32'h39cbc8a3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bada48),
	.w1(32'hb9b8c7c0),
	.w2(32'hb84e22a9),
	.w3(32'h3a4f000d),
	.w4(32'h3a387a91),
	.w5(32'hb9de2a57),
	.w6(32'h3a742060),
	.w7(32'h3acfb96f),
	.w8(32'h3a916108),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55575c),
	.w1(32'hbaf75a4f),
	.w2(32'h3a24d214),
	.w3(32'hbaceaee2),
	.w4(32'hb9e5222b),
	.w5(32'hba25db74),
	.w6(32'h3a9bd2ed),
	.w7(32'hb9ca4aad),
	.w8(32'h3ac6fff6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e6ced),
	.w1(32'h37f16428),
	.w2(32'h3b02d6e9),
	.w3(32'hb89acd92),
	.w4(32'h3abe8e7f),
	.w5(32'hb9d750cc),
	.w6(32'h3b12dc00),
	.w7(32'h3ae24406),
	.w8(32'h3aa14f8e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6914a4),
	.w1(32'hbb17c6e4),
	.w2(32'hbb229d47),
	.w3(32'h39aa389b),
	.w4(32'hb9eede8d),
	.w5(32'hb8a60894),
	.w6(32'h3b30872a),
	.w7(32'hbae9591b),
	.w8(32'hba80f1de),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e54bf),
	.w1(32'hba9a14f0),
	.w2(32'hbaca1b92),
	.w3(32'hba64a41d),
	.w4(32'h3a048153),
	.w5(32'h3aa9a407),
	.w6(32'hbaea334c),
	.w7(32'hbad07a62),
	.w8(32'hb98cfd85),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60264f),
	.w1(32'hbab50af9),
	.w2(32'h3af37298),
	.w3(32'h3a3842a6),
	.w4(32'h3b509ebf),
	.w5(32'hba891210),
	.w6(32'h3a1e3aaf),
	.w7(32'h3af7c193),
	.w8(32'h3ad6eddf),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2abe08),
	.w1(32'h3aef5b22),
	.w2(32'h3b8a841e),
	.w3(32'h37b2f3dc),
	.w4(32'h3a089bd0),
	.w5(32'h3a406792),
	.w6(32'h3b46800e),
	.w7(32'h3baaf69c),
	.w8(32'h3a1fc750),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bfe30),
	.w1(32'h3ab5ee39),
	.w2(32'h3acaa245),
	.w3(32'h3a883fe6),
	.w4(32'h3a9accec),
	.w5(32'h3b173204),
	.w6(32'h3aaf1644),
	.w7(32'h3a919c8c),
	.w8(32'h39fc1ebd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa05686),
	.w1(32'hba008536),
	.w2(32'hba7755ed),
	.w3(32'h3b1112bf),
	.w4(32'hba9d42fc),
	.w5(32'h3ad30dce),
	.w6(32'h39ddb5ab),
	.w7(32'hbb12d72c),
	.w8(32'h3b08b13f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcc7f0),
	.w1(32'h3a84d7b3),
	.w2(32'h3a816e87),
	.w3(32'h39c15ac1),
	.w4(32'h3a9ff596),
	.w5(32'h3ad1005f),
	.w6(32'h3a3352c3),
	.w7(32'h3a77fa7c),
	.w8(32'h3a7f0f67),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bad6a5),
	.w1(32'h389439f0),
	.w2(32'hba21fb0e),
	.w3(32'h3afac0b3),
	.w4(32'hb9cfe3bd),
	.w5(32'h3b62ca05),
	.w6(32'h3ab7c13d),
	.w7(32'hbac0c356),
	.w8(32'h387c150c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4cd66),
	.w1(32'h3a7915cc),
	.w2(32'hb9e260ed),
	.w3(32'h3a9082e8),
	.w4(32'h39266d12),
	.w5(32'h3aa2e5c1),
	.w6(32'h3a85b2a6),
	.w7(32'hba22057e),
	.w8(32'h3aa94bef),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6548),
	.w1(32'h3ae23034),
	.w2(32'h3a80e613),
	.w3(32'h39fc74e3),
	.w4(32'hba00eb27),
	.w5(32'h3b0a73eb),
	.w6(32'hb899c0dd),
	.w7(32'hb9e1a8c7),
	.w8(32'h3aeab347),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada833b),
	.w1(32'hba2b07a1),
	.w2(32'hbac7a7e3),
	.w3(32'h3a79aad9),
	.w4(32'h3921186b),
	.w5(32'h3a32c340),
	.w6(32'hb90706ae),
	.w7(32'hba9f9820),
	.w8(32'hbaf0a473),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a3b05),
	.w1(32'hbaf59ad3),
	.w2(32'hb95bca03),
	.w3(32'h3acfd20f),
	.w4(32'h3b10fe24),
	.w5(32'hba0fb656),
	.w6(32'hb9debf0f),
	.w7(32'hba7ffdd2),
	.w8(32'h3aa2be3a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bebf18),
	.w1(32'hb92b32e9),
	.w2(32'hbaffaee0),
	.w3(32'h3982b031),
	.w4(32'hbaf1cf24),
	.w5(32'h3ab99c20),
	.w6(32'h3a88b6f5),
	.w7(32'hb9129b84),
	.w8(32'h39f63bed),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a51344),
	.w1(32'hba7b6ce9),
	.w2(32'hbb878dfa),
	.w3(32'h3ab2726b),
	.w4(32'hbb397500),
	.w5(32'h3832e7c3),
	.w6(32'h382b7217),
	.w7(32'hbb85ee31),
	.w8(32'h39cc261c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39533a8a),
	.w1(32'h39e029c4),
	.w2(32'h3a63769a),
	.w3(32'h39b84c7d),
	.w4(32'h3a37dc2c),
	.w5(32'hba4b980e),
	.w6(32'h3a25701b),
	.w7(32'h3a6d0adb),
	.w8(32'hba89d29b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95029f8),
	.w1(32'h390d20a8),
	.w2(32'h3a2172c3),
	.w3(32'hba29518c),
	.w4(32'hb9e76f9b),
	.w5(32'hb9900f83),
	.w6(32'hbaadc765),
	.w7(32'hba25cde5),
	.w8(32'hb990e2b1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383fecd2),
	.w1(32'h39e87a46),
	.w2(32'h39dd0723),
	.w3(32'h38ba2675),
	.w4(32'h3a001bb2),
	.w5(32'h3b14ff3b),
	.w6(32'h399ac3d6),
	.w7(32'h39eba918),
	.w8(32'h3b09d37e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af99b87),
	.w1(32'h3b35b187),
	.w2(32'h3b3e3eb5),
	.w3(32'h3b242dad),
	.w4(32'h3ad51770),
	.w5(32'hb9359100),
	.w6(32'h3b4a532e),
	.w7(32'h3b3454b9),
	.w8(32'hb9ee2a81),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa657ff),
	.w1(32'hba618b8b),
	.w2(32'h3a9e6f35),
	.w3(32'hb95ff826),
	.w4(32'h38cfea83),
	.w5(32'h3a7c5e53),
	.w6(32'h38dda121),
	.w7(32'h39edade9),
	.w8(32'h3a58a200),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fc1f0),
	.w1(32'h38f5bee9),
	.w2(32'h3a316603),
	.w3(32'h3831d3fb),
	.w4(32'h3a575bbd),
	.w5(32'hba8b54e8),
	.w6(32'hb9d40fac),
	.w7(32'h39e991db),
	.w8(32'hb99a6500),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12a0be),
	.w1(32'hb9f77bce),
	.w2(32'hba30d31a),
	.w3(32'hba547c7b),
	.w4(32'hba96a5b2),
	.w5(32'hb9f23347),
	.w6(32'h37816357),
	.w7(32'hba05c8cf),
	.w8(32'hb9b62650),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39e478),
	.w1(32'hb988f339),
	.w2(32'hb9da2091),
	.w3(32'hb96c885f),
	.w4(32'hb9d8dacd),
	.w5(32'hba37610f),
	.w6(32'hb9076043),
	.w7(32'hb9fa56be),
	.w8(32'hba3a538e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba731aeb),
	.w1(32'hbaa5559c),
	.w2(32'hbaa5eeaa),
	.w3(32'hba3ac931),
	.w4(32'hba51ca3c),
	.w5(32'h3900b997),
	.w6(32'hba983b4f),
	.w7(32'hbad3d33a),
	.w8(32'hb8fd9543),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba064d57),
	.w1(32'h394a5541),
	.w2(32'h39ad6347),
	.w3(32'h39a2209e),
	.w4(32'h3a0c81fa),
	.w5(32'h3a63cd9f),
	.w6(32'h39dd9304),
	.w7(32'h3a12df73),
	.w8(32'h3aced3fe),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31230),
	.w1(32'h3ada09e4),
	.w2(32'h3af210b6),
	.w3(32'h3ab7796a),
	.w4(32'h3ae976a0),
	.w5(32'hb94a4473),
	.w6(32'h3af8830e),
	.w7(32'h3b0cc222),
	.w8(32'hb97a216e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4cffc),
	.w1(32'hb9990a64),
	.w2(32'hb9c00451),
	.w3(32'hb9d5df8e),
	.w4(32'hb9d3e073),
	.w5(32'hba20dabc),
	.w6(32'hb9d705b4),
	.w7(32'hb9c88b44),
	.w8(32'hb98ec079),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d4f3b),
	.w1(32'hb9fded61),
	.w2(32'hba42934d),
	.w3(32'hba5f68ca),
	.w4(32'hba5d9502),
	.w5(32'h3a6916de),
	.w6(32'hba1ee561),
	.w7(32'hba807ac8),
	.w8(32'h3a8deab6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ffbfb),
	.w1(32'h3aceaad9),
	.w2(32'h3a1963c5),
	.w3(32'h398a8575),
	.w4(32'h395e57ef),
	.w5(32'hb999991c),
	.w6(32'h3a00a967),
	.w7(32'h39cfbf30),
	.w8(32'hb9d49bc8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c9263),
	.w1(32'h39c7d14c),
	.w2(32'h39282665),
	.w3(32'hb92de172),
	.w4(32'hb9612244),
	.w5(32'hba194993),
	.w6(32'h3984d6c6),
	.w7(32'h39a3fcb5),
	.w8(32'h386081dc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dea21b),
	.w1(32'h3a9c70f2),
	.w2(32'h3a8ba0fd),
	.w3(32'h3a3d0434),
	.w4(32'h39f93228),
	.w5(32'hb9d73712),
	.w6(32'h3abc8b0f),
	.w7(32'h3a0ea2b0),
	.w8(32'hba910c55),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ee525),
	.w1(32'hba3c8230),
	.w2(32'hba89a9ea),
	.w3(32'hb96f7680),
	.w4(32'hba2fcb87),
	.w5(32'h3aaa03c2),
	.w6(32'hb9bf86c2),
	.w7(32'hba4d3167),
	.w8(32'h3a95f255),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a567a),
	.w1(32'h3ac0a154),
	.w2(32'h3a2c68ee),
	.w3(32'h3a91a276),
	.w4(32'h392a3ad7),
	.w5(32'h3a911682),
	.w6(32'h3ac65a37),
	.w7(32'h3a676568),
	.w8(32'h3a748218),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a690b14),
	.w1(32'h3a6f96d3),
	.w2(32'h3a87da14),
	.w3(32'h3a8cd39d),
	.w4(32'h3a8fefa2),
	.w5(32'hba803a7e),
	.w6(32'h3a6b4e1f),
	.w7(32'h3a855d7f),
	.w8(32'hba870dc8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba764c7d),
	.w1(32'hba9469ee),
	.w2(32'hba9355f8),
	.w3(32'hbaae124b),
	.w4(32'hba93467a),
	.w5(32'hbadfa016),
	.w6(32'hba94b574),
	.w7(32'hbaaeb155),
	.w8(32'hbaac6330),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5212bc),
	.w1(32'hba2d6532),
	.w2(32'hba0f8731),
	.w3(32'hbab5dbf7),
	.w4(32'hba7c9789),
	.w5(32'hba48fd06),
	.w6(32'hba8950aa),
	.w7(32'hba13a6db),
	.w8(32'hb8b77d26),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba312aac),
	.w1(32'h39384854),
	.w2(32'h3a0c9128),
	.w3(32'hb8b8ae8d),
	.w4(32'h39d26193),
	.w5(32'h3a916be6),
	.w6(32'h3a0adba8),
	.w7(32'h3a39c711),
	.w8(32'h39ea45a8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38622325),
	.w1(32'h3a5159d8),
	.w2(32'h3a8be151),
	.w3(32'h3ad8ea31),
	.w4(32'h3ad76158),
	.w5(32'h38451354),
	.w6(32'h3aa9481f),
	.w7(32'h3adb6be5),
	.w8(32'hb9cadcfb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98957fb),
	.w1(32'hba55a886),
	.w2(32'hb90b2a43),
	.w3(32'hba06ba33),
	.w4(32'h37ef968f),
	.w5(32'hb98c5d55),
	.w6(32'hba8cc6e1),
	.w7(32'h37ca205b),
	.w8(32'hb9efc0ed),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391069b8),
	.w1(32'h39d36070),
	.w2(32'h395bf78e),
	.w3(32'hba53d5e7),
	.w4(32'hba65c15f),
	.w5(32'hb9aff8c3),
	.w6(32'hba117b64),
	.w7(32'hb98b5ab4),
	.w8(32'hba769297),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e8a0),
	.w1(32'hba6a5afd),
	.w2(32'hba1808cb),
	.w3(32'hb9307911),
	.w4(32'h39aa0c0a),
	.w5(32'hb98b68f4),
	.w6(32'hba575eb2),
	.w7(32'hb9affc46),
	.w8(32'hba7cc2b0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94830e5),
	.w1(32'h3946e13e),
	.w2(32'hb8b6b4eb),
	.w3(32'hba05d5b5),
	.w4(32'hba0fd478),
	.w5(32'h3900b865),
	.w6(32'hbaa260c5),
	.w7(32'hba5d9f5d),
	.w8(32'h399b574c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c41d3),
	.w1(32'h3b0fa3e8),
	.w2(32'h3ae2cb83),
	.w3(32'h3aa78915),
	.w4(32'h3ae2f068),
	.w5(32'h3a086a5f),
	.w6(32'h3aba88a1),
	.w7(32'h3abd5d15),
	.w8(32'hb89801a1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783b0f4),
	.w1(32'hb8617c94),
	.w2(32'hb95996e8),
	.w3(32'hb9c7f2ea),
	.w4(32'hb9982d74),
	.w5(32'hba306ec2),
	.w6(32'hb9d92a53),
	.w7(32'hb9daf6c6),
	.w8(32'hba19ded2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96e40f),
	.w1(32'hbaca09e2),
	.w2(32'hbab735cc),
	.w3(32'hba571869),
	.w4(32'hba793de2),
	.w5(32'h3973ff77),
	.w6(32'h35f4debf),
	.w7(32'hb988dae7),
	.w8(32'h399020dc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule