module layer_6_featuremap_115(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd61027),
	.w1(32'h3b8b7fbb),
	.w2(32'h3b8dd486),
	.w3(32'hba0d1561),
	.w4(32'h39be8a25),
	.w5(32'h3a2184ef),
	.w6(32'h3b45326e),
	.w7(32'h3b0dbaf4),
	.w8(32'h39980580),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9c8f9),
	.w1(32'h3a72d30d),
	.w2(32'hb92e6e0f),
	.w3(32'hbbe93892),
	.w4(32'hbbfe1938),
	.w5(32'hbbff68b1),
	.w6(32'h3bd62353),
	.w7(32'h3c13b22a),
	.w8(32'h3c1d05ad),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6c3df),
	.w1(32'h3c4af48f),
	.w2(32'hbbc3656e),
	.w3(32'hbc5aa57a),
	.w4(32'hbc074d24),
	.w5(32'h3c01c677),
	.w6(32'hbc4ca9fa),
	.w7(32'hbc9f8974),
	.w8(32'hbb1e36eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7f5d1),
	.w1(32'hbb14d838),
	.w2(32'hbb55d24e),
	.w3(32'hb98b301a),
	.w4(32'h3ad43c14),
	.w5(32'h3abcea2e),
	.w6(32'h3a1a54fe),
	.w7(32'h3ae8b80e),
	.w8(32'h3b2283da),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cdbf1),
	.w1(32'h3d0ad89b),
	.w2(32'h3d613ae1),
	.w3(32'hbce40d34),
	.w4(32'hbd428390),
	.w5(32'hbc1aa2e8),
	.w6(32'h3c1c218c),
	.w7(32'hbd13bfcb),
	.w8(32'hbd323005),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f1106),
	.w1(32'h39d3325a),
	.w2(32'hb8e90ee1),
	.w3(32'hbc38cbbf),
	.w4(32'hbc1170c5),
	.w5(32'hbb8eb849),
	.w6(32'hbbd3000a),
	.w7(32'hbc16a87d),
	.w8(32'hbc0c0720),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2c344),
	.w1(32'hbcded263),
	.w2(32'hbce7903c),
	.w3(32'hbb9ddecf),
	.w4(32'h38964f17),
	.w5(32'hbc074552),
	.w6(32'hbc905467),
	.w7(32'hbb49d530),
	.w8(32'hbb80b8e3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575479),
	.w1(32'h3c55433e),
	.w2(32'hbbf77939),
	.w3(32'hbc495294),
	.w4(32'hbc867de3),
	.w5(32'hbc1ece72),
	.w6(32'hbcdf7357),
	.w7(32'hbd25ad9c),
	.w8(32'hbca05215),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc942b0b),
	.w1(32'h3aec9dcb),
	.w2(32'h3d25dfd9),
	.w3(32'h3bb95a71),
	.w4(32'hbd01b8a8),
	.w5(32'hbd19f947),
	.w6(32'h3ce5cb9f),
	.w7(32'h3d5f5889),
	.w8(32'h3c62bdc7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa18e4),
	.w1(32'h3a3198eb),
	.w2(32'h3b73b1fd),
	.w3(32'hbb9507de),
	.w4(32'hbbd0c6d1),
	.w5(32'hbc197e50),
	.w6(32'h39ed2279),
	.w7(32'hba8324a5),
	.w8(32'hbc119345),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213c7b),
	.w1(32'h3a2afb86),
	.w2(32'hbb3d181f),
	.w3(32'hbbb39794),
	.w4(32'hbb8dd9cf),
	.w5(32'hbc254fe9),
	.w6(32'hbc176c48),
	.w7(32'h3acf9467),
	.w8(32'hbc1143c3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ecb2),
	.w1(32'h3b425488),
	.w2(32'h3c87f7b6),
	.w3(32'h3b9cf50a),
	.w4(32'h3bcf07ae),
	.w5(32'hbbe7a193),
	.w6(32'h3c77aa89),
	.w7(32'h3c5e3837),
	.w8(32'hbb9ff7bd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5283f9),
	.w1(32'hbb2af1ac),
	.w2(32'h3adf2d5f),
	.w3(32'hbb2d5472),
	.w4(32'h3bdb8f8a),
	.w5(32'hbaabac4e),
	.w6(32'hb9323a62),
	.w7(32'h3bd51056),
	.w8(32'hbb005bc8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc244e2a),
	.w1(32'hbc1023a2),
	.w2(32'hbc248b64),
	.w3(32'hbbe7a0ff),
	.w4(32'h3ac1dcca),
	.w5(32'hbc172d1f),
	.w6(32'hbc85e26c),
	.w7(32'h3ba19ede),
	.w8(32'hbcb1f5b5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b4d3d),
	.w1(32'h3b4047d2),
	.w2(32'hbac919e2),
	.w3(32'hbc1a6106),
	.w4(32'hbc32be7f),
	.w5(32'hbc2febb2),
	.w6(32'h3616a1f1),
	.w7(32'hbafa5eb4),
	.w8(32'hbc3437d5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb874c8),
	.w1(32'h3aabaefa),
	.w2(32'h39d7b00a),
	.w3(32'hbb6eab24),
	.w4(32'hbaa6d23b),
	.w5(32'hbb1e5513),
	.w6(32'hba6b24ea),
	.w7(32'hb9a0fc27),
	.w8(32'h3b05b3f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a991d97),
	.w1(32'h3c6ffc36),
	.w2(32'h3c13e6a1),
	.w3(32'h3bda12f5),
	.w4(32'h3b1c2c03),
	.w5(32'h3c013876),
	.w6(32'h3c52ff41),
	.w7(32'hba37318a),
	.w8(32'h3b978e22),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1626),
	.w1(32'h3a701b48),
	.w2(32'h3b68a04e),
	.w3(32'hba8ee2ff),
	.w4(32'hb8ce3e6e),
	.w5(32'hbb74c1cc),
	.w6(32'hbab13dc9),
	.w7(32'h3b3db62b),
	.w8(32'hbaf8e607),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3723ece2),
	.w1(32'hbac6fc5d),
	.w2(32'hbaa3af5c),
	.w3(32'h3a59469d),
	.w4(32'h3ad20f81),
	.w5(32'h3b62f0ef),
	.w6(32'hbb60fc2c),
	.w7(32'hbb958b44),
	.w8(32'hbb0a8d2d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922735),
	.w1(32'hbc00dbb8),
	.w2(32'h3cb4e2a1),
	.w3(32'h3a915889),
	.w4(32'hbb1fd480),
	.w5(32'hbc12df31),
	.w6(32'h3c3c2284),
	.w7(32'h3cb0cd4e),
	.w8(32'h3aaa2dee),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c177d6b),
	.w1(32'hba9983ce),
	.w2(32'hbacee38f),
	.w3(32'h39924bdc),
	.w4(32'hba3eb299),
	.w5(32'hb999b811),
	.w6(32'hba9ae826),
	.w7(32'h3aad0064),
	.w8(32'h3aa55334),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d32f2),
	.w1(32'h3c28dd99),
	.w2(32'h3c5d544f),
	.w3(32'h3c091d9d),
	.w4(32'h3c031d7b),
	.w5(32'h3c36e4d5),
	.w6(32'h3c9232a2),
	.w7(32'h3c7b7edf),
	.w8(32'h3c8a9118),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47aa0f),
	.w1(32'hbb56f25d),
	.w2(32'hbc373a28),
	.w3(32'hbbc20703),
	.w4(32'h3c9c3165),
	.w5(32'h3cc03a42),
	.w6(32'hbccfaf49),
	.w7(32'hbccd76f4),
	.w8(32'hbc826c53),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb87da9),
	.w1(32'hbcc10b66),
	.w2(32'hbc71b439),
	.w3(32'h3d06ad4a),
	.w4(32'h3cfdf2f5),
	.w5(32'h3c092ae9),
	.w6(32'h3cd8f2ea),
	.w7(32'h3d34696d),
	.w8(32'h3cf704fd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45b509),
	.w1(32'h3c24ae25),
	.w2(32'h3cb6c6e3),
	.w3(32'hbc95fc37),
	.w4(32'hbc80a085),
	.w5(32'hbc1e2410),
	.w6(32'h3ca79cea),
	.w7(32'h3c8e7670),
	.w8(32'h3bbb61d2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4bafd),
	.w1(32'hbc556888),
	.w2(32'hbc27be1a),
	.w3(32'hbc3dd765),
	.w4(32'hbc5f0bf9),
	.w5(32'hbc6310b3),
	.w6(32'hbbf4b50d),
	.w7(32'hbbd146f6),
	.w8(32'hbc11167f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946875),
	.w1(32'h3bf900e2),
	.w2(32'h3b998f32),
	.w3(32'h3c15f2d4),
	.w4(32'h3ba88f90),
	.w5(32'h3ba28a23),
	.w6(32'h3be2bd17),
	.w7(32'h3c05f625),
	.w8(32'h3ba83d8d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88c06),
	.w1(32'hbbcb0382),
	.w2(32'hbb871b5e),
	.w3(32'h3b53166b),
	.w4(32'h3bb5c3a1),
	.w5(32'h3a553e21),
	.w6(32'hbb83efba),
	.w7(32'h3b894d58),
	.w8(32'h3ba82d0f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d5d2c),
	.w1(32'hbb8f86c2),
	.w2(32'hbb502630),
	.w3(32'hbafc4050),
	.w4(32'hbb90b597),
	.w5(32'hbbeace53),
	.w6(32'hbb2fdc8b),
	.w7(32'hbb29e906),
	.w8(32'hbb4c1f0e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29cd9d),
	.w1(32'hbc5a6cf9),
	.w2(32'h39ca4155),
	.w3(32'hbb1467d4),
	.w4(32'hbc05978e),
	.w5(32'hbc88b1f8),
	.w6(32'h3c0ea5d5),
	.w7(32'h3ca6a660),
	.w8(32'h3bcd6a8b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c506ed2),
	.w1(32'h3c35ad99),
	.w2(32'hbc2d95d0),
	.w3(32'hbcb10e29),
	.w4(32'hbc0ee979),
	.w5(32'h3cd3549f),
	.w6(32'hbd069215),
	.w7(32'hbd0cd80f),
	.w8(32'h3c0d227e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca60391),
	.w1(32'h3c9f2514),
	.w2(32'h3d01c309),
	.w3(32'hbcee3eda),
	.w4(32'hbcd79222),
	.w5(32'hbc552788),
	.w6(32'h3ad52cf2),
	.w7(32'hbbd1c0fd),
	.w8(32'hbc85b11a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf08890),
	.w1(32'hbaa3e8f3),
	.w2(32'hbbfc1c51),
	.w3(32'h3b33b889),
	.w4(32'h3bd8d174),
	.w5(32'hb9001071),
	.w6(32'h3b7d6b5c),
	.w7(32'h3ca378d6),
	.w8(32'h3c8fd6eb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a6737),
	.w1(32'hbc1629ad),
	.w2(32'hbc62fa74),
	.w3(32'hbbb87c7f),
	.w4(32'hbbce7cbc),
	.w5(32'hbb8d1c68),
	.w6(32'hbc1d6983),
	.w7(32'hbbe6203c),
	.w8(32'hbcaef152),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc726a38),
	.w1(32'h3bf47f23),
	.w2(32'h3a1b25fd),
	.w3(32'hbb349894),
	.w4(32'hbba24af2),
	.w5(32'hbb357f57),
	.w6(32'h3b8b46ee),
	.w7(32'hbb825bb3),
	.w8(32'hbbda2749),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9806f37),
	.w1(32'hbad9058c),
	.w2(32'hbb7160c0),
	.w3(32'h3b94146e),
	.w4(32'h3c776560),
	.w5(32'h3c2a1043),
	.w6(32'hbab251ee),
	.w7(32'hbb056c41),
	.w8(32'h3ac2d646),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb792572),
	.w1(32'h3a6d742d),
	.w2(32'h3b5302e3),
	.w3(32'hbbac9ba6),
	.w4(32'hbb8e88ac),
	.w5(32'hba0974ee),
	.w6(32'hbb9997d3),
	.w7(32'hbbe255a2),
	.w8(32'hbbd7c964),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb875f5f),
	.w1(32'hbbdfb54b),
	.w2(32'hbbd85723),
	.w3(32'hbb8fdeba),
	.w4(32'hbbceb50b),
	.w5(32'hbc206817),
	.w6(32'hba75054f),
	.w7(32'hbb198b7f),
	.w8(32'hbb96eccc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b929),
	.w1(32'hbc0a959a),
	.w2(32'hbc678967),
	.w3(32'hbbcd6057),
	.w4(32'hbc1ed065),
	.w5(32'hbc2b4e50),
	.w6(32'hbc061377),
	.w7(32'hbbe9b074),
	.w8(32'hbbbe4655),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88e3b9),
	.w1(32'h3a20ca65),
	.w2(32'h3ccbc9c3),
	.w3(32'h3c7e981d),
	.w4(32'hbc26b57c),
	.w5(32'hbcfe7e42),
	.w6(32'h3d03cbfb),
	.w7(32'h3cf13378),
	.w8(32'h3c99c458),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c961752),
	.w1(32'h3c382837),
	.w2(32'h3cb88507),
	.w3(32'hbd14c790),
	.w4(32'hbd43e891),
	.w5(32'hbd43e080),
	.w6(32'hbc20edfd),
	.w7(32'hbc8cf2f2),
	.w8(32'hbce15645),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e0581),
	.w1(32'hbbaa977a),
	.w2(32'hbbabe508),
	.w3(32'h3807f101),
	.w4(32'h3b350923),
	.w5(32'h3a3c1e5a),
	.w6(32'hbb7eda93),
	.w7(32'h3a329ffe),
	.w8(32'h3ae9aef2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fcdf4),
	.w1(32'h3b33a89f),
	.w2(32'h3a568e1d),
	.w3(32'h3b0870e2),
	.w4(32'h3bcefc39),
	.w5(32'h3b839559),
	.w6(32'h3b39d599),
	.w7(32'h3ad6a7e3),
	.w8(32'hb9354e3d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a8f4f),
	.w1(32'h3a1f3416),
	.w2(32'hb9faf50d),
	.w3(32'hbaaf0a93),
	.w4(32'h3b704d83),
	.w5(32'h3c010502),
	.w6(32'h3acbb058),
	.w7(32'h393a0d9c),
	.w8(32'h3c08672f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6f2a),
	.w1(32'h3b1ba750),
	.w2(32'h3b06dc99),
	.w3(32'hb9286b08),
	.w4(32'h3a98dbbe),
	.w5(32'hba9f701d),
	.w6(32'h3b007fc7),
	.w7(32'h3b5350f7),
	.w8(32'h3b5e1246),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd413aa),
	.w1(32'hbc4e6ee6),
	.w2(32'hbcdc3472),
	.w3(32'hbc948c43),
	.w4(32'hbc530749),
	.w5(32'hbc8ccce7),
	.w6(32'hbcb60fd7),
	.w7(32'hbca3ea79),
	.w8(32'hbbbc18cf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb10991),
	.w1(32'h3ad5617f),
	.w2(32'hbc2c5c9f),
	.w3(32'hbc2bfdcf),
	.w4(32'hbb82deb8),
	.w5(32'hbc675df0),
	.w6(32'hba9477b1),
	.w7(32'h3bea7be0),
	.w8(32'h3c38cc08),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b120e56),
	.w1(32'hbc3112f4),
	.w2(32'hbc29591c),
	.w3(32'hbc4578b6),
	.w4(32'hbb507e9e),
	.w5(32'hbc4a9888),
	.w6(32'hbca2b11c),
	.w7(32'hbc232884),
	.w8(32'hbc68b4ac),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a539),
	.w1(32'h3b4b839f),
	.w2(32'hbada107a),
	.w3(32'hbad60fdd),
	.w4(32'hba71bd85),
	.w5(32'hb92ddc03),
	.w6(32'hbb1323e6),
	.w7(32'hbb56c7df),
	.w8(32'hbae7650d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cc76a),
	.w1(32'h3ba5a7b0),
	.w2(32'hbcd7a9bf),
	.w3(32'hbbca6fef),
	.w4(32'h3cd006bb),
	.w5(32'h3cf44a07),
	.w6(32'hbcebf3ed),
	.w7(32'hbcd37f29),
	.w8(32'hbbf3c1b0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca59a08),
	.w1(32'hbbe3b24e),
	.w2(32'hbc45f020),
	.w3(32'hbb74a4aa),
	.w4(32'h39d93073),
	.w5(32'hbb9c8a11),
	.w6(32'hbbf84933),
	.w7(32'hbacbd191),
	.w8(32'hbb848d90),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8950),
	.w1(32'hbb94edea),
	.w2(32'hbbdd02b6),
	.w3(32'h3a9d6045),
	.w4(32'hba42db50),
	.w5(32'h38fbbdda),
	.w6(32'hbb7d1ce8),
	.w7(32'hbad85b0a),
	.w8(32'hba45edef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ac9a2),
	.w1(32'hbba08411),
	.w2(32'hbbb263f6),
	.w3(32'h3aeab69c),
	.w4(32'h3b9a6db3),
	.w5(32'h3b5f8c36),
	.w6(32'hbb995e62),
	.w7(32'h3b2acaf0),
	.w8(32'h3c02b30b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a5505),
	.w1(32'hbc6b1f4a),
	.w2(32'hbbf8f021),
	.w3(32'hbb418022),
	.w4(32'h3ae74560),
	.w5(32'hbbe543cd),
	.w6(32'hbb80057f),
	.w7(32'h3c1faa60),
	.w8(32'h3c6e7756),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d7292),
	.w1(32'hbc24fce3),
	.w2(32'hbc4d8e1f),
	.w3(32'hbb4cbcd5),
	.w4(32'hba393341),
	.w5(32'hbbadf35a),
	.w6(32'h3b333b38),
	.w7(32'h3c112eed),
	.w8(32'h3baba6cf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7404e),
	.w1(32'hbc331d99),
	.w2(32'hbc77e413),
	.w3(32'h3cbb527f),
	.w4(32'h3cee66ff),
	.w5(32'h3c133d8c),
	.w6(32'h3c47a0cc),
	.w7(32'hb9f662ea),
	.w8(32'hbc30df33),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6756b),
	.w1(32'hbb7019d0),
	.w2(32'hbb554bc5),
	.w3(32'hbb12dd18),
	.w4(32'hbb65bfdd),
	.w5(32'hbb6583ff),
	.w6(32'hbb165eda),
	.w7(32'hbaf5056d),
	.w8(32'hbb9583ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9700bc),
	.w1(32'h3b98e7c4),
	.w2(32'hbbb19b54),
	.w3(32'h3c40c591),
	.w4(32'h3b52e96e),
	.w5(32'hba6025c2),
	.w6(32'h3c1a2b45),
	.w7(32'h3bc3d6f5),
	.w8(32'h3a1ccbb7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08827),
	.w1(32'h3b472983),
	.w2(32'h3b5e001a),
	.w3(32'h3b7ad227),
	.w4(32'h3b44c668),
	.w5(32'h3a7c9d53),
	.w6(32'h3b8f1bc8),
	.w7(32'h3b721387),
	.w8(32'h3b3592da),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97b172),
	.w1(32'hbba57a11),
	.w2(32'h3c615d45),
	.w3(32'h3c18efcb),
	.w4(32'h3a5c90a1),
	.w5(32'hbca61eb1),
	.w6(32'hbc285797),
	.w7(32'hbbd24b1d),
	.w8(32'hbc45d46c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6292ff),
	.w1(32'hbb748c4b),
	.w2(32'hbc80d456),
	.w3(32'h3ba00d1f),
	.w4(32'hbba768a7),
	.w5(32'hbc67b6ad),
	.w6(32'hbb69064e),
	.w7(32'hbbf7488d),
	.w8(32'hbc78883b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6d97),
	.w1(32'h3c9dc124),
	.w2(32'h3c6b41c7),
	.w3(32'h3bb4f840),
	.w4(32'hbb898142),
	.w5(32'h3c427279),
	.w6(32'h3c6f743f),
	.w7(32'h3bc8e540),
	.w8(32'h3c16a26c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51f2f1),
	.w1(32'h3c886305),
	.w2(32'h3cd9c32a),
	.w3(32'hb95ade32),
	.w4(32'h3be8745f),
	.w5(32'h3c753712),
	.w6(32'h3ce2eeea),
	.w7(32'h3d21bdaf),
	.w8(32'h3c9390b3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf613c0),
	.w1(32'hb8ee3a82),
	.w2(32'hba8710cf),
	.w3(32'h3bba72c1),
	.w4(32'h3c299be3),
	.w5(32'h3c159372),
	.w6(32'h3aa232c8),
	.w7(32'h3b5e9e2a),
	.w8(32'h3b8cf1b3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule