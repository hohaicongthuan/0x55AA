module layer_8_featuremap_180(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56fca8),
	.w1(32'h3c2f31da),
	.w2(32'h3ce7986c),
	.w3(32'hb9e3448c),
	.w4(32'h3bdb44f0),
	.w5(32'h3c9d1d35),
	.w6(32'h3ba081fb),
	.w7(32'h3afec374),
	.w8(32'h3bb58160),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b2f9),
	.w1(32'hbb69e9f6),
	.w2(32'hbb4c4e5a),
	.w3(32'hbb3abad0),
	.w4(32'h3a1686d4),
	.w5(32'hbb07db1a),
	.w6(32'hba426c8b),
	.w7(32'hbab0e560),
	.w8(32'h3b948052),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b958),
	.w1(32'hbcafaead),
	.w2(32'hbc2ce3f1),
	.w3(32'hba22f48a),
	.w4(32'hbadcb357),
	.w5(32'hbbd5879d),
	.w6(32'hbc0f7244),
	.w7(32'hbc89b68e),
	.w8(32'hbc1bcaaa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b857822),
	.w1(32'hbbffd89a),
	.w2(32'hbb871078),
	.w3(32'hb982fe8c),
	.w4(32'hbc6641f2),
	.w5(32'h3b564c61),
	.w6(32'h3aebb2bd),
	.w7(32'hbc236eee),
	.w8(32'hbcb66a0c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c14e),
	.w1(32'h3a7608ee),
	.w2(32'h386175b9),
	.w3(32'h3bd0392f),
	.w4(32'hbb13a5ee),
	.w5(32'hba37fe59),
	.w6(32'hba0efbfc),
	.w7(32'h3a1c4370),
	.w8(32'hbb980c3f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ffcd8),
	.w1(32'hbbfe728f),
	.w2(32'h3b69592b),
	.w3(32'h3bc79f2c),
	.w4(32'hbb269ff6),
	.w5(32'h3c2d9705),
	.w6(32'hbc91841f),
	.w7(32'hbc96a39a),
	.w8(32'h3c13a064),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc51655),
	.w1(32'h3b06d9de),
	.w2(32'hbb0abec1),
	.w3(32'hbb9aa64d),
	.w4(32'hbb957803),
	.w5(32'hbb84237b),
	.w6(32'h3af9508a),
	.w7(32'h39a993e5),
	.w8(32'hbbb28bed),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdf4e8),
	.w1(32'h3c4d17b6),
	.w2(32'h3a436e49),
	.w3(32'h3ac62be1),
	.w4(32'h3ad43f7f),
	.w5(32'hbc3fd106),
	.w6(32'h3a2d74ac),
	.w7(32'h3b1a7be2),
	.w8(32'hbb9b16b4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2589),
	.w1(32'hbb50ee77),
	.w2(32'hbbe6e6fb),
	.w3(32'hbb351d52),
	.w4(32'hbbd3e9f1),
	.w5(32'hbb232606),
	.w6(32'h3a973a0a),
	.w7(32'hbaa2cdd9),
	.w8(32'hbc170b3b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb468b43),
	.w1(32'h3ca08a65),
	.w2(32'h3c9996fa),
	.w3(32'h3c878f9b),
	.w4(32'h3c50146f),
	.w5(32'h3c2637f1),
	.w6(32'h3b2faab8),
	.w7(32'h3c1f194d),
	.w8(32'h3a9f53dd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc036f3),
	.w1(32'h387bdd2b),
	.w2(32'hbc94e1b4),
	.w3(32'hbc15d21f),
	.w4(32'hbb3b9c36),
	.w5(32'hbc2bf2cf),
	.w6(32'h3b7cf3f2),
	.w7(32'hbc100fbf),
	.w8(32'h3bca9cea),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6315),
	.w1(32'h3bc49731),
	.w2(32'h3c17eab6),
	.w3(32'hbba3cdad),
	.w4(32'hb8bdabad),
	.w5(32'hbaa058a9),
	.w6(32'hba32b5d4),
	.w7(32'hbb0eede5),
	.w8(32'h3ba8d4c0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a205c9b),
	.w1(32'hbb2a3f8e),
	.w2(32'h3b943c49),
	.w3(32'hbca93dfa),
	.w4(32'hbbc1bd74),
	.w5(32'hbb7aee95),
	.w6(32'hba2c1c8d),
	.w7(32'hb7fb91a4),
	.w8(32'hbc845d57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e19c7),
	.w1(32'h3bb0271f),
	.w2(32'h38c60eef),
	.w3(32'hbb421205),
	.w4(32'h3b460606),
	.w5(32'h3bfbdf3e),
	.w6(32'hbc14e153),
	.w7(32'h3ae543c8),
	.w8(32'h3c2ebc15),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1dccf),
	.w1(32'h3b417193),
	.w2(32'hbb7a276f),
	.w3(32'hbac5bf52),
	.w4(32'hbb9b3e2c),
	.w5(32'hbb846b6f),
	.w6(32'h3b682cb9),
	.w7(32'h3a9a63b5),
	.w8(32'hbbbd0d4c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a461),
	.w1(32'hbc2080eb),
	.w2(32'hbba7373b),
	.w3(32'h3b526260),
	.w4(32'hbac571f8),
	.w5(32'h3b73453f),
	.w6(32'hbbbd50b6),
	.w7(32'hbc8d4ea5),
	.w8(32'h3b4b5ca9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2959c),
	.w1(32'hbaba139a),
	.w2(32'hba3a7af4),
	.w3(32'hbb564685),
	.w4(32'hbb3efd48),
	.w5(32'hbb340227),
	.w6(32'hbb893ced),
	.w7(32'hbb75932c),
	.w8(32'hbbbc68b7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73c2e),
	.w1(32'hbb830483),
	.w2(32'hbbe374c3),
	.w3(32'hba62a1ab),
	.w4(32'hbb94657b),
	.w5(32'h3a0432b6),
	.w6(32'hbb3df1ff),
	.w7(32'hbb958d52),
	.w8(32'h3c373c1f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98329b),
	.w1(32'hbb975b9d),
	.w2(32'h3c5e4739),
	.w3(32'hbc0b4695),
	.w4(32'h3beda737),
	.w5(32'h3d0c53ab),
	.w6(32'hbca89635),
	.w7(32'hbd3f8aa0),
	.w8(32'hbbf3fa15),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb6c9a),
	.w1(32'h3be513df),
	.w2(32'h3c17b6b2),
	.w3(32'hbb370202),
	.w4(32'hbb9953a0),
	.w5(32'hbb240f26),
	.w6(32'h3b5c666a),
	.w7(32'h3b534a63),
	.w8(32'h3969128a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810af2),
	.w1(32'h3b680262),
	.w2(32'h3b99dc94),
	.w3(32'hbaa085cd),
	.w4(32'hbb43e625),
	.w5(32'hbb8ce0a5),
	.w6(32'hbb2586b3),
	.w7(32'hbb822ef5),
	.w8(32'hbc36d437),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac914),
	.w1(32'hbc34c917),
	.w2(32'hbba0afc2),
	.w3(32'h3c08c080),
	.w4(32'hbb333cc0),
	.w5(32'h3bc09f4a),
	.w6(32'hbb83b491),
	.w7(32'h3b88d12e),
	.w8(32'h3c9f823f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b622b),
	.w1(32'h3b2e08cd),
	.w2(32'h3d5aa922),
	.w3(32'hbc6dee28),
	.w4(32'h3ca15076),
	.w5(32'h3d240453),
	.w6(32'hbbe7946e),
	.w7(32'hbbb2228d),
	.w8(32'h3d10a242),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa5ffd),
	.w1(32'hbb181a8d),
	.w2(32'h3a5eb054),
	.w3(32'hbc47f659),
	.w4(32'hbb96d5f1),
	.w5(32'hbc0b1252),
	.w6(32'hbbf95406),
	.w7(32'hbc4056dc),
	.w8(32'h3bd82331),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fcd20),
	.w1(32'hbc0affc2),
	.w2(32'h3c3b7474),
	.w3(32'hbbf3a513),
	.w4(32'h3b9686f0),
	.w5(32'h3bcde73f),
	.w6(32'hbc5ab7a2),
	.w7(32'hbc6aab0b),
	.w8(32'h3bb87d24),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74ad11),
	.w1(32'h3b11f260),
	.w2(32'hbc1d9f54),
	.w3(32'h3b9d3edf),
	.w4(32'hbb310140),
	.w5(32'h39ae357e),
	.w6(32'h39676cc2),
	.w7(32'hba52b8cd),
	.w8(32'hb9e78e4f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19eebb),
	.w1(32'hbcd47e8c),
	.w2(32'hbca95734),
	.w3(32'h3a5fa179),
	.w4(32'hbc3b7e6e),
	.w5(32'hbb1030d2),
	.w6(32'hbc155f7f),
	.w7(32'hbcbb454a),
	.w8(32'hbb1505ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed801c),
	.w1(32'hbc981691),
	.w2(32'h3d78527e),
	.w3(32'hbd1be918),
	.w4(32'hbd07759d),
	.w5(32'h3ca79255),
	.w6(32'h3d315c22),
	.w7(32'hbbfb65eb),
	.w8(32'hbd2fac32),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc6ad),
	.w1(32'h3bcb2cae),
	.w2(32'h3c118dbc),
	.w3(32'h3b8dac15),
	.w4(32'h3b41df33),
	.w5(32'hbc1fc406),
	.w6(32'hb6c2931a),
	.w7(32'h3c0b034e),
	.w8(32'h3a97c7bd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd044),
	.w1(32'hbaf1d181),
	.w2(32'hb9a7b7ca),
	.w3(32'hbca70fba),
	.w4(32'h3c26f800),
	.w5(32'h3c1c059c),
	.w6(32'hbace590f),
	.w7(32'h3b4a7515),
	.w8(32'h3be39569),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd025b),
	.w1(32'h3c0687eb),
	.w2(32'h3c2d7346),
	.w3(32'h3c886be3),
	.w4(32'h3b54a756),
	.w5(32'hbc034167),
	.w6(32'hba983b20),
	.w7(32'h3bcda1a5),
	.w8(32'h3a114420),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc846a82),
	.w1(32'hbb5c4a65),
	.w2(32'hbc8dc2de),
	.w3(32'hbc8cddbd),
	.w4(32'h3ba0b4e2),
	.w5(32'hbb87564e),
	.w6(32'h3905e063),
	.w7(32'hbc30b18a),
	.w8(32'h3b7ab518),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037eeb),
	.w1(32'hbb75ca55),
	.w2(32'hba909739),
	.w3(32'hbb062d68),
	.w4(32'hb82e07a9),
	.w5(32'hbbe5911f),
	.w6(32'h3af9da57),
	.w7(32'h3b432d3c),
	.w8(32'h3c66d7fb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f1c13),
	.w1(32'hbc203c08),
	.w2(32'hbbcc94a7),
	.w3(32'hbc682d3b),
	.w4(32'hbaf9b0fc),
	.w5(32'hbc31d6d0),
	.w6(32'hbb1367ee),
	.w7(32'hba340fdb),
	.w8(32'hbb63b6f1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cf066),
	.w1(32'h3c89c194),
	.w2(32'h3c3403f8),
	.w3(32'hbb9def8a),
	.w4(32'h3bcc2439),
	.w5(32'hbadb0aa0),
	.w6(32'h3c8032f3),
	.w7(32'h3c96002a),
	.w8(32'h3c1cd6bc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca99b78),
	.w1(32'h3ba22940),
	.w2(32'h3c00da3f),
	.w3(32'hbc966651),
	.w4(32'h3b4814a0),
	.w5(32'h3b8c98b4),
	.w6(32'h398c069f),
	.w7(32'hbbaa7aa1),
	.w8(32'h3b380996),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39af0),
	.w1(32'hbb9999e8),
	.w2(32'h3bad22f8),
	.w3(32'hbb7b07d7),
	.w4(32'hbc1de520),
	.w5(32'hbba29431),
	.w6(32'h39cf6930),
	.w7(32'h3c0679b6),
	.w8(32'h3c06b8ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c126224),
	.w1(32'h39ba5079),
	.w2(32'hbb62ca14),
	.w3(32'h393068e8),
	.w4(32'hbbc8c8d2),
	.w5(32'hbbbde99d),
	.w6(32'h3b10cc1f),
	.w7(32'h3aaefe58),
	.w8(32'hbc12c116),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6943a),
	.w1(32'h39107421),
	.w2(32'hbb9d94b6),
	.w3(32'h3bb2b3db),
	.w4(32'hbb6e25aa),
	.w5(32'hba9c473d),
	.w6(32'h38c9bd1a),
	.w7(32'hbbc52028),
	.w8(32'h3bf8da4d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd84cb8),
	.w1(32'hb994adef),
	.w2(32'hbba17efa),
	.w3(32'hbaaf64d9),
	.w4(32'hbb106097),
	.w5(32'hbb993c16),
	.w6(32'hbbc1de30),
	.w7(32'hbbbfeb3d),
	.w8(32'hba9f15ec),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d968),
	.w1(32'h3cabeec2),
	.w2(32'h3ce9bb50),
	.w3(32'h3c461566),
	.w4(32'h3c6af8c2),
	.w5(32'h3cc480cb),
	.w6(32'h3c126c80),
	.w7(32'h3b89246a),
	.w8(32'hbb2f493f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeafee2),
	.w1(32'hbc6de438),
	.w2(32'hbae625d2),
	.w3(32'hb9da60e3),
	.w4(32'hbb27dc39),
	.w5(32'h3c423674),
	.w6(32'hbbf297b6),
	.w7(32'hbc93ba0b),
	.w8(32'h3b09f617),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03dd7f),
	.w1(32'hbb86b76c),
	.w2(32'h3bd1136a),
	.w3(32'h3b844669),
	.w4(32'hbb3ea9e1),
	.w5(32'hbc27b84a),
	.w6(32'hbab83ad3),
	.w7(32'h3c01feaf),
	.w8(32'h3ca1986b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ed3d7),
	.w1(32'hbaf7b74a),
	.w2(32'h3b29aa40),
	.w3(32'hbbec2594),
	.w4(32'h3bd94bac),
	.w5(32'h3bb88370),
	.w6(32'hbc16b55a),
	.w7(32'h3b051d6d),
	.w8(32'h3c397649),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd03885),
	.w1(32'hbb841af4),
	.w2(32'hbb137ea3),
	.w3(32'hbc308647),
	.w4(32'h3b499754),
	.w5(32'h3bd54895),
	.w6(32'hbc01d3ea),
	.w7(32'hbc25713c),
	.w8(32'hbb828cf6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f1e5e),
	.w1(32'hbb8530a2),
	.w2(32'hbbac2a8e),
	.w3(32'hbc267952),
	.w4(32'hbb17eb7b),
	.w5(32'h36e73c90),
	.w6(32'h3a292694),
	.w7(32'hbadf82b9),
	.w8(32'h3b6233e4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaea3eb),
	.w1(32'hbc2190e1),
	.w2(32'hbba895a2),
	.w3(32'h3af3b192),
	.w4(32'hbb15a2d2),
	.w5(32'hbbbe9bfb),
	.w6(32'hbc2f802b),
	.w7(32'hbbfedf23),
	.w8(32'hbb8a040d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc828795),
	.w1(32'hbc2feaac),
	.w2(32'hbb96cc2c),
	.w3(32'hbc0f273f),
	.w4(32'hbba46a6c),
	.w5(32'hbb3f5e48),
	.w6(32'hbbd8d6c1),
	.w7(32'hbc33eb55),
	.w8(32'h3b4f2bd3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07471f),
	.w1(32'hbb803553),
	.w2(32'h3c316a3d),
	.w3(32'hbb7f00f0),
	.w4(32'h3afac2ac),
	.w5(32'h3ad0d5ea),
	.w6(32'h3a8aed6f),
	.w7(32'hbb4be5c9),
	.w8(32'h3be85178),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f1348),
	.w1(32'hbb9551d9),
	.w2(32'h3b9a4d61),
	.w3(32'hbbe175b0),
	.w4(32'h3b909f76),
	.w5(32'h3c066a4b),
	.w6(32'h3af7fd95),
	.w7(32'h3955c451),
	.w8(32'hbb9241da),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46d6dd),
	.w1(32'h3b1a2c69),
	.w2(32'h3bb7cc9f),
	.w3(32'h3c7fdb95),
	.w4(32'h39b5578b),
	.w5(32'h3bab9d41),
	.w6(32'h3bbc929c),
	.w7(32'h3baf8370),
	.w8(32'hbad977b9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67d738),
	.w1(32'hba40ebfe),
	.w2(32'h3bd39aac),
	.w3(32'h3a7b9846),
	.w4(32'h3cd920d0),
	.w5(32'h3d2297e2),
	.w6(32'hbc21c57d),
	.w7(32'hbc9f1b59),
	.w8(32'hbbac0a9d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75d23),
	.w1(32'h3b556068),
	.w2(32'hbb27316a),
	.w3(32'h3c704397),
	.w4(32'h3afac651),
	.w5(32'hb984dd68),
	.w6(32'hbaf94542),
	.w7(32'hb81625a4),
	.w8(32'hbb534be0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb97c4),
	.w1(32'h3c869f3a),
	.w2(32'h3c1d525a),
	.w3(32'h3b82c8a9),
	.w4(32'h3c1e01ac),
	.w5(32'hbabf65a5),
	.w6(32'hba1a7615),
	.w7(32'h3c41d9e4),
	.w8(32'h3b460dcd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adedd47),
	.w1(32'hbc3739a7),
	.w2(32'h3a295631),
	.w3(32'hbbd98cc5),
	.w4(32'hbb63bc82),
	.w5(32'hbbbc22bd),
	.w6(32'hbb9e0d23),
	.w7(32'hbb51efa5),
	.w8(32'h3c28a6c5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2ce5),
	.w1(32'h3b62a400),
	.w2(32'h3ca40990),
	.w3(32'hbbf2e018),
	.w4(32'h3c4e4406),
	.w5(32'h3c8a565f),
	.w6(32'h3c57b1ff),
	.w7(32'h3c893460),
	.w8(32'h3c91ae25),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc6518),
	.w1(32'h3c817fff),
	.w2(32'h3ad5d654),
	.w3(32'h39047db0),
	.w4(32'h3a4549ea),
	.w5(32'hbd274437),
	.w6(32'hbb3f8cf6),
	.w7(32'h3cea17cf),
	.w8(32'h3cc5f98a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9eb46),
	.w1(32'hbae02ace),
	.w2(32'h3b961e2b),
	.w3(32'hbce311c3),
	.w4(32'hbb1dbb35),
	.w5(32'hbb8ed482),
	.w6(32'h3bbcdfc6),
	.w7(32'h3c340b5a),
	.w8(32'h3c359530),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02bd70),
	.w1(32'hb9d2e789),
	.w2(32'h3b09b5d9),
	.w3(32'hbc3f23be),
	.w4(32'h3b887df6),
	.w5(32'h3b2bb7ba),
	.w6(32'hbb4b5d6d),
	.w7(32'hbaf362a4),
	.w8(32'h3bbbeba2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0bba2),
	.w1(32'hbb59d987),
	.w2(32'h3c3c0f75),
	.w3(32'hbb824b07),
	.w4(32'h3bdbf6ae),
	.w5(32'h3b803458),
	.w6(32'hbbf28de5),
	.w7(32'h3b1208c3),
	.w8(32'h3c400378),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d667),
	.w1(32'hbc7730fe),
	.w2(32'hba99f749),
	.w3(32'hbbd6318c),
	.w4(32'hbb98237a),
	.w5(32'h392765a9),
	.w6(32'hbc803b18),
	.w7(32'hbc8a07db),
	.w8(32'h3ab4515f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c224096),
	.w1(32'hbc86234b),
	.w2(32'hbb8bd1b8),
	.w3(32'h3b9db471),
	.w4(32'hbc7ff554),
	.w5(32'h3ba0d299),
	.w6(32'h3bd905c5),
	.w7(32'h3a8c022d),
	.w8(32'h3b94f6a2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d5da3),
	.w1(32'h3c8d6485),
	.w2(32'h3c8e6b7a),
	.w3(32'h3d03cd1d),
	.w4(32'h3c3a297d),
	.w5(32'h3c92a993),
	.w6(32'h3b786588),
	.w7(32'hbad19752),
	.w8(32'hbba53f4d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387b25ad),
	.w1(32'h3bba3191),
	.w2(32'h3c215ff5),
	.w3(32'h3b868da2),
	.w4(32'h3c128681),
	.w5(32'h3c0b0f79),
	.w6(32'h3a1beae4),
	.w7(32'h3c216803),
	.w8(32'h3c50b495),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c035c86),
	.w1(32'h3b10e5ec),
	.w2(32'h3b8cc9b1),
	.w3(32'h3af006af),
	.w4(32'h3b9e72ce),
	.w5(32'h3baea728),
	.w6(32'h39fd6fb9),
	.w7(32'h3b8bb3d6),
	.w8(32'h3c227e6a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133dcc),
	.w1(32'hbbef491e),
	.w2(32'hbba4e4ac),
	.w3(32'hbbf96c65),
	.w4(32'hbbff8eb4),
	.w5(32'h3b04d220),
	.w6(32'hbb4b7ce9),
	.w7(32'hbb2ab132),
	.w8(32'hbb8608c6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0e462),
	.w1(32'hbc5196cb),
	.w2(32'h3b8342c1),
	.w3(32'hbbd853f9),
	.w4(32'h3c0fa0cd),
	.w5(32'h3c605f90),
	.w6(32'hbc276720),
	.w7(32'hbba993c4),
	.w8(32'h3c5ff730),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4bd21),
	.w1(32'h3b215daf),
	.w2(32'h3bc6d87b),
	.w3(32'hbbc50fd1),
	.w4(32'h3b2c752e),
	.w5(32'h3c012999),
	.w6(32'hbaa4cf08),
	.w7(32'h3aa10297),
	.w8(32'hbb99568f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d5baa),
	.w1(32'hbc5f2050),
	.w2(32'hbbaf8971),
	.w3(32'h3c81caf7),
	.w4(32'hbbc2f985),
	.w5(32'hbbb01c43),
	.w6(32'hbc29793d),
	.w7(32'hbc09d772),
	.w8(32'h3a5640ee),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c8a6),
	.w1(32'hbc80cbb1),
	.w2(32'hbb4cd937),
	.w3(32'hbc4009c3),
	.w4(32'hbb68cb4c),
	.w5(32'h3c8c54e1),
	.w6(32'hbc3969d1),
	.w7(32'h3a37985f),
	.w8(32'h3c106ca4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c832389),
	.w1(32'h3b482dfc),
	.w2(32'hbc4d4d17),
	.w3(32'h3be81320),
	.w4(32'h3b9f766c),
	.w5(32'h3c4df9d3),
	.w6(32'h3bb58e1a),
	.w7(32'hbcd70885),
	.w8(32'hbcd411e6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be87d),
	.w1(32'h3bed2cd7),
	.w2(32'h3ba3421d),
	.w3(32'h3ca39483),
	.w4(32'h3bdc1ccf),
	.w5(32'h3aa490b4),
	.w6(32'h3a41a09b),
	.w7(32'h3be4d19a),
	.w8(32'h3bb4f71e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf350),
	.w1(32'hba8f5645),
	.w2(32'h3bdf7eec),
	.w3(32'hbc033d78),
	.w4(32'h3b10d3ad),
	.w5(32'hb98322b8),
	.w6(32'hbc191446),
	.w7(32'hbb9a3b4f),
	.w8(32'h3b456fb3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33d20c),
	.w1(32'h3c6ff721),
	.w2(32'h3c84bfcf),
	.w3(32'h39e1a215),
	.w4(32'h3ba9c2b6),
	.w5(32'h3a9405cd),
	.w6(32'h3c338d46),
	.w7(32'h3c2f36da),
	.w8(32'h3af6b994),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f3c8b),
	.w1(32'hbc8dd7f6),
	.w2(32'hbb38edef),
	.w3(32'hbbf5ca7c),
	.w4(32'hbbd2dd49),
	.w5(32'h3b8c4f1e),
	.w6(32'hbc6dca8a),
	.w7(32'hbcce2a17),
	.w8(32'hbaaeb293),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c429521),
	.w1(32'h3bb158fd),
	.w2(32'h3b054402),
	.w3(32'h3c607621),
	.w4(32'h3bae78ef),
	.w5(32'h3bcedb2e),
	.w6(32'hbaa4ba4b),
	.w7(32'hbbc6d22e),
	.w8(32'hbae0719b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d3635),
	.w1(32'h3be8eb96),
	.w2(32'h3b63ed9c),
	.w3(32'hbb0817c9),
	.w4(32'hbb3ac813),
	.w5(32'hbc867135),
	.w6(32'h3b042ca3),
	.w7(32'h3b670c89),
	.w8(32'h3bc30c83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fb2e3),
	.w1(32'h3aa75678),
	.w2(32'h3c54f9f1),
	.w3(32'hbcc4d810),
	.w4(32'hbb0bdd59),
	.w5(32'hb8cbefe0),
	.w6(32'h3b8ab795),
	.w7(32'h3b96b240),
	.w8(32'h3a91dca0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2526fe),
	.w1(32'hbae7e52e),
	.w2(32'h3c517eba),
	.w3(32'hbb9f16b0),
	.w4(32'h3c3dcb1a),
	.w5(32'h3ca0b10b),
	.w6(32'hbb83caab),
	.w7(32'hbc964033),
	.w8(32'hbcc2728f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cd32d),
	.w1(32'h3bb820c1),
	.w2(32'hba7c79be),
	.w3(32'h3adfdab2),
	.w4(32'h3b561c39),
	.w5(32'h3b49a5cb),
	.w6(32'h3bafa549),
	.w7(32'h3be49d60),
	.w8(32'h3bc4e595),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4927ed),
	.w1(32'hbb0e2674),
	.w2(32'hbc175e99),
	.w3(32'h3b4a575a),
	.w4(32'hbb4e599d),
	.w5(32'hbb7fbb79),
	.w6(32'hbc322c22),
	.w7(32'hbbb7385b),
	.w8(32'h3a9ffaa9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19591a),
	.w1(32'hbc123e23),
	.w2(32'hbc198ee5),
	.w3(32'hbbffc063),
	.w4(32'hbae44bbd),
	.w5(32'hbb502c85),
	.w6(32'hbb7e10f8),
	.w7(32'hbbdfa85e),
	.w8(32'h3aa9a0a5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd416b),
	.w1(32'hbc52e319),
	.w2(32'hbb849708),
	.w3(32'hbc1d895a),
	.w4(32'hbbb4a3b0),
	.w5(32'h3be643b4),
	.w6(32'hbc786c69),
	.w7(32'hbc27104c),
	.w8(32'h3bcfba60),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf61732),
	.w1(32'h3c881a2d),
	.w2(32'h3c6e9dd8),
	.w3(32'h3d0b46df),
	.w4(32'h3c3a5fbc),
	.w5(32'h3c172026),
	.w6(32'h3c4511ac),
	.w7(32'hbb959a06),
	.w8(32'h3b75ea53),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6bc1f),
	.w1(32'h3ae7471e),
	.w2(32'h3b4dcc49),
	.w3(32'hbbca57e1),
	.w4(32'h3abacbbc),
	.w5(32'hbba41efb),
	.w6(32'hbc02948c),
	.w7(32'hbc991435),
	.w8(32'hbc01a821),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42deae),
	.w1(32'h3cb92657),
	.w2(32'h3d129f3d),
	.w3(32'hbbe82d12),
	.w4(32'h3c6fa5ff),
	.w5(32'h3d07b099),
	.w6(32'h3b89861d),
	.w7(32'h3c8188dd),
	.w8(32'h3caf9f27),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab50fc),
	.w1(32'h3c7dde38),
	.w2(32'h3a100d94),
	.w3(32'h3b9769cc),
	.w4(32'h3c6b2130),
	.w5(32'h3be54f11),
	.w6(32'h3c0b2b88),
	.w7(32'h3add2d59),
	.w8(32'hbc47fe94),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cc706),
	.w1(32'hbc6a9228),
	.w2(32'h3b8d307c),
	.w3(32'hbb14cf0f),
	.w4(32'hbba4d339),
	.w5(32'h3b8e1af2),
	.w6(32'hbb9f0e21),
	.w7(32'h3a579153),
	.w8(32'h3c20d1fa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93d5fe),
	.w1(32'h3c736370),
	.w2(32'h3b00b887),
	.w3(32'h3bf32b14),
	.w4(32'h3c104af5),
	.w5(32'hbabb2fdf),
	.w6(32'h3a622a49),
	.w7(32'h39b86516),
	.w8(32'hbc161bed),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc975e3e),
	.w1(32'hbc26a73b),
	.w2(32'hbaf6969d),
	.w3(32'hbc5eeee2),
	.w4(32'hbc1362b4),
	.w5(32'hbba443e5),
	.w6(32'hbc700859),
	.w7(32'hbc189dfb),
	.w8(32'hbbb6cadc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d93be),
	.w1(32'h3c2ab60b),
	.w2(32'h3bb8dfcd),
	.w3(32'hbc19eb9f),
	.w4(32'h3bb0ab4d),
	.w5(32'hbae3b8d8),
	.w6(32'hb99839b4),
	.w7(32'h3b63b489),
	.w8(32'h3b6f4f97),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39bb8e),
	.w1(32'hb88c43a0),
	.w2(32'h3b64ea82),
	.w3(32'h3adbdef9),
	.w4(32'hbb0c7d46),
	.w5(32'hbc1c5be4),
	.w6(32'hbc0282f8),
	.w7(32'hbae0e927),
	.w8(32'hbb1efea9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c7f6),
	.w1(32'hbaac9363),
	.w2(32'hbb911907),
	.w3(32'h3a7cc32e),
	.w4(32'hbac175fc),
	.w5(32'hbbbeda8b),
	.w6(32'h3a29904a),
	.w7(32'hbab860f8),
	.w8(32'hbb0beca6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910e43),
	.w1(32'hbb9c6a6f),
	.w2(32'h3ac9b597),
	.w3(32'hbc10243f),
	.w4(32'hbab368cf),
	.w5(32'h391fe107),
	.w6(32'hbbd73cc2),
	.w7(32'hbbc45e0c),
	.w8(32'h3b751d6f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6cced),
	.w1(32'h3be5c12a),
	.w2(32'h3c5f985c),
	.w3(32'hbbe04899),
	.w4(32'hba5f1863),
	.w5(32'hbb58fb6a),
	.w6(32'h3c04c8d2),
	.w7(32'h3c04aaff),
	.w8(32'h3c293dae),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cfa8c),
	.w1(32'h3c051d97),
	.w2(32'hbaabf8b7),
	.w3(32'hbc8448e7),
	.w4(32'hb9331002),
	.w5(32'hbc28210a),
	.w6(32'h3c0010b6),
	.w7(32'h3bf70f38),
	.w8(32'hbb627190),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d863),
	.w1(32'h3bca66c2),
	.w2(32'hb9920b0c),
	.w3(32'hbc5d94c5),
	.w4(32'hbbd330bb),
	.w5(32'hbc3329a4),
	.w6(32'hbc15887f),
	.w7(32'h3b653d4e),
	.w8(32'h3abc3792),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e88863),
	.w1(32'hbc2b58e4),
	.w2(32'hbafe9316),
	.w3(32'hbc589469),
	.w4(32'hbb4a4671),
	.w5(32'hbaf76486),
	.w6(32'hbb03b7a0),
	.w7(32'h3b3d8bb0),
	.w8(32'hb9ab0038),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd2bcd),
	.w1(32'hbb46530d),
	.w2(32'h3a6031f4),
	.w3(32'hbbd804f7),
	.w4(32'hbbd63341),
	.w5(32'hbbf46b7f),
	.w6(32'hbb9f8e9d),
	.w7(32'h3bead870),
	.w8(32'h3bafe110),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb945),
	.w1(32'h395ff062),
	.w2(32'h3ce49587),
	.w3(32'hbc31e571),
	.w4(32'h3a883727),
	.w5(32'hbb4e4089),
	.w6(32'hbc976300),
	.w7(32'h3cb7b2c7),
	.w8(32'h3d1b9a5d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0750b),
	.w1(32'hba8f9afa),
	.w2(32'h3b0e7e71),
	.w3(32'hbc700008),
	.w4(32'h3bf95353),
	.w5(32'h3b29ec23),
	.w6(32'hbb620db3),
	.w7(32'hbb86ea6d),
	.w8(32'hbb809312),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd1b71),
	.w1(32'h3b2d593a),
	.w2(32'hbc0286be),
	.w3(32'hb97a373a),
	.w4(32'h3b05aaf4),
	.w5(32'hbb84b8af),
	.w6(32'h3bcec31f),
	.w7(32'h3adbda3f),
	.w8(32'hbbdb5ef2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98883c),
	.w1(32'h3b8500e1),
	.w2(32'hba88c66b),
	.w3(32'h3bee646c),
	.w4(32'h3bcfb32c),
	.w5(32'h3b8790d6),
	.w6(32'h3aa0af81),
	.w7(32'hbb708068),
	.w8(32'h3b58603d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a62d8a),
	.w1(32'h3c915f10),
	.w2(32'hbca637da),
	.w3(32'hbc27321c),
	.w4(32'hbc0131e5),
	.w5(32'hbc194a00),
	.w6(32'h3bc4c049),
	.w7(32'h3b9d969c),
	.w8(32'hbb8dff38),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a008),
	.w1(32'hbbb6a193),
	.w2(32'hbbc7c47b),
	.w3(32'h3c732e21),
	.w4(32'hba95e770),
	.w5(32'h3b41f7bd),
	.w6(32'h3aba6b5c),
	.w7(32'hbba9815f),
	.w8(32'h3c071d4e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92366f5),
	.w1(32'hba77e0d5),
	.w2(32'hbb910c0a),
	.w3(32'h3b59ea9b),
	.w4(32'h3a3628f4),
	.w5(32'h3ba2a5bd),
	.w6(32'h3b5bb644),
	.w7(32'hbbaa9997),
	.w8(32'hb99d597a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9dfba),
	.w1(32'h3bf62f89),
	.w2(32'h3c1b67d0),
	.w3(32'hbabaead7),
	.w4(32'h3b476954),
	.w5(32'hba9a92ab),
	.w6(32'hbbc5b04a),
	.w7(32'h3ab7c5a0),
	.w8(32'hbb0c961a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb55dd8),
	.w1(32'hbcae9787),
	.w2(32'h3bfcd08f),
	.w3(32'hbc86d2e2),
	.w4(32'hbcb9b0c6),
	.w5(32'hbc47f237),
	.w6(32'hbbdd21d9),
	.w7(32'h3bd7717a),
	.w8(32'h3c261419),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7ad72),
	.w1(32'h3be9a3f6),
	.w2(32'h3b8d36f4),
	.w3(32'h3bf1e9bb),
	.w4(32'h376429fa),
	.w5(32'h3bf23efe),
	.w6(32'h3b92e1b6),
	.w7(32'h3bc03c41),
	.w8(32'hbae18afb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb77bf7),
	.w1(32'hbb0be350),
	.w2(32'hbaedfdc9),
	.w3(32'h3bf7bf4c),
	.w4(32'hb9eefce1),
	.w5(32'h3a32b73d),
	.w6(32'hbb3be952),
	.w7(32'hbb502c14),
	.w8(32'h3ac1d54e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6f5e),
	.w1(32'h3b4c13bf),
	.w2(32'h3bfa9543),
	.w3(32'h39a14e3e),
	.w4(32'h3be38861),
	.w5(32'h3b5db81c),
	.w6(32'h39b934ba),
	.w7(32'h3b50fd5b),
	.w8(32'h3bb336bb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31e583),
	.w1(32'hbb9a1ab8),
	.w2(32'hbba262b8),
	.w3(32'h3b8dc19f),
	.w4(32'hbb41970d),
	.w5(32'hbb496a33),
	.w6(32'hba1e694d),
	.w7(32'hbb68f2f8),
	.w8(32'h3ba0a8c3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c6738),
	.w1(32'h3bc55dd0),
	.w2(32'hbaf4a7dc),
	.w3(32'hbbe69f95),
	.w4(32'hb9a17889),
	.w5(32'h3b5c914e),
	.w6(32'h3ad592f5),
	.w7(32'h3a91100c),
	.w8(32'h3c0f0262),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7147),
	.w1(32'hbc177cd7),
	.w2(32'hbbf18c54),
	.w3(32'h3c1e2c62),
	.w4(32'hbc13836b),
	.w5(32'hbc061501),
	.w6(32'hbc20b0a6),
	.w7(32'hbb86f125),
	.w8(32'h3c3ad3eb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d7ef),
	.w1(32'h3c31937b),
	.w2(32'h3b02cb80),
	.w3(32'hbc4877f1),
	.w4(32'h3c4f7b46),
	.w5(32'h3c62ed6a),
	.w6(32'hbae46d95),
	.w7(32'hbc48a961),
	.w8(32'hbc848b45),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b711),
	.w1(32'h3a725891),
	.w2(32'h3b090a96),
	.w3(32'h3b0efb86),
	.w4(32'h3b67cc83),
	.w5(32'h3b64294b),
	.w6(32'hba8c2383),
	.w7(32'h3b0847b9),
	.w8(32'h3b81102a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b35d9),
	.w1(32'hbc0bd3ca),
	.w2(32'hbbb58057),
	.w3(32'hbb525ec1),
	.w4(32'hbb7a8173),
	.w5(32'h3c2b61b1),
	.w6(32'hbbe8a015),
	.w7(32'hbc581859),
	.w8(32'hbbe4f01b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60dfb6),
	.w1(32'hba15844b),
	.w2(32'h3ba9c37d),
	.w3(32'h3d1e4a62),
	.w4(32'h3b547024),
	.w5(32'h3bbe0402),
	.w6(32'h3b2d0d24),
	.w7(32'h3a6ed1d7),
	.w8(32'h3aa06396),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78627),
	.w1(32'hbb0cac8f),
	.w2(32'hbbb21104),
	.w3(32'h3bf71558),
	.w4(32'hbafe1206),
	.w5(32'hbb4f6e72),
	.w6(32'hbb1111c5),
	.w7(32'hbbb9e25d),
	.w8(32'hbc083ed9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c7d6c),
	.w1(32'hbc1e83ad),
	.w2(32'hbb7e4f62),
	.w3(32'hbc898889),
	.w4(32'hb8ead4dd),
	.w5(32'h3ba1eaee),
	.w6(32'hbb8506a9),
	.w7(32'hbc325928),
	.w8(32'h3a3f288f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae0a3),
	.w1(32'hbb93b269),
	.w2(32'hbbf8adb8),
	.w3(32'h3c41843c),
	.w4(32'h3bc135c7),
	.w5(32'hbac2cb8d),
	.w6(32'h3b536f1b),
	.w7(32'hbaa4cc2b),
	.w8(32'h3b625574),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc721e8c),
	.w1(32'h39ec5628),
	.w2(32'h3b711456),
	.w3(32'hbc492c69),
	.w4(32'hbbe0b970),
	.w5(32'hbaab1ded),
	.w6(32'hbb6e1a54),
	.w7(32'hbbb8708f),
	.w8(32'h3bc8d1cf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2066d5),
	.w1(32'hbac640db),
	.w2(32'h3a9f40ef),
	.w3(32'hbc4c4792),
	.w4(32'h3ba08063),
	.w5(32'h3b111fa3),
	.w6(32'hbb27acf4),
	.w7(32'h3a05ce79),
	.w8(32'h3bf0808a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51ff68),
	.w1(32'hbafebef2),
	.w2(32'h3b02d1a6),
	.w3(32'hba9a3eee),
	.w4(32'hbb1d33dd),
	.w5(32'hba8f7ea2),
	.w6(32'hb91f5d04),
	.w7(32'h3aac3a86),
	.w8(32'hbb489db0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70953b),
	.w1(32'h3a884aea),
	.w2(32'hbba8289e),
	.w3(32'hb9ac0eed),
	.w4(32'hba596f6d),
	.w5(32'hbbf2a6b3),
	.w6(32'hbb9d06d6),
	.w7(32'hbbcf7242),
	.w8(32'hbc0affee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194306),
	.w1(32'hbc2585ba),
	.w2(32'hb8bd6d9e),
	.w3(32'hbb1b06dd),
	.w4(32'h3af29efb),
	.w5(32'hbc0c38d4),
	.w6(32'hbbe1fefa),
	.w7(32'hbc0471a4),
	.w8(32'h3c39d431),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af135e4),
	.w1(32'hba2b0bde),
	.w2(32'h3a7aa3cd),
	.w3(32'hbbe3549f),
	.w4(32'hba8591af),
	.w5(32'h3993b221),
	.w6(32'h3a84d30a),
	.w7(32'hba918813),
	.w8(32'h39f4b931),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb961),
	.w1(32'h3b44c378),
	.w2(32'h3c93583a),
	.w3(32'hbbb78431),
	.w4(32'h3bb33772),
	.w5(32'h3cb723df),
	.w6(32'hba9359de),
	.w7(32'h3bccc249),
	.w8(32'h3b98517d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule