module layer_10_featuremap_399(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec25b),
	.w1(32'hba193b8f),
	.w2(32'h3b75e453),
	.w3(32'hba952946),
	.w4(32'hbb9373e8),
	.w5(32'hbac67edb),
	.w6(32'hbacc08b5),
	.w7(32'hbbff1494),
	.w8(32'hbc96823b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbf237),
	.w1(32'hbbd102cd),
	.w2(32'hbc08f8fe),
	.w3(32'hbc14d074),
	.w4(32'hbc0b079d),
	.w5(32'hbb4a63cf),
	.w6(32'hbc1a6f49),
	.w7(32'hbaeba026),
	.w8(32'h3bca62d0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1b1f),
	.w1(32'h3acc95ff),
	.w2(32'h3b82fd07),
	.w3(32'hbbc733fe),
	.w4(32'hbbb3ba5c),
	.w5(32'h3b9596b9),
	.w6(32'hba5dbb6f),
	.w7(32'h3b6f0314),
	.w8(32'h3b65d9a5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149044),
	.w1(32'h3af64bf3),
	.w2(32'hbbb66bd1),
	.w3(32'h3b383f73),
	.w4(32'h3b9e30cf),
	.w5(32'hbb1aca43),
	.w6(32'h3bb2f0f4),
	.w7(32'hbb11c968),
	.w8(32'h3c1769ad),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd0c7),
	.w1(32'hbc079b18),
	.w2(32'h3afdd5be),
	.w3(32'h3a27e3c3),
	.w4(32'hbc12ee82),
	.w5(32'hbb5945e0),
	.w6(32'h3c078fb0),
	.w7(32'hbc51fd2a),
	.w8(32'hbc2f7210),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf4707),
	.w1(32'h3bbc0212),
	.w2(32'h3a8d5dfa),
	.w3(32'hbc565335),
	.w4(32'h3b28c921),
	.w5(32'hbaf43c54),
	.w6(32'hbc84342f),
	.w7(32'hbc329e8b),
	.w8(32'hbcb0d007),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c48f1),
	.w1(32'h3946b452),
	.w2(32'h3b0c570f),
	.w3(32'h3a73405a),
	.w4(32'hbb8e5869),
	.w5(32'hbc305e3f),
	.w6(32'hbc2e1c28),
	.w7(32'h3a1dc0f5),
	.w8(32'h3badc7f3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1b617),
	.w1(32'h3b5703d5),
	.w2(32'h3c1ca715),
	.w3(32'hbc0d5a21),
	.w4(32'h3c1021aa),
	.w5(32'h3c873204),
	.w6(32'hbb00469e),
	.w7(32'h3c12440e),
	.w8(32'hbabb25ac),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17569d),
	.w1(32'h3bd66aa0),
	.w2(32'hbbc54367),
	.w3(32'h3a699744),
	.w4(32'h3b9e821a),
	.w5(32'hbb4d9064),
	.w6(32'h3b9c97bd),
	.w7(32'h3ac847c1),
	.w8(32'h3bbc04aa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c80f9),
	.w1(32'hbc83f1d9),
	.w2(32'hbca18b42),
	.w3(32'hbab7f44a),
	.w4(32'hbc8c6ed6),
	.w5(32'hbcb5843c),
	.w6(32'h3bdd7441),
	.w7(32'hbc42d65b),
	.w8(32'hbc98bc65),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc907e56),
	.w1(32'hbc545869),
	.w2(32'hbc6879c7),
	.w3(32'hbc2ac1eb),
	.w4(32'hbb44cea9),
	.w5(32'hbb92918b),
	.w6(32'hbc1df32a),
	.w7(32'hbae3a8cc),
	.w8(32'h3b0afaa5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d03cd),
	.w1(32'hbb01613f),
	.w2(32'h3b82e4e3),
	.w3(32'hbb9faeb6),
	.w4(32'hbbea8d86),
	.w5(32'h3a9a0d0e),
	.w6(32'h3ae0be71),
	.w7(32'hbba81770),
	.w8(32'hbadf2f45),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc596b7),
	.w1(32'h3ba07306),
	.w2(32'hbbc732b9),
	.w3(32'hbae595cc),
	.w4(32'hbb957ec7),
	.w5(32'hba53b558),
	.w6(32'hbc1c407c),
	.w7(32'h3a4c0f78),
	.w8(32'h3be2d3ed),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5ed21),
	.w1(32'hbb674ff5),
	.w2(32'hbb5040d2),
	.w3(32'h3a9ee799),
	.w4(32'hbba01b94),
	.w5(32'hbb390cac),
	.w6(32'h39a4e02e),
	.w7(32'h3a98a172),
	.w8(32'h3bcb4e4c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9517e),
	.w1(32'hbadde529),
	.w2(32'hbc01665c),
	.w3(32'hbad3d974),
	.w4(32'hbb0426d4),
	.w5(32'hbb4ebb80),
	.w6(32'hb8fb0c3a),
	.w7(32'h3a82231b),
	.w8(32'h3c78aa24),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e100),
	.w1(32'h3bcbe361),
	.w2(32'h3b8cd0b6),
	.w3(32'hbb8518ab),
	.w4(32'hbabbf88c),
	.w5(32'h3b9b6c74),
	.w6(32'hbb0d5856),
	.w7(32'hbbb79e36),
	.w8(32'h3bb5c855),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae299e6),
	.w1(32'hbb90e89d),
	.w2(32'hbc1a998f),
	.w3(32'hbb45d755),
	.w4(32'hbc062316),
	.w5(32'hbc93386e),
	.w6(32'hbb0a3ab2),
	.w7(32'h3943dd6c),
	.w8(32'hba5dc7b9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6292f),
	.w1(32'h3bcfda0d),
	.w2(32'h3c30787d),
	.w3(32'hbc0acc16),
	.w4(32'hba131057),
	.w5(32'h3a41e70c),
	.w6(32'hbb2408ea),
	.w7(32'hbab88df1),
	.w8(32'hbb942528),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a862ca6),
	.w1(32'h3ab85309),
	.w2(32'hbb0698ca),
	.w3(32'hbb8e35f4),
	.w4(32'h3c02f153),
	.w5(32'h3b3843ad),
	.w6(32'h390088c1),
	.w7(32'h3a8df84b),
	.w8(32'h3bb67187),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc334),
	.w1(32'h3a433262),
	.w2(32'hbb42fe6c),
	.w3(32'hbbac7d45),
	.w4(32'h3be68708),
	.w5(32'hbb2bee00),
	.w6(32'hba5ade24),
	.w7(32'h3b27a34f),
	.w8(32'hbc6c7d2c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa07acf),
	.w1(32'h3c475fe6),
	.w2(32'h3c664203),
	.w3(32'hbb3c9699),
	.w4(32'h3996b20b),
	.w5(32'h3bde66b0),
	.w6(32'hbb125260),
	.w7(32'hbbba4cdb),
	.w8(32'hbb983016),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa15f4),
	.w1(32'h3c3e4971),
	.w2(32'hbc098960),
	.w3(32'h3c0259b4),
	.w4(32'h3b87ebe9),
	.w5(32'h3b663b4e),
	.w6(32'h3983418f),
	.w7(32'hbae0c9a9),
	.w8(32'h3c5496bd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86950d),
	.w1(32'hbb881731),
	.w2(32'hba76edad),
	.w3(32'hbbb20d4f),
	.w4(32'hbbfa9ff5),
	.w5(32'hbbaa75d9),
	.w6(32'hbc411cea),
	.w7(32'hbbaaecf9),
	.w8(32'hbc1defc5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc861947),
	.w1(32'h3c1f9036),
	.w2(32'h3c5cf76c),
	.w3(32'hb8005f78),
	.w4(32'hbc431292),
	.w5(32'hbc4b1822),
	.w6(32'hbc04d259),
	.w7(32'hbc57cda3),
	.w8(32'hbc2e474c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7581c2),
	.w1(32'h3c0e5574),
	.w2(32'hbc1e877e),
	.w3(32'hbc021c45),
	.w4(32'h39d6cccd),
	.w5(32'h3b60af8e),
	.w6(32'hbc71caf0),
	.w7(32'hbac66334),
	.w8(32'h3c414652),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5776a9),
	.w1(32'h3bec753a),
	.w2(32'h3c5e12b7),
	.w3(32'hba5426ab),
	.w4(32'hbc05710a),
	.w5(32'hbbadead6),
	.w6(32'hbaf79c50),
	.w7(32'hbc855ab9),
	.w8(32'hbc9e31e4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886b7e),
	.w1(32'hbb92172f),
	.w2(32'hbc080039),
	.w3(32'hbbd4c1fc),
	.w4(32'h3ab8894e),
	.w5(32'hbb5ae7ae),
	.w6(32'hbc17d072),
	.w7(32'h3b709db2),
	.w8(32'hbbf60cde),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac56cae),
	.w1(32'hb9b9f052),
	.w2(32'hbb60c450),
	.w3(32'hbb1aeff9),
	.w4(32'hbba0360c),
	.w5(32'hbbb836d3),
	.w6(32'hbc2d3f1d),
	.w7(32'hbc80d2a4),
	.w8(32'h3b1497fc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56939d),
	.w1(32'hbc2155fd),
	.w2(32'hbc43e0c4),
	.w3(32'hbb39f8d7),
	.w4(32'hbbcb40c5),
	.w5(32'hbbabf759),
	.w6(32'h39d0d763),
	.w7(32'hba8575e9),
	.w8(32'hbc31557f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44e057),
	.w1(32'h3b9242f4),
	.w2(32'h3b9d388d),
	.w3(32'hba49cf35),
	.w4(32'h3b26dffe),
	.w5(32'h3b8139f3),
	.w6(32'hbbea4e22),
	.w7(32'hbc1eac2e),
	.w8(32'hbc36fd02),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba7dd2),
	.w1(32'hbc07c386),
	.w2(32'hbbdf6352),
	.w3(32'h3bb49c03),
	.w4(32'hba155dda),
	.w5(32'hbb800a6e),
	.w6(32'hbb285c91),
	.w7(32'h3a5497e6),
	.w8(32'hba4f59fe),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc480c20),
	.w1(32'hbad6db0a),
	.w2(32'hbbedaa5b),
	.w3(32'hbaffb9c2),
	.w4(32'hbbb50d10),
	.w5(32'hbc1312d6),
	.w6(32'h3b8d2902),
	.w7(32'h3a4b713d),
	.w8(32'hba426ca8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b6a1a),
	.w1(32'hbc380323),
	.w2(32'hbc719659),
	.w3(32'hba792cf6),
	.w4(32'hbc173504),
	.w5(32'hbc16b0a5),
	.w6(32'hb9947709),
	.w7(32'hbbb994d8),
	.w8(32'hbc2d0c90),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33ba25),
	.w1(32'hbbb22b6e),
	.w2(32'hb995497e),
	.w3(32'hbbf1d90e),
	.w4(32'hbc2be45b),
	.w5(32'hbc0233f1),
	.w6(32'hbc2d6271),
	.w7(32'hbbb4160b),
	.w8(32'hbbdb821c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4196),
	.w1(32'h3b622a05),
	.w2(32'h3bcb2488),
	.w3(32'hbbc65f9e),
	.w4(32'h3c4b7145),
	.w5(32'h3ca614e5),
	.w6(32'hbb9f88e5),
	.w7(32'h3b85f2e7),
	.w8(32'h3ba426a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79312),
	.w1(32'h3b3b6bfa),
	.w2(32'hbb1279a5),
	.w3(32'h3b896fe5),
	.w4(32'hba80f3bb),
	.w5(32'hbbc53c7a),
	.w6(32'h3bbed6a8),
	.w7(32'hba7824ed),
	.w8(32'hbac86664),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeae1a),
	.w1(32'hbbd9b237),
	.w2(32'hbc6e420f),
	.w3(32'hbc0638e2),
	.w4(32'hbaa6da0a),
	.w5(32'h37ae7571),
	.w6(32'hb996ac95),
	.w7(32'hba775b32),
	.w8(32'h3bbb10dc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4f5f4),
	.w1(32'h3b094f74),
	.w2(32'hbc2c9c58),
	.w3(32'hbae3f941),
	.w4(32'hb9dde7a6),
	.w5(32'hbb9f05b6),
	.w6(32'hbb993f7f),
	.w7(32'h3b5f9024),
	.w8(32'h3a7beccd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0584ba),
	.w1(32'h3c97da08),
	.w2(32'h3be5a1c9),
	.w3(32'hbb380033),
	.w4(32'h3b970eed),
	.w5(32'h3b99c993),
	.w6(32'hbb0d5c4e),
	.w7(32'h39dcbed5),
	.w8(32'hbac13710),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaf2ff),
	.w1(32'h3c351465),
	.w2(32'h3c4b7d0f),
	.w3(32'h3ab4ceb9),
	.w4(32'h399a69a7),
	.w5(32'h3ac3cd5e),
	.w6(32'h3bbd2a24),
	.w7(32'hbc0dcc59),
	.w8(32'hbc189cd2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4419),
	.w1(32'h3b5e0a8c),
	.w2(32'h3c1a7637),
	.w3(32'h3aae8253),
	.w4(32'h393cd7e6),
	.w5(32'hbc13c98a),
	.w6(32'hbb2d1786),
	.w7(32'h3be451e5),
	.w8(32'h3bd179f4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c071cb),
	.w1(32'hba01403e),
	.w2(32'hbbb3af1b),
	.w3(32'hbafda9af),
	.w4(32'hb9b0a81f),
	.w5(32'h3b45d488),
	.w6(32'h3bb12b46),
	.w7(32'h3b926b7a),
	.w8(32'h3c2414fd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c0706),
	.w1(32'hbb795e51),
	.w2(32'h3ba7f154),
	.w3(32'h3b4e32ce),
	.w4(32'hbb8fe0e3),
	.w5(32'hbb89760a),
	.w6(32'h3a9518dc),
	.w7(32'hbbcee209),
	.w8(32'hbc4c7512),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a913),
	.w1(32'h3c5532af),
	.w2(32'h3ca0c1f5),
	.w3(32'hb8bff4af),
	.w4(32'h3b6c94b1),
	.w5(32'h3ba8412b),
	.w6(32'hbbf60ab9),
	.w7(32'hbaa86686),
	.w8(32'hbbe73bbc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a948b),
	.w1(32'hbbe969d9),
	.w2(32'hbc3fd66f),
	.w3(32'h3a676d09),
	.w4(32'hbbb20dc4),
	.w5(32'hbc41d3f7),
	.w6(32'h3a7362e7),
	.w7(32'hbc17706d),
	.w8(32'hbc54e1c7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25db3d),
	.w1(32'hbb9f41f1),
	.w2(32'hbbea95f8),
	.w3(32'hbbf390ca),
	.w4(32'h3aaae3b0),
	.w5(32'h3b62a41c),
	.w6(32'hbb47c283),
	.w7(32'hb9bec8e6),
	.w8(32'h3b9ec852),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69930),
	.w1(32'h3b2b7d7c),
	.w2(32'hba1b6d5f),
	.w3(32'hbba12461),
	.w4(32'hbb17aec4),
	.w5(32'hbb8b1283),
	.w6(32'hba5c9bf1),
	.w7(32'h3c2a47f6),
	.w8(32'h3c95a414),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf594bd),
	.w1(32'hbaf62a05),
	.w2(32'hbb80add1),
	.w3(32'hbb3fc1e4),
	.w4(32'hbc024ec0),
	.w5(32'h3b4c12f2),
	.w6(32'h3c38e763),
	.w7(32'hbb0b6f6f),
	.w8(32'h3bdffaba),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc005d),
	.w1(32'h39ca69b0),
	.w2(32'hbbfe8956),
	.w3(32'h3acdbb91),
	.w4(32'h3be1dd1e),
	.w5(32'hbc043757),
	.w6(32'h3b919b7a),
	.w7(32'h3b1c9860),
	.w8(32'h3b292917),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec7f3),
	.w1(32'h3ba4dc6e),
	.w2(32'h3b14979e),
	.w3(32'hbc0072a4),
	.w4(32'hbaec6531),
	.w5(32'hba789e05),
	.w6(32'h3ad7e514),
	.w7(32'h3bb9afd9),
	.w8(32'h3bd7511a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0baec),
	.w1(32'hbaf23705),
	.w2(32'h3af74d4f),
	.w3(32'hb98dc2d5),
	.w4(32'hbb9aa3e5),
	.w5(32'h3b505080),
	.w6(32'h3b4b2d9c),
	.w7(32'h38305f88),
	.w8(32'h3b8c9df6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc638f3),
	.w1(32'hbc5c7c68),
	.w2(32'hbcc6f856),
	.w3(32'hbb363683),
	.w4(32'hbaf3cff2),
	.w5(32'hbbad2984),
	.w6(32'hbb62d61a),
	.w7(32'h3b851022),
	.w8(32'h3c308465),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72d39b),
	.w1(32'h3c616292),
	.w2(32'h3c4eeb85),
	.w3(32'h3b14adbd),
	.w4(32'h3b4d5c97),
	.w5(32'h3b5ad12a),
	.w6(32'hbb9e6979),
	.w7(32'hbb59dc98),
	.w8(32'hbbb3dc22),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b550995),
	.w1(32'h3b7925e9),
	.w2(32'h3bfb70bb),
	.w3(32'hbb95813e),
	.w4(32'h3b982c6c),
	.w5(32'h3cb0d529),
	.w6(32'hbbc69464),
	.w7(32'hbb40672c),
	.w8(32'hbb739ced),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a699acd),
	.w1(32'h3c03f955),
	.w2(32'hbc15bef8),
	.w3(32'h3941cd3b),
	.w4(32'h3b662241),
	.w5(32'hbc694656),
	.w6(32'hbb8d0705),
	.w7(32'hbb2b222d),
	.w8(32'hbc1259ca),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41ff80),
	.w1(32'hbb297063),
	.w2(32'hb8b8ad4a),
	.w3(32'hb9ca7156),
	.w4(32'hbb993b56),
	.w5(32'hbbf85d66),
	.w6(32'h3c48b497),
	.w7(32'h3b3ebdd7),
	.w8(32'hbb82fd33),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3410e8),
	.w1(32'hb998f77b),
	.w2(32'h3bae7198),
	.w3(32'hbb224fc6),
	.w4(32'hbb7b18dc),
	.w5(32'hba70f9b4),
	.w6(32'hbba37d47),
	.w7(32'hbc6dd620),
	.w8(32'hbc800942),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399134cf),
	.w1(32'hbb794caf),
	.w2(32'h3b927ee0),
	.w3(32'hbbf9d763),
	.w4(32'h3b7b4d47),
	.w5(32'hba96d975),
	.w6(32'hbbfeb939),
	.w7(32'hbacd761f),
	.w8(32'h3aec6253),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b5508),
	.w1(32'h3c00d52f),
	.w2(32'h3c25c8b6),
	.w3(32'h3b8d7116),
	.w4(32'h3bcfec66),
	.w5(32'h3b6016cb),
	.w6(32'hbc3a780b),
	.w7(32'h3c122820),
	.w8(32'h3b31bc8e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd229e0),
	.w1(32'h3b25811f),
	.w2(32'hbb45c833),
	.w3(32'h3c336ef2),
	.w4(32'h3b508ccd),
	.w5(32'hbbc36549),
	.w6(32'h3c1ea15e),
	.w7(32'h3c251e69),
	.w8(32'hbbb40308),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8427c5),
	.w1(32'hbbddc46f),
	.w2(32'hbb3f2cfc),
	.w3(32'hbc2c4412),
	.w4(32'hbc3bed93),
	.w5(32'hbc30f09e),
	.w6(32'h3b4a7a7e),
	.w7(32'hbba9d5e0),
	.w8(32'hbc83e19e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b08d),
	.w1(32'h3bd2a356),
	.w2(32'h3b96d307),
	.w3(32'hbc39dee9),
	.w4(32'h3b85c391),
	.w5(32'h3baba479),
	.w6(32'hbbd49c3b),
	.w7(32'hbb9e79e6),
	.w8(32'hbb621a13),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba276857),
	.w1(32'h39918dc8),
	.w2(32'hb9bc899a),
	.w3(32'h3abb31dd),
	.w4(32'h3a5ae928),
	.w5(32'h3abec210),
	.w6(32'h3bb7570b),
	.w7(32'h3c01eb6f),
	.w8(32'h3bf05ce7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f34b),
	.w1(32'hbb95f871),
	.w2(32'h3b991610),
	.w3(32'h3bade126),
	.w4(32'hbb88b097),
	.w5(32'h3ad4e156),
	.w6(32'h3c0f8676),
	.w7(32'hbbdeb11d),
	.w8(32'hbc32312b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38b2ae),
	.w1(32'h3c32066b),
	.w2(32'h3c6c19f5),
	.w3(32'hbb648b55),
	.w4(32'hba6577bd),
	.w5(32'hbb1e9469),
	.w6(32'hbbded29a),
	.w7(32'hbb7ba359),
	.w8(32'hbc1b924d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b899246),
	.w1(32'h3beb8c42),
	.w2(32'h3be6ad11),
	.w3(32'hbbd9da1d),
	.w4(32'hb9f85228),
	.w5(32'hbad0a5e6),
	.w6(32'hbc2c2ceb),
	.w7(32'hbbf2fd3c),
	.w8(32'hbc89fc9c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b055d77),
	.w1(32'hbb086e88),
	.w2(32'h3ae4296d),
	.w3(32'hbb7bd7f9),
	.w4(32'hbbb834a2),
	.w5(32'hb9c5968c),
	.w6(32'hbc2d0037),
	.w7(32'hbb707df0),
	.w8(32'hbc424267),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a372549),
	.w1(32'hbc4befd8),
	.w2(32'hbc4eafb6),
	.w3(32'hbbbc5614),
	.w4(32'hbc10e073),
	.w5(32'h3b116c55),
	.w6(32'hbb46799b),
	.w7(32'h3b7818ee),
	.w8(32'h3b8eb14e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2b67),
	.w1(32'hbc4b21b8),
	.w2(32'hbc2688e7),
	.w3(32'hbc18a35d),
	.w4(32'hbbb23a19),
	.w5(32'h3b86af29),
	.w6(32'hbb9bcf9e),
	.w7(32'h3c053110),
	.w8(32'h3c6cc57e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2fbf),
	.w1(32'h3819b70e),
	.w2(32'h38049a6f),
	.w3(32'h3bb0e0a1),
	.w4(32'h37747e1b),
	.w5(32'h37d654c4),
	.w6(32'h3b923079),
	.w7(32'h37caec6b),
	.w8(32'h38285fdf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d6d355),
	.w1(32'hb70c4126),
	.w2(32'hb60e7ae7),
	.w3(32'hb685165b),
	.w4(32'hb75a46f6),
	.w5(32'h37352483),
	.w6(32'hb34656f8),
	.w7(32'h36c41fa1),
	.w8(32'h36c83e0a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cc3b5c),
	.w1(32'hb7f9530b),
	.w2(32'hb764d480),
	.w3(32'hb7785bd0),
	.w4(32'hb708e1f3),
	.w5(32'hb7929a38),
	.w6(32'hb709572f),
	.w7(32'hb7bb46a9),
	.w8(32'hb674e014),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76f0fc4),
	.w1(32'h36583f73),
	.w2(32'hb63428b0),
	.w3(32'h37f329bc),
	.w4(32'hb71c0551),
	.w5(32'hb782278d),
	.w6(32'h366d5210),
	.w7(32'h35ff75d0),
	.w8(32'hb7daefcc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c875d2),
	.w1(32'hb2804fb5),
	.w2(32'hb7333935),
	.w3(32'h36f48f35),
	.w4(32'h36a5b0eb),
	.w5(32'hb69b44b4),
	.w6(32'h378dea4a),
	.w7(32'h378aa548),
	.w8(32'hb702f957),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372b5d44),
	.w1(32'h37cdece2),
	.w2(32'h37b68b95),
	.w3(32'h37703281),
	.w4(32'h3802d99d),
	.w5(32'h3794698c),
	.w6(32'h35fb55ec),
	.w7(32'h37228ff0),
	.w8(32'hb7730f80),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63565e6),
	.w1(32'hb7513329),
	.w2(32'hb7d40134),
	.w3(32'h3741a8df),
	.w4(32'h362cbfa3),
	.w5(32'hb788e39b),
	.w6(32'hb846cb6e),
	.w7(32'h36b628d2),
	.w8(32'hb6983525),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7058e87),
	.w1(32'hb6c07a5a),
	.w2(32'h3713bf9a),
	.w3(32'hb6e56980),
	.w4(32'hb738a421),
	.w5(32'hb4817df8),
	.w6(32'hb7fe5743),
	.w7(32'hb70c12ea),
	.w8(32'hb73e817f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3623bef4),
	.w1(32'h37492fbc),
	.w2(32'h3780a917),
	.w3(32'h37914829),
	.w4(32'hb7c1d5cf),
	.w5(32'hb31d1f23),
	.w6(32'hb6a71713),
	.w7(32'hb6c41e80),
	.w8(32'h37cf8064),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb650dbb8),
	.w1(32'hb6c0ed43),
	.w2(32'h3793f869),
	.w3(32'h37e6e570),
	.w4(32'hb701ecf9),
	.w5(32'h3686eab0),
	.w6(32'h38112018),
	.w7(32'hb78eea71),
	.w8(32'h362fb972),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74eec9c),
	.w1(32'hb5dc6659),
	.w2(32'h3653366c),
	.w3(32'h36d600c0),
	.w4(32'hb6c47274),
	.w5(32'hb6a6206f),
	.w6(32'hb783cbf3),
	.w7(32'hb6d1e1fe),
	.w8(32'h36d9f7be),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57b8b4e),
	.w1(32'hb7a457b6),
	.w2(32'h376afae3),
	.w3(32'hb74a4ed4),
	.w4(32'hb7ed6eb4),
	.w5(32'h36b277a2),
	.w6(32'hb6b1c795),
	.w7(32'hb769f460),
	.w8(32'h363832dd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371240ac),
	.w1(32'hb77a4bb3),
	.w2(32'hb6ae1019),
	.w3(32'h3702ce45),
	.w4(32'hb791bdea),
	.w5(32'hb5cb8adb),
	.w6(32'hb6f8e4a0),
	.w7(32'h371a7aa9),
	.w8(32'h3731090d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b5066a),
	.w1(32'hb8082da7),
	.w2(32'h3582f5a5),
	.w3(32'h35c5b86d),
	.w4(32'hb7d383d1),
	.w5(32'h37019d9f),
	.w6(32'h36b76db1),
	.w7(32'hb7b6d636),
	.w8(32'h377759e8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78cf944),
	.w1(32'hb6bbe389),
	.w2(32'hb7de4b82),
	.w3(32'hb744f5d0),
	.w4(32'hb7a3f9df),
	.w5(32'hb5ca5faf),
	.w6(32'h3694f39b),
	.w7(32'h36dae579),
	.w8(32'hb70e4e44),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba4398),
	.w1(32'h36ea0b94),
	.w2(32'hb6da59d6),
	.w3(32'h35cc7352),
	.w4(32'hb76f07e0),
	.w5(32'hb7a23308),
	.w6(32'hb8758947),
	.w7(32'h36a71aee),
	.w8(32'hb71606f9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3505c41a),
	.w1(32'hb79cb612),
	.w2(32'h37443409),
	.w3(32'h367719f5),
	.w4(32'h38163221),
	.w5(32'h370b3a90),
	.w6(32'h36b5e08b),
	.w7(32'hb623bd07),
	.w8(32'hb64e0570),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803e1e3),
	.w1(32'h3791b0a7),
	.w2(32'hb711d239),
	.w3(32'h3805f22e),
	.w4(32'hb6a0a82d),
	.w5(32'hb7efc32f),
	.w6(32'h386de720),
	.w7(32'hb6c735e7),
	.w8(32'h37069208),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3628fd94),
	.w1(32'hb5b4b42f),
	.w2(32'hb70ef153),
	.w3(32'hb7b7e903),
	.w4(32'hb38bb05c),
	.w5(32'h37b13a99),
	.w6(32'hb67d6dce),
	.w7(32'hb7f384d9),
	.w8(32'h37540835),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38074bca),
	.w1(32'h373d8cc5),
	.w2(32'h37404cb7),
	.w3(32'h35c39deb),
	.w4(32'h32401792),
	.w5(32'hb78c10c4),
	.w6(32'h3773784e),
	.w7(32'h376eaacb),
	.w8(32'hb72c8ac7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716bff3),
	.w1(32'hb6c3c621),
	.w2(32'hb80273db),
	.w3(32'h37996523),
	.w4(32'hb6915d2b),
	.w5(32'hb71abbe5),
	.w6(32'hb826ed18),
	.w7(32'h376e16eb),
	.w8(32'h36df9203),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e9aae),
	.w1(32'h36e6bc98),
	.w2(32'h36006056),
	.w3(32'h36773e8d),
	.w4(32'h3690303f),
	.w5(32'hb5117682),
	.w6(32'h376dd954),
	.w7(32'h37df7985),
	.w8(32'h377748d8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a99e3f),
	.w1(32'h373c2de6),
	.w2(32'h377fd29e),
	.w3(32'h36f235fc),
	.w4(32'h37271aba),
	.w5(32'h37db1cfc),
	.w6(32'h37cf328a),
	.w7(32'h366bc0d6),
	.w8(32'h377dd99f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ef1958),
	.w1(32'hb770a0be),
	.w2(32'h373993f1),
	.w3(32'hb7b19462),
	.w4(32'hb6863ddd),
	.w5(32'h37d092bb),
	.w6(32'hb60d86cd),
	.w7(32'hb76441f6),
	.w8(32'h377e75aa),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ae6194),
	.w1(32'h3766b727),
	.w2(32'h37f54193),
	.w3(32'h37ca843d),
	.w4(32'h3802d806),
	.w5(32'h37de7327),
	.w6(32'h364c1047),
	.w7(32'h382c118c),
	.w8(32'h380f1701),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772657b),
	.w1(32'h3768d305),
	.w2(32'h379a30a0),
	.w3(32'hb6baac04),
	.w4(32'h3717d771),
	.w5(32'h3759ab0c),
	.w6(32'hb79ca4c1),
	.w7(32'hb7ae344b),
	.w8(32'hb762e11c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f69aad),
	.w1(32'h36d64c5f),
	.w2(32'hb70c1b1e),
	.w3(32'h37bc7901),
	.w4(32'h36b27a98),
	.w5(32'hb698df9d),
	.w6(32'h3655c619),
	.w7(32'hb64f9861),
	.w8(32'hb870f17a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3590759c),
	.w1(32'hb79ffc9a),
	.w2(32'hb7c4842b),
	.w3(32'h380566a4),
	.w4(32'hb718f45c),
	.w5(32'hb6000ace),
	.w6(32'hb5c24409),
	.w7(32'hb4600c0d),
	.w8(32'h368f7cfc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b50f7),
	.w1(32'h377a49e9),
	.w2(32'h37aadfd5),
	.w3(32'h380aa8d6),
	.w4(32'hb6e25c94),
	.w5(32'hb5c9576a),
	.w6(32'h384c047c),
	.w7(32'h378cc5c2),
	.w8(32'h374a9c05),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58571d0),
	.w1(32'h37174f10),
	.w2(32'hb7a89caf),
	.w3(32'h368a8095),
	.w4(32'hb6aa91ba),
	.w5(32'hb738a34f),
	.w6(32'h372c226a),
	.w7(32'h36312f5b),
	.w8(32'hb60ad117),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f4a8e3),
	.w1(32'h37941aee),
	.w2(32'h36b5146b),
	.w3(32'hb830869a),
	.w4(32'hb6244fe7),
	.w5(32'h35246f4f),
	.w6(32'hb6b7f517),
	.w7(32'h382243d0),
	.w8(32'h37c89bba),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6866cd7),
	.w1(32'h371f6a4c),
	.w2(32'h37a172d6),
	.w3(32'h37c4509c),
	.w4(32'h3780240e),
	.w5(32'h378801d0),
	.w6(32'hb7f98dc9),
	.w7(32'hb75173b5),
	.w8(32'h3796b8ae),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837200b),
	.w1(32'h37ccdd8d),
	.w2(32'h37db0252),
	.w3(32'h384b27d3),
	.w4(32'h371094d1),
	.w5(32'h37cc182f),
	.w6(32'h35ff11fc),
	.w7(32'h36e621a0),
	.w8(32'h35e8b619),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb630eeb1),
	.w1(32'hb74e39e1),
	.w2(32'h37c0b9ad),
	.w3(32'h374cd190),
	.w4(32'hb7d66c34),
	.w5(32'h3760b219),
	.w6(32'hb709816c),
	.w7(32'hb712c784),
	.w8(32'h383378ae),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374c91b5),
	.w1(32'h37d49e84),
	.w2(32'h36368dd4),
	.w3(32'hb633456b),
	.w4(32'hb7637de8),
	.w5(32'hb7bbd932),
	.w6(32'h38098f92),
	.w7(32'h36eeb9d8),
	.w8(32'hb66d026e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72a064d),
	.w1(32'hb7ed0352),
	.w2(32'hb704304c),
	.w3(32'h37bb2dae),
	.w4(32'h36c59b15),
	.w5(32'h37a3fd4d),
	.w6(32'h37dedfcf),
	.w7(32'h37819058),
	.w8(32'h37a94791),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d83fcc),
	.w1(32'hb787a5a3),
	.w2(32'h34520385),
	.w3(32'h354ad4c0),
	.w4(32'hb6b13351),
	.w5(32'h3684d8e1),
	.w6(32'h359ac8bf),
	.w7(32'hb4d8ad7c),
	.w8(32'hb5b1cd58),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78823eb),
	.w1(32'hb7795502),
	.w2(32'h36c62802),
	.w3(32'hb7761147),
	.w4(32'hb74db79b),
	.w5(32'h378374e4),
	.w6(32'hb6702eb4),
	.w7(32'hb7350108),
	.w8(32'h373dafaa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3725cf0c),
	.w1(32'hb66eca36),
	.w2(32'h359f1096),
	.w3(32'h3784c2f8),
	.w4(32'hb7801d55),
	.w5(32'h3581dedf),
	.w6(32'h375f8b32),
	.w7(32'hb68b1ad3),
	.w8(32'h361fccb3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f1d63),
	.w1(32'h373bac2b),
	.w2(32'h371549df),
	.w3(32'h37f845af),
	.w4(32'h381acb65),
	.w5(32'h37d96da6),
	.w6(32'h382691c6),
	.w7(32'h382f6b97),
	.w8(32'h3803d989),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c67ef9),
	.w1(32'h3715c492),
	.w2(32'h368c3771),
	.w3(32'h3865805f),
	.w4(32'h370f796e),
	.w5(32'h379ed280),
	.w6(32'h3811120f),
	.w7(32'h38263346),
	.w8(32'h3765fcc6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70d7f5c),
	.w1(32'hb78ff548),
	.w2(32'h3711a8f4),
	.w3(32'h3739c4ce),
	.w4(32'hb562955a),
	.w5(32'h35187e82),
	.w6(32'h3664429b),
	.w7(32'hb7928ddd),
	.w8(32'h36d3e12b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5d013),
	.w1(32'hb742374c),
	.w2(32'hb6fc6e31),
	.w3(32'h38013085),
	.w4(32'hb75f5a4c),
	.w5(32'h36cb3240),
	.w6(32'h37c875d7),
	.w7(32'h33734ee2),
	.w8(32'hb709d9f2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb786b2f3),
	.w1(32'h3679009b),
	.w2(32'h37d97c0d),
	.w3(32'hb70f33d5),
	.w4(32'hb7094d74),
	.w5(32'hb6eeffdc),
	.w6(32'hb72ef202),
	.w7(32'hb5a354e2),
	.w8(32'h365d5693),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373fa388),
	.w1(32'h36e8661b),
	.w2(32'hb7a3159e),
	.w3(32'hb7b59f3b),
	.w4(32'h36e78bb8),
	.w5(32'hb74ba6ed),
	.w6(32'h374e84c7),
	.w7(32'h378632d3),
	.w8(32'hb7887673),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37149b33),
	.w1(32'hb780a5a0),
	.w2(32'h37c0c92f),
	.w3(32'h373affa1),
	.w4(32'hb79c1b2d),
	.w5(32'hb6ed4bd5),
	.w6(32'hb81afb26),
	.w7(32'hb75f1ba7),
	.w8(32'h36ef751c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7272dfa),
	.w1(32'hb53df3de),
	.w2(32'h357a336b),
	.w3(32'hb786d5ef),
	.w4(32'hb668b5be),
	.w5(32'h3622436f),
	.w6(32'hb7fcbbd3),
	.w7(32'h3761e445),
	.w8(32'h34dc779b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bccfe3),
	.w1(32'hb7cc2dfc),
	.w2(32'h377000df),
	.w3(32'hb53925bf),
	.w4(32'h37194a66),
	.w5(32'h3791b9af),
	.w6(32'h3657ad46),
	.w7(32'h3768fc8c),
	.w8(32'h3679453a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377951ea),
	.w1(32'hb7c0a12f),
	.w2(32'h36f5894c),
	.w3(32'h3751b4b7),
	.w4(32'h376d830e),
	.w5(32'h3770ac3a),
	.w6(32'hb7b20640),
	.w7(32'h37ef798d),
	.w8(32'h367c6362),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c40c2c),
	.w1(32'h3710c256),
	.w2(32'h36949dbc),
	.w3(32'h351e3939),
	.w4(32'hb66cfab1),
	.w5(32'h3570bfd9),
	.w6(32'hb735521f),
	.w7(32'hb7c30575),
	.w8(32'hb6da94c5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb56d7490),
	.w1(32'hb70c4154),
	.w2(32'h382deed3),
	.w3(32'h37857599),
	.w4(32'hb8234411),
	.w5(32'h36d49bc2),
	.w6(32'h37197b22),
	.w7(32'hb806f243),
	.w8(32'hb71f2de2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3781e871),
	.w1(32'h3691030d),
	.w2(32'h36a235a5),
	.w3(32'hb6b941ee),
	.w4(32'h3704668f),
	.w5(32'h36a17a4e),
	.w6(32'hb69cc002),
	.w7(32'h3798b786),
	.w8(32'h350685d3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb746e28e),
	.w1(32'h371af354),
	.w2(32'hb7d87b73),
	.w3(32'h37175db9),
	.w4(32'hb73beded),
	.w5(32'hb750ba6b),
	.w6(32'hb7d6cdcc),
	.w7(32'h367c39ad),
	.w8(32'h37244e94),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6abed41),
	.w1(32'hb7d61c90),
	.w2(32'h36f154dc),
	.w3(32'hb7e0c5c1),
	.w4(32'hb6c8c52d),
	.w5(32'hb68fd330),
	.w6(32'hb7cd25ab),
	.w7(32'hb657304e),
	.w8(32'hb63eec58),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37924dbb),
	.w1(32'hb799865c),
	.w2(32'hb7959fa0),
	.w3(32'hb80325a3),
	.w4(32'hb7afbfd4),
	.w5(32'h36357bc8),
	.w6(32'hb727de95),
	.w7(32'hb7a9d55c),
	.w8(32'hb7c44a69),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ad0896),
	.w1(32'hb7e12f19),
	.w2(32'hb73be4e9),
	.w3(32'hb6665f1a),
	.w4(32'h370e326f),
	.w5(32'h37033b7f),
	.w6(32'hb7e2eee9),
	.w7(32'h373d12bb),
	.w8(32'hb71af3a8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eea51e),
	.w1(32'hb803c8cf),
	.w2(32'hb71905ef),
	.w3(32'h38091e38),
	.w4(32'hb4f1b1e6),
	.w5(32'h362800ca),
	.w6(32'hb795d3ab),
	.w7(32'h378f52e6),
	.w8(32'hb63bff6f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fd53a6),
	.w1(32'h3754c5be),
	.w2(32'hb6b1f0c0),
	.w3(32'h371f92b3),
	.w4(32'hb6c239c0),
	.w5(32'hb792fe3f),
	.w6(32'hb704d9c7),
	.w7(32'h3741ca4c),
	.w8(32'h372aa3b6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64f002e),
	.w1(32'hb7abc259),
	.w2(32'hb7c6a39b),
	.w3(32'hb8034ae7),
	.w4(32'hb52c48a3),
	.w5(32'h35a2ccea),
	.w6(32'h36e02c8c),
	.w7(32'h359076f8),
	.w8(32'h366200cf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363f7ea5),
	.w1(32'h38092a02),
	.w2(32'h37c9e9de),
	.w3(32'h366048f7),
	.w4(32'hb62cbfbb),
	.w5(32'hb72b9e59),
	.w6(32'h3782a91d),
	.w7(32'hb605d76c),
	.w8(32'hb681e861),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b22c75),
	.w1(32'hb6ac9de0),
	.w2(32'hb6f3e02e),
	.w3(32'hb68593d2),
	.w4(32'hb669084c),
	.w5(32'hb789d1f8),
	.w6(32'hb6927e10),
	.w7(32'hb796e723),
	.w8(32'hb6532075),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7723b83),
	.w1(32'hb7bdcb88),
	.w2(32'hb73f850e),
	.w3(32'hb6c184d2),
	.w4(32'hb7df069e),
	.w5(32'hb78655ed),
	.w6(32'h33ff3170),
	.w7(32'h365c2c35),
	.w8(32'hb7978617),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5f8d9),
	.w1(32'h36df1785),
	.w2(32'hb6a59fcd),
	.w3(32'h36e78243),
	.w4(32'h382c696b),
	.w5(32'hb7867cfe),
	.w6(32'hb7281442),
	.w7(32'h37819b9d),
	.w8(32'h364e6a41),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ed7508),
	.w1(32'h36bf8fec),
	.w2(32'h359786d7),
	.w3(32'h36f25bb5),
	.w4(32'h35f0eaca),
	.w5(32'h370c5629),
	.w6(32'h3703c5b0),
	.w7(32'hb624f8ce),
	.w8(32'h36d17f62),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fc855c),
	.w1(32'hb7bc353e),
	.w2(32'hb75296ec),
	.w3(32'h37471e5d),
	.w4(32'hb74f00a4),
	.w5(32'hb5ca7fc7),
	.w6(32'h372ea913),
	.w7(32'hb5e36ebb),
	.w8(32'hb6898916),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7935c1d),
	.w1(32'hb742b535),
	.w2(32'hb74771cc),
	.w3(32'hb6aead37),
	.w4(32'hb689f939),
	.w5(32'h36fca818),
	.w6(32'hb72fb357),
	.w7(32'h37ebc3c8),
	.w8(32'h369d4676),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b191a0),
	.w1(32'hb6585711),
	.w2(32'h376dcb35),
	.w3(32'h38147648),
	.w4(32'h3764697a),
	.w5(32'h376dd710),
	.w6(32'h38115ddf),
	.w7(32'h37378e67),
	.w8(32'h3790d37e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710a0d1),
	.w1(32'h35886e75),
	.w2(32'hb7e85ecf),
	.w3(32'hb7297842),
	.w4(32'h374ea5ae),
	.w5(32'hb7af73f9),
	.w6(32'h371abcba),
	.w7(32'h37ee85d8),
	.w8(32'hb7ec5181),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787e381),
	.w1(32'hb62de4c6),
	.w2(32'hb4844d0c),
	.w3(32'h381c9309),
	.w4(32'h37697445),
	.w5(32'h371af28c),
	.w6(32'hb646f271),
	.w7(32'h3764e650),
	.w8(32'h35d41de8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3706e8bd),
	.w1(32'hb48b54ba),
	.w2(32'hb72a93a5),
	.w3(32'h372eb567),
	.w4(32'h37c27272),
	.w5(32'h373eeed8),
	.w6(32'hb6cce49d),
	.w7(32'h3796bd09),
	.w8(32'h3784c288),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a5191a),
	.w1(32'hb715a66f),
	.w2(32'hb7279d57),
	.w3(32'h377331a9),
	.w4(32'hb79f7ab3),
	.w5(32'hb6fda342),
	.w6(32'h378687c7),
	.w7(32'h35bdf0c4),
	.w8(32'h362d328f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5564b52),
	.w1(32'hb80b3abe),
	.w2(32'hb72bf4bc),
	.w3(32'hb6cdcb7d),
	.w4(32'h3541ae66),
	.w5(32'h37583277),
	.w6(32'hb70fbcd4),
	.w7(32'hb7268797),
	.w8(32'h37636db6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b15317),
	.w1(32'hb65a95a7),
	.w2(32'h370f1995),
	.w3(32'h36cd3412),
	.w4(32'h36ab27ec),
	.w5(32'hb6837908),
	.w6(32'h3698f2fe),
	.w7(32'h37599aa0),
	.w8(32'h37945518),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb40b7912),
	.w1(32'hb6f553c2),
	.w2(32'h371d4097),
	.w3(32'hb66a71fc),
	.w4(32'hb787cfb5),
	.w5(32'hb5bc0e44),
	.w6(32'h37fec4b1),
	.w7(32'h35da8d81),
	.w8(32'hb79b8047),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378bfde3),
	.w1(32'h36b431d7),
	.w2(32'h379ae710),
	.w3(32'h36ac161a),
	.w4(32'hb64981d6),
	.w5(32'h37a415f5),
	.w6(32'hb7b1b5a5),
	.w7(32'hb5b3c05e),
	.w8(32'h3763f2fb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c798bf),
	.w1(32'hb68b7046),
	.w2(32'h3610ff37),
	.w3(32'hb7b39eef),
	.w4(32'hb7d5997d),
	.w5(32'hb77d406b),
	.w6(32'hb7772457),
	.w7(32'h35588f1f),
	.w8(32'hb6c4ebb5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67ec95f),
	.w1(32'h37b50395),
	.w2(32'h380aacb9),
	.w3(32'hb795ffb6),
	.w4(32'h37750b99),
	.w5(32'h378b7408),
	.w6(32'h3727bf38),
	.w7(32'hb6ac5680),
	.w8(32'hb7218dc1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722a0c5),
	.w1(32'h369830f5),
	.w2(32'hb60c300e),
	.w3(32'h37072aa0),
	.w4(32'hb73d8ad2),
	.w5(32'hb6340954),
	.w6(32'h3721f319),
	.w7(32'h36aef520),
	.w8(32'hb62803d9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cd8f75),
	.w1(32'h379b55d9),
	.w2(32'h3785674e),
	.w3(32'h37c11ea4),
	.w4(32'h3789825d),
	.w5(32'h36f43825),
	.w6(32'h37313863),
	.w7(32'h37e4062f),
	.w8(32'h37b592bd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb724c3ee),
	.w1(32'hb69661c2),
	.w2(32'h37080a28),
	.w3(32'hb7ca06cc),
	.w4(32'hb67dfbed),
	.w5(32'h37e087c2),
	.w6(32'hb734f5e4),
	.w7(32'hb736bd8f),
	.w8(32'h3738c95c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a1e38),
	.w1(32'h35969df1),
	.w2(32'h36a10417),
	.w3(32'h370e1c6b),
	.w4(32'hb742b3c7),
	.w5(32'h36411a09),
	.w6(32'h36ede8ff),
	.w7(32'hb6356461),
	.w8(32'h37e8524f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3786bb84),
	.w1(32'h3732b31f),
	.w2(32'h373a1196),
	.w3(32'h373d45dc),
	.w4(32'h36da9b5e),
	.w5(32'h378b59e0),
	.w6(32'h381d791e),
	.w7(32'h37c2365c),
	.w8(32'h37cb8676),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c9c835),
	.w1(32'h36b17e70),
	.w2(32'h3789fbe5),
	.w3(32'h37a9377e),
	.w4(32'h35099aae),
	.w5(32'h369662b6),
	.w6(32'hb6f438c9),
	.w7(32'hb752cc9e),
	.w8(32'hb781f813),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cd8565),
	.w1(32'hb698d5f8),
	.w2(32'hb741216c),
	.w3(32'h37ac1d06),
	.w4(32'h34c153f5),
	.w5(32'hb71f0261),
	.w6(32'hb74aacfe),
	.w7(32'h37eb60e5),
	.w8(32'h363c9e67),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38095780),
	.w1(32'hb7249f6d),
	.w2(32'hb72a7252),
	.w3(32'h36e6ed01),
	.w4(32'hb78f9694),
	.w5(32'h359f0e27),
	.w6(32'h3821aeb1),
	.w7(32'hb787ece0),
	.w8(32'h3494ff09),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8060cfc),
	.w1(32'hb62aa3cd),
	.w2(32'h37711969),
	.w3(32'hb7c39e38),
	.w4(32'hb7a69d73),
	.w5(32'h379a4bb3),
	.w6(32'hb706b8d8),
	.w7(32'hb7db49df),
	.w8(32'h37d59e96),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37175a6f),
	.w1(32'h34207f5e),
	.w2(32'h37228990),
	.w3(32'h375892b9),
	.w4(32'hb796cb45),
	.w5(32'hb6479d12),
	.w6(32'h3845d550),
	.w7(32'hb617edc7),
	.w8(32'hb7934967),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362ff2ce),
	.w1(32'h361bb636),
	.w2(32'hb7bb96b2),
	.w3(32'hb681955c),
	.w4(32'hb78e5a91),
	.w5(32'hb7b9800d),
	.w6(32'hb6e4b684),
	.w7(32'hb79b7725),
	.w8(32'hb78c3d98),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5050b),
	.w1(32'hb7721ddc),
	.w2(32'hb788ee97),
	.w3(32'h3579afee),
	.w4(32'hb7c8ce30),
	.w5(32'hb70f330b),
	.w6(32'hb74b207e),
	.w7(32'hb75909f2),
	.w8(32'hb67ccefb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb784c2fd),
	.w1(32'hb5e95efa),
	.w2(32'h36cd37b6),
	.w3(32'hb5cc3d98),
	.w4(32'hb6a4ef8e),
	.w5(32'hb65fe56a),
	.w6(32'hb547eff6),
	.w7(32'h36f9ea96),
	.w8(32'hb748b053),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728f4e4),
	.w1(32'hb7d34255),
	.w2(32'h375f4a0d),
	.w3(32'h37759500),
	.w4(32'hb8010e7f),
	.w5(32'h36056f90),
	.w6(32'h369ccd29),
	.w7(32'hb7dd5b6e),
	.w8(32'hb61276b4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37328227),
	.w1(32'hb686c0cc),
	.w2(32'hb8004dd1),
	.w3(32'h355b924d),
	.w4(32'h35fa610a),
	.w5(32'hb668739f),
	.w6(32'hb6880fff),
	.w7(32'h38188b1a),
	.w8(32'h383efcd8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792fb5c),
	.w1(32'hb5cfbe87),
	.w2(32'h36cea234),
	.w3(32'hb6e44e3b),
	.w4(32'hb7196071),
	.w5(32'hb707e0e7),
	.w6(32'h36fc70b9),
	.w7(32'h37b4c29b),
	.w8(32'h3663e3e3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736f2d1),
	.w1(32'hb7592159),
	.w2(32'hb7812320),
	.w3(32'h371c7450),
	.w4(32'hb75b0555),
	.w5(32'hb690e58e),
	.w6(32'h36f1c1cb),
	.w7(32'hb758d4ed),
	.w8(32'h37ae57dd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da78fd),
	.w1(32'hb706af2e),
	.w2(32'h377ad0b3),
	.w3(32'hb791737b),
	.w4(32'hb767697f),
	.w5(32'h3541a895),
	.w6(32'h38157066),
	.w7(32'hb79fe47c),
	.w8(32'hb6b1b2c5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71289dc),
	.w1(32'h372a6c28),
	.w2(32'hb6afc86d),
	.w3(32'h364bdf4b),
	.w4(32'h369a7930),
	.w5(32'h3743e319),
	.w6(32'hb75c92c6),
	.w7(32'hb7419b71),
	.w8(32'h35f90758),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3703b58a),
	.w1(32'hb73c516b),
	.w2(32'hb6ba5a7b),
	.w3(32'h37b37beb),
	.w4(32'hb795d217),
	.w5(32'hb7a911f6),
	.w6(32'h3601938f),
	.w7(32'hb749e931),
	.w8(32'h37017e79),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b9cc2b),
	.w1(32'h371459e4),
	.w2(32'h36fb8a9a),
	.w3(32'hb780c44e),
	.w4(32'hb6c4c113),
	.w5(32'hb66dc788),
	.w6(32'hb738f44a),
	.w7(32'hb6187f83),
	.w8(32'hb7debe92),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c3918),
	.w1(32'hb6f2877a),
	.w2(32'h36408948),
	.w3(32'h35e3e83b),
	.w4(32'hb7295571),
	.w5(32'hb7874d4d),
	.w6(32'hb5ea0177),
	.w7(32'hb6d9d8a3),
	.w8(32'h37494cb2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb784aab0),
	.w1(32'hb716bd9f),
	.w2(32'h37c1128b),
	.w3(32'hb80cb53e),
	.w4(32'hb75c3c31),
	.w5(32'hb712bce6),
	.w6(32'hb704f7a1),
	.w7(32'hb7c13cc6),
	.w8(32'h36d401a4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ba317),
	.w1(32'hb5fc929a),
	.w2(32'h37eb3a4f),
	.w3(32'hb7a4e140),
	.w4(32'hb725660b),
	.w5(32'h37403b00),
	.w6(32'h356c75c8),
	.w7(32'hb7308ec5),
	.w8(32'hb69b50da),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f19e16),
	.w1(32'hb71f8c25),
	.w2(32'hb616fdd1),
	.w3(32'h35e54d74),
	.w4(32'hb65607b6),
	.w5(32'hb68ea8f5),
	.w6(32'hb7898828),
	.w7(32'hb7969d68),
	.w8(32'hb5aca670),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f1ae6d),
	.w1(32'h37e2f5dd),
	.w2(32'h374d81c7),
	.w3(32'hb6e5cb8b),
	.w4(32'h375e0a75),
	.w5(32'hb6f6f8a1),
	.w6(32'hb79bc024),
	.w7(32'h36a524f9),
	.w8(32'hb6f4c0b8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a9c66a),
	.w1(32'h3795da22),
	.w2(32'h3794505a),
	.w3(32'h363908b6),
	.w4(32'h352dc046),
	.w5(32'h37205444),
	.w6(32'h36625723),
	.w7(32'h370e4f7a),
	.w8(32'hb6c1b790),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38050054),
	.w1(32'h37885215),
	.w2(32'h37eed8f9),
	.w3(32'h37927051),
	.w4(32'hb793c1b2),
	.w5(32'h37fe0bd3),
	.w6(32'hb7643565),
	.w7(32'hb7573d24),
	.w8(32'h3745eee8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6842a15),
	.w1(32'hb82bf055),
	.w2(32'h379d5b04),
	.w3(32'hb79e056d),
	.w4(32'hb7939243),
	.w5(32'h3765d2a4),
	.w6(32'h3657c19e),
	.w7(32'h36678101),
	.w8(32'h3726de91),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36db7c1e),
	.w1(32'hb78b9366),
	.w2(32'h354ce21b),
	.w3(32'hb780d995),
	.w4(32'hb6fbcd00),
	.w5(32'h35f9a2b5),
	.w6(32'h37f2a5b5),
	.w7(32'hb7363511),
	.w8(32'hb43ab7c2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0dd4c),
	.w1(32'hb7b06020),
	.w2(32'hb829bba8),
	.w3(32'hb76bdf92),
	.w4(32'hb75314c1),
	.w5(32'hb7c93865),
	.w6(32'hb7184ae8),
	.w7(32'hb7a51352),
	.w8(32'hb7ea4c40),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7867fb9),
	.w1(32'hb7aaa002),
	.w2(32'h37e84d11),
	.w3(32'h36cdb1f6),
	.w4(32'hb80d0022),
	.w5(32'h3790da59),
	.w6(32'hb6cdeb08),
	.w7(32'hb8480a8a),
	.w8(32'hb6cef2ea),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6298dea),
	.w1(32'hb7902c6e),
	.w2(32'h36a8c562),
	.w3(32'hb7724c20),
	.w4(32'hb72a6ea9),
	.w5(32'hb6a66b12),
	.w6(32'hb80e74a0),
	.w7(32'hb6a47ac1),
	.w8(32'hb7219a2e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab6781),
	.w1(32'h366f832b),
	.w2(32'h36c02988),
	.w3(32'hb51aa3bb),
	.w4(32'hb7ed95fb),
	.w5(32'hb7a46801),
	.w6(32'hb76c0e4b),
	.w7(32'hb8106754),
	.w8(32'hb4193ca2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b180b2),
	.w1(32'h35a65a7f),
	.w2(32'h3758dfe5),
	.w3(32'hb65f4d5b),
	.w4(32'hb6fa23f1),
	.w5(32'hb6321fbc),
	.w6(32'h378cde41),
	.w7(32'hb55986d3),
	.w8(32'h376e3853),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78aefc3),
	.w1(32'h35d09c4f),
	.w2(32'h369933e3),
	.w3(32'hb723baba),
	.w4(32'hb7015068),
	.w5(32'hb789e2ec),
	.w6(32'h371cc3ee),
	.w7(32'hb68a5a18),
	.w8(32'h37ffd817),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710edac),
	.w1(32'h3719ee1d),
	.w2(32'hb7845baf),
	.w3(32'hb56d447a),
	.w4(32'hb64831e9),
	.w5(32'hb6af69e4),
	.w6(32'h385ab8d8),
	.w7(32'hb733cd96),
	.w8(32'h37976153),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78df63a),
	.w1(32'h37a6cb0f),
	.w2(32'hb7ab8432),
	.w3(32'hb7600878),
	.w4(32'h374d0a67),
	.w5(32'hb7c73d92),
	.w6(32'h37843ebd),
	.w7(32'h37979ead),
	.w8(32'h36a3a710),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79febb0),
	.w1(32'hb6bf26b2),
	.w2(32'hb62cb355),
	.w3(32'hb66ea8bc),
	.w4(32'hb700b634),
	.w5(32'h372beaef),
	.w6(32'hb6a2d886),
	.w7(32'h3610af4a),
	.w8(32'h3601ccf8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370bbab1),
	.w1(32'hb4517d7e),
	.w2(32'hb7cf087f),
	.w3(32'h38018e2c),
	.w4(32'hb787476e),
	.w5(32'hb7913703),
	.w6(32'h356238a2),
	.w7(32'h3695dff2),
	.w8(32'hb73ad4b3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e3d280),
	.w1(32'h37d91434),
	.w2(32'hb7dbcdf9),
	.w3(32'h37d1f3fa),
	.w4(32'h36bc8b5c),
	.w5(32'hb7b95fdc),
	.w6(32'h37e41955),
	.w7(32'hb6d9614c),
	.w8(32'h34bbef05),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dcd2e8),
	.w1(32'h36cc1e27),
	.w2(32'hb78389b0),
	.w3(32'h381062b9),
	.w4(32'hb70b23fb),
	.w5(32'h36ff5780),
	.w6(32'h381b539c),
	.w7(32'hb735589b),
	.w8(32'h37963595),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37231b32),
	.w1(32'hb76509f5),
	.w2(32'h35db0835),
	.w3(32'h34914944),
	.w4(32'hb752b89a),
	.w5(32'h36df47d0),
	.w6(32'h37d9f562),
	.w7(32'hb80eb55a),
	.w8(32'hb6b77acc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3683179f),
	.w1(32'hb6ff71fe),
	.w2(32'h3547de9c),
	.w3(32'h377341a0),
	.w4(32'hb721668f),
	.w5(32'hb613d490),
	.w6(32'h368b3d2b),
	.w7(32'h3783a34e),
	.w8(32'hb71cc0ee),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c7e32e),
	.w1(32'hb66325a1),
	.w2(32'h367078ea),
	.w3(32'h3721339c),
	.w4(32'hb74ee2dc),
	.w5(32'hb7180399),
	.w6(32'hb6919df1),
	.w7(32'hb80083d4),
	.w8(32'h355418c8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3750e613),
	.w1(32'h364a4f2e),
	.w2(32'h37750a5d),
	.w3(32'h36937234),
	.w4(32'hb64bcd0d),
	.w5(32'hb5c90cb9),
	.w6(32'h377ba8a0),
	.w7(32'h36c3dd60),
	.w8(32'hb519d9fa),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a1f176),
	.w1(32'hb7a399c5),
	.w2(32'h36ae1fcb),
	.w3(32'hb6cb8a71),
	.w4(32'hb726c4ad),
	.w5(32'h3690e907),
	.w6(32'hb6a65de6),
	.w7(32'hb6f9ff28),
	.w8(32'hb6d15be7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ac29f),
	.w1(32'hb53e7d51),
	.w2(32'hb7e17605),
	.w3(32'h373ceab4),
	.w4(32'hb75131c1),
	.w5(32'hb71ecd24),
	.w6(32'hb746d08e),
	.w7(32'hb60b2ee6),
	.w8(32'hb74f8e9d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7459ee6),
	.w1(32'hb6e5e043),
	.w2(32'h363e6d64),
	.w3(32'hb622fbda),
	.w4(32'hb6909910),
	.w5(32'h360ceb3a),
	.w6(32'hb79ea722),
	.w7(32'h37a9110c),
	.w8(32'h38096ccc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359e4faa),
	.w1(32'hb792c164),
	.w2(32'hb6d57d4a),
	.w3(32'hb625f3f8),
	.w4(32'hb74b0369),
	.w5(32'h37b73d7b),
	.w6(32'h383805b3),
	.w7(32'hb66602ce),
	.w8(32'hb4971d0e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f65459),
	.w1(32'h379546ad),
	.w2(32'hb79f061a),
	.w3(32'hb73e23f9),
	.w4(32'h362324c9),
	.w5(32'hb810ba03),
	.w6(32'h371b24ce),
	.w7(32'h3627b988),
	.w8(32'hb4bf6fd4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a9b70c),
	.w1(32'h39b75c53),
	.w2(32'hbb93edf2),
	.w3(32'h37e6d460),
	.w4(32'hbae68448),
	.w5(32'h3a849c54),
	.w6(32'h380aae37),
	.w7(32'h39c810ef),
	.w8(32'hb97056b2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba858),
	.w1(32'hba4fba61),
	.w2(32'hbb209b13),
	.w3(32'h3b92a23b),
	.w4(32'h3a014f6a),
	.w5(32'h3b65640b),
	.w6(32'hba0363dd),
	.w7(32'hba4ba327),
	.w8(32'hbb35ae5d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804bf9),
	.w1(32'hbab28c33),
	.w2(32'hbb28f615),
	.w3(32'hbb869300),
	.w4(32'h396b4459),
	.w5(32'hbb908509),
	.w6(32'hbbb52083),
	.w7(32'h3b2e0ec6),
	.w8(32'h3b2049d2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acc81),
	.w1(32'h3aaed52e),
	.w2(32'hbbc0d36e),
	.w3(32'h3b543fd7),
	.w4(32'h3b83a911),
	.w5(32'hbc113f6c),
	.w6(32'h3bafa398),
	.w7(32'h3ade1079),
	.w8(32'hbbe493a8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fffbc),
	.w1(32'h3aede9ff),
	.w2(32'h392f0a42),
	.w3(32'hba803eb3),
	.w4(32'h3b38057a),
	.w5(32'h3a92f204),
	.w6(32'h3aa3142b),
	.w7(32'h3a1c8a50),
	.w8(32'hb9bf9519),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae87775),
	.w1(32'hba5fa885),
	.w2(32'hb839bba7),
	.w3(32'hbb069e93),
	.w4(32'h3ac78ee2),
	.w5(32'h3a29f395),
	.w6(32'hbb1d82c2),
	.w7(32'h3b89f6dc),
	.w8(32'h3b5f0e96),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7af2),
	.w1(32'hba1e76c7),
	.w2(32'h3aa3354b),
	.w3(32'h37f4afc5),
	.w4(32'h3acc0747),
	.w5(32'h3b085701),
	.w6(32'h3b98c128),
	.w7(32'h3b2ceea1),
	.w8(32'h3b961675),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62f370),
	.w1(32'hbb052ff2),
	.w2(32'hbba91999),
	.w3(32'h3b34e6ca),
	.w4(32'h3a3d749b),
	.w5(32'hbbb43ad7),
	.w6(32'h3b834a30),
	.w7(32'hbb20f010),
	.w8(32'hbbb3d33e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd860a9),
	.w1(32'hbbb87bf3),
	.w2(32'hbc23e196),
	.w3(32'hbaf199b5),
	.w4(32'hbb2b14b5),
	.w5(32'hbafb5427),
	.w6(32'hbc0598d1),
	.w7(32'hbb30c685),
	.w8(32'hbb83b2d0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b15cb),
	.w1(32'hbaec58c4),
	.w2(32'h3b15dd66),
	.w3(32'hbc26ce78),
	.w4(32'hba318d73),
	.w5(32'h3b833247),
	.w6(32'hbc05a970),
	.w7(32'hbb81e02d),
	.w8(32'h3a21a579),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b224681),
	.w1(32'h3a8c7a15),
	.w2(32'hbaae2d51),
	.w3(32'h3a83866c),
	.w4(32'hba657681),
	.w5(32'h3abb9df0),
	.w6(32'hbb21d5d1),
	.w7(32'hba8e0b8d),
	.w8(32'h3933bdcb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40397a),
	.w1(32'h3b78054f),
	.w2(32'h3bd3c390),
	.w3(32'h3aa5b150),
	.w4(32'h3baea262),
	.w5(32'h3bb25fa5),
	.w6(32'hbb522aa2),
	.w7(32'h3a8fb513),
	.w8(32'h3bd22a06),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6924c4),
	.w1(32'hbb8763dd),
	.w2(32'h394420ab),
	.w3(32'h3b0cdb46),
	.w4(32'hbbfd74bc),
	.w5(32'h3c6c787e),
	.w6(32'hb89ca2f9),
	.w7(32'hbb91c987),
	.w8(32'h3bc1ab28),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b827b11),
	.w1(32'hbaba62a9),
	.w2(32'hb995e45c),
	.w3(32'h3c0adcd6),
	.w4(32'hb9f21406),
	.w5(32'hbb23d33c),
	.w6(32'h3b876a6d),
	.w7(32'hbb914069),
	.w8(32'hbb8da87d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8feddb),
	.w1(32'hbb875f6c),
	.w2(32'hbba4c29f),
	.w3(32'hbb84d7ba),
	.w4(32'hbb120da8),
	.w5(32'hbaf466de),
	.w6(32'hbb8e2f5d),
	.w7(32'hbba08fb7),
	.w8(32'hbb766312),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb768380),
	.w1(32'hbb8bf704),
	.w2(32'hbb4c1064),
	.w3(32'hbc25ccd6),
	.w4(32'hbb1a7fd5),
	.w5(32'h3b9b8acc),
	.w6(32'hbc0410fb),
	.w7(32'h383d80be),
	.w8(32'h3a6d21c3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf8d40),
	.w1(32'h3b666e96),
	.w2(32'hbb8e2552),
	.w3(32'hbb9adbeb),
	.w4(32'h3b63aad8),
	.w5(32'hbb4e1287),
	.w6(32'hbb66e181),
	.w7(32'h3b4d08b2),
	.w8(32'hbc0d840f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe57c1),
	.w1(32'hbbb96c71),
	.w2(32'hbbf4d4ba),
	.w3(32'hbc2104ba),
	.w4(32'hbbfcfc1e),
	.w5(32'hbc26a9ec),
	.w6(32'hbb04275d),
	.w7(32'hbbd1fb09),
	.w8(32'hbb8604ac),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade443),
	.w1(32'h3a27dc46),
	.w2(32'hbaea4dc6),
	.w3(32'hbaf7b2f1),
	.w4(32'hbb02c56a),
	.w5(32'hbb69ced9),
	.w6(32'hbbc3a0ee),
	.w7(32'hba704e8a),
	.w8(32'h3a7a9c85),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16790),
	.w1(32'h3b3d5b35),
	.w2(32'h3b304d57),
	.w3(32'h3b8c164d),
	.w4(32'h3b3835e9),
	.w5(32'h3c4bd675),
	.w6(32'h3b32a2a2),
	.w7(32'hbb5a47df),
	.w8(32'h3bf6ac39),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18f466),
	.w1(32'hbb1763a8),
	.w2(32'h3a936847),
	.w3(32'h3ba33fe7),
	.w4(32'hbb74cf2e),
	.w5(32'h3b8c2d95),
	.w6(32'hb9e9d5ca),
	.w7(32'hbbedb26b),
	.w8(32'hbb56499f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b5253),
	.w1(32'h3aea3231),
	.w2(32'h3bd4631a),
	.w3(32'hbb8154f6),
	.w4(32'hbaa93140),
	.w5(32'h3c28a786),
	.w6(32'hbb30eccb),
	.w7(32'hba9cc735),
	.w8(32'h3b764584),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1dfc9),
	.w1(32'h3a75fe86),
	.w2(32'hba18eef0),
	.w3(32'hbb6c41e3),
	.w4(32'h3ae25794),
	.w5(32'h3b474af1),
	.w6(32'hbbbd28ed),
	.w7(32'h3b8180cc),
	.w8(32'h3bfb11ab),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac432c0),
	.w1(32'hbb8a98f9),
	.w2(32'hbac88236),
	.w3(32'hbab83873),
	.w4(32'hbbc5b1cc),
	.w5(32'hbbfa8089),
	.w6(32'h3c027747),
	.w7(32'h3baf312d),
	.w8(32'h3b59e64c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ad075),
	.w1(32'h3b30d531),
	.w2(32'h3acd576a),
	.w3(32'hbb8507a3),
	.w4(32'h3af8f809),
	.w5(32'hba4869ac),
	.w6(32'h3ad16729),
	.w7(32'h3b90fd63),
	.w8(32'h3b630309),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b255bab),
	.w1(32'h3a48c47f),
	.w2(32'h3b138a51),
	.w3(32'hbb902752),
	.w4(32'hbbc7d8fd),
	.w5(32'hbafd5f5d),
	.w6(32'h3b58c323),
	.w7(32'h3b847ac1),
	.w8(32'h3a35e8d8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0665dc),
	.w1(32'h3b2f2a59),
	.w2(32'h3a8abe90),
	.w3(32'hbae4f257),
	.w4(32'h3b6eefa2),
	.w5(32'h3b68f092),
	.w6(32'hbb5f33b4),
	.w7(32'h3c04c1f0),
	.w8(32'hbbc03449),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156789),
	.w1(32'hbb935eb2),
	.w2(32'hbb4ee20c),
	.w3(32'hbc534330),
	.w4(32'hbbdafc25),
	.w5(32'h3c152fb4),
	.w6(32'hbc372c7c),
	.w7(32'hbba0fba6),
	.w8(32'hbb4dbb28),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13bbc8),
	.w1(32'h38fa4c29),
	.w2(32'h3a8c7ab8),
	.w3(32'hbb9f3985),
	.w4(32'hbba0cc07),
	.w5(32'hbaac13af),
	.w6(32'hbafc1a43),
	.w7(32'hbabdea15),
	.w8(32'hba4f9894),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11ac93),
	.w1(32'h3b798fd4),
	.w2(32'h3bbaf476),
	.w3(32'hbaa4d092),
	.w4(32'h3996a33b),
	.w5(32'hbbbe37b0),
	.w6(32'hbb84f74e),
	.w7(32'hbb71c010),
	.w8(32'hbb90a37d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb27eb),
	.w1(32'h3b24bdac),
	.w2(32'h3b311064),
	.w3(32'hbbe405c5),
	.w4(32'hbb39f408),
	.w5(32'hbb615840),
	.w6(32'hbb7f7664),
	.w7(32'hbc0411ae),
	.w8(32'hbbe1ee7c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86762),
	.w1(32'h3a9fd9e0),
	.w2(32'h3ae4998a),
	.w3(32'hbbfff2f8),
	.w4(32'hbbac80ff),
	.w5(32'hb97250dd),
	.w6(32'hbb98954c),
	.w7(32'hbb69afa4),
	.w8(32'h39f434ef),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c0d4d),
	.w1(32'hbbb1824e),
	.w2(32'hbbd7b4b1),
	.w3(32'hbaa92e11),
	.w4(32'hbb6af6d4),
	.w5(32'h3abe86f7),
	.w6(32'hbb187911),
	.w7(32'hbb033b2b),
	.w8(32'hbb8b6f8f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba436240),
	.w1(32'hb8b8970e),
	.w2(32'h3a3d029a),
	.w3(32'hba2ffca6),
	.w4(32'hbb04a362),
	.w5(32'h3b857cd8),
	.w6(32'hbb826c91),
	.w7(32'h3b5f7429),
	.w8(32'hba03c2f0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6413f),
	.w1(32'hbbd3f6d4),
	.w2(32'h3b1e75b2),
	.w3(32'h3b95af6c),
	.w4(32'hbbf8ec76),
	.w5(32'h3bc11261),
	.w6(32'h3bbf6fe7),
	.w7(32'hbbb8b652),
	.w8(32'h3902a9f8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb41f),
	.w1(32'hba4ecb8d),
	.w2(32'h39d78596),
	.w3(32'h3b83b560),
	.w4(32'hbbe60c2a),
	.w5(32'hbbabcd1e),
	.w6(32'h3b154514),
	.w7(32'hbb7d16f4),
	.w8(32'h3ae3ad14),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dba995),
	.w1(32'h3b212e62),
	.w2(32'h3b6d34e4),
	.w3(32'hbad4f6e4),
	.w4(32'hbacdc215),
	.w5(32'h3b5328e4),
	.w6(32'h3ab2673f),
	.w7(32'hbaae107a),
	.w8(32'h3b3c90ce),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be71ff4),
	.w1(32'hba4edfeb),
	.w2(32'h3b3adac8),
	.w3(32'h3be0601f),
	.w4(32'h3a10e0a6),
	.w5(32'h3c532930),
	.w6(32'h3b9ea837),
	.w7(32'hbab20e9d),
	.w8(32'hb97d79c3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8752e),
	.w1(32'hbbfdaf0b),
	.w2(32'hbbe8efbe),
	.w3(32'h39f77086),
	.w4(32'hbc03df24),
	.w5(32'h3aa51aff),
	.w6(32'hbb25d18c),
	.w7(32'hbc552e5e),
	.w8(32'hbb9c24e9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca9e96),
	.w1(32'h3b84b902),
	.w2(32'h3abcb317),
	.w3(32'hbba8b884),
	.w4(32'h3aa8d9a9),
	.w5(32'hbb384bb7),
	.w6(32'hbb72fb8f),
	.w7(32'hbbc62517),
	.w8(32'hbb370b6b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b811ccb),
	.w1(32'h39063959),
	.w2(32'hbb4aebf7),
	.w3(32'h37071302),
	.w4(32'hbb11d660),
	.w5(32'hbc2b140e),
	.w6(32'hbb265fdc),
	.w7(32'h39e3c3d3),
	.w8(32'hba810867),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cdc5),
	.w1(32'hbab2badd),
	.w2(32'hba035864),
	.w3(32'h3aefa57e),
	.w4(32'hbb417057),
	.w5(32'h3ba8c2b2),
	.w6(32'hb906ec8b),
	.w7(32'hba974a17),
	.w8(32'hb9f1ceef),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa81c),
	.w1(32'hbabe2c17),
	.w2(32'hbb8e60d3),
	.w3(32'h3b1b710a),
	.w4(32'hbb4f25ef),
	.w5(32'h38bb22f5),
	.w6(32'h3be30a44),
	.w7(32'hbba57a50),
	.w8(32'hbbb0e7e5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0ee1),
	.w1(32'h3b262c0d),
	.w2(32'h3b1665e7),
	.w3(32'hbb2abfb0),
	.w4(32'h3ac68527),
	.w5(32'h3bf0ad01),
	.w6(32'hbb99bca8),
	.w7(32'hba3fbebc),
	.w8(32'h3b184b01),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba971472),
	.w1(32'h3a673cab),
	.w2(32'hba170e59),
	.w3(32'hbb249333),
	.w4(32'hbb850d9b),
	.w5(32'h3bf0cc6a),
	.w6(32'hbafc012a),
	.w7(32'h38fb1a7b),
	.w8(32'h3c10b801),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93578ca),
	.w1(32'h3c318b48),
	.w2(32'hbac6cbab),
	.w3(32'h3a00287e),
	.w4(32'h3c5a00fd),
	.w5(32'hbc3ecb09),
	.w6(32'hbb9d1cf7),
	.w7(32'h3ba43f57),
	.w8(32'hba428db1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972ad3),
	.w1(32'hbad1ac85),
	.w2(32'hbba4eded),
	.w3(32'h3bfbb7e4),
	.w4(32'hbb168ca0),
	.w5(32'h3b255b95),
	.w6(32'h3b1ff66e),
	.w7(32'hbb08bb5f),
	.w8(32'hbabacb6e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940696),
	.w1(32'h3a094d33),
	.w2(32'hbb6fce5f),
	.w3(32'hbbbe096d),
	.w4(32'h3b6c8088),
	.w5(32'hbb933e6d),
	.w6(32'hbbb38529),
	.w7(32'h3b22bcb5),
	.w8(32'hbaeb09fb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105f8e),
	.w1(32'h3b0905b5),
	.w2(32'h3bdca71b),
	.w3(32'h39bd38f3),
	.w4(32'hb9d1d8fe),
	.w5(32'h3b24f973),
	.w6(32'hbae4ee3c),
	.w7(32'h3bd1bcf4),
	.w8(32'h3bfc7835),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103f9f),
	.w1(32'hbb0527c2),
	.w2(32'hbb49f9d1),
	.w3(32'h3b216e4d),
	.w4(32'hbb230bba),
	.w5(32'hbba873a0),
	.w6(32'h3b3aa0ec),
	.w7(32'h3aa10a27),
	.w8(32'h3ab0dfd0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0158c),
	.w1(32'hbb444192),
	.w2(32'hbbd96265),
	.w3(32'hbbd879ed),
	.w4(32'hbbcc61f1),
	.w5(32'hbbca5cc1),
	.w6(32'h3b7a3a29),
	.w7(32'hbc3d42ee),
	.w8(32'hbc1970eb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393982f1),
	.w1(32'h39bca278),
	.w2(32'h3a8b2f20),
	.w3(32'h3b5657da),
	.w4(32'h3c1feffd),
	.w5(32'h3bc10dea),
	.w6(32'h3ba39ce5),
	.w7(32'h3b89323f),
	.w8(32'h3b9b8786),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d41f),
	.w1(32'hbb7db1d8),
	.w2(32'hba999edd),
	.w3(32'h3c103187),
	.w4(32'hbbafbbb8),
	.w5(32'h3b9f3278),
	.w6(32'hb9b6e658),
	.w7(32'hbc252f43),
	.w8(32'h3b9febbb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad89b4),
	.w1(32'hba5dbc66),
	.w2(32'hbb13f2a7),
	.w3(32'hbb592334),
	.w4(32'hba8fe7b0),
	.w5(32'h3bd22e32),
	.w6(32'h3b20c9c1),
	.w7(32'hb9ed3bcf),
	.w8(32'hbab4dc96),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf06050),
	.w1(32'hbb876c88),
	.w2(32'h38a80612),
	.w3(32'hbba90ed6),
	.w4(32'hbb91da8d),
	.w5(32'h3c3aa022),
	.w6(32'hbbf29c16),
	.w7(32'hbb70c7c3),
	.w8(32'hbad3f63c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43722d),
	.w1(32'hbb958e56),
	.w2(32'hba7b94c8),
	.w3(32'hb7099d35),
	.w4(32'hbba1b1fc),
	.w5(32'hbb8c35ae),
	.w6(32'hba077d69),
	.w7(32'h3b7b32dd),
	.w8(32'hba930b75),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042f6a),
	.w1(32'hbaff20d3),
	.w2(32'hbb5dfdde),
	.w3(32'hb9bd2d6b),
	.w4(32'hbb41a728),
	.w5(32'h399653f9),
	.w6(32'hba59cf4d),
	.w7(32'hbb02b5ef),
	.w8(32'h3a644301),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12f441),
	.w1(32'h3b291041),
	.w2(32'h3a8f183d),
	.w3(32'h3bcdfd90),
	.w4(32'h3bb08db5),
	.w5(32'h3abe1997),
	.w6(32'h3b320231),
	.w7(32'h3be41876),
	.w8(32'h3bb49a89),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4974c2),
	.w1(32'h3af7df1c),
	.w2(32'hb9fe16e4),
	.w3(32'hbb53d852),
	.w4(32'h3b4a0729),
	.w5(32'h3b6228b5),
	.w6(32'h3b23a4f1),
	.w7(32'h3a7ac73b),
	.w8(32'hb90d47f3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule