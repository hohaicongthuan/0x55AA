module layer_8_featuremap_188(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a0466),
	.w1(32'hbb9bf880),
	.w2(32'hbd0d4c8a),
	.w3(32'h3cbe6504),
	.w4(32'h3c9e9656),
	.w5(32'hbc78b8cc),
	.w6(32'h3cf04109),
	.w7(32'h3b81a217),
	.w8(32'hbc922f4a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2486d),
	.w1(32'hb9523acd),
	.w2(32'h3b7ef52f),
	.w3(32'hbcad64f8),
	.w4(32'h3b9e7865),
	.w5(32'h3c2c6250),
	.w6(32'h3ba87f0d),
	.w7(32'hbb08854f),
	.w8(32'h3b3724d4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dbde5),
	.w1(32'h3962ee1c),
	.w2(32'hbc079d7c),
	.w3(32'h3bc2a26a),
	.w4(32'hbc3b9f83),
	.w5(32'hbd0e22f5),
	.w6(32'h3cca815f),
	.w7(32'h3c3a2e79),
	.w8(32'h3c4bdd23),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2716),
	.w1(32'h3bd39637),
	.w2(32'h3bbfd824),
	.w3(32'hbcb32498),
	.w4(32'h3b8d206d),
	.w5(32'hbcee5470),
	.w6(32'h3cd9249c),
	.w7(32'h3c507d1d),
	.w8(32'h3ca3d8e2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9069d13),
	.w1(32'h3acf9986),
	.w2(32'h3b3e03fc),
	.w3(32'hbc8db16b),
	.w4(32'h3c01eaec),
	.w5(32'h3c56644e),
	.w6(32'h3c092afb),
	.w7(32'h3b7d83fc),
	.w8(32'h3ba63525),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a39de),
	.w1(32'hbc2f273a),
	.w2(32'h3c407cf6),
	.w3(32'hbc551e16),
	.w4(32'hbb289816),
	.w5(32'h3c1c3ad3),
	.w6(32'hbc4ac586),
	.w7(32'hbc30af4b),
	.w8(32'h3c59715d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb055f0),
	.w1(32'h3b52f149),
	.w2(32'h3b932727),
	.w3(32'hbcc42709),
	.w4(32'h39ebb4f0),
	.w5(32'h3b8bfe00),
	.w6(32'h3ab3e887),
	.w7(32'h3ba90903),
	.w8(32'h3b539431),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab470cd),
	.w1(32'hbc340554),
	.w2(32'hbb590010),
	.w3(32'h3c1de274),
	.w4(32'hbc4fdc4a),
	.w5(32'hbc13f8fd),
	.w6(32'h3c20d028),
	.w7(32'h3b828f6b),
	.w8(32'h3bae39a2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a93fa),
	.w1(32'hba4043c5),
	.w2(32'hbb63b083),
	.w3(32'h3cbcb280),
	.w4(32'h3c509d7d),
	.w5(32'h3c2cb057),
	.w6(32'h3c522e13),
	.w7(32'hbaf30eb4),
	.w8(32'hbbbeb04a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994eefa),
	.w1(32'hbc38873b),
	.w2(32'hbd4cae23),
	.w3(32'h3ca18919),
	.w4(32'hbc909b35),
	.w5(32'hbd352f20),
	.w6(32'h3cfcba7f),
	.w7(32'h3b82ca51),
	.w8(32'hbaede80a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf9e1a),
	.w1(32'hbc403f15),
	.w2(32'hb88facfe),
	.w3(32'hbc306e54),
	.w4(32'hbaf19df6),
	.w5(32'h3c05ea66),
	.w6(32'h3c7d68db),
	.w7(32'h3c133f10),
	.w8(32'hbb82e84e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4953c5),
	.w1(32'hbb399967),
	.w2(32'hbc72ec63),
	.w3(32'h3cc328f7),
	.w4(32'hb9dc9646),
	.w5(32'hbc10040d),
	.w6(32'h3c647a89),
	.w7(32'hbbd6613b),
	.w8(32'h3afc29a0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18468f),
	.w1(32'hbb0178c8),
	.w2(32'h3b15fbfd),
	.w3(32'h3a9db7e0),
	.w4(32'h3a6cdcca),
	.w5(32'h39ccf725),
	.w6(32'hb9aa84b5),
	.w7(32'hbad7ba5d),
	.w8(32'h3bdae9a5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb502eab),
	.w1(32'h3c8675a5),
	.w2(32'hbaa86a36),
	.w3(32'hbc3da522),
	.w4(32'h3bd57829),
	.w5(32'hbd032d20),
	.w6(32'h3cce4f2d),
	.w7(32'h3cc9c3f8),
	.w8(32'h3c3bb24f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0906),
	.w1(32'hbb01f630),
	.w2(32'hbbad365b),
	.w3(32'hbccf80f3),
	.w4(32'hbb8b91c9),
	.w5(32'hbbcdd69e),
	.w6(32'hba33e54f),
	.w7(32'hbae88a13),
	.w8(32'hb90f0208),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783c284),
	.w1(32'h3c339505),
	.w2(32'h3c0f3391),
	.w3(32'hbb41d002),
	.w4(32'h3c918f8f),
	.w5(32'h3cd0a117),
	.w6(32'hbbe457d5),
	.w7(32'hbba96a84),
	.w8(32'hbc122b03),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083a0e),
	.w1(32'h3b728b7c),
	.w2(32'hbc8b61df),
	.w3(32'hbbf3f4fa),
	.w4(32'hbb82953a),
	.w5(32'hbc8c08ec),
	.w6(32'h3b172e41),
	.w7(32'hbb95489e),
	.w8(32'hbb4296cf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc9ced),
	.w1(32'hbbaeb52e),
	.w2(32'hbb13b877),
	.w3(32'hbbadf797),
	.w4(32'h3a7249aa),
	.w5(32'h3bc5bc54),
	.w6(32'h3c325aa8),
	.w7(32'h3ba19537),
	.w8(32'h3cd5340f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccf6c1),
	.w1(32'hbd16e210),
	.w2(32'hbd4b8591),
	.w3(32'h3d578647),
	.w4(32'h3ba6d4ee),
	.w5(32'hbbf73aaa),
	.w6(32'h3d342960),
	.w7(32'hbc72c14c),
	.w8(32'hbd3708fc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c912a5b),
	.w1(32'hbc685836),
	.w2(32'hbc10c8d5),
	.w3(32'h3d0e5605),
	.w4(32'hbae6f9eb),
	.w5(32'hbaf716a9),
	.w6(32'h3cecb2e6),
	.w7(32'h3c5d5a7b),
	.w8(32'h3c28be5f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cbd43),
	.w1(32'hbc7feb65),
	.w2(32'hbc163c78),
	.w3(32'h3970060a),
	.w4(32'hbbe240ce),
	.w5(32'h3988802e),
	.w6(32'hbcdb20ef),
	.w7(32'hbbe50b9c),
	.w8(32'hb9b43f39),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e3bf),
	.w1(32'h3c2bd006),
	.w2(32'h3c05f218),
	.w3(32'hbbbdb8c5),
	.w4(32'h3b4293b0),
	.w5(32'hbc1a7f28),
	.w6(32'h3c32ce3b),
	.w7(32'h3c2fdd68),
	.w8(32'h3c462b18),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c68d9),
	.w1(32'hbbffb47b),
	.w2(32'hbd87b8dc),
	.w3(32'h3d39e217),
	.w4(32'h3c86f69e),
	.w5(32'hbd4b2fd6),
	.w6(32'h3d559fbb),
	.w7(32'h3b7eec59),
	.w8(32'hbc8b9c49),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38ac16),
	.w1(32'hbb38aa8a),
	.w2(32'hb9e23252),
	.w3(32'h3c12ca80),
	.w4(32'h38b6adb8),
	.w5(32'hbc4475ef),
	.w6(32'h3c51edad),
	.w7(32'h3c333ba6),
	.w8(32'h3c1fce6e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5ab4),
	.w1(32'hbb318ff8),
	.w2(32'hbc74d9dd),
	.w3(32'hbbc317a4),
	.w4(32'hbbb1699b),
	.w5(32'hbc9e58c3),
	.w6(32'h3bb69b4c),
	.w7(32'hbaed9ba0),
	.w8(32'hbaa6ce3b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147f26),
	.w1(32'h3aebb8e3),
	.w2(32'hbcccc8e7),
	.w3(32'h3ca71752),
	.w4(32'h3cb58876),
	.w5(32'hbbcc6999),
	.w6(32'h3d01946c),
	.w7(32'h3bb67b2e),
	.w8(32'hbb5db5a7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9fde1),
	.w1(32'h3a775596),
	.w2(32'h3bb58549),
	.w3(32'hbbfa8810),
	.w4(32'hbbd0b4ca),
	.w5(32'hbcf01526),
	.w6(32'hbb2ebd16),
	.w7(32'h3b3e9a05),
	.w8(32'h3ba55b7b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86193d),
	.w1(32'hbd588d8f),
	.w2(32'hbda1ebd6),
	.w3(32'h3d91d682),
	.w4(32'hbc55e5e1),
	.w5(32'h3c62e022),
	.w6(32'h3db68a52),
	.w7(32'h3d2ce099),
	.w8(32'h3b3dd05c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c661c60),
	.w1(32'hbbc54560),
	.w2(32'hbc82b7d4),
	.w3(32'h3d135e08),
	.w4(32'h3bb7972a),
	.w5(32'hbc21cd02),
	.w6(32'h3c8d3b37),
	.w7(32'h3ba8eabe),
	.w8(32'h3b67c5c6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4d6db),
	.w1(32'hba447a43),
	.w2(32'h3b422727),
	.w3(32'h3b016918),
	.w4(32'h3cc6138c),
	.w5(32'h3cbe9d86),
	.w6(32'h3b36ebc0),
	.w7(32'h3b8f8637),
	.w8(32'hbaf331d1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f38b),
	.w1(32'h3b62fb15),
	.w2(32'hbc606b6f),
	.w3(32'h3c5a43a3),
	.w4(32'hbb5e4c53),
	.w5(32'hbc2ffbed),
	.w6(32'h3b73daee),
	.w7(32'hb9fe90c7),
	.w8(32'hba926898),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2540bc),
	.w1(32'hbb2ba233),
	.w2(32'h3ba085f2),
	.w3(32'hbbba790c),
	.w4(32'h3b19cd34),
	.w5(32'h3c42ecb6),
	.w6(32'hbadc99e9),
	.w7(32'hb8ba84ea),
	.w8(32'h3bcd8423),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37f4dd),
	.w1(32'h3b74f75c),
	.w2(32'h3ba49976),
	.w3(32'h3b36052e),
	.w4(32'h3a67304a),
	.w5(32'hbafbe015),
	.w6(32'h3b44b50b),
	.w7(32'hbb0f7403),
	.w8(32'hbb5126ff),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40458c),
	.w1(32'h3c3ab4d1),
	.w2(32'h3b9c1892),
	.w3(32'h3aac8f32),
	.w4(32'h3bfb7b40),
	.w5(32'h3c07c259),
	.w6(32'h3bd1a09f),
	.w7(32'h3c659280),
	.w8(32'h3b106daa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35eb52),
	.w1(32'h3c086c35),
	.w2(32'h3bf9a05d),
	.w3(32'hbc1a4835),
	.w4(32'h3a1d6f66),
	.w5(32'h3bc08041),
	.w6(32'hbb8c55c5),
	.w7(32'hbbdd4a58),
	.w8(32'hbac72709),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb174c9),
	.w1(32'hbb8c7b5d),
	.w2(32'hbca0fc33),
	.w3(32'h3c2edeb4),
	.w4(32'hbbdc8f4d),
	.w5(32'hbc9ceab4),
	.w6(32'h3c073014),
	.w7(32'hbbdd76da),
	.w8(32'hbc62f8ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f6dd3),
	.w1(32'h3b7b67b5),
	.w2(32'h3bbeca50),
	.w3(32'hbc2bd9be),
	.w4(32'h3b69dd5f),
	.w5(32'h3b9febd4),
	.w6(32'h3ab4a6ac),
	.w7(32'h3b84dc7f),
	.w8(32'h3bea467a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9842),
	.w1(32'h3bbffcfb),
	.w2(32'h3bf89a80),
	.w3(32'h3c288832),
	.w4(32'h3bc96228),
	.w5(32'h3bfd3d90),
	.w6(32'h3c2dbc9d),
	.w7(32'h3ba7b26b),
	.w8(32'h3c018119),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b590d08),
	.w1(32'h3b83f7ea),
	.w2(32'h3bba3063),
	.w3(32'h3ba6c5fb),
	.w4(32'h3be0b508),
	.w5(32'h3c76875b),
	.w6(32'hb9adbd3d),
	.w7(32'hbab520cb),
	.w8(32'h3c1482dc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fff15),
	.w1(32'h3bd7105a),
	.w2(32'hba6a6b06),
	.w3(32'h3ab429e5),
	.w4(32'h3b47a080),
	.w5(32'hbad39c15),
	.w6(32'h3b300291),
	.w7(32'h3bde0021),
	.w8(32'h3c35c73b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d030302),
	.w1(32'hbc077041),
	.w2(32'hbc029dd1),
	.w3(32'h3d82888b),
	.w4(32'h3cbdde13),
	.w5(32'h3ca4f8a4),
	.w6(32'h3d7ef19c),
	.w7(32'h3ca4255f),
	.w8(32'h3cfc1549),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9edf39),
	.w1(32'hbad83951),
	.w2(32'h3b64f058),
	.w3(32'h3bf916cf),
	.w4(32'h3c05ab3a),
	.w5(32'h3c88360e),
	.w6(32'hbb57831f),
	.w7(32'hbc03bb00),
	.w8(32'hbc23f64e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc6b9e),
	.w1(32'hbab314ae),
	.w2(32'h3ab80394),
	.w3(32'h3c432f70),
	.w4(32'hba440184),
	.w5(32'h3b4f26b6),
	.w6(32'hbb15305a),
	.w7(32'h3b2d0a31),
	.w8(32'h3b2a6667),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca08c),
	.w1(32'hba800f08),
	.w2(32'hbace97a5),
	.w3(32'h3c7e3357),
	.w4(32'h38b83526),
	.w5(32'h3c562241),
	.w6(32'h3c6a7321),
	.w7(32'h3baf842e),
	.w8(32'h3bb19c0a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5011),
	.w1(32'hbcb6383b),
	.w2(32'hbd364cf4),
	.w3(32'h3ce7db55),
	.w4(32'hbc0d4727),
	.w5(32'hbd02e798),
	.w6(32'h3cb672a3),
	.w7(32'hbc31c951),
	.w8(32'hbcb3722a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3acf73),
	.w1(32'hbc202e07),
	.w2(32'hbc1a0172),
	.w3(32'h3aa30c14),
	.w4(32'hbbb147be),
	.w5(32'hbb9f3aae),
	.w6(32'h3b69aaab),
	.w7(32'hbbb067f7),
	.w8(32'hbc0e26bc),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad943d2),
	.w1(32'hbbc7401f),
	.w2(32'hbc3c43ea),
	.w3(32'h3ac61bfb),
	.w4(32'hbb9f8875),
	.w5(32'hbc62565f),
	.w6(32'hbb2805b6),
	.w7(32'h3b21e234),
	.w8(32'h3b76f3cb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f67bf),
	.w1(32'h3a4cb344),
	.w2(32'hbca99560),
	.w3(32'h3b60310e),
	.w4(32'h3ae301e3),
	.w5(32'hbc34a595),
	.w6(32'h3cb0351b),
	.w7(32'h3bdf5622),
	.w8(32'hbc1576ad),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4563c),
	.w1(32'hba70646d),
	.w2(32'hbc47590e),
	.w3(32'h3c0a7c2e),
	.w4(32'hbb44a2ae),
	.w5(32'hbc3d0ee3),
	.w6(32'h3c3a5487),
	.w7(32'h3be7b3b5),
	.w8(32'h3be191f5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04549f),
	.w1(32'h3b3daa9d),
	.w2(32'h3c34d3c9),
	.w3(32'hbbb4ea1f),
	.w4(32'h3cc3a26a),
	.w5(32'h3ce8f062),
	.w6(32'h3c4aee1c),
	.w7(32'h3c43d0b7),
	.w8(32'h3c99b8d0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd76bc9),
	.w1(32'h3c1cefd5),
	.w2(32'h3c7ff215),
	.w3(32'h3cd761b4),
	.w4(32'hbb78060b),
	.w5(32'h3c5f1448),
	.w6(32'h3b6de820),
	.w7(32'hbc617574),
	.w8(32'h3c52a4b3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff8de7),
	.w1(32'hbce8f8c1),
	.w2(32'hbcfcfc9f),
	.w3(32'h3d2c006a),
	.w4(32'hbbdad020),
	.w5(32'hbc8785f2),
	.w6(32'h3d681987),
	.w7(32'h3c90c85b),
	.w8(32'hbb11b1a0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00481d),
	.w1(32'hbb21579b),
	.w2(32'hbc0c160b),
	.w3(32'h3c9f1ac2),
	.w4(32'h3bf6b5a5),
	.w5(32'hbaa83057),
	.w6(32'h3cc91b68),
	.w7(32'h3c169c2d),
	.w8(32'h3b1a8074),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c532d42),
	.w1(32'hbb3b7281),
	.w2(32'hbc38712e),
	.w3(32'h3ccf543b),
	.w4(32'h3ba27a8e),
	.w5(32'hbc14efa8),
	.w6(32'h3c462126),
	.w7(32'h3a85df17),
	.w8(32'hbbd92f8b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babb5cf),
	.w1(32'hbb2be8e9),
	.w2(32'h3c4a25e2),
	.w3(32'h3c871b4f),
	.w4(32'h3aaf762c),
	.w5(32'h3c3ab421),
	.w6(32'h3bde104f),
	.w7(32'h3bf74b8f),
	.w8(32'h3c072a9b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf53c3d),
	.w1(32'h3bb4c892),
	.w2(32'hbc10c3dd),
	.w3(32'h3d036e8c),
	.w4(32'hbbe5424e),
	.w5(32'hbc5cd3f1),
	.w6(32'h3cb79a54),
	.w7(32'h3b7dfd61),
	.w8(32'hbc902280),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4178c9),
	.w1(32'h3be23c51),
	.w2(32'hbc7df916),
	.w3(32'h3c26f5b4),
	.w4(32'hbb065a0e),
	.w5(32'hbc78176b),
	.w6(32'h3c0ba632),
	.w7(32'h3bc1c9e5),
	.w8(32'h3c2ae51c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4b29b),
	.w1(32'hbc11dc17),
	.w2(32'hbbced80f),
	.w3(32'h3cbea6d7),
	.w4(32'h3a87f21a),
	.w5(32'h3a8ba000),
	.w6(32'h3c8a2c08),
	.w7(32'h3b668e67),
	.w8(32'h3b52fb3e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43f08),
	.w1(32'hbb041b86),
	.w2(32'hbc4ab6b0),
	.w3(32'h3c59bfe8),
	.w4(32'hba9b6be0),
	.w5(32'hbbbe496d),
	.w6(32'h3b3d6f39),
	.w7(32'h3771d8b0),
	.w8(32'hbbca43d7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff113d),
	.w1(32'h3bba7569),
	.w2(32'hbbad03e9),
	.w3(32'h3bbd4ce8),
	.w4(32'h3c1ce5c5),
	.w5(32'hbbb0c434),
	.w6(32'h3c4b325a),
	.w7(32'h3c710579),
	.w8(32'h3c8b10ab),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5004d4),
	.w1(32'hb9b33572),
	.w2(32'h3b83bd81),
	.w3(32'hbc192a90),
	.w4(32'hb91a09ea),
	.w5(32'hbc90a760),
	.w6(32'h3b8d4254),
	.w7(32'h3c09948f),
	.w8(32'h3c7aed82),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7266f),
	.w1(32'hbaf2c782),
	.w2(32'hbbd34805),
	.w3(32'hbc3fbbfe),
	.w4(32'h3ba60ae9),
	.w5(32'h3b8d6433),
	.w6(32'hbb8bc225),
	.w7(32'hbc31fad3),
	.w8(32'hbb56a4f9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9955a3),
	.w1(32'hbb36cc46),
	.w2(32'h3bc090b2),
	.w3(32'h3d1fd096),
	.w4(32'h3c15023b),
	.w5(32'h3c87376e),
	.w6(32'h3d1aa96d),
	.w7(32'h3bf208d2),
	.w8(32'h3c09402f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42288a),
	.w1(32'hbc2f7478),
	.w2(32'hbc60525d),
	.w3(32'h3c2bc65a),
	.w4(32'hbc8042fc),
	.w5(32'hbcc0ebcf),
	.w6(32'h3a6878fd),
	.w7(32'hbb8aed2d),
	.w8(32'hbb5f1f12),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb72f3),
	.w1(32'h3ba6bba3),
	.w2(32'h3b388513),
	.w3(32'hbc45ed0f),
	.w4(32'h3bf4e775),
	.w5(32'h3b83a8b3),
	.w6(32'h3baea6e7),
	.w7(32'h3b41d02d),
	.w8(32'h3b6dc61c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3c10),
	.w1(32'hbb52fc2c),
	.w2(32'hba6a2b38),
	.w3(32'h3bb07dee),
	.w4(32'h3b42f09b),
	.w5(32'hbb8b859f),
	.w6(32'h3c3d4fad),
	.w7(32'h3c014957),
	.w8(32'h3b4e0c5b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b6cf7),
	.w1(32'hbc391df1),
	.w2(32'hbc9acb88),
	.w3(32'h3c140b2d),
	.w4(32'hbc40155a),
	.w5(32'hbcac296e),
	.w6(32'hbb3ea791),
	.w7(32'hbbb7f9fe),
	.w8(32'hbbbd721e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795201),
	.w1(32'hbb43fdf7),
	.w2(32'hbc017062),
	.w3(32'hbc923fc4),
	.w4(32'hbba60938),
	.w5(32'hbc404b88),
	.w6(32'hbadec3d7),
	.w7(32'hbb153adb),
	.w8(32'hbaf93783),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52b5c),
	.w1(32'h3c6fea16),
	.w2(32'h37330fca),
	.w3(32'h3b9f1549),
	.w4(32'h3af0061e),
	.w5(32'hbb54f9d4),
	.w6(32'h3c82c5ea),
	.w7(32'h3c3d4248),
	.w8(32'h3b2a8ec2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52a225),
	.w1(32'h3bc8200f),
	.w2(32'hbd2842bb),
	.w3(32'h3c8e7486),
	.w4(32'h3bb78ed3),
	.w5(32'hbd134b3a),
	.w6(32'h3d49f3a2),
	.w7(32'h3d1399b4),
	.w8(32'h3b7b9c76),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a4fb),
	.w1(32'hbc0910de),
	.w2(32'h3aba1cb0),
	.w3(32'hbc8e3f6c),
	.w4(32'hbc63df79),
	.w5(32'hba9877d5),
	.w6(32'hbb19b3d2),
	.w7(32'hbb331629),
	.w8(32'hbb61696b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aeb93),
	.w1(32'hbb98eef4),
	.w2(32'hbcfa7249),
	.w3(32'h3c9c7ef5),
	.w4(32'hba86e882),
	.w5(32'hbcb1d8f4),
	.w6(32'h3cbf8d94),
	.w7(32'h3bf4f98d),
	.w8(32'h3b938965),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c3127),
	.w1(32'hbc2dacb2),
	.w2(32'hbce25204),
	.w3(32'hbcdaf9b2),
	.w4(32'hbc84f0b3),
	.w5(32'hbd12ae0a),
	.w6(32'hbab5fd1e),
	.w7(32'hbbaa978e),
	.w8(32'hbb45958b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44aa69),
	.w1(32'h357a2f60),
	.w2(32'h3b9d091a),
	.w3(32'hbcaf971b),
	.w4(32'h3c52b62f),
	.w5(32'h3bd4f265),
	.w6(32'h3c94f0ea),
	.w7(32'h3c49481d),
	.w8(32'h3c61f666),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9242288),
	.w1(32'hbb32c214),
	.w2(32'hbb41675b),
	.w3(32'hb828a547),
	.w4(32'h3a5be4b8),
	.w5(32'h3be2231e),
	.w6(32'hba7b84f4),
	.w7(32'h39a08d96),
	.w8(32'hbb8c9342),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9523a),
	.w1(32'h3bdb87de),
	.w2(32'hb918c935),
	.w3(32'h3c6d8ecb),
	.w4(32'h3cc4fe88),
	.w5(32'h3ca98136),
	.w6(32'h3ba52509),
	.w7(32'h3c44f0f4),
	.w8(32'h3c4c6bbf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199b7e),
	.w1(32'h39b756d5),
	.w2(32'hbb163b47),
	.w3(32'h3c868986),
	.w4(32'h3a552a5f),
	.w5(32'h3b1006e6),
	.w6(32'h3a9c68a5),
	.w7(32'hbab792a3),
	.w8(32'h3b9df604),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79d259),
	.w1(32'hbc167a78),
	.w2(32'hbc4c1a1e),
	.w3(32'h3d16c4a8),
	.w4(32'h3bc80841),
	.w5(32'hb91706d5),
	.w6(32'h3cc41e47),
	.w7(32'h3b60ff05),
	.w8(32'hbbb0dc8b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc0bf6),
	.w1(32'hbb899889),
	.w2(32'hbca7b73b),
	.w3(32'h3c575325),
	.w4(32'hbb9330b2),
	.w5(32'hbcaf37a4),
	.w6(32'h3c267a41),
	.w7(32'hbb5c4fc5),
	.w8(32'hbc85e6d6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d250e),
	.w1(32'h3bdd2df6),
	.w2(32'h3c18e8cc),
	.w3(32'hb95d121e),
	.w4(32'hbaf08077),
	.w5(32'h3b61b8c5),
	.w6(32'h3bc53b08),
	.w7(32'h3c27a55e),
	.w8(32'h3bf0f4af),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d87e8),
	.w1(32'h3bb691ca),
	.w2(32'hbc26a574),
	.w3(32'h3c467878),
	.w4(32'hbaf432c4),
	.w5(32'hbcb4bc40),
	.w6(32'h3c920300),
	.w7(32'h3bff2ca1),
	.w8(32'h3af1d57f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65e67d),
	.w1(32'h3c42d9cb),
	.w2(32'hbbcadc62),
	.w3(32'hbc8831f8),
	.w4(32'h3c9692dd),
	.w5(32'hbab9a032),
	.w6(32'h3cb6b637),
	.w7(32'h3c9b6aa7),
	.w8(32'h3c5ad925),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb31d59),
	.w1(32'hbc965820),
	.w2(32'hbc80d961),
	.w3(32'h3ca2e274),
	.w4(32'h3a884ea1),
	.w5(32'h3a7ed874),
	.w6(32'h3ccd30f4),
	.w7(32'h3b2c6eec),
	.w8(32'h3ae03ab1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d352ea7),
	.w1(32'h3a5239d6),
	.w2(32'h3c9ed966),
	.w3(32'h3d42654f),
	.w4(32'h3c1ec954),
	.w5(32'h3c734d80),
	.w6(32'h3d26cb9e),
	.w7(32'h3cf30986),
	.w8(32'h3d04f104),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b7c1b),
	.w1(32'hbb892d6f),
	.w2(32'hbd100369),
	.w3(32'h3d38dac7),
	.w4(32'h3c4c4c99),
	.w5(32'hbd17ced1),
	.w6(32'h3da6d115),
	.w7(32'h3d0fd5f2),
	.w8(32'h3c84b50d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c432fc8),
	.w1(32'h3c5c6a95),
	.w2(32'h3ca229cc),
	.w3(32'hba061779),
	.w4(32'h3c16beb1),
	.w5(32'hbc3cad7d),
	.w6(32'h3ce0fb25),
	.w7(32'h3d0b6fed),
	.w8(32'h3ca381a7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b49d9),
	.w1(32'hba0ecf0a),
	.w2(32'hbb128fe4),
	.w3(32'hbccc9e26),
	.w4(32'h3b41e2e2),
	.w5(32'h3bd3425e),
	.w6(32'hb98b1453),
	.w7(32'h3b0623f9),
	.w8(32'hbbe97d60),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94136d),
	.w1(32'h3a6b4811),
	.w2(32'h399a7bf0),
	.w3(32'h3a1496aa),
	.w4(32'hba6e0b63),
	.w5(32'hbb2db2c7),
	.w6(32'h3a188b1a),
	.w7(32'h3ac9e280),
	.w8(32'h3baa8695),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2bf6a),
	.w1(32'h3ab3565c),
	.w2(32'hbbe8b70d),
	.w3(32'h39c46ad5),
	.w4(32'hbb8753ef),
	.w5(32'hbc583310),
	.w6(32'h3bc7cdec),
	.w7(32'h3b8a20cc),
	.w8(32'hba24f414),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00ddd),
	.w1(32'h3a13f237),
	.w2(32'hbd0aea40),
	.w3(32'hbc1693d3),
	.w4(32'hbab178f1),
	.w5(32'hbd1867d2),
	.w6(32'h3c9668a4),
	.w7(32'h3c52683e),
	.w8(32'h3c474904),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9d19a),
	.w1(32'hbc3b2730),
	.w2(32'hbca86cdb),
	.w3(32'hbcac5f5b),
	.w4(32'hbbf1063b),
	.w5(32'hbc917cc3),
	.w6(32'h3c3d1736),
	.w7(32'hbb63ff4c),
	.w8(32'h3ba2b4c2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1acb0a),
	.w1(32'h3c7cad84),
	.w2(32'h3c866879),
	.w3(32'hbce06c9e),
	.w4(32'h3c36492a),
	.w5(32'h3bee8e94),
	.w6(32'h3be2572b),
	.w7(32'h3c2b065b),
	.w8(32'h3bac1cc6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8803f0),
	.w1(32'hbc2a3ffb),
	.w2(32'hba9ea523),
	.w3(32'h3bf85356),
	.w4(32'h3a9b1912),
	.w5(32'h3c328353),
	.w6(32'h3b2d9d66),
	.w7(32'h39e5273c),
	.w8(32'h3b8c8dfe),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda67ee),
	.w1(32'hbba57c23),
	.w2(32'hbbd2d5e9),
	.w3(32'h3c9a1cc5),
	.w4(32'h3b835d45),
	.w5(32'h3b129b53),
	.w6(32'h3c32d9d1),
	.w7(32'h3b432127),
	.w8(32'h3b5c4831),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81136e),
	.w1(32'h3b5a08bc),
	.w2(32'h3be405ef),
	.w3(32'hbab4b4b3),
	.w4(32'h3c05f9f3),
	.w5(32'h3c635213),
	.w6(32'hba580509),
	.w7(32'h3865f9d2),
	.w8(32'hbb04b013),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1b588),
	.w1(32'hbc1b4ec3),
	.w2(32'hbc843d91),
	.w3(32'h3c527ed4),
	.w4(32'hb996378f),
	.w5(32'hbc0b94b3),
	.w6(32'h3c483975),
	.w7(32'h3aed1049),
	.w8(32'hbb8705d2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c15e),
	.w1(32'hbb3b8563),
	.w2(32'hbc960d46),
	.w3(32'h3d09b56c),
	.w4(32'h3cd404c5),
	.w5(32'h3aaac4c7),
	.w6(32'h3d2984bd),
	.w7(32'h3c8d3fc5),
	.w8(32'h3c272e7c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17236e),
	.w1(32'hba378fd5),
	.w2(32'h3b3e408c),
	.w3(32'h3c2d2219),
	.w4(32'h3be7ced1),
	.w5(32'h3c3ab0ad),
	.w6(32'h39c24af6),
	.w7(32'hbab137dd),
	.w8(32'h3c1b3119),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b198ec9),
	.w1(32'h3b145c99),
	.w2(32'hbaab99d6),
	.w3(32'h3c2c205d),
	.w4(32'h3c0b1886),
	.w5(32'h3b691758),
	.w6(32'hbb22b18e),
	.w7(32'h3ad1159b),
	.w8(32'h3c46d093),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae08745),
	.w1(32'h3b543eff),
	.w2(32'hbb033fba),
	.w3(32'h3be5334f),
	.w4(32'hbc1d45c5),
	.w5(32'hbc722d41),
	.w6(32'h3c079fe4),
	.w7(32'h3bf6bedc),
	.w8(32'h3b34d11a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6fce),
	.w1(32'hbb4d3f0d),
	.w2(32'h3b4cdfdb),
	.w3(32'h3a94f8b4),
	.w4(32'hbc20281c),
	.w5(32'hbb878568),
	.w6(32'hbb23c092),
	.w7(32'h3c25e0b5),
	.w8(32'h3c3ffd0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9e87e),
	.w1(32'hbc88bdeb),
	.w2(32'hbc8a5599),
	.w3(32'h3ca4f5a8),
	.w4(32'hbb9dbb09),
	.w5(32'h3bf71a87),
	.w6(32'hbc2a5f5c),
	.w7(32'hbc9040a1),
	.w8(32'hbbf8570c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81dd64),
	.w1(32'h3c32db53),
	.w2(32'h3c027cc0),
	.w3(32'hba12d840),
	.w4(32'h3c26512e),
	.w5(32'hbb57fc06),
	.w6(32'h3bd0bae1),
	.w7(32'h3c28b5b5),
	.w8(32'h3b85fd56),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caadb8a),
	.w1(32'hbc8664d8),
	.w2(32'hbd052701),
	.w3(32'h3919b969),
	.w4(32'hbcbb2298),
	.w5(32'hbcdfdb0d),
	.w6(32'h3c837fac),
	.w7(32'h3a69eca5),
	.w8(32'hbb26ae3b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22319d),
	.w1(32'hbbba7a26),
	.w2(32'hbb8b58ba),
	.w3(32'hbc277b1f),
	.w4(32'h3b58d099),
	.w5(32'h3a2231c8),
	.w6(32'hbc579b9f),
	.w7(32'hbc90fbda),
	.w8(32'hbc53001d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9e570),
	.w1(32'hbc3bb8a7),
	.w2(32'hbcdd318e),
	.w3(32'h3c18ef08),
	.w4(32'h3ad01709),
	.w5(32'hbc38856f),
	.w6(32'h3ce063b4),
	.w7(32'h3c385ed0),
	.w8(32'hbb9186f0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ecb48),
	.w1(32'h3c3286b2),
	.w2(32'hbc428ded),
	.w3(32'h3c53a375),
	.w4(32'h3c3c0d6c),
	.w5(32'hbc4bb0c2),
	.w6(32'h3ca82eda),
	.w7(32'h3c7da902),
	.w8(32'h3bb9e095),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb61e9),
	.w1(32'h3b2e61f3),
	.w2(32'hbb64956c),
	.w3(32'hbbb49c48),
	.w4(32'h3be3d60b),
	.w5(32'h3b8910fa),
	.w6(32'h3bfda1c1),
	.w7(32'h390827c8),
	.w8(32'h3c7d15a6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1be27),
	.w1(32'hba3e8f65),
	.w2(32'h3c366257),
	.w3(32'hbbf7d126),
	.w4(32'h3907747e),
	.w5(32'h3c87f9a9),
	.w6(32'hbbded609),
	.w7(32'hbae29c4b),
	.w8(32'h3b6cbc86),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e60c),
	.w1(32'h3a95681a),
	.w2(32'h3acff44a),
	.w3(32'h3c76f0c8),
	.w4(32'h3c23e379),
	.w5(32'h3bcb09ef),
	.w6(32'h3c1ec630),
	.w7(32'h3b595c1e),
	.w8(32'h3b281c8a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29cf82),
	.w1(32'h3c22ffd0),
	.w2(32'h3be5a3bd),
	.w3(32'h3c415d5c),
	.w4(32'h3c732d0f),
	.w5(32'hb98e425a),
	.w6(32'h3ca2e9ef),
	.w7(32'h3c42958f),
	.w8(32'h3aeec237),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c542c62),
	.w1(32'hbb6d0151),
	.w2(32'h3b9cc039),
	.w3(32'h3b103719),
	.w4(32'h3b64e16c),
	.w5(32'h3c705dab),
	.w6(32'h3b8449d2),
	.w7(32'hbb96fb21),
	.w8(32'h3ba7f526),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2e8a6),
	.w1(32'hbb9c8f14),
	.w2(32'h3c62763a),
	.w3(32'hb99c50f0),
	.w4(32'hbc2734ac),
	.w5(32'h3bd7b0af),
	.w6(32'hbb5a578d),
	.w7(32'hba374fa2),
	.w8(32'hba051c7a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afffc53),
	.w1(32'hbc95006f),
	.w2(32'hbd386a82),
	.w3(32'hbb7683a3),
	.w4(32'hbca188d7),
	.w5(32'hbd055035),
	.w6(32'hbbcc8bb2),
	.w7(32'hbc485daa),
	.w8(32'hbb84f3d4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd92a06),
	.w1(32'h3bd75076),
	.w2(32'h3a81799c),
	.w3(32'hbc9237e5),
	.w4(32'h3c15fcb3),
	.w5(32'h3a4a7782),
	.w6(32'h3c01e681),
	.w7(32'h3c2443a3),
	.w8(32'h3b3a14f5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23cf56),
	.w1(32'h3a1e1f76),
	.w2(32'h3abd0712),
	.w3(32'hbb8c2887),
	.w4(32'h3bad4a60),
	.w5(32'h3b8e18ef),
	.w6(32'h3b11b837),
	.w7(32'hba33aa6b),
	.w8(32'hba8545c0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838d17),
	.w1(32'h3c022027),
	.w2(32'h3c2a2bce),
	.w3(32'h3b84c56c),
	.w4(32'h3c68ef18),
	.w5(32'h3c806833),
	.w6(32'h3b28aacd),
	.w7(32'h3adcb656),
	.w8(32'h3c1e8427),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3674),
	.w1(32'hbaa49f07),
	.w2(32'h3c1e7ff9),
	.w3(32'h3cadac12),
	.w4(32'h3acc52fd),
	.w5(32'h3bc6d824),
	.w6(32'h3c422def),
	.w7(32'hbbba295b),
	.w8(32'h3ac266fb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e688f),
	.w1(32'h3bc29a8a),
	.w2(32'hbc141d8a),
	.w3(32'hbbb10319),
	.w4(32'h3bb00c1b),
	.w5(32'hbc2feda0),
	.w6(32'h3c2aa13a),
	.w7(32'h393fa415),
	.w8(32'hbb515dee),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b381a),
	.w1(32'hbbe85312),
	.w2(32'hbc122f70),
	.w3(32'hbc6af072),
	.w4(32'hbbdac96e),
	.w5(32'hbbaa5532),
	.w6(32'hb9c7a8c8),
	.w7(32'hbbdb4e97),
	.w8(32'hbb90c809),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1290a0),
	.w1(32'h3aabf210),
	.w2(32'hbc13d325),
	.w3(32'h3ca24efa),
	.w4(32'h3bfc7c7a),
	.w5(32'hbc188e84),
	.w6(32'h3c801e8e),
	.w7(32'h3c461b29),
	.w8(32'h3b2dfdf3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108e0e),
	.w1(32'hbbb47919),
	.w2(32'hbbe4fcc4),
	.w3(32'hbb9828c7),
	.w4(32'hbada16c0),
	.w5(32'hbc8a6517),
	.w6(32'h3bab61aa),
	.w7(32'h3a3ee2d6),
	.w8(32'hbbd3b7f8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b861b),
	.w1(32'hbb326712),
	.w2(32'hba518a47),
	.w3(32'hbbaf7ea7),
	.w4(32'hb8ff9aa8),
	.w5(32'h3a9c88fd),
	.w6(32'hbb9a752f),
	.w7(32'hbbb2cbc1),
	.w8(32'hbba9b2c2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c647c),
	.w1(32'h3b9b4310),
	.w2(32'h3c55eb74),
	.w3(32'hbc25848f),
	.w4(32'hbb3cae2e),
	.w5(32'h3a4c674b),
	.w6(32'hbc191f4a),
	.w7(32'hbb452300),
	.w8(32'hbab035fe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6198),
	.w1(32'h3a88618e),
	.w2(32'hbc8acd78),
	.w3(32'h3b5f0792),
	.w4(32'h3bbef59b),
	.w5(32'hbcbbe6f8),
	.w6(32'h3c232660),
	.w7(32'hba08dad3),
	.w8(32'h3b185293),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9df22),
	.w1(32'hbac9db46),
	.w2(32'h3a1f3c56),
	.w3(32'hbcfeec75),
	.w4(32'hbbee7485),
	.w5(32'hbbb144a6),
	.w6(32'h3bc1d5f2),
	.w7(32'h3bc06a5b),
	.w8(32'h3a335883),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4839),
	.w1(32'hbb880cc8),
	.w2(32'hbbaa038f),
	.w3(32'h3ba1419e),
	.w4(32'hbb298d9b),
	.w5(32'hbb58f49b),
	.w6(32'h3aabeb07),
	.w7(32'hbbeeff8c),
	.w8(32'hbbc3ebb7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99650da),
	.w1(32'h39537fce),
	.w2(32'hbbb8c72a),
	.w3(32'h3b659326),
	.w4(32'h3bcbc0b1),
	.w5(32'h390aa9f1),
	.w6(32'h3b39097f),
	.w7(32'hb9c4bce0),
	.w8(32'hbbebfe42),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule