module layer_8_featuremap_46(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a18cd),
	.w1(32'h39b0150b),
	.w2(32'h3814a765),
	.w3(32'h3bb80e96),
	.w4(32'h3ada4109),
	.w5(32'hba5b8292),
	.w6(32'h3bf82089),
	.w7(32'h3b9a0311),
	.w8(32'h3b06e797),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad364e2),
	.w1(32'hbb1cc510),
	.w2(32'hbb821fe0),
	.w3(32'h3a01cc1c),
	.w4(32'hb9cacd07),
	.w5(32'hbac9cc9a),
	.w6(32'h3a5ec3c9),
	.w7(32'h397d7a52),
	.w8(32'h39463274),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e4ce),
	.w1(32'hba24d0b7),
	.w2(32'hb80932da),
	.w3(32'hbac39d80),
	.w4(32'h38365b9f),
	.w5(32'h3a42ed7a),
	.w6(32'hbadcf082),
	.w7(32'hba420d78),
	.w8(32'h3ab9cc8f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff678f),
	.w1(32'hba91f4a3),
	.w2(32'hba53e77c),
	.w3(32'h38fedc13),
	.w4(32'hb909b760),
	.w5(32'hbae4479e),
	.w6(32'h3a48b5be),
	.w7(32'h39eaa20e),
	.w8(32'hba1ae566),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24e9f5),
	.w1(32'hbc0644b8),
	.w2(32'hbbb9f2a6),
	.w3(32'hba83d974),
	.w4(32'hbb8ab963),
	.w5(32'hbb84e740),
	.w6(32'h3b04d7fa),
	.w7(32'hba91a90f),
	.w8(32'hbaf4329c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00ef79),
	.w1(32'h3b360d4d),
	.w2(32'h3b267ffb),
	.w3(32'hba9fade5),
	.w4(32'h3b0a8217),
	.w5(32'h3b513b67),
	.w6(32'hbb4d9234),
	.w7(32'hba7b2305),
	.w8(32'h37b7f267),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba234eee),
	.w1(32'hba1e701b),
	.w2(32'h36863b7d),
	.w3(32'hb9b8f5b3),
	.w4(32'hb9d22d76),
	.w5(32'hb934b4d2),
	.w6(32'hb74277e0),
	.w7(32'hb9ba5596),
	.w8(32'h37bf7ebd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b43ad),
	.w1(32'hbac6ce34),
	.w2(32'hbba5a1dc),
	.w3(32'h38cc8368),
	.w4(32'hbb2d56f8),
	.w5(32'hbbb721ef),
	.w6(32'h3b3308b3),
	.w7(32'hb988ae4f),
	.w8(32'hbb8f9af8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb136dd2),
	.w1(32'hbb8b90eb),
	.w2(32'hbb5755b8),
	.w3(32'h3af9b1b7),
	.w4(32'hbab6cd98),
	.w5(32'hbafb94c4),
	.w6(32'h3b6fb989),
	.w7(32'h3adbae4a),
	.w8(32'h3b1402d0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de1cd0),
	.w1(32'h3859340d),
	.w2(32'hbaf6c534),
	.w3(32'h3ac639c6),
	.w4(32'h3a3c5e55),
	.w5(32'hb9b0408f),
	.w6(32'h3a2dbb04),
	.w7(32'h3a9036ad),
	.w8(32'h3ade8e67),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9af871),
	.w1(32'hbb778937),
	.w2(32'hbb0c0571),
	.w3(32'h3b71737e),
	.w4(32'hb9781e85),
	.w5(32'hbb69657a),
	.w6(32'h3be98d8f),
	.w7(32'h3b84328b),
	.w8(32'hba8fe079),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906db71),
	.w1(32'hba4bc4e5),
	.w2(32'hba9ca09a),
	.w3(32'hb9e7fa9f),
	.w4(32'h39ae871d),
	.w5(32'hba637509),
	.w6(32'h3a4c70ce),
	.w7(32'h3b028b03),
	.w8(32'h3ad3a9bc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952fa3),
	.w1(32'hbb133c52),
	.w2(32'hbb7219f7),
	.w3(32'hbb40d7a1),
	.w4(32'hba7c73d5),
	.w5(32'hba4113ba),
	.w6(32'hbb55d06d),
	.w7(32'hbb031b72),
	.w8(32'h3a1004a7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f34ed),
	.w1(32'h3a39baf3),
	.w2(32'h3a6c525c),
	.w3(32'hba9a6ff3),
	.w4(32'hb984e889),
	.w5(32'h3a1088ed),
	.w6(32'hbaabe79f),
	.w7(32'hb9bbae13),
	.w8(32'h39ced63d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b09c28),
	.w1(32'hb9743935),
	.w2(32'hb94c3c33),
	.w3(32'hb99e6c85),
	.w4(32'hb9568643),
	.w5(32'hb90aa1a9),
	.w6(32'hb9a43f8d),
	.w7(32'hb94cea28),
	.w8(32'hb93da1d1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30ef1a),
	.w1(32'hb9d209f8),
	.w2(32'hb9119c05),
	.w3(32'hb98b4882),
	.w4(32'hba1b2fe1),
	.w5(32'hba639ca1),
	.w6(32'hb9d5dc49),
	.w7(32'hba9989e1),
	.w8(32'hba1739b3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0c3f),
	.w1(32'h3b81821c),
	.w2(32'h3b2e6fe9),
	.w3(32'h3b85af2a),
	.w4(32'h3b24ff61),
	.w5(32'h3abbd3fd),
	.w6(32'h3b2ef5fe),
	.w7(32'h3a2526d6),
	.w8(32'hb9b6a7dd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca8ad),
	.w1(32'hbb9005d3),
	.w2(32'hbb8c6a9d),
	.w3(32'hbaf00f6f),
	.w4(32'hbb06dac8),
	.w5(32'hba2e61f0),
	.w6(32'hbb0f744b),
	.w7(32'hbb06b9ce),
	.w8(32'h3aba6253),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee474),
	.w1(32'hbc38d339),
	.w2(32'hbb379f01),
	.w3(32'hbad6e072),
	.w4(32'hbc05acd7),
	.w5(32'hbc538b08),
	.w6(32'h3c681b90),
	.w7(32'h3a32f3a5),
	.w8(32'hbba4af36),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04a7dc),
	.w1(32'hbc88a064),
	.w2(32'hbc4ab5ab),
	.w3(32'hbb8dbf75),
	.w4(32'hbc13faa8),
	.w5(32'hbba8356b),
	.w6(32'h3ae6bdf5),
	.w7(32'hbb23a561),
	.w8(32'hbbb4aa7c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd45f7),
	.w1(32'h38d86a2f),
	.w2(32'h3ae44fc1),
	.w3(32'h3a22d018),
	.w4(32'h3b35bf5a),
	.w5(32'h3b8e1d16),
	.w6(32'hbaa9feb8),
	.w7(32'h3aea1183),
	.w8(32'h39d839d8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1471c7),
	.w1(32'hbaf1a6a6),
	.w2(32'hbbb5f690),
	.w3(32'hbc43fd53),
	.w4(32'hbb8239df),
	.w5(32'hba383c5e),
	.w6(32'hbc0ce624),
	.w7(32'hbb489090),
	.w8(32'hba2bfb78),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca76751),
	.w1(32'hba7413c8),
	.w2(32'hb90d9814),
	.w3(32'h3cb9608e),
	.w4(32'h3b9500de),
	.w5(32'hba592471),
	.w6(32'h3d053535),
	.w7(32'h3cbb545b),
	.w8(32'h3c23ccfb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164949),
	.w1(32'hbba413a4),
	.w2(32'hbbcee248),
	.w3(32'hba3fb404),
	.w4(32'hbb244cb2),
	.w5(32'hbb513f64),
	.w6(32'hb9a7a0b4),
	.w7(32'hbaef7b31),
	.w8(32'hbb3574ec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c680f32),
	.w1(32'h3c4f3785),
	.w2(32'h3c17150b),
	.w3(32'h3c46a7ee),
	.w4(32'h3c10158d),
	.w5(32'h3bfcef11),
	.w6(32'h3befd7d4),
	.w7(32'h3bb7c584),
	.w8(32'h3bcef306),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb38f60),
	.w1(32'hbbc46988),
	.w2(32'hbc0b60c5),
	.w3(32'h3bffd4c1),
	.w4(32'hbaf132e0),
	.w5(32'hbbd92258),
	.w6(32'h3c4eabb7),
	.w7(32'h3bf5e9b9),
	.w8(32'h39e6a8b8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f5a26),
	.w1(32'hb9409372),
	.w2(32'hba7e399c),
	.w3(32'h3a929d7f),
	.w4(32'hb82f95f2),
	.w5(32'hba93eb50),
	.w6(32'h3a68a0bb),
	.w7(32'h383ad158),
	.w8(32'hb9d2c365),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71a547),
	.w1(32'hbc1ac3c1),
	.w2(32'hbc6610d5),
	.w3(32'h3c0b679a),
	.w4(32'h3cd7c7fa),
	.w5(32'hbc2028c5),
	.w6(32'h3d5d6b23),
	.w7(32'h3da73247),
	.w8(32'h3bf98a03),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea5636),
	.w1(32'hbb115de9),
	.w2(32'hbb38a27c),
	.w3(32'h3b1341f5),
	.w4(32'hba167ec6),
	.w5(32'hbb10bada),
	.w6(32'h3b91ffe0),
	.w7(32'h3b6214a3),
	.w8(32'h3aa5d734),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d43d0),
	.w1(32'hba384a24),
	.w2(32'hb7f218a1),
	.w3(32'hba0ce6a0),
	.w4(32'hb8def287),
	.w5(32'h39b71901),
	.w6(32'hb9735642),
	.w7(32'hb8873dcf),
	.w8(32'hb9ad82f8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b8a9),
	.w1(32'h3a80aea1),
	.w2(32'h3ab8f793),
	.w3(32'hbb078f0b),
	.w4(32'h3811c59d),
	.w5(32'hb90769d8),
	.w6(32'hbbb24e17),
	.w7(32'hbb4fe5d8),
	.w8(32'hbb099519),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe6895),
	.w1(32'hbb0d1675),
	.w2(32'hbaeb4d17),
	.w3(32'hb99d7a1a),
	.w4(32'hbaed9f54),
	.w5(32'hbb084b77),
	.w6(32'h3ade1a71),
	.w7(32'hb8355f34),
	.w8(32'hba748340),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399afb48),
	.w1(32'h3911269c),
	.w2(32'h38c49b05),
	.w3(32'h39a885d0),
	.w4(32'h395a672c),
	.w5(32'h38e772b6),
	.w6(32'h39986136),
	.w7(32'h386c9107),
	.w8(32'hb8cf7c0b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcbcc7),
	.w1(32'hb907969e),
	.w2(32'hb8ba507d),
	.w3(32'hb8def6d0),
	.w4(32'hb9065713),
	.w5(32'hb89b8f81),
	.w6(32'h3636ca7f),
	.w7(32'hb860151b),
	.w8(32'hb6c4eebc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066519),
	.w1(32'hba987de5),
	.w2(32'hbab5c8d9),
	.w3(32'hbb21423f),
	.w4(32'hba9f5b01),
	.w5(32'h39ca5b55),
	.w6(32'hbbc60f54),
	.w7(32'hbba88630),
	.w8(32'hbb707030),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd245e5),
	.w1(32'h3a42a298),
	.w2(32'hbb870d52),
	.w3(32'h3bf5adbf),
	.w4(32'h3b332642),
	.w5(32'hbb7c53e7),
	.w6(32'h3bc649ae),
	.w7(32'h3b2891a8),
	.w8(32'hbb352835),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f08599),
	.w1(32'h399dd111),
	.w2(32'h3a8c4f9d),
	.w3(32'hb84537b1),
	.w4(32'h389a36f9),
	.w5(32'h3a8a67e3),
	.w6(32'h39607759),
	.w7(32'h39276f14),
	.w8(32'h3a944247),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44e8d8),
	.w1(32'hbb7d5f81),
	.w2(32'hbb5f5c6d),
	.w3(32'h381dc624),
	.w4(32'h38b6cd6b),
	.w5(32'h3a1c18d1),
	.w6(32'h3b1435c6),
	.w7(32'h3b74baeb),
	.w8(32'h3b854544),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed2559),
	.w1(32'hb94406ab),
	.w2(32'h38a0200e),
	.w3(32'h39108c4a),
	.w4(32'hb9b443e1),
	.w5(32'hb8baee64),
	.w6(32'hb9e70510),
	.w7(32'hb9d99fc7),
	.w8(32'hb9116214),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3d25),
	.w1(32'h3a4116d3),
	.w2(32'h3a5304a1),
	.w3(32'h3a32c045),
	.w4(32'h39db100d),
	.w5(32'h3a0e0fca),
	.w6(32'h391c433e),
	.w7(32'h39e151a8),
	.w8(32'h3a583605),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4577e1),
	.w1(32'hba8cf2d3),
	.w2(32'hbb8cf207),
	.w3(32'h3be75c4d),
	.w4(32'h3bb5913e),
	.w5(32'hb91c2471),
	.w6(32'h3b951f72),
	.w7(32'h3bdbd98c),
	.w8(32'h3b23a492),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14dd5f),
	.w1(32'hbb294aca),
	.w2(32'hbae2c03a),
	.w3(32'hbb0537d6),
	.w4(32'hbb427066),
	.w5(32'hbb74fc32),
	.w6(32'hbadec473),
	.w7(32'hbab504a2),
	.w8(32'hbb7c6f91),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233874),
	.w1(32'hba8a8aaf),
	.w2(32'hb9809206),
	.w3(32'hbb23ea68),
	.w4(32'hba27229b),
	.w5(32'hba8c3df7),
	.w6(32'h3965bd79),
	.w7(32'hb9995cd1),
	.w8(32'hba7697f5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38874c),
	.w1(32'h38f18844),
	.w2(32'hb83c8ea2),
	.w3(32'h3b56061b),
	.w4(32'h3ab95ee8),
	.w5(32'hba356014),
	.w6(32'h3b8df7c3),
	.w7(32'h3b58b262),
	.w8(32'h3a673304),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1a16),
	.w1(32'hbc283392),
	.w2(32'hbbd63dc6),
	.w3(32'hbc107d38),
	.w4(32'hbc3865a9),
	.w5(32'hbc2d4f3d),
	.w6(32'hb9ba9347),
	.w7(32'hbb639beb),
	.w8(32'hbc08988d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87002e),
	.w1(32'h3a986b75),
	.w2(32'h3a42aacd),
	.w3(32'h38d07a71),
	.w4(32'hb8d5cf50),
	.w5(32'hbac2e9bb),
	.w6(32'h3a3550c8),
	.w7(32'h3a573a2d),
	.w8(32'hbb1c28a5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9572a7),
	.w1(32'h3a8740bd),
	.w2(32'hbae61cd2),
	.w3(32'hbad1d1ab),
	.w4(32'h3a0d6f56),
	.w5(32'h3a5720ce),
	.w6(32'hbb04beca),
	.w7(32'hbac98442),
	.w8(32'hb98d1113),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fada7),
	.w1(32'hbc283201),
	.w2(32'hbb9431d2),
	.w3(32'hbb802f76),
	.w4(32'hbc04d902),
	.w5(32'hbc0360a4),
	.w6(32'h3b866ebf),
	.w7(32'h3aada907),
	.w8(32'hbaea1b9f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba406393),
	.w1(32'hb95c6aa1),
	.w2(32'hb8831d24),
	.w3(32'hb9f76d97),
	.w4(32'hb822412e),
	.w5(32'hb9ab95a3),
	.w6(32'h396297be),
	.w7(32'h3a042b1d),
	.w8(32'hba38a519),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb068f6),
	.w1(32'hbbd6c939),
	.w2(32'hbb873bb7),
	.w3(32'hbb94bb4a),
	.w4(32'hbb9a3a64),
	.w5(32'hbba3a096),
	.w6(32'hbabfb84e),
	.w7(32'hb9c8e295),
	.w8(32'hbb241f01),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78a2f3),
	.w1(32'hbacb1dd1),
	.w2(32'hbab2dbe3),
	.w3(32'hbb1662a4),
	.w4(32'h377914b0),
	.w5(32'h3ad8da28),
	.w6(32'h3988f2c4),
	.w7(32'h3b674779),
	.w8(32'h3bb58fb8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18a00a),
	.w1(32'hbc2cee44),
	.w2(32'hbb1e1c22),
	.w3(32'hbc1bb878),
	.w4(32'hbc9c6202),
	.w5(32'hbc387ea0),
	.w6(32'h3ac1cbb6),
	.w7(32'hbbb8c147),
	.w8(32'hbc251ed3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8e70),
	.w1(32'hbabb1dce),
	.w2(32'hbb2ac850),
	.w3(32'h3b098ef8),
	.w4(32'hbb01248b),
	.w5(32'hbaf99436),
	.w6(32'h3c26fb34),
	.w7(32'h3b5f7c4b),
	.w8(32'h3a3ff31e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9096dd7),
	.w1(32'hba19f55e),
	.w2(32'hbaf33be4),
	.w3(32'h3a93affc),
	.w4(32'h3a9a41c4),
	.w5(32'hbabf89f0),
	.w6(32'hb83056c6),
	.w7(32'hba02c0c9),
	.w8(32'hba894fd6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a257ef8),
	.w1(32'hba52cc8d),
	.w2(32'hbb0832ba),
	.w3(32'h38e05a8d),
	.w4(32'h3a137d7f),
	.w5(32'hba78de4a),
	.w6(32'h38ce7854),
	.w7(32'hbacad66f),
	.w8(32'hbaa34e9d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750c32),
	.w1(32'hbbe2d833),
	.w2(32'hbbbe735e),
	.w3(32'hba5ef5bc),
	.w4(32'hbbf7b8a6),
	.w5(32'hbc2fe109),
	.w6(32'h3b784d0b),
	.w7(32'h3ad6e475),
	.w8(32'hba694bca),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6de733),
	.w1(32'h3ad9e366),
	.w2(32'hb95130cd),
	.w3(32'h3a175a3f),
	.w4(32'h3a369875),
	.w5(32'h3a8a76b0),
	.w6(32'hba534e8f),
	.w7(32'hbaf73097),
	.w8(32'hb82d91b8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9864ae),
	.w1(32'h3aadf7a4),
	.w2(32'h3a848e37),
	.w3(32'h3b048fd9),
	.w4(32'hba5f4710),
	.w5(32'hbb25be11),
	.w6(32'h3b61d72e),
	.w7(32'hba8f8173),
	.w8(32'hbb878546),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e8363a),
	.w1(32'hbae7bae8),
	.w2(32'h3a2a8a28),
	.w3(32'hb8810e3c),
	.w4(32'hbab493c9),
	.w5(32'hba4f3c9c),
	.w6(32'h3b4b7623),
	.w7(32'h3b5cd4f1),
	.w8(32'hb9ffff5a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25976f),
	.w1(32'hb71de518),
	.w2(32'hb9007c3f),
	.w3(32'h3ab23bb0),
	.w4(32'h39d7bad7),
	.w5(32'h3ae5bad6),
	.w6(32'h3b054ce2),
	.w7(32'h39431ee4),
	.w8(32'h3aaec86f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a9f4b),
	.w1(32'h3b797ecb),
	.w2(32'hba8d8de3),
	.w3(32'h3acd042a),
	.w4(32'h3ab3d74a),
	.w5(32'h3ab30c03),
	.w6(32'h3b0a06b6),
	.w7(32'h3a3fd085),
	.w8(32'h3a9ce754),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac818fd),
	.w1(32'hbab10a45),
	.w2(32'hb9665618),
	.w3(32'hba46e6ef),
	.w4(32'hba6ee56c),
	.w5(32'hba20a333),
	.w6(32'hbaa63a4d),
	.w7(32'hba01f890),
	.w8(32'h36d138f4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59e6b),
	.w1(32'hbb5d6932),
	.w2(32'hbbdd8ea3),
	.w3(32'h3b7d3fe8),
	.w4(32'hba34e84b),
	.w5(32'hbbb89c60),
	.w6(32'h3bbd6b3e),
	.w7(32'h3b98af62),
	.w8(32'hb91b119a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972994e),
	.w1(32'hbb0071db),
	.w2(32'h3aaa1810),
	.w3(32'hbb40410b),
	.w4(32'hbb6df1e9),
	.w5(32'hbab5d170),
	.w6(32'h3a7c87c1),
	.w7(32'hbada027a),
	.w8(32'hbb11b3d0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca42d),
	.w1(32'h3b2c0056),
	.w2(32'h3b062312),
	.w3(32'h3b7db198),
	.w4(32'h3b015be0),
	.w5(32'h3abed58b),
	.w6(32'h3b808f4c),
	.w7(32'h3b496ee9),
	.w8(32'h3b13f8f7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d9846),
	.w1(32'h3978c83f),
	.w2(32'hba893db2),
	.w3(32'h3b64ada3),
	.w4(32'hba25043b),
	.w5(32'hbb3a22e7),
	.w6(32'h3b3754b6),
	.w7(32'h3a1f7f27),
	.w8(32'hbafbfd12),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695a21),
	.w1(32'hbb4a52a5),
	.w2(32'hbb5cb5f0),
	.w3(32'hbaae75f7),
	.w4(32'hba472e83),
	.w5(32'h3ac1d528),
	.w6(32'hbaa8b3df),
	.w7(32'hba7dc43b),
	.w8(32'hb97b2769),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bded0),
	.w1(32'h3a15b5db),
	.w2(32'hb8ec822b),
	.w3(32'h3a62bb08),
	.w4(32'h3a71e4ed),
	.w5(32'hba9af42c),
	.w6(32'h3ad1c10d),
	.w7(32'hba609046),
	.w8(32'h3a6b66c1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa644b6),
	.w1(32'hba89b49b),
	.w2(32'hbb2cf88b),
	.w3(32'h39724d4e),
	.w4(32'hbae18bb5),
	.w5(32'hbb3bc22c),
	.w6(32'hb9c43256),
	.w7(32'hbac4f6bf),
	.w8(32'hbb18320d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c9f73),
	.w1(32'h3aa1ca8c),
	.w2(32'h3b75bb2b),
	.w3(32'h3c39d970),
	.w4(32'h3b5e56d0),
	.w5(32'hbb0ec8df),
	.w6(32'h3ca61fb2),
	.w7(32'h3c511300),
	.w8(32'h3a3e8e59),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab84e36),
	.w1(32'h3a5f0abf),
	.w2(32'h3a1dcfe8),
	.w3(32'h3a4dfe79),
	.w4(32'h38897288),
	.w5(32'hb9db37ea),
	.w6(32'h38f948ea),
	.w7(32'h37e581b7),
	.w8(32'hb93ac8d3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae76c96),
	.w1(32'hbc066189),
	.w2(32'hbc0413cc),
	.w3(32'h378a343e),
	.w4(32'hbbc76e44),
	.w5(32'hbbc901a6),
	.w6(32'h3b1e1f16),
	.w7(32'hba947b2d),
	.w8(32'hbb90402d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfdbdc),
	.w1(32'hba35fd76),
	.w2(32'hb78d01c7),
	.w3(32'h37952ae2),
	.w4(32'hbaac4718),
	.w5(32'hba49af36),
	.w6(32'hb9b449b6),
	.w7(32'h3982afe0),
	.w8(32'h392d54fa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9efc88),
	.w1(32'hbb7374b7),
	.w2(32'hbbddba51),
	.w3(32'h3b91c8a2),
	.w4(32'hba41633b),
	.w5(32'hbb62a712),
	.w6(32'h3beaac59),
	.w7(32'h3b830101),
	.w8(32'h3b424520),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898fba8),
	.w1(32'hb90d0a0d),
	.w2(32'hb90f894b),
	.w3(32'hb8a3c4d4),
	.w4(32'hb9d948ec),
	.w5(32'hba17144c),
	.w6(32'hb9087fa2),
	.w7(32'hb8d63240),
	.w8(32'hb9a96b50),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc99bc0),
	.w1(32'h3b0e7d65),
	.w2(32'h3b1b7daa),
	.w3(32'h3c021294),
	.w4(32'h3b2caa31),
	.w5(32'h3afe9da8),
	.w6(32'h3be6eb60),
	.w7(32'h3ba5c825),
	.w8(32'h3b4a092c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b434d),
	.w1(32'hb9c9db54),
	.w2(32'hb9e45a72),
	.w3(32'hb98cb3c2),
	.w4(32'hba38149f),
	.w5(32'hba59099b),
	.w6(32'hb9d8404e),
	.w7(32'hb993c2b1),
	.w8(32'hb8f258e0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55573d),
	.w1(32'hbad4a3aa),
	.w2(32'hbaa4473e),
	.w3(32'h3ba04164),
	.w4(32'hb85a023a),
	.w5(32'hbb4e6251),
	.w6(32'h3c15d817),
	.w7(32'h3bbc5660),
	.w8(32'hb73c3c4e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3309b4),
	.w1(32'hb69cf07e),
	.w2(32'hbb8ab3d7),
	.w3(32'h3b578dbb),
	.w4(32'hba9f1b26),
	.w5(32'hbb6a8e07),
	.w6(32'h3b8d5de1),
	.w7(32'h395dc8d1),
	.w8(32'hbb5ca9fa),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05b540),
	.w1(32'h3b39c95e),
	.w2(32'h3b3214c9),
	.w3(32'h3b1a353c),
	.w4(32'h3b044c1a),
	.w5(32'h3b16cb04),
	.w6(32'h3b01b555),
	.w7(32'h3b07b20f),
	.w8(32'h3ab5831a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0e8dd),
	.w1(32'hba1cf47a),
	.w2(32'hbab0f52f),
	.w3(32'hbad18944),
	.w4(32'h39e241d3),
	.w5(32'h39d91b09),
	.w6(32'hb92efe19),
	.w7(32'hba4f20e8),
	.w8(32'hb99477de),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde4877),
	.w1(32'hbbea0a71),
	.w2(32'hbb0a2e90),
	.w3(32'hbae24d5a),
	.w4(32'hbb19fbf0),
	.w5(32'h3a9886fd),
	.w6(32'hb9ff6132),
	.w7(32'hbaad6204),
	.w8(32'hba0b25d2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb119f1),
	.w1(32'hbc29d395),
	.w2(32'hbbde9b6a),
	.w3(32'hbb686eb2),
	.w4(32'hbc01faec),
	.w5(32'hbbf0cf7e),
	.w6(32'h3ab1fdca),
	.w7(32'h3a0c95e1),
	.w8(32'hbaa282cd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2a46f),
	.w1(32'hbbe04183),
	.w2(32'hbc265c4c),
	.w3(32'hbb68f844),
	.w4(32'hbba4a3ac),
	.w5(32'hbbb0444f),
	.w6(32'h3a9a042a),
	.w7(32'h39fec018),
	.w8(32'hba5b5a1b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88296),
	.w1(32'hbc0d39f6),
	.w2(32'hbbffd77d),
	.w3(32'h3bf6edbc),
	.w4(32'hbb2f8baa),
	.w5(32'hbc09ec8e),
	.w6(32'h3c99f214),
	.w7(32'h3c31e4ed),
	.w8(32'h3a8d08ae),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dcaf9),
	.w1(32'hbb94be79),
	.w2(32'hbbbe7d2a),
	.w3(32'h3c1017f8),
	.w4(32'hbb7d4b6e),
	.w5(32'hbbf75500),
	.w6(32'h3c048e0e),
	.w7(32'h3b0d94bd),
	.w8(32'hbb54ef25),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15e234),
	.w1(32'hba7b4100),
	.w2(32'hb8abcd07),
	.w3(32'hba86aea2),
	.w4(32'hba50aa04),
	.w5(32'h398fd44a),
	.w6(32'hb9898737),
	.w7(32'hb7c1f8b6),
	.w8(32'hb9bd3c83),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e229ed),
	.w1(32'hb92148e1),
	.w2(32'h38fc5e9e),
	.w3(32'hb78009a2),
	.w4(32'hb98d955e),
	.w5(32'h39823749),
	.w6(32'hb94fefd9),
	.w7(32'h38fdb331),
	.w8(32'hb9cff8f8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e184),
	.w1(32'hbae86389),
	.w2(32'hba996028),
	.w3(32'hbb2379d5),
	.w4(32'hbb23bd4a),
	.w5(32'hbaf68556),
	.w6(32'hba6ce46c),
	.w7(32'hbb14aff3),
	.w8(32'hba5fc1bc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bbada),
	.w1(32'hba9049bb),
	.w2(32'hba92980f),
	.w3(32'h3b4a9b78),
	.w4(32'hb9faf81a),
	.w5(32'h38c237ee),
	.w6(32'h3ba36b87),
	.w7(32'h3ac5bb02),
	.w8(32'h39d24ca8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a2e88),
	.w1(32'hbb291aef),
	.w2(32'hba06388d),
	.w3(32'hbb5fd665),
	.w4(32'hbb26281c),
	.w5(32'hb9183351),
	.w6(32'hb9b28d6c),
	.w7(32'h39725b26),
	.w8(32'hba8dcac3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4500),
	.w1(32'h3a654881),
	.w2(32'h39953e8f),
	.w3(32'h3a769fc2),
	.w4(32'h39eebfab),
	.w5(32'hba4bb844),
	.w6(32'hba4dbdee),
	.w7(32'hb9a3f295),
	.w8(32'hba7f03f4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bcb23),
	.w1(32'hbaba25b4),
	.w2(32'h3b458c93),
	.w3(32'hba8ca783),
	.w4(32'h3a23e8ae),
	.w5(32'h3b951e2d),
	.w6(32'hba531acb),
	.w7(32'hba221f0a),
	.w8(32'hb71d453c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0783e8),
	.w1(32'hbc13a1ce),
	.w2(32'hbbbb9699),
	.w3(32'hbbdb5dbe),
	.w4(32'hbc135c5c),
	.w5(32'hbbcf4064),
	.w6(32'hbb755860),
	.w7(32'hbb55f8f5),
	.w8(32'hbb968a6b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50b821),
	.w1(32'hbc235ee0),
	.w2(32'hbc1956c5),
	.w3(32'hbc44f4a7),
	.w4(32'hbc1b3888),
	.w5(32'hbbc68402),
	.w6(32'hbbde3b55),
	.w7(32'hbc0fc046),
	.w8(32'hbbb557a0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bd139),
	.w1(32'h3a9c94dd),
	.w2(32'h3a7a40b9),
	.w3(32'h3b6dbd94),
	.w4(32'h39923476),
	.w5(32'hbb1c4a2c),
	.w6(32'h3ae36355),
	.w7(32'h3b08f156),
	.w8(32'hba5c7c65),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71dd12),
	.w1(32'hbc18dd6f),
	.w2(32'hbb3cfa68),
	.w3(32'hb9a9ffd8),
	.w4(32'hbbcd8fc2),
	.w5(32'hbafd7960),
	.w6(32'h3c1efd0d),
	.w7(32'h3ba84b23),
	.w8(32'h3b76dd5f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192fc4),
	.w1(32'h39ccbcf1),
	.w2(32'hba982263),
	.w3(32'hbad389b4),
	.w4(32'hb9ce874d),
	.w5(32'h3a00ee0e),
	.w6(32'hba98ce08),
	.w7(32'hbb134dec),
	.w8(32'h39b7f6e4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396845de),
	.w1(32'h3a236ae2),
	.w2(32'h3a719dc3),
	.w3(32'h3a252a09),
	.w4(32'h3a21a9be),
	.w5(32'h3a126a4a),
	.w6(32'h3a7e236e),
	.w7(32'h3aa598f4),
	.w8(32'h38c4314d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9307b),
	.w1(32'h383973f5),
	.w2(32'h393abf4a),
	.w3(32'h3979fcb3),
	.w4(32'hb9a214dc),
	.w5(32'h36f92f11),
	.w6(32'hb8fa311c),
	.w7(32'h396903a6),
	.w8(32'hb9ee7c95),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6303),
	.w1(32'hba388de8),
	.w2(32'hbb153329),
	.w3(32'hbad2d7b3),
	.w4(32'hbab76040),
	.w5(32'hbada2d4b),
	.w6(32'hbab0332b),
	.w7(32'hbae696fc),
	.w8(32'hbaa043d6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012a21),
	.w1(32'hbbc51b39),
	.w2(32'hbbca654b),
	.w3(32'hbbbf7971),
	.w4(32'hbbb48e25),
	.w5(32'hbba0ce08),
	.w6(32'hbb89087c),
	.w7(32'hba98dbf9),
	.w8(32'hbaf3acbc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcce623),
	.w1(32'h3c01d84a),
	.w2(32'h3b4656e1),
	.w3(32'h3babd477),
	.w4(32'h3bb0e2fe),
	.w5(32'h3acf0e15),
	.w6(32'h3bbe1350),
	.w7(32'h3bdf6cae),
	.w8(32'h391c7e86),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acbb0),
	.w1(32'hbb48bf5f),
	.w2(32'hbaccc66d),
	.w3(32'hbacaa269),
	.w4(32'h3a17939c),
	.w5(32'h3b42d707),
	.w6(32'hba98695b),
	.w7(32'hba8ae605),
	.w8(32'hb9b8cb2b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5d696),
	.w1(32'hbae17375),
	.w2(32'hbad80a96),
	.w3(32'hbaf58f0a),
	.w4(32'hbaa17978),
	.w5(32'hba4195cf),
	.w6(32'hbb22803a),
	.w7(32'hbb0b059e),
	.w8(32'hba537eff),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29e53b),
	.w1(32'h39a9e681),
	.w2(32'h3ac37505),
	.w3(32'h3c0566e7),
	.w4(32'hba1ffbeb),
	.w5(32'hbae99b4f),
	.w6(32'h3c74b06e),
	.w7(32'h3be1910b),
	.w8(32'h3a931543),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00b25b),
	.w1(32'hbbbead96),
	.w2(32'hb8a96abe),
	.w3(32'h390f17b0),
	.w4(32'hbb73efa3),
	.w5(32'hbb120b16),
	.w6(32'h39a66587),
	.w7(32'h3b4ad8bc),
	.w8(32'h3b6a783d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbedb89),
	.w1(32'hbbb58e18),
	.w2(32'hbb840a56),
	.w3(32'hbbce3bf8),
	.w4(32'hbba5fa54),
	.w5(32'hbb244c04),
	.w6(32'hbb8e6771),
	.w7(32'hbb8b88c2),
	.w8(32'hbb797652),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8572dd),
	.w1(32'hbabb80e2),
	.w2(32'hbaa158ad),
	.w3(32'hbb511334),
	.w4(32'hba9499a9),
	.w5(32'h38ee4fdd),
	.w6(32'hbb5e0e6b),
	.w7(32'hbb3eee55),
	.w8(32'hbb3d0ad7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe55195),
	.w1(32'hbbc42b53),
	.w2(32'hbb0b0631),
	.w3(32'hbb661452),
	.w4(32'hba927b83),
	.w5(32'hba9dd4bc),
	.w6(32'h3af1c576),
	.w7(32'h3abf21f6),
	.w8(32'h3ad84baf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b01cf),
	.w1(32'hbbcd248c),
	.w2(32'hbaef451b),
	.w3(32'h3a8abe35),
	.w4(32'hbb470e69),
	.w5(32'hbaad3958),
	.w6(32'h3b4ed1d9),
	.w7(32'h3b1b2af0),
	.w8(32'hba3090bd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff2cb2),
	.w1(32'hba94a45e),
	.w2(32'hbb0d5926),
	.w3(32'hbb95f82d),
	.w4(32'hba70f1f6),
	.w5(32'hbb38c3b9),
	.w6(32'hb93f8124),
	.w7(32'hba7e4dd9),
	.w8(32'h37aa95e6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89574a),
	.w1(32'h3b338043),
	.w2(32'h3b85fac1),
	.w3(32'hba27e1a7),
	.w4(32'hba8f7ff8),
	.w5(32'h3b3acfff),
	.w6(32'hbb80f14e),
	.w7(32'hbb8e4675),
	.w8(32'hbafa21a4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83768c),
	.w1(32'h3a43cf03),
	.w2(32'h37f3cadb),
	.w3(32'hba95f3f3),
	.w4(32'h39ba8a4b),
	.w5(32'hb8afe365),
	.w6(32'h39d13269),
	.w7(32'hba1d53af),
	.w8(32'h3908e80e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd7077),
	.w1(32'hba2f3377),
	.w2(32'hba1183fc),
	.w3(32'hb9d53dde),
	.w4(32'hb7deb15a),
	.w5(32'hb91a0773),
	.w6(32'h3a6648d1),
	.w7(32'h39c507d7),
	.w8(32'h3a80cbfd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274241),
	.w1(32'h3b7b5654),
	.w2(32'h3b62b99a),
	.w3(32'h3b9715a3),
	.w4(32'h3bb0a564),
	.w5(32'h3b9e466f),
	.w6(32'h3bde1882),
	.w7(32'h3bc03b95),
	.w8(32'h3b791e45),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cb1be),
	.w1(32'h3ba27ac8),
	.w2(32'hba5095b8),
	.w3(32'h3b1f87c3),
	.w4(32'h3bcfd120),
	.w5(32'h3a863774),
	.w6(32'hb9d2d6ca),
	.w7(32'hba17110c),
	.w8(32'h3b592977),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38bea6),
	.w1(32'h3b0b3adb),
	.w2(32'h3b7076f5),
	.w3(32'h3b0c4c7b),
	.w4(32'h3b0d3604),
	.w5(32'h3b42b5be),
	.w6(32'h3b73dda8),
	.w7(32'h3b34e91a),
	.w8(32'hbaa6b719),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3877cb45),
	.w1(32'h3a411d4b),
	.w2(32'hba442ea9),
	.w3(32'h3adf2cfd),
	.w4(32'hbad49d3b),
	.w5(32'hbb112317),
	.w6(32'h3a882356),
	.w7(32'h3ac1dbd6),
	.w8(32'hba78205e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbbe8),
	.w1(32'h3b6d384f),
	.w2(32'h3b50fae1),
	.w3(32'hbb0ffec6),
	.w4(32'h3a118c94),
	.w5(32'h3a8216b7),
	.w6(32'h3ad740f3),
	.w7(32'hb97d606c),
	.w8(32'h3a152604),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0ca0),
	.w1(32'hbb7ca06f),
	.w2(32'h3a9cd7aa),
	.w3(32'h3b2cacd3),
	.w4(32'h3aca10d4),
	.w5(32'h3a7db1cd),
	.w6(32'hbace50f8),
	.w7(32'hb9a95020),
	.w8(32'hbb26f261),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d811),
	.w1(32'h3b1470b4),
	.w2(32'hbaa1b138),
	.w3(32'h3b4f99d7),
	.w4(32'h3b1e977b),
	.w5(32'hba68e808),
	.w6(32'h3b5c4fe5),
	.w7(32'h3b8160a3),
	.w8(32'h3b259a31),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e9053),
	.w1(32'h37b6c0dd),
	.w2(32'h3a0117ac),
	.w3(32'hb954fdcd),
	.w4(32'hb9580463),
	.w5(32'hba635428),
	.w6(32'hbb1b3c56),
	.w7(32'hbab1f184),
	.w8(32'hbbad482f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aff59),
	.w1(32'h3acc1e8c),
	.w2(32'hbaef117e),
	.w3(32'hba928715),
	.w4(32'hbab916e1),
	.w5(32'hbad8c2a4),
	.w6(32'hbbda0a45),
	.w7(32'hbbea4674),
	.w8(32'hba9f2da5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9962f8),
	.w1(32'hbb6d3049),
	.w2(32'h3b69031e),
	.w3(32'hbb2e4078),
	.w4(32'h3994b913),
	.w5(32'hba7ae58b),
	.w6(32'hbbc1ff50),
	.w7(32'hb840de63),
	.w8(32'hba3df69f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0928),
	.w1(32'h37a4b7a4),
	.w2(32'h3a6aeb7b),
	.w3(32'hbb6fa42e),
	.w4(32'hbab0b2d1),
	.w5(32'hbb15fc20),
	.w6(32'h3abe3a5e),
	.w7(32'hba8ea480),
	.w8(32'h3a2f123b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeae31),
	.w1(32'h3a805f22),
	.w2(32'h3b13f5b4),
	.w3(32'h3b436491),
	.w4(32'h3b73a7e9),
	.w5(32'h3b92cf17),
	.w6(32'h3b1759ee),
	.w7(32'h3b4ca8b6),
	.w8(32'h3babcb5e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a5b68),
	.w1(32'h3c006869),
	.w2(32'h3bc9796a),
	.w3(32'h3b64f221),
	.w4(32'h3c0a1696),
	.w5(32'h3c128d01),
	.w6(32'h3b78e193),
	.w7(32'h3afc9dab),
	.w8(32'h3b738551),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule