module layer_10_featuremap_24(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcdd38),
	.w1(32'h3b9c0b59),
	.w2(32'hbc5295f4),
	.w3(32'h3ba0c5d7),
	.w4(32'h3b5b613a),
	.w5(32'hbb4588d8),
	.w6(32'hbc56e282),
	.w7(32'hbbcecb5e),
	.w8(32'hba3708fa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c228504),
	.w1(32'h3c6aac9b),
	.w2(32'hbc1df155),
	.w3(32'h3c76615a),
	.w4(32'h3c67b164),
	.w5(32'hbbe44382),
	.w6(32'h3b44b2e3),
	.w7(32'h3c157fb0),
	.w8(32'hbb5c848c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc698bd1),
	.w1(32'hbb93951e),
	.w2(32'h3c0fb0eb),
	.w3(32'hbc448ce9),
	.w4(32'hbc1bcd5f),
	.w5(32'h3c9dda0f),
	.w6(32'hbc43dc3c),
	.w7(32'hbbce5fc9),
	.w8(32'h3c658984),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d0ef5),
	.w1(32'h3b033bc3),
	.w2(32'h3c8f2ce2),
	.w3(32'h3d1e9301),
	.w4(32'h3cafaacb),
	.w5(32'h3ca67f8a),
	.w6(32'h3cc6f65b),
	.w7(32'h3c9d5ca1),
	.w8(32'h3bc2dea8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c520f93),
	.w1(32'h3a8fae0a),
	.w2(32'hbc2c280a),
	.w3(32'h3c91ae80),
	.w4(32'h3c60291b),
	.w5(32'hbd3fd4b9),
	.w6(32'h3c56a4ed),
	.w7(32'h3c93aa83),
	.w8(32'hbd14207c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd79dcc),
	.w1(32'hbc80b1d9),
	.w2(32'h3b363050),
	.w3(32'hbd5413a4),
	.w4(32'hbc55b373),
	.w5(32'h39a8e5cf),
	.w6(32'hbcffe2f0),
	.w7(32'hbc4f81bc),
	.w8(32'hb99b7bf3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dd16c),
	.w1(32'h3a880b1d),
	.w2(32'h3b4592ad),
	.w3(32'h3b66284c),
	.w4(32'hbabc1bf5),
	.w5(32'h3abc0ff0),
	.w6(32'h3b38157a),
	.w7(32'hbac1e3fb),
	.w8(32'h3bb3e72c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6ada7),
	.w1(32'h3ad330ad),
	.w2(32'h3bbfbc7b),
	.w3(32'h3c2a209c),
	.w4(32'h3b019ff7),
	.w5(32'hbbd26bac),
	.w6(32'h3bf9e314),
	.w7(32'h3c0e30cf),
	.w8(32'hbb7de3f3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9507c7),
	.w1(32'h3b8b3797),
	.w2(32'h3a30e5ce),
	.w3(32'h3b404c7e),
	.w4(32'hbb23fb09),
	.w5(32'hbb92f62a),
	.w6(32'hbab4cdc5),
	.w7(32'hbb771d4e),
	.w8(32'hbb5baaf7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977984),
	.w1(32'h3b5dcdc0),
	.w2(32'hbb8d6189),
	.w3(32'h3ba89134),
	.w4(32'h3bb1747f),
	.w5(32'hbba8dc70),
	.w6(32'h3ad6e4f4),
	.w7(32'h3c011ae9),
	.w8(32'hbb65cb9b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf87f8),
	.w1(32'hbb823cfd),
	.w2(32'hbadae165),
	.w3(32'hbbc7d07e),
	.w4(32'hbb16e397),
	.w5(32'h3c00ce75),
	.w6(32'hbb833801),
	.w7(32'hbb7d25c3),
	.w8(32'h3b4acae7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380307),
	.w1(32'h3b95418d),
	.w2(32'h3b532609),
	.w3(32'h3cbf1ea3),
	.w4(32'h3c5e45db),
	.w5(32'hbb39a385),
	.w6(32'h3cc0e192),
	.w7(32'h3c3371ab),
	.w8(32'hba72ec57),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8abeb),
	.w1(32'h3bc2941c),
	.w2(32'h3b869c69),
	.w3(32'h3bb6cc9f),
	.w4(32'h3bc67957),
	.w5(32'h3b4a8e9e),
	.w6(32'h3ba968cd),
	.w7(32'h3b98f585),
	.w8(32'h3b821145),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4a53c),
	.w1(32'hbb050bb7),
	.w2(32'h3c134744),
	.w3(32'h3c1f0587),
	.w4(32'h3af6e35c),
	.w5(32'hbb8a82d5),
	.w6(32'h3c13002d),
	.w7(32'h3a80f1ef),
	.w8(32'hbc090801),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fcd53),
	.w1(32'hbb76b9ea),
	.w2(32'hbad12ed9),
	.w3(32'hbc83784d),
	.w4(32'hbc554812),
	.w5(32'hbb88efc1),
	.w6(32'hbc3a6d18),
	.w7(32'hbc12676f),
	.w8(32'hbbcbc50c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a971218),
	.w1(32'h3a050dbe),
	.w2(32'hbb137088),
	.w3(32'h39b87900),
	.w4(32'hbb25e078),
	.w5(32'hbb973b58),
	.w6(32'hbb2ec026),
	.w7(32'h3a8ced96),
	.w8(32'hbb6f05ba),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91af20),
	.w1(32'hb9a6dd14),
	.w2(32'h3b85b588),
	.w3(32'hbb67e5e2),
	.w4(32'hbb036e52),
	.w5(32'h3adff73c),
	.w6(32'hbb474999),
	.w7(32'hbb1c3fa9),
	.w8(32'h3c3ccb39),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a942d),
	.w1(32'h3bdb39fc),
	.w2(32'hba86c32b),
	.w3(32'h3903a39b),
	.w4(32'h3bac47dd),
	.w5(32'h3b8aa4ba),
	.w6(32'h3c296c26),
	.w7(32'h3c421ea9),
	.w8(32'hb9f8e61c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d14e8f),
	.w1(32'hbb3f8eb9),
	.w2(32'h3b859605),
	.w3(32'h3c03bea1),
	.w4(32'h3b3b300d),
	.w5(32'h3bf2def8),
	.w6(32'h3bbb3930),
	.w7(32'h3b9d8685),
	.w8(32'h3bfd34db),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f761),
	.w1(32'h3bc2b2ca),
	.w2(32'hbb241748),
	.w3(32'h3c836879),
	.w4(32'h3b21182c),
	.w5(32'h3b3532c2),
	.w6(32'h3ba10f16),
	.w7(32'hbb740eea),
	.w8(32'hbaefa66d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9184d4),
	.w1(32'hbb887324),
	.w2(32'h3c8488d4),
	.w3(32'h3ac20457),
	.w4(32'hba9129b7),
	.w5(32'h3c914885),
	.w6(32'hba63ba2f),
	.w7(32'hbb68fcc1),
	.w8(32'h3c8a6079),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caba610),
	.w1(32'h3c9c97e3),
	.w2(32'h3c0f15ad),
	.w3(32'h3d0204c5),
	.w4(32'h3c92a0b4),
	.w5(32'h3b9152d5),
	.w6(32'h3c6f577c),
	.w7(32'h3c7fda53),
	.w8(32'hbc04c690),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21dd04),
	.w1(32'h3c22e468),
	.w2(32'h38e5c670),
	.w3(32'h3c94f3b7),
	.w4(32'h3c7781b1),
	.w5(32'hbaaefed6),
	.w6(32'h3ba1bd88),
	.w7(32'h3bb69701),
	.w8(32'hb99cc154),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee189),
	.w1(32'h3b9d6ada),
	.w2(32'h3b6154bc),
	.w3(32'h3b76272a),
	.w4(32'h3c03f3f7),
	.w5(32'h3c0d657c),
	.w6(32'h3b8aefd1),
	.w7(32'h3bbfd717),
	.w8(32'h3b74544c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c848),
	.w1(32'h3b9469e4),
	.w2(32'h3b9b04c3),
	.w3(32'h3c5b711d),
	.w4(32'h3bac67d0),
	.w5(32'h39a7f8b7),
	.w6(32'h3c580a20),
	.w7(32'h3b809d4f),
	.w8(32'h3bcbc36b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45d01a),
	.w1(32'h3b361f9e),
	.w2(32'h3be1e5bc),
	.w3(32'h3b44fb3a),
	.w4(32'hb9d6eb71),
	.w5(32'h3cfbc052),
	.w6(32'h3ba6b536),
	.w7(32'hb9816657),
	.w8(32'h3cb6e02d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dbf1b),
	.w1(32'h3c492a60),
	.w2(32'hba66be3c),
	.w3(32'h3d19592a),
	.w4(32'h3cd5f448),
	.w5(32'hbb765bea),
	.w6(32'h3cf6820a),
	.w7(32'h3caad0f9),
	.w8(32'h3a2347e7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa3adb),
	.w1(32'hbade376f),
	.w2(32'h3c2148a1),
	.w3(32'hbb1ac16a),
	.w4(32'hbb98ae9b),
	.w5(32'hbbcb6d46),
	.w6(32'h3aa2f0f1),
	.w7(32'hb9924112),
	.w8(32'hb9ee696d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9507bd),
	.w1(32'h3c6328ff),
	.w2(32'hbc04b6f3),
	.w3(32'hbaa82266),
	.w4(32'h39995f5b),
	.w5(32'hbb85ffc9),
	.w6(32'h3aaa073c),
	.w7(32'h3b6fcb37),
	.w8(32'hbc89ae07),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481b8c),
	.w1(32'hbb9e6ce3),
	.w2(32'hba9a40b5),
	.w3(32'hbbed43c3),
	.w4(32'hbbabee7f),
	.w5(32'hbbed1a6f),
	.w6(32'hbc3c853e),
	.w7(32'hbc64e2cc),
	.w8(32'h39dfa44e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b502dbd),
	.w1(32'h3aec0f75),
	.w2(32'hbc48cb15),
	.w3(32'hbb821a4e),
	.w4(32'hbb80a06f),
	.w5(32'h3be52b31),
	.w6(32'h3b6d2bb0),
	.w7(32'h3b59e8c9),
	.w8(32'hbb585a76),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bfb3a),
	.w1(32'hbc06bcc6),
	.w2(32'hbca572f6),
	.w3(32'h3c5236c6),
	.w4(32'h3c064486),
	.w5(32'h3ccc2f5e),
	.w6(32'h3b1958e4),
	.w7(32'h3bccfac9),
	.w8(32'hba117537),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e1ef0),
	.w1(32'hbbdd4348),
	.w2(32'hbb655e63),
	.w3(32'h3cbac436),
	.w4(32'h3c5c9181),
	.w5(32'hba108655),
	.w6(32'h3b37156d),
	.w7(32'h3c357034),
	.w8(32'hbb2f9ada),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9894),
	.w1(32'hbb8f8829),
	.w2(32'hbbd52027),
	.w3(32'h3ab819e8),
	.w4(32'hba99b8d8),
	.w5(32'h3b41c9c4),
	.w6(32'hbb4cb208),
	.w7(32'hbb2a5f73),
	.w8(32'h3c10d33c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98e6a5),
	.w1(32'hbb8c11e4),
	.w2(32'h3af3a758),
	.w3(32'hbc69075d),
	.w4(32'h3b578e49),
	.w5(32'h3b1d622d),
	.w6(32'hb93c6d8c),
	.w7(32'h3b32bb78),
	.w8(32'hbb7ef401),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957fbe9),
	.w1(32'hbaf25c92),
	.w2(32'hbc7e7079),
	.w3(32'h3b325ba5),
	.w4(32'h3a826f36),
	.w5(32'h3b56708f),
	.w6(32'hbb9d1a4d),
	.w7(32'hbbc92bc2),
	.w8(32'hbc120c42),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc912bd0),
	.w1(32'hbca524b8),
	.w2(32'h3a40ef8f),
	.w3(32'h3c5caafd),
	.w4(32'h3c5065fa),
	.w5(32'hbc1300f5),
	.w6(32'hbc324fdf),
	.w7(32'hbc738df1),
	.w8(32'hba8c8191),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d806d),
	.w1(32'h3c119541),
	.w2(32'h3c8e7315),
	.w3(32'hba41fa66),
	.w4(32'hbb8be9e7),
	.w5(32'hbcdb3dd9),
	.w6(32'h3b7bc8f1),
	.w7(32'h3a25ba7f),
	.w8(32'h3c54a816),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfcf889),
	.w1(32'h3cd95829),
	.w2(32'hbb37dab3),
	.w3(32'hbd00d700),
	.w4(32'hbca3e1d0),
	.w5(32'h3bfcef39),
	.w6(32'h3c5e6fd8),
	.w7(32'h3b6e7d75),
	.w8(32'hbbaf1455),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f6329),
	.w1(32'h3b9a25b2),
	.w2(32'h3c1dc6e4),
	.w3(32'h3bac81a0),
	.w4(32'h3b051312),
	.w5(32'h3b4e4d33),
	.w6(32'h3c28dbed),
	.w7(32'h3c6affff),
	.w8(32'h3b56b0bf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1681de),
	.w1(32'h3b1f5d63),
	.w2(32'hbbda300c),
	.w3(32'hba7a29f2),
	.w4(32'hbab1d2a0),
	.w5(32'hbbec6e96),
	.w6(32'h3bb2f493),
	.w7(32'h3a8db4e9),
	.w8(32'h3b461385),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9c59),
	.w1(32'h3b126178),
	.w2(32'h3bc855c8),
	.w3(32'hbc18cb90),
	.w4(32'hbaa61302),
	.w5(32'hbbd7230a),
	.w6(32'h3c81dfbf),
	.w7(32'h3c8c42f3),
	.w8(32'h3b18f838),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217c78),
	.w1(32'hbb952502),
	.w2(32'h3ad52c46),
	.w3(32'hbb43827f),
	.w4(32'h3b9b48b9),
	.w5(32'hba9b17c8),
	.w6(32'hbbed666d),
	.w7(32'hbb7cfb62),
	.w8(32'hbb8c1167),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa474ab),
	.w1(32'h3b81d0dc),
	.w2(32'hbb9e186a),
	.w3(32'h3a79e834),
	.w4(32'h3abe9a2e),
	.w5(32'hbc2d271a),
	.w6(32'hbb9c09f1),
	.w7(32'hbba69545),
	.w8(32'hbc347d2c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901e72),
	.w1(32'hbbc2af57),
	.w2(32'hbb7a21c9),
	.w3(32'hbbb4ecf7),
	.w4(32'hbc183048),
	.w5(32'h3b47704f),
	.w6(32'hbad1a6d3),
	.w7(32'hbbf665d0),
	.w8(32'h3b848bca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5906),
	.w1(32'h3b563322),
	.w2(32'h3bace8c5),
	.w3(32'hbc35fb80),
	.w4(32'hbae43751),
	.w5(32'hbb48ddc1),
	.w6(32'hba275b43),
	.w7(32'h3b109ce1),
	.w8(32'h3bc50a38),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4643cd),
	.w1(32'h3b817979),
	.w2(32'h3baa5961),
	.w3(32'h3adf2810),
	.w4(32'hbb8b9d37),
	.w5(32'h3899f2b1),
	.w6(32'h3c0cc50f),
	.w7(32'h3bd217d4),
	.w8(32'h3c07bcf1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9179c),
	.w1(32'h3ac8813f),
	.w2(32'h3ba39554),
	.w3(32'hbb2b1dd2),
	.w4(32'h3a47e170),
	.w5(32'h3b11fb71),
	.w6(32'h3b13aa20),
	.w7(32'h3be1c34d),
	.w8(32'h3ae72528),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850391),
	.w1(32'h3b553b5c),
	.w2(32'hbb8d7c86),
	.w3(32'h3a38b01e),
	.w4(32'hba85b0de),
	.w5(32'h3bed5371),
	.w6(32'h3a120f69),
	.w7(32'hbb3b6b58),
	.w8(32'hbc021dc0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23fea9),
	.w1(32'hbbfd64e4),
	.w2(32'hba0bfdc6),
	.w3(32'h3c0736ad),
	.w4(32'h3c003f3d),
	.w5(32'hbad0a228),
	.w6(32'hbc55299b),
	.w7(32'hbbdc0cae),
	.w8(32'h3bcbd14f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b89b11),
	.w1(32'h3c314c31),
	.w2(32'h3a4343f4),
	.w3(32'hbbe560ea),
	.w4(32'hbbb0e871),
	.w5(32'hbbc99947),
	.w6(32'h3bbb3264),
	.w7(32'h3c15e2dd),
	.w8(32'hbbf2fb89),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03f331),
	.w1(32'h3b77f0c1),
	.w2(32'h3b22c251),
	.w3(32'hbc2a393e),
	.w4(32'hbb572f00),
	.w5(32'h3bf1d4e5),
	.w6(32'hbad0c87c),
	.w7(32'h3bd00f47),
	.w8(32'h3c0c4efa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c475ddd),
	.w1(32'h3c8b890c),
	.w2(32'hbba6ff7c),
	.w3(32'hbc0a8ec1),
	.w4(32'h3aa2ca65),
	.w5(32'h3aa0821c),
	.w6(32'h3c4734d1),
	.w7(32'h3bbf3655),
	.w8(32'h3ba29df2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41e1f5),
	.w1(32'hbc193d9e),
	.w2(32'h3c174b2f),
	.w3(32'hbbb6be74),
	.w4(32'hbac133fd),
	.w5(32'hbcab4fc1),
	.w6(32'h3a4b682f),
	.w7(32'h3b16490a),
	.w8(32'hbbb44f43),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23d48a),
	.w1(32'h3c163087),
	.w2(32'hbbf01569),
	.w3(32'hbcf4430f),
	.w4(32'hbc823cd9),
	.w5(32'h3d3aa27d),
	.w6(32'hbc046675),
	.w7(32'hbb178515),
	.w8(32'h3b908178),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df16a),
	.w1(32'hbbefc367),
	.w2(32'hbbac26f4),
	.w3(32'h3d3bb05b),
	.w4(32'h3cd53a52),
	.w5(32'h3abe6f80),
	.w6(32'h3c247be3),
	.w7(32'h3c43f269),
	.w8(32'h3a4c83c8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd6c5),
	.w1(32'hbb04c036),
	.w2(32'h3c248205),
	.w3(32'hb922debc),
	.w4(32'h38b9a781),
	.w5(32'hba9192b5),
	.w6(32'hbb83c83c),
	.w7(32'h3bace63b),
	.w8(32'h38bc6740),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7088ac),
	.w1(32'h3c24eb6b),
	.w2(32'hba9eff0d),
	.w3(32'h3964ebbe),
	.w4(32'h3b9c0ab3),
	.w5(32'hbad1e214),
	.w6(32'h3bb443f7),
	.w7(32'h3b9cbb5a),
	.w8(32'h3c4261a8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944e8ef),
	.w1(32'hbb874a8b),
	.w2(32'h3b1e8730),
	.w3(32'hbaf20e4d),
	.w4(32'hbbbd3a90),
	.w5(32'hb89e9069),
	.w6(32'h3c61d7b4),
	.w7(32'h3c324b95),
	.w8(32'hbc01efa7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18fd0f),
	.w1(32'h3b448574),
	.w2(32'h3c15ab0c),
	.w3(32'hbb04bb20),
	.w4(32'h3b4daf16),
	.w5(32'hbca11fe9),
	.w6(32'hbaaeb2c3),
	.w7(32'hb9d0456d),
	.w8(32'h3b931970),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c957436),
	.w1(32'h3c31fbcc),
	.w2(32'hbb3f3078),
	.w3(32'hbca97800),
	.w4(32'hbc706ef1),
	.w5(32'hbc0d2b4d),
	.w6(32'h3c505647),
	.w7(32'h3c15f090),
	.w8(32'hbb04ba35),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8e64c),
	.w1(32'hbb63d3be),
	.w2(32'h3b8a2797),
	.w3(32'hbb863dde),
	.w4(32'h3b26e22f),
	.w5(32'hbc53a6e0),
	.w6(32'h3a442f7b),
	.w7(32'h3bcc5870),
	.w8(32'hbb716aae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac930cb),
	.w1(32'hbbc6b3b0),
	.w2(32'hbafb3054),
	.w3(32'h39dd5713),
	.w4(32'h3b5fc683),
	.w5(32'hbb409278),
	.w6(32'hbc6a3de2),
	.w7(32'h3b4d9798),
	.w8(32'h39f4f774),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba7a1),
	.w1(32'hbc04979b),
	.w2(32'hbb82e14f),
	.w3(32'hbb12e527),
	.w4(32'hbb87a64e),
	.w5(32'h3bb977b7),
	.w6(32'hba4b1489),
	.w7(32'hbb75b241),
	.w8(32'hbbcde2ab),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1b708),
	.w1(32'hbc526b8d),
	.w2(32'hbb3cfb33),
	.w3(32'h3c72ea48),
	.w4(32'h3c4ea0e4),
	.w5(32'hbb1c5823),
	.w6(32'hbc358469),
	.w7(32'hbb220492),
	.w8(32'h3985e1c3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142c19),
	.w1(32'h3a8e25d4),
	.w2(32'h3b963efa),
	.w3(32'hbbc49389),
	.w4(32'hbb96a72d),
	.w5(32'h3ad304c6),
	.w6(32'hbaf86fb9),
	.w7(32'hbb397973),
	.w8(32'h3b3b0f73),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004dc9),
	.w1(32'h3c3d8ce7),
	.w2(32'h3a8ed14c),
	.w3(32'h3bea0f73),
	.w4(32'h3c0504c2),
	.w5(32'hba8acb0d),
	.w6(32'h3bd61c04),
	.w7(32'h3c12f924),
	.w8(32'h3bce1ed3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93f1e7),
	.w1(32'h3b053c23),
	.w2(32'hb9aa128a),
	.w3(32'hbb947065),
	.w4(32'hbc25b67e),
	.w5(32'hbac98719),
	.w6(32'h3beaca5a),
	.w7(32'h3b1acf31),
	.w8(32'hbb972f94),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bc672),
	.w1(32'h3a69f7a9),
	.w2(32'h3b1d37be),
	.w3(32'hbc0868cb),
	.w4(32'hbae5e4a2),
	.w5(32'hba0e989a),
	.w6(32'hbc14fc00),
	.w7(32'hbbee21d5),
	.w8(32'h3b75582f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b662b02),
	.w1(32'h3b635ca6),
	.w2(32'h3bad2bae),
	.w3(32'hb9cfdd84),
	.w4(32'h39fe66e8),
	.w5(32'h3b1f0e62),
	.w6(32'h3b6fce7d),
	.w7(32'h3b8f3905),
	.w8(32'hbb071374),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49cd10),
	.w1(32'h3c45454c),
	.w2(32'hba5e948a),
	.w3(32'h3b999834),
	.w4(32'h3b47dfa8),
	.w5(32'h3a3a8bf6),
	.w6(32'h3bb1e298),
	.w7(32'h3c20dc7d),
	.w8(32'h3c30307c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d263),
	.w1(32'h3c07111a),
	.w2(32'h3b3a4064),
	.w3(32'hbb91734e),
	.w4(32'hbb316ac0),
	.w5(32'hba762f51),
	.w6(32'h3bf64b73),
	.w7(32'h3b0cfe06),
	.w8(32'hbc11f227),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc35c4),
	.w1(32'hbaf1614e),
	.w2(32'h38359d27),
	.w3(32'hbba724b1),
	.w4(32'hbc1f3e3a),
	.w5(32'h3b495a96),
	.w6(32'h3b5fa057),
	.w7(32'h3968d029),
	.w8(32'hbb97e701),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9475033),
	.w1(32'h3b0ae2ca),
	.w2(32'h3903a9fd),
	.w3(32'h3be52ebd),
	.w4(32'h3bd115bf),
	.w5(32'hbb224af5),
	.w6(32'hbbfb3dc0),
	.w7(32'hbb961424),
	.w8(32'h3b04bad2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f45418),
	.w1(32'hbb52f9e0),
	.w2(32'h3b8e7c0f),
	.w3(32'hbb1fe2a6),
	.w4(32'hbbb841cd),
	.w5(32'hbb0136c7),
	.w6(32'h3a81ccaf),
	.w7(32'hbadcf478),
	.w8(32'hbba5bac6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cef8bd),
	.w1(32'hbb8c0cdb),
	.w2(32'h3aa4da1c),
	.w3(32'hbb39a38b),
	.w4(32'hbc199cbb),
	.w5(32'h3ad6d0d5),
	.w6(32'hbc51444e),
	.w7(32'hbc3d8a8a),
	.w8(32'h3b01f4b2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba055322),
	.w1(32'h3bc0a400),
	.w2(32'hbbea7ed7),
	.w3(32'h3b57bb2c),
	.w4(32'h3b196ea4),
	.w5(32'h3c20de5d),
	.w6(32'hbc04baca),
	.w7(32'h3adea7ea),
	.w8(32'hbc642cf2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a4bd4),
	.w1(32'hbbf105d5),
	.w2(32'h3c01454f),
	.w3(32'h3a86490d),
	.w4(32'hbb52e25e),
	.w5(32'hbac5e7da),
	.w6(32'hbc6f0290),
	.w7(32'hbba60e1b),
	.w8(32'h3c7d876c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a9e3),
	.w1(32'h3b9aedc9),
	.w2(32'hba8d9463),
	.w3(32'hbbd71022),
	.w4(32'h3a16fbb8),
	.w5(32'hbc266052),
	.w6(32'h3bf25b55),
	.w7(32'h3b47166a),
	.w8(32'h3a0b3e9f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d0b6),
	.w1(32'hbae56d1e),
	.w2(32'hbb1e862b),
	.w3(32'hbc27800a),
	.w4(32'hbc210c21),
	.w5(32'hbbb13760),
	.w6(32'h39971521),
	.w7(32'h39b05c80),
	.w8(32'h3a53eb71),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dea53),
	.w1(32'hbaa15e2d),
	.w2(32'hbb237cfa),
	.w3(32'hbbb99d6f),
	.w4(32'hbbf14360),
	.w5(32'hbbf10ba9),
	.w6(32'h3b6defe9),
	.w7(32'h3a5f8708),
	.w8(32'hb9938d12),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1d503),
	.w1(32'hbb3db4f9),
	.w2(32'h3aa44ce4),
	.w3(32'hbb62bdb6),
	.w4(32'hbbeb53d8),
	.w5(32'hbbc24743),
	.w6(32'h3b00e024),
	.w7(32'h3a301271),
	.w8(32'hbaeb1dd6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066413),
	.w1(32'hbbd918d6),
	.w2(32'h3c7049a8),
	.w3(32'hbc553997),
	.w4(32'hbc36cf0b),
	.w5(32'hba81e739),
	.w6(32'hbb6e81e2),
	.w7(32'h3b35d8f2),
	.w8(32'h3c48414f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bb4d4),
	.w1(32'h3ba5c5ef),
	.w2(32'h3c4df852),
	.w3(32'h3b3cf8a9),
	.w4(32'h3bf99fa5),
	.w5(32'hbb698629),
	.w6(32'h3c73cd41),
	.w7(32'h3c37a1ea),
	.w8(32'hba111d19),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ddbc),
	.w1(32'h3a433644),
	.w2(32'h3b0b6eb6),
	.w3(32'hbb9e6079),
	.w4(32'h3aa90070),
	.w5(32'h3aaa08c1),
	.w6(32'h3b0af435),
	.w7(32'h3c3ff3e8),
	.w8(32'h3b6d1b00),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14b200),
	.w1(32'hbade61b3),
	.w2(32'h3a87cdda),
	.w3(32'hbc168292),
	.w4(32'hbb0dea22),
	.w5(32'h3b4baa1c),
	.w6(32'h3c1021d7),
	.w7(32'hb9d71ac3),
	.w8(32'h3b61fb32),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974c995),
	.w1(32'h3aefcd50),
	.w2(32'h3b7e73d0),
	.w3(32'hbaa4b4aa),
	.w4(32'hb9ec4d98),
	.w5(32'hb97bfb26),
	.w6(32'h3ad980ff),
	.w7(32'h3b2b4f25),
	.w8(32'hb9f4abab),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4620c),
	.w1(32'h3b5520a2),
	.w2(32'h3bc421a3),
	.w3(32'h39736ea3),
	.w4(32'h3ae38132),
	.w5(32'h3bfb389b),
	.w6(32'hba2beaae),
	.w7(32'h3aa46829),
	.w8(32'h3bf15f46),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58837d),
	.w1(32'h3c1031ac),
	.w2(32'hbc037211),
	.w3(32'h3b413f4e),
	.w4(32'hbb0d3f7d),
	.w5(32'hbbc62f9b),
	.w6(32'h3c105998),
	.w7(32'h3c02b669),
	.w8(32'h3b7c186c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ef59c),
	.w1(32'hba05fb9b),
	.w2(32'hbaf8efd7),
	.w3(32'hbbe7093d),
	.w4(32'h3bcdbcac),
	.w5(32'h3b20ad8b),
	.w6(32'h3bbc024c),
	.w7(32'hbb0011d5),
	.w8(32'h3ad8ab58),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0502c4),
	.w1(32'h3b0a059e),
	.w2(32'h3c2cee38),
	.w3(32'h3a8293ee),
	.w4(32'hba27e210),
	.w5(32'h3a0cf639),
	.w6(32'h37efc440),
	.w7(32'h3b1a6128),
	.w8(32'h3c291424),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba5442),
	.w1(32'h3caa00c5),
	.w2(32'h3c536a1e),
	.w3(32'h3bc91535),
	.w4(32'h3c0270cc),
	.w5(32'h3be02be8),
	.w6(32'h3c97b0b6),
	.w7(32'h3c5f81bc),
	.w8(32'h3bc831f9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d54c3),
	.w1(32'h3c4f23e9),
	.w2(32'h3b9b57b4),
	.w3(32'h3c13c786),
	.w4(32'h3c1829c2),
	.w5(32'hbb2381de),
	.w6(32'h3b8e6a3c),
	.w7(32'h3bd0e06d),
	.w8(32'hbac3bed0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0352e8),
	.w1(32'h3c0690f7),
	.w2(32'h3b8bb66d),
	.w3(32'hba2db194),
	.w4(32'h3ad348a1),
	.w5(32'hba0719c0),
	.w6(32'h3b2d55e5),
	.w7(32'h3b79ef31),
	.w8(32'hbb402ff6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba163c89),
	.w1(32'h3b8a5254),
	.w2(32'hbbc54b3a),
	.w3(32'hbc119ff7),
	.w4(32'hbb6da575),
	.w5(32'hbb84bd57),
	.w6(32'hbb676007),
	.w7(32'hbb11be11),
	.w8(32'h394c9728),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27fd92),
	.w1(32'hbb9f3f13),
	.w2(32'h3bac2948),
	.w3(32'hbbd6d6db),
	.w4(32'h3b4834c4),
	.w5(32'h3b4a2001),
	.w6(32'hbc195aa8),
	.w7(32'hbc470cee),
	.w8(32'hbb651013),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0673c3),
	.w1(32'h3a7c6e60),
	.w2(32'h3bdbd290),
	.w3(32'h3c6abda2),
	.w4(32'h3c4f4d4a),
	.w5(32'h3af1d64f),
	.w6(32'hbc25970c),
	.w7(32'hbb58e7d8),
	.w8(32'h3bebf2af),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd023),
	.w1(32'h385c7571),
	.w2(32'hbb642778),
	.w3(32'h3c1f0784),
	.w4(32'h3c68970e),
	.w5(32'h3b8a742e),
	.w6(32'hbba06aaf),
	.w7(32'h3bc97dfc),
	.w8(32'hbc07b8ed),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc549c00),
	.w1(32'hbc000092),
	.w2(32'h3c08919b),
	.w3(32'hbbce9372),
	.w4(32'h3b8ad02f),
	.w5(32'hba83b20c),
	.w6(32'hbb309536),
	.w7(32'h3b187b58),
	.w8(32'h3be8808c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ec6f7),
	.w1(32'h3c982156),
	.w2(32'hbbdef0a2),
	.w3(32'hba61b908),
	.w4(32'h3b89d534),
	.w5(32'h3b53d3b5),
	.w6(32'h3b013cc5),
	.w7(32'h3bd8daac),
	.w8(32'hbc3f4c42),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba705d2),
	.w1(32'hbc8d6e6f),
	.w2(32'hbc270583),
	.w3(32'h3cbc4c11),
	.w4(32'h3c9e090e),
	.w5(32'h3c0bdc8c),
	.w6(32'hbc772a52),
	.w7(32'hbc71ac1c),
	.w8(32'hbc8a3025),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e7fb4),
	.w1(32'hbc9b7bf7),
	.w2(32'hbbd71482),
	.w3(32'h3cb45382),
	.w4(32'h3c64fea2),
	.w5(32'hbbc94a5a),
	.w6(32'hbc82e998),
	.w7(32'hbc9891e0),
	.w8(32'hbb897cd3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0496da),
	.w1(32'hbc2f2790),
	.w2(32'hbb5fa708),
	.w3(32'hbb06aa5f),
	.w4(32'hb824bfe6),
	.w5(32'hbb36ed9c),
	.w6(32'hbaba9281),
	.w7(32'hbb33d860),
	.w8(32'hbb0da057),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2846f4),
	.w1(32'hbc4b31c0),
	.w2(32'h3b6996c2),
	.w3(32'hbc18392f),
	.w4(32'hbb55cfa8),
	.w5(32'h3909caa1),
	.w6(32'hbb9f1982),
	.w7(32'h3bbc6354),
	.w8(32'h3c5b30dc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1811e),
	.w1(32'h3b905d23),
	.w2(32'h3b1ca2ac),
	.w3(32'hbb5ec803),
	.w4(32'hbb2887bb),
	.w5(32'h3aa59184),
	.w6(32'h3c37e298),
	.w7(32'h3c94e3ae),
	.w8(32'hb957a4b4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d04ad),
	.w1(32'hb9718a99),
	.w2(32'h3bd095e9),
	.w3(32'hbaeda3d2),
	.w4(32'h3b48a0f7),
	.w5(32'h3bc3044d),
	.w6(32'h3b0d685d),
	.w7(32'hb88d5e89),
	.w8(32'h3be9dfa2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cdae7),
	.w1(32'h3a026c0d),
	.w2(32'hbc752334),
	.w3(32'hbabffbf1),
	.w4(32'h3aebce55),
	.w5(32'hbb8742ff),
	.w6(32'h3b818a0d),
	.w7(32'h3b298d14),
	.w8(32'h3af4867f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc542597),
	.w1(32'hbc094b99),
	.w2(32'h3be0776a),
	.w3(32'hbb8a4c33),
	.w4(32'h399e4fc1),
	.w5(32'hbc08aacd),
	.w6(32'h39ca3323),
	.w7(32'hbbc10456),
	.w8(32'hbb757d93),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb457a6),
	.w1(32'hbaa3c4df),
	.w2(32'hbc526fa9),
	.w3(32'h3a09c9f9),
	.w4(32'hbbc0fcfd),
	.w5(32'h3c2bc6d5),
	.w6(32'hba136c2e),
	.w7(32'hbbd37579),
	.w8(32'hbc0fb8ef),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc498d98),
	.w1(32'hbc628c2c),
	.w2(32'h3c549269),
	.w3(32'h3c819bee),
	.w4(32'h3c61d834),
	.w5(32'hbab29c38),
	.w6(32'hbc7a0357),
	.w7(32'hbbe9dc7b),
	.w8(32'h3b2b4c86),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18870d),
	.w1(32'h3a3a1f61),
	.w2(32'h3962b832),
	.w3(32'h3c438676),
	.w4(32'h3c9e41ec),
	.w5(32'hbc3e0698),
	.w6(32'hbbdff593),
	.w7(32'h3b4beef0),
	.w8(32'hb9a9b158),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c275b13),
	.w1(32'h3c272a64),
	.w2(32'h3b4e0560),
	.w3(32'hbc6600e1),
	.w4(32'hbc5aba61),
	.w5(32'h3b3fc6f5),
	.w6(32'h3baefa2a),
	.w7(32'h3ac8853d),
	.w8(32'h3c0408ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab44a58),
	.w1(32'h3bbee7aa),
	.w2(32'hbcb18b7a),
	.w3(32'h3b13443a),
	.w4(32'h3b8dcbf4),
	.w5(32'hbc0c4623),
	.w6(32'hb9f0a9f3),
	.w7(32'h3b3babee),
	.w8(32'hbb45b086),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e0703),
	.w1(32'hbca998c0),
	.w2(32'hbbe1329f),
	.w3(32'hbafeece2),
	.w4(32'hba2d44e7),
	.w5(32'h3cd2025d),
	.w6(32'hbb8fe862),
	.w7(32'hbc3e1bf2),
	.w8(32'hba118c1a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ff55c),
	.w1(32'hbc79b72c),
	.w2(32'h38b442b4),
	.w3(32'h3d056900),
	.w4(32'h3cbe69f4),
	.w5(32'hba2f521c),
	.w6(32'h3bcd46f6),
	.w7(32'h3ba88636),
	.w8(32'h3b6b1543),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031601),
	.w1(32'h3ab73ad5),
	.w2(32'h3b957100),
	.w3(32'hbaf95506),
	.w4(32'hbacb4eb3),
	.w5(32'hba1850e2),
	.w6(32'h3aff64d3),
	.w7(32'h3aaa3f2c),
	.w8(32'h3c0c130c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59e8cf),
	.w1(32'h3c308ee4),
	.w2(32'hbbe1fff0),
	.w3(32'hbbc5e699),
	.w4(32'h3a519b98),
	.w5(32'hbb8694eb),
	.w6(32'h3bc0b424),
	.w7(32'h3c05ecd9),
	.w8(32'h3bc12b3b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00cf50),
	.w1(32'hbbcc99e1),
	.w2(32'hbb211522),
	.w3(32'hbb9cd440),
	.w4(32'hbb38d8e9),
	.w5(32'hbc04abe5),
	.w6(32'h3bf67e57),
	.w7(32'h3b8c6cc5),
	.w8(32'hbbb2f0b7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ba58),
	.w1(32'hbc28a9fd),
	.w2(32'hbc13e2f7),
	.w3(32'h3b4b0988),
	.w4(32'h3bbb8e33),
	.w5(32'h3bf3c920),
	.w6(32'hbc037466),
	.w7(32'hbc27f02b),
	.w8(32'hbc7bca24),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c72bf),
	.w1(32'hbc8fe205),
	.w2(32'hb8fe1685),
	.w3(32'h3cd4e5d7),
	.w4(32'h3c948772),
	.w5(32'h3adef810),
	.w6(32'hbc897a67),
	.w7(32'hbc545d24),
	.w8(32'hbc4d5f42),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf032),
	.w1(32'hbb1a237c),
	.w2(32'h37fb8e9b),
	.w3(32'h3a73f183),
	.w4(32'h39a5b6b4),
	.w5(32'hb9d4979a),
	.w6(32'hbc56ea88),
	.w7(32'hbbbe04f3),
	.w8(32'hb92dcfdb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e4ef3),
	.w1(32'hb82a09ea),
	.w2(32'hb9ee7a43),
	.w3(32'hbb51b36d),
	.w4(32'hb9921b62),
	.w5(32'hbb21a21e),
	.w6(32'h39223a6c),
	.w7(32'hba19ab53),
	.w8(32'hbb3c6fbe),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab739f7),
	.w1(32'hb90a5b4e),
	.w2(32'h3c32cc47),
	.w3(32'hba74aa6c),
	.w4(32'hbaf3c469),
	.w5(32'h3b96ed3e),
	.w6(32'hbb1af591),
	.w7(32'hbafbaa2c),
	.w8(32'h3b730c31),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbed5cc),
	.w1(32'hbc488992),
	.w2(32'h3b24763d),
	.w3(32'hb91dc703),
	.w4(32'hbc2b80ca),
	.w5(32'h39829db6),
	.w6(32'hbbf8107a),
	.w7(32'hbc65cc4d),
	.w8(32'h3ab4dce9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1030c),
	.w1(32'h3afcfb98),
	.w2(32'hbb3c9afc),
	.w3(32'hbade70de),
	.w4(32'h3ab83870),
	.w5(32'hba25f48f),
	.w6(32'h3adc82d2),
	.w7(32'h3ba744e3),
	.w8(32'h3ae5343a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6091b9),
	.w1(32'h3b826f6b),
	.w2(32'hba84c465),
	.w3(32'h397b23e9),
	.w4(32'hbbb1fd19),
	.w5(32'hbaa63ea0),
	.w6(32'h3bc4c466),
	.w7(32'hbaf4b60d),
	.w8(32'h3b76d78e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a738bb2),
	.w1(32'h3aa00526),
	.w2(32'hba03afd9),
	.w3(32'hbb660787),
	.w4(32'hbbec2edf),
	.w5(32'hbb4b67d0),
	.w6(32'h3bc62b91),
	.w7(32'h3bd467bd),
	.w8(32'h3b0aae9d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b130008),
	.w1(32'hbb64d63a),
	.w2(32'hbc30f40d),
	.w3(32'h3a98a0d7),
	.w4(32'hbc1b0595),
	.w5(32'hbb3dca61),
	.w6(32'h3ba53748),
	.w7(32'hbb401c0e),
	.w8(32'h3b684480),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e98c0),
	.w1(32'hbb10fee5),
	.w2(32'hbc886acd),
	.w3(32'hbb1eb5b9),
	.w4(32'hbc5037b1),
	.w5(32'h3bb86c18),
	.w6(32'h3b4be0ea),
	.w7(32'h3bddc753),
	.w8(32'hbc9015e0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc948beb),
	.w1(32'hbc2584f9),
	.w2(32'hbb6f8afb),
	.w3(32'h3c768740),
	.w4(32'h3c58c341),
	.w5(32'hbb7902df),
	.w6(32'hbc8c1c76),
	.w7(32'hbc480932),
	.w8(32'h3bf0fe46),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a140a),
	.w1(32'h3bfbc031),
	.w2(32'h3b4df68f),
	.w3(32'h3aa5e92a),
	.w4(32'hb89e159a),
	.w5(32'hbafc7565),
	.w6(32'h3c82371f),
	.w7(32'h3c080975),
	.w8(32'hbb54c5ae),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e897f),
	.w1(32'hbbc93f3f),
	.w2(32'h3ca98e9c),
	.w3(32'h3c800db2),
	.w4(32'h3ca076e0),
	.w5(32'h3c40f9ce),
	.w6(32'hbc4458c1),
	.w7(32'hbc5fb2b7),
	.w8(32'h3c1d7061),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf6a2c),
	.w1(32'h3ca4e431),
	.w2(32'h3bb61dce),
	.w3(32'hba5736d0),
	.w4(32'hbba810d0),
	.w5(32'hbb21934d),
	.w6(32'h3b95144b),
	.w7(32'h3c33a081),
	.w8(32'h3bfa0881),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3eeda),
	.w1(32'hbb283c3b),
	.w2(32'h39badd13),
	.w3(32'hbc26afa3),
	.w4(32'hbb8b35a3),
	.w5(32'hbbcf889c),
	.w6(32'h3bfa2cbd),
	.w7(32'h3b00d77c),
	.w8(32'hbb404a8d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec632c),
	.w1(32'hb9ab12eb),
	.w2(32'hbbdc7ec4),
	.w3(32'hbb2ac6da),
	.w4(32'hbb7d1302),
	.w5(32'h3adf933a),
	.w6(32'hbb1528f2),
	.w7(32'hbaced032),
	.w8(32'hbb2e79a0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e527e),
	.w1(32'hbc6d465f),
	.w2(32'hbc17b884),
	.w3(32'h3afa1fcc),
	.w4(32'h3af91842),
	.w5(32'hbab04f48),
	.w6(32'hbbfbe16b),
	.w7(32'hbb408da2),
	.w8(32'h3ba82a4a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c04f2),
	.w1(32'hbb7cb24d),
	.w2(32'h3c32e85a),
	.w3(32'hbc86c1bc),
	.w4(32'hbba2cfd7),
	.w5(32'h3c557596),
	.w6(32'hbb4813fe),
	.w7(32'hbc361e4a),
	.w8(32'hbbca3b0b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c229fcf),
	.w1(32'h3c03081c),
	.w2(32'hbaa2ba6f),
	.w3(32'h3c820fe2),
	.w4(32'h3c33ef76),
	.w5(32'hbb67f969),
	.w6(32'hbc209313),
	.w7(32'hbbb7f752),
	.w8(32'hba74529b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118814),
	.w1(32'h3b042194),
	.w2(32'hbc6c36f5),
	.w3(32'hba9bebaa),
	.w4(32'hbab45e88),
	.w5(32'h3cb61e8f),
	.w6(32'h3a7d9e93),
	.w7(32'h3b30cd00),
	.w8(32'hbc18f76a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc471ed7),
	.w1(32'hbbaa1f9f),
	.w2(32'h3b54081f),
	.w3(32'h3cce37da),
	.w4(32'h3c1c07a0),
	.w5(32'hb91918db),
	.w6(32'hbc62d2d7),
	.w7(32'hbadec0ab),
	.w8(32'h39d525ef),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba20a4b),
	.w1(32'h3b9f2a53),
	.w2(32'h3b4181d4),
	.w3(32'h3a26a5d2),
	.w4(32'h39fc9706),
	.w5(32'hbbb58ed0),
	.w6(32'h3ac9e610),
	.w7(32'h3aa29607),
	.w8(32'h3b5f8d15),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc0795),
	.w1(32'h3b997c68),
	.w2(32'h3cfe5ec1),
	.w3(32'hbb1572a0),
	.w4(32'h3b9872b5),
	.w5(32'h3b7beb7b),
	.w6(32'h3afeec34),
	.w7(32'h3b3419d7),
	.w8(32'h3c65b75d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0757c5),
	.w1(32'h3d0836d6),
	.w2(32'hbb9a6886),
	.w3(32'h3a2c93fc),
	.w4(32'h3c67fadd),
	.w5(32'hbbc64705),
	.w6(32'h3ccf5a8f),
	.w7(32'h3c58f9b9),
	.w8(32'h3b82a77d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39fd82),
	.w1(32'h3955e5dc),
	.w2(32'h37b9ae74),
	.w3(32'hbc03c00a),
	.w4(32'hbba2c968),
	.w5(32'hbbb2d957),
	.w6(32'h3bcb6f3e),
	.w7(32'h3b358276),
	.w8(32'h3924ba24),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ceaae),
	.w1(32'h3b54307b),
	.w2(32'hbb45974d),
	.w3(32'hbb31abc9),
	.w4(32'hbb07068b),
	.w5(32'hbb8d017d),
	.w6(32'h3b65d90a),
	.w7(32'h3b8ac773),
	.w8(32'h3bb271b3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad13a),
	.w1(32'hbaf0cee8),
	.w2(32'h3c1accd4),
	.w3(32'hba5d71c1),
	.w4(32'hba8fa68b),
	.w5(32'h3b85a86c),
	.w6(32'h3bcf02b8),
	.w7(32'h3c115a9e),
	.w8(32'h38dd873b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19e262),
	.w1(32'h3b2ebb2b),
	.w2(32'hbb177cfc),
	.w3(32'h3b182e62),
	.w4(32'h39e97156),
	.w5(32'hbc17e119),
	.w6(32'h3b0ca223),
	.w7(32'h3bfb87a7),
	.w8(32'hbb92d31a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4baab),
	.w1(32'hbbb4e38f),
	.w2(32'h39db5995),
	.w3(32'h3bfc8601),
	.w4(32'h3c664b5b),
	.w5(32'hbba9ff73),
	.w6(32'hbc431f2b),
	.w7(32'hbc3a978d),
	.w8(32'hbaa49333),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cb45),
	.w1(32'hbb0aef1f),
	.w2(32'h3c61c41a),
	.w3(32'hbbe78735),
	.w4(32'hbb9596a5),
	.w5(32'h3b030b08),
	.w6(32'hba458317),
	.w7(32'h3b89e1bf),
	.w8(32'h3bf0258d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf855a),
	.w1(32'h3bad09de),
	.w2(32'hbb4d51ed),
	.w3(32'hba5ade01),
	.w4(32'h3a82875c),
	.w5(32'hbb323ddc),
	.w6(32'h3baec41b),
	.w7(32'h3c186372),
	.w8(32'hbb88c78b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ec4de),
	.w1(32'hbb74c2c6),
	.w2(32'h3b56e69c),
	.w3(32'hbb3f3535),
	.w4(32'hba7ffa8a),
	.w5(32'hbafc43e6),
	.w6(32'hbbde73d3),
	.w7(32'hbb438453),
	.w8(32'hbb0a4266),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812987),
	.w1(32'h3b512315),
	.w2(32'h3b4a8462),
	.w3(32'h3a6af31d),
	.w4(32'h3aa6300f),
	.w5(32'hb8900367),
	.w6(32'hba829275),
	.w7(32'hba119caa),
	.w8(32'h3b1c33c1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba93cb9),
	.w1(32'h3b9dbaab),
	.w2(32'h3ce0e4ca),
	.w3(32'h3b3e2c1d),
	.w4(32'hbb48b17b),
	.w5(32'hbcb6364a),
	.w6(32'hba60ec10),
	.w7(32'h3bdff4c3),
	.w8(32'h3c90c4fc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d18e71e),
	.w1(32'h3c6807ce),
	.w2(32'hbaeec90a),
	.w3(32'hbca7cbe9),
	.w4(32'hbb120adf),
	.w5(32'h3c8f6272),
	.w6(32'h3c12d184),
	.w7(32'hbbdde1ef),
	.w8(32'hbbb50262),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75ec49),
	.w1(32'h3b01fea0),
	.w2(32'hb9bf9694),
	.w3(32'h39da105a),
	.w4(32'h3bd8f4ae),
	.w5(32'h3b4e253e),
	.w6(32'hbbc4b8b7),
	.w7(32'hbb70b8ab),
	.w8(32'hb979c3f0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e29dfc),
	.w1(32'hb9124bd3),
	.w2(32'h3ac42f86),
	.w3(32'h3ab54b54),
	.w4(32'h3b3c96cf),
	.w5(32'h3b0daf8f),
	.w6(32'hba3ae975),
	.w7(32'hba32758b),
	.w8(32'hbaccac2a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5980),
	.w1(32'h3ab07947),
	.w2(32'h3c28d0b2),
	.w3(32'h3b8625b8),
	.w4(32'h3c187157),
	.w5(32'h3c82c139),
	.w6(32'h3b9690a6),
	.w7(32'h3c72f6ea),
	.w8(32'hba2349a1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c345380),
	.w1(32'h3c781ce8),
	.w2(32'hb8e6f357),
	.w3(32'h3c991bb4),
	.w4(32'h3c77559c),
	.w5(32'h39bf2d40),
	.w6(32'h3c34edf8),
	.w7(32'h3c85ecd4),
	.w8(32'h3b89025b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd1c1),
	.w1(32'h3b5b1028),
	.w2(32'hbca47382),
	.w3(32'hbb858629),
	.w4(32'hbb8a72ba),
	.w5(32'hbc357967),
	.w6(32'h3a064157),
	.w7(32'hbb046cd7),
	.w8(32'hbbb451f5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c5f6b),
	.w1(32'hbbac1532),
	.w2(32'h3c144c77),
	.w3(32'hbc6eca73),
	.w4(32'hbb458016),
	.w5(32'h3c3f8409),
	.w6(32'hbb9f8a73),
	.w7(32'hbb2affbc),
	.w8(32'h3b90cf33),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e540c),
	.w1(32'h3a39ded2),
	.w2(32'hba81ef5e),
	.w3(32'h3c908fe1),
	.w4(32'h3c70ef56),
	.w5(32'hba936fb9),
	.w6(32'h3c4fd09e),
	.w7(32'h3cb2de73),
	.w8(32'h3ae22cb3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1beb91),
	.w1(32'h3ad1f2ac),
	.w2(32'hbc4b1e8b),
	.w3(32'hbc023c6b),
	.w4(32'hbb8674c9),
	.w5(32'hbca15e4b),
	.w6(32'hba6073f0),
	.w7(32'hbba6a21e),
	.w8(32'hbc86c961),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9397b7),
	.w1(32'hbbe90359),
	.w2(32'hbb91c03f),
	.w3(32'hbcdb7108),
	.w4(32'hbca52022),
	.w5(32'hbb097542),
	.w6(32'hbc867c95),
	.w7(32'hbcbd6ffc),
	.w8(32'hbb3e3b01),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a7c0),
	.w1(32'h3adee35d),
	.w2(32'hbb43cc89),
	.w3(32'hba532360),
	.w4(32'h3ae38b1a),
	.w5(32'h3b929bd9),
	.w6(32'h3a887210),
	.w7(32'h3afdcc9b),
	.w8(32'hbaf6f312),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bd5ad),
	.w1(32'hbb8a7562),
	.w2(32'hba99e47d),
	.w3(32'hbb7c1184),
	.w4(32'hbbf85d49),
	.w5(32'h3b2824be),
	.w6(32'h3b7cb44e),
	.w7(32'hbaa8aa47),
	.w8(32'h3ab0eee1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e78ae),
	.w1(32'h3b3b8b1a),
	.w2(32'hbad83abc),
	.w3(32'h3ad9e0e7),
	.w4(32'h39984310),
	.w5(32'hba67936d),
	.w6(32'h3b9e862b),
	.w7(32'h3a73708e),
	.w8(32'hbb490e75),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd9b2),
	.w1(32'h3bde96f0),
	.w2(32'hbae584cf),
	.w3(32'h3af86ca8),
	.w4(32'h3ab8e022),
	.w5(32'h3a77ea68),
	.w6(32'h3bbe3943),
	.w7(32'hbae1ced8),
	.w8(32'h3c2d3143),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6346354),
	.w1(32'h3957ba97),
	.w2(32'h39c63f33),
	.w3(32'hbadbda8e),
	.w4(32'hba68ccc5),
	.w5(32'hbb98f917),
	.w6(32'h3ba68c1c),
	.w7(32'h3c121cb6),
	.w8(32'hba7d36d1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b839b),
	.w1(32'h3c10731d),
	.w2(32'hbc564b9a),
	.w3(32'hb9c194b5),
	.w4(32'h3aee522c),
	.w5(32'hbb02c7b8),
	.w6(32'hbb8e71c3),
	.w7(32'h3ae776a3),
	.w8(32'hb6b8c467),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc93398),
	.w1(32'hba1d4370),
	.w2(32'h3d12e5a0),
	.w3(32'h3bf97f29),
	.w4(32'h3ab1884e),
	.w5(32'h3d1939de),
	.w6(32'h3ac720c1),
	.w7(32'hbb62ad96),
	.w8(32'h3c894145),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1f633f),
	.w1(32'h3cda1499),
	.w2(32'hbb28ba6c),
	.w3(32'h3d5c7650),
	.w4(32'h3d42241c),
	.w5(32'hbacf692f),
	.w6(32'h3d1a37e7),
	.w7(32'h3d30005c),
	.w8(32'hbb58e826),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac5257),
	.w1(32'h3a9359a9),
	.w2(32'hbbb846d4),
	.w3(32'h3b4ddb59),
	.w4(32'h3ba2aafb),
	.w5(32'hbc7b72c9),
	.w6(32'hba2c2420),
	.w7(32'h3af79c73),
	.w8(32'hbc33bf91),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1bfa),
	.w1(32'h3bdea7da),
	.w2(32'h3be518ad),
	.w3(32'hbc82b7cf),
	.w4(32'hbb9a5556),
	.w5(32'hbbbdb0ab),
	.w6(32'hbca7427a),
	.w7(32'hbc349513),
	.w8(32'hbc7a84ee),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd8b7),
	.w1(32'hbc147f3e),
	.w2(32'hbcc8887b),
	.w3(32'hbc50d838),
	.w4(32'hbcbb61ec),
	.w5(32'hbc95bae1),
	.w6(32'hbc0de95d),
	.w7(32'hbc8c6674),
	.w8(32'h3a25bbd4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78d9ad),
	.w1(32'h3babaeda),
	.w2(32'hbab501ff),
	.w3(32'hbcf43718),
	.w4(32'hbc99231e),
	.w5(32'hba4c7f77),
	.w6(32'hbc7e831f),
	.w7(32'hbccd2487),
	.w8(32'h3bf4365c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e27a7),
	.w1(32'h3aec1d79),
	.w2(32'hbb458040),
	.w3(32'hba369892),
	.w4(32'hbc60f283),
	.w5(32'h3b014717),
	.w6(32'hbb85d680),
	.w7(32'hbb9ed757),
	.w8(32'hb9082198),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab580ae),
	.w1(32'hbb23202e),
	.w2(32'h3be04873),
	.w3(32'h3bc678e6),
	.w4(32'h3b8e254f),
	.w5(32'h3b956b89),
	.w6(32'h3b3bca57),
	.w7(32'h3b972702),
	.w8(32'hba42207a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4cc9),
	.w1(32'h3bf1bc9f),
	.w2(32'hbb27bb6d),
	.w3(32'h3bf4259d),
	.w4(32'h3c34b44d),
	.w5(32'hbc72077c),
	.w6(32'h3b88c107),
	.w7(32'h3a94e9d8),
	.w8(32'hbc6fbee3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16e52d),
	.w1(32'hbc4c1dac),
	.w2(32'hbcadfe30),
	.w3(32'hbc355117),
	.w4(32'hbc76ffba),
	.w5(32'hbcb67221),
	.w6(32'hbc71c30d),
	.w7(32'hbc5691df),
	.w8(32'hbc29bc3b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bd61d),
	.w1(32'hbbe07333),
	.w2(32'hbbd8875d),
	.w3(32'hbd18a850),
	.w4(32'hbcc97782),
	.w5(32'hbc205155),
	.w6(32'hbcc5fe2a),
	.w7(32'hbcd07397),
	.w8(32'hbbf3dea2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba945c5),
	.w1(32'hbb868516),
	.w2(32'h3a33d270),
	.w3(32'h3b0d38ef),
	.w4(32'h3b042ee4),
	.w5(32'hbbabd400),
	.w6(32'h3a3c1dd3),
	.w7(32'h391307dd),
	.w8(32'hbbc1a8ee),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85da7d),
	.w1(32'hbb29a59d),
	.w2(32'h3be89eab),
	.w3(32'hbb11da66),
	.w4(32'hba8f98d2),
	.w5(32'h3bea2308),
	.w6(32'hba939e50),
	.w7(32'h3c20517a),
	.w8(32'hbbeb1f71),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27fa42),
	.w1(32'h3c158b5d),
	.w2(32'hba4c08c8),
	.w3(32'hba33633a),
	.w4(32'h3b853a81),
	.w5(32'hbc5bb6ce),
	.w6(32'hbb0771e0),
	.w7(32'h3c607ea0),
	.w8(32'h3be32cc0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9d181),
	.w1(32'h3a8341e7),
	.w2(32'h3ba54140),
	.w3(32'hbc333aa5),
	.w4(32'h3af36b07),
	.w5(32'h3bfdca40),
	.w6(32'hbc0e1a2c),
	.w7(32'hbb3df09c),
	.w8(32'hbaab8be4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb966af),
	.w1(32'h3c36ca42),
	.w2(32'h3abed74f),
	.w3(32'h3bb3b6cb),
	.w4(32'h3b83ee28),
	.w5(32'hbaed2e0f),
	.w6(32'hba07d76b),
	.w7(32'h3c14234d),
	.w8(32'hba047cc3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8eca6),
	.w1(32'hbbbd7cc0),
	.w2(32'h392faeac),
	.w3(32'hbbf50072),
	.w4(32'hbb3cb551),
	.w5(32'h3b5a2012),
	.w6(32'hbbb0215d),
	.w7(32'hba36e90b),
	.w8(32'h3ba9753b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46abfa),
	.w1(32'h3c37f0ad),
	.w2(32'h3ad8c2f0),
	.w3(32'h3ab80ce0),
	.w4(32'h3c683880),
	.w5(32'hba9ee3e5),
	.w6(32'h3bfa522d),
	.w7(32'h3c8c41ce),
	.w8(32'hbb66a847),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca9e95),
	.w1(32'h3b8c3e09),
	.w2(32'hbba3b2af),
	.w3(32'hba52727d),
	.w4(32'hbb0fe379),
	.w5(32'hbb89025a),
	.w6(32'hbae2cf9b),
	.w7(32'h3b2256ca),
	.w8(32'h3a902d19),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99bd63),
	.w1(32'hbbf95d6a),
	.w2(32'hba36a689),
	.w3(32'hbab79e46),
	.w4(32'hba921e0b),
	.w5(32'h3bde3f3d),
	.w6(32'h3b0f2865),
	.w7(32'hba93fa2b),
	.w8(32'h3b0bd63d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8041),
	.w1(32'h3c08b8fb),
	.w2(32'hbc55fd4d),
	.w3(32'h3be32278),
	.w4(32'h3bb3a780),
	.w5(32'hbca596cf),
	.w6(32'h3b5605a6),
	.w7(32'hbb1ba27f),
	.w8(32'hbc41eecd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe24af),
	.w1(32'hbc49ff05),
	.w2(32'hbbe89638),
	.w3(32'hbd03e631),
	.w4(32'hbd05ace4),
	.w5(32'hbadbf223),
	.w6(32'hbcea63b6),
	.w7(32'hbcc51579),
	.w8(32'hb9ccdcc2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe84b6),
	.w1(32'hba75bb66),
	.w2(32'h3ac6285d),
	.w3(32'hbc3f0257),
	.w4(32'hbc2df8b0),
	.w5(32'hbb69b3cf),
	.w6(32'hbc135a29),
	.w7(32'hbc3093a2),
	.w8(32'h3c173934),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7d035),
	.w1(32'h3afba429),
	.w2(32'h3b6d4eac),
	.w3(32'hbc2f10a0),
	.w4(32'hba4fb388),
	.w5(32'h3a022726),
	.w6(32'hbbb9f153),
	.w7(32'hbb9f5afc),
	.w8(32'h3bca0b7e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c220b),
	.w1(32'h39ffe404),
	.w2(32'hbb447d9e),
	.w3(32'h3b3a98ff),
	.w4(32'h3a559b50),
	.w5(32'hbae09383),
	.w6(32'h3c1bc14a),
	.w7(32'h3c18c8f3),
	.w8(32'hba42a818),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba216f94),
	.w1(32'hba910333),
	.w2(32'h3a6cd45c),
	.w3(32'hb9be6c40),
	.w4(32'h3a777263),
	.w5(32'h3af14f1f),
	.w6(32'hb97acba9),
	.w7(32'hba151a6c),
	.w8(32'h3bd19b5c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67db3b),
	.w1(32'h3b69af72),
	.w2(32'hbb816247),
	.w3(32'h3bec8d19),
	.w4(32'h3b46a572),
	.w5(32'hbba3b4ce),
	.w6(32'h3c34d930),
	.w7(32'h3c2d7787),
	.w8(32'hbc2adf5e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe16d9),
	.w1(32'hbc0fd8f6),
	.w2(32'h3bf7609a),
	.w3(32'hbaf2f614),
	.w4(32'h3b1cf6a9),
	.w5(32'h3c08d835),
	.w6(32'hbb08f12b),
	.w7(32'hbb1713a9),
	.w8(32'h3bdae3c2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfff9d),
	.w1(32'h3bc7f486),
	.w2(32'hbc05d4e7),
	.w3(32'h3c2bc472),
	.w4(32'h3c01a988),
	.w5(32'hbb8d08d0),
	.w6(32'h3c06f4a5),
	.w7(32'h3c0ac533),
	.w8(32'hbab5abf9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861ed35),
	.w1(32'h3b652e35),
	.w2(32'h3ac7865e),
	.w3(32'hbbb2e9e9),
	.w4(32'h3b17a6b8),
	.w5(32'h3b9c82f4),
	.w6(32'hbc1cfd40),
	.w7(32'hbb7a3939),
	.w8(32'h3a0e5c02),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5251),
	.w1(32'hbb674ecd),
	.w2(32'hbc64d2fe),
	.w3(32'h3bd9d413),
	.w4(32'hb9c5d850),
	.w5(32'hbbc82e52),
	.w6(32'hbb3476a2),
	.w7(32'h3ae14ed7),
	.w8(32'h3c25319e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc784df9),
	.w1(32'h3bb62e52),
	.w2(32'hbc09511d),
	.w3(32'hbc8f1724),
	.w4(32'hbc35c35b),
	.w5(32'hbc884835),
	.w6(32'hb8a99e2f),
	.w7(32'hbc35a1b7),
	.w8(32'hbc703cb9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd75711),
	.w1(32'hbb81c9c0),
	.w2(32'hbbe32f5d),
	.w3(32'hbc5c28ac),
	.w4(32'hbbd5f858),
	.w5(32'hbb1c8320),
	.w6(32'hbc842498),
	.w7(32'hbc3b04ce),
	.w8(32'hbbb2cfe8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb630176),
	.w1(32'h3895bd5c),
	.w2(32'hbc466088),
	.w3(32'h3a9cbf2c),
	.w4(32'h3a2953b9),
	.w5(32'hbc015783),
	.w6(32'hbb8136ed),
	.w7(32'hbb27f8d0),
	.w8(32'hbb5c6568),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0efff2),
	.w1(32'hbb843f80),
	.w2(32'h3c7b29ea),
	.w3(32'hbc038893),
	.w4(32'hbb020a70),
	.w5(32'h3cf3a47e),
	.w6(32'hbbaee7d2),
	.w7(32'hbab7004b),
	.w8(32'h3c9e1b10),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc49d87),
	.w1(32'h3c7b85ed),
	.w2(32'h3a3d0ca6),
	.w3(32'h3d026623),
	.w4(32'h3cadb956),
	.w5(32'hbbc56b57),
	.w6(32'h3cf4efc1),
	.w7(32'h3c75aee7),
	.w8(32'h3b01125d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718e3c),
	.w1(32'h3abc6ff9),
	.w2(32'h3b0a1e37),
	.w3(32'hbb3896dd),
	.w4(32'hbba3f089),
	.w5(32'h3bcb0dbc),
	.w6(32'hbac72783),
	.w7(32'hbc3aeb4c),
	.w8(32'h3b455f10),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8fdd7),
	.w1(32'h3b37d125),
	.w2(32'h39eac159),
	.w3(32'h3c3f0bc2),
	.w4(32'h3bfdcf77),
	.w5(32'h3b8e8c35),
	.w6(32'h3bb46fe4),
	.w7(32'h3888049e),
	.w8(32'h3ae27fb5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18546d),
	.w1(32'hb900dd17),
	.w2(32'h3c2c4144),
	.w3(32'h3b98f97c),
	.w4(32'h3bffaaf1),
	.w5(32'h3c046aab),
	.w6(32'h3798fb29),
	.w7(32'h38c4d6f1),
	.w8(32'h3c3e22e4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6e174),
	.w1(32'h3bd4998a),
	.w2(32'hbb59ca27),
	.w3(32'h3b6652d1),
	.w4(32'h3b7ff8f6),
	.w5(32'hba1428ac),
	.w6(32'h3bdaff7c),
	.w7(32'h3b9ee2b6),
	.w8(32'h3b10374c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af24bb7),
	.w1(32'h3b97d9ae),
	.w2(32'hbbed5827),
	.w3(32'hba6e2495),
	.w4(32'h3a7a99e4),
	.w5(32'hbc1ee349),
	.w6(32'h394eceab),
	.w7(32'hbb866e13),
	.w8(32'hbb630340),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d5c63),
	.w1(32'hbb65439a),
	.w2(32'h3c13f300),
	.w3(32'hbc9030df),
	.w4(32'hbc670612),
	.w5(32'h3ae5ca4c),
	.w6(32'hbc237fac),
	.w7(32'hbbae6dc1),
	.w8(32'h3aae9af2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50e60),
	.w1(32'h3b895a02),
	.w2(32'hbcbb2db5),
	.w3(32'h3a212036),
	.w4(32'hba763bda),
	.w5(32'hbc9fa101),
	.w6(32'hbb85f4d7),
	.w7(32'hbc23b21f),
	.w8(32'hbb7849f9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9af9e4),
	.w1(32'h3ac70c7b),
	.w2(32'hbc6c50a6),
	.w3(32'hbce79e2b),
	.w4(32'hbc95b9c9),
	.w5(32'hbc829995),
	.w6(32'hbcccb3bd),
	.w7(32'hbccdb86e),
	.w8(32'hbb901f3f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f87a3),
	.w1(32'hbbd039ed),
	.w2(32'h3a820de3),
	.w3(32'hbcc09b7d),
	.w4(32'hbc7757c6),
	.w5(32'hba1ac9ca),
	.w6(32'hbc910829),
	.w7(32'hbca0b1ca),
	.w8(32'h3c02c83b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d529),
	.w1(32'hba6d9bd9),
	.w2(32'hba80674e),
	.w3(32'hbbd3a5db),
	.w4(32'hb9ae7140),
	.w5(32'h3ae81927),
	.w6(32'hbb131e5e),
	.w7(32'h3a3fc959),
	.w8(32'h3ba62240),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d70de0),
	.w1(32'h3b42c410),
	.w2(32'hbbd7bf7d),
	.w3(32'h3b216a81),
	.w4(32'h3b65af01),
	.w5(32'hbc32ed05),
	.w6(32'h3b9b83a0),
	.w7(32'h3b82d1b9),
	.w8(32'hbc1e3ffd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc395ae8),
	.w1(32'hbb9e12ae),
	.w2(32'hbc78c9bd),
	.w3(32'hbc7a189c),
	.w4(32'hbc98436c),
	.w5(32'hbb5acf17),
	.w6(32'hbc54365e),
	.w7(32'hbbddadb3),
	.w8(32'h3b85ea26),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb580596),
	.w1(32'hbb35a278),
	.w2(32'h3b076511),
	.w3(32'hbb8f19e0),
	.w4(32'hba33c15f),
	.w5(32'h3bcbf8db),
	.w6(32'h3b3825e3),
	.w7(32'h3b1a11df),
	.w8(32'h3b488f47),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad57b4d),
	.w1(32'hbb3ad59a),
	.w2(32'h3aabcac7),
	.w3(32'h3b78aca5),
	.w4(32'hbb04170a),
	.w5(32'h3b15812c),
	.w6(32'h3c0ee961),
	.w7(32'h3b91a847),
	.w8(32'hbbe8b81d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb4e23),
	.w1(32'hbb8d4c12),
	.w2(32'hbb476dc7),
	.w3(32'h3c224043),
	.w4(32'h3b542b97),
	.w5(32'hbb3e1353),
	.w6(32'h39d938ac),
	.w7(32'hb9adcbd8),
	.w8(32'hbbd4f6a2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c188a),
	.w1(32'hbb2d2470),
	.w2(32'h396e9227),
	.w3(32'hbb09b8fc),
	.w4(32'hb9dd1c78),
	.w5(32'h3a10fb85),
	.w6(32'hbac88301),
	.w7(32'h3a6a7bee),
	.w8(32'h3b1a43d6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71d1e0),
	.w1(32'h3b1a7ec8),
	.w2(32'h3b926f55),
	.w3(32'h3b35979f),
	.w4(32'h3bc0fdb2),
	.w5(32'h3b9d9d2d),
	.w6(32'h3b04ec1d),
	.w7(32'h3b393a41),
	.w8(32'h39804444),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd171b),
	.w1(32'hbc066e8d),
	.w2(32'hbba4a281),
	.w3(32'h3c013629),
	.w4(32'h3bb977b6),
	.w5(32'hbaa2861b),
	.w6(32'h3a9fd9e1),
	.w7(32'h3bc72ae1),
	.w8(32'h3c375a93),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd62f08),
	.w1(32'hbc2c4a3c),
	.w2(32'h3a0d9ac0),
	.w3(32'hbc2082fc),
	.w4(32'hbc429a27),
	.w5(32'h391c3cfd),
	.w6(32'hba8ccfcc),
	.w7(32'hbab3e686),
	.w8(32'hbac2ca8f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91474f),
	.w1(32'h393e9d91),
	.w2(32'h3c14d934),
	.w3(32'hbb9d8bfc),
	.w4(32'hbbcb3655),
	.w5(32'h398562a9),
	.w6(32'hbc1c97b6),
	.w7(32'hbb8b4486),
	.w8(32'hbb9730b2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24ce97),
	.w1(32'h38b30f33),
	.w2(32'hbcb42d1e),
	.w3(32'hbaddeebd),
	.w4(32'hba925c6c),
	.w5(32'hbd327760),
	.w6(32'hbc0ed758),
	.w7(32'hbc584c2c),
	.w8(32'hbc9f0fdd),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfb0af),
	.w1(32'hbc61a046),
	.w2(32'h3b789ea3),
	.w3(32'hbd7d2c1b),
	.w4(32'hbd37ca24),
	.w5(32'h3be06a89),
	.w6(32'hbd185198),
	.w7(32'hbd18b182),
	.w8(32'hbb6503e1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e826),
	.w1(32'h393840ef),
	.w2(32'hbc981a4e),
	.w3(32'h3acddd2c),
	.w4(32'h3afa58e0),
	.w5(32'hbca5a14f),
	.w6(32'hbbaab555),
	.w7(32'hbb10d6cd),
	.w8(32'hbadfd181),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb01365),
	.w1(32'hbb849c3a),
	.w2(32'hbcd44ee7),
	.w3(32'hbcf63126),
	.w4(32'hbcb7eea6),
	.w5(32'hbcd2f636),
	.w6(32'hbbae121a),
	.w7(32'hbc6825da),
	.w8(32'hbc23d009),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca930f1),
	.w1(32'hbac0c7e3),
	.w2(32'hbc4d19ee),
	.w3(32'hbd3ae959),
	.w4(32'hbca13528),
	.w5(32'hbbc1a7f9),
	.w6(32'hbccf7da6),
	.w7(32'hbd09d988),
	.w8(32'h3b63c6d7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddfb9c),
	.w1(32'h3b71d6d0),
	.w2(32'hbbc0b8eb),
	.w3(32'hbc0f7d31),
	.w4(32'hbbd95f38),
	.w5(32'hbbfc981e),
	.w6(32'hbbffc61b),
	.w7(32'hbb6997dd),
	.w8(32'h3bc5e9b5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba724cb),
	.w1(32'h3b804710),
	.w2(32'hbc988e70),
	.w3(32'hbc995667),
	.w4(32'hbc283bce),
	.w5(32'hbcbdc608),
	.w6(32'hbc0de2d5),
	.w7(32'hbbd29e3e),
	.w8(32'hbc53580a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd7e38),
	.w1(32'hbb8c5e15),
	.w2(32'hbb3b6d82),
	.w3(32'hbd32b839),
	.w4(32'hbce830b4),
	.w5(32'hbbc1b201),
	.w6(32'hbd1a2253),
	.w7(32'hbd101bbb),
	.w8(32'h3bdb6107),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94385a),
	.w1(32'h3b92a4be),
	.w2(32'h3a934776),
	.w3(32'hbc1ce129),
	.w4(32'hbb6831c7),
	.w5(32'hbad56b24),
	.w6(32'hbbf18ea7),
	.w7(32'hb9aa319f),
	.w8(32'h3be9f098),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a94be),
	.w1(32'h3bb229e7),
	.w2(32'h3a8dcf70),
	.w3(32'hbb19c431),
	.w4(32'h3b19a899),
	.w5(32'h3c0eaada),
	.w6(32'hbb6ecd7f),
	.w7(32'h3be659b8),
	.w8(32'hbc040eff),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa309),
	.w1(32'hbba92dba),
	.w2(32'hbc6bdad6),
	.w3(32'h3c5fc1a7),
	.w4(32'h3c1b1bc9),
	.w5(32'hbc73332d),
	.w6(32'h3b3ea39c),
	.w7(32'h3ba2e1fa),
	.w8(32'hbb3fc33b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe36c30),
	.w1(32'h3a03f78b),
	.w2(32'hb9f37d12),
	.w3(32'hbc8322c0),
	.w4(32'hbc06df86),
	.w5(32'h3c103624),
	.w6(32'hbc1a9e1e),
	.w7(32'hbc018d69),
	.w8(32'h3a8b3f52),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97c0e8),
	.w1(32'hbbf4afd3),
	.w2(32'h3cb60002),
	.w3(32'h3ae4082b),
	.w4(32'h3b48ff7d),
	.w5(32'h3c9e4743),
	.w6(32'h39e8fd55),
	.w7(32'h3b8e6af5),
	.w8(32'h3c151e1c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00fe52),
	.w1(32'h3c8903a4),
	.w2(32'hbbeda7e9),
	.w3(32'h3cf23a72),
	.w4(32'h3ce8896f),
	.w5(32'hbc772c39),
	.w6(32'h3c5fd23e),
	.w7(32'h3c77964e),
	.w8(32'h3ad91506),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4edd42),
	.w1(32'hbaf4c4ed),
	.w2(32'hbba39424),
	.w3(32'hbce2838b),
	.w4(32'hbcbd4c75),
	.w5(32'hbc2d5389),
	.w6(32'hbcbc9c38),
	.w7(32'hbcd8b3c8),
	.w8(32'hbc4d1a5d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa19c0),
	.w1(32'hbbc4e4f9),
	.w2(32'h3ca1e322),
	.w3(32'hbc3efccd),
	.w4(32'hbc316da1),
	.w5(32'h3d10d442),
	.w6(32'hbc35f79e),
	.w7(32'hbc51d20d),
	.w8(32'h3c814b46),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca25d22),
	.w1(32'h3c63ffbd),
	.w2(32'hb9fa81bf),
	.w3(32'h3d4660ee),
	.w4(32'h3d2182b0),
	.w5(32'hbbafa093),
	.w6(32'h3d15b0f0),
	.w7(32'h3d2f6cde),
	.w8(32'h3b0bb852),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa33906),
	.w1(32'h3aad1550),
	.w2(32'h3b9be05d),
	.w3(32'hbc3bbbed),
	.w4(32'hbbc3505a),
	.w5(32'h3b191f85),
	.w6(32'hbbcf2687),
	.w7(32'hbba828e3),
	.w8(32'hbbf2aa18),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be503a6),
	.w1(32'h3be3d052),
	.w2(32'hbbbfa327),
	.w3(32'h3bf8d94e),
	.w4(32'h3c0f02bb),
	.w5(32'h3b85fb17),
	.w6(32'hb9e37f52),
	.w7(32'h3ac68934),
	.w8(32'h3bab1560),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16856e),
	.w1(32'hbb8e7810),
	.w2(32'hbb731b97),
	.w3(32'h3b8bb674),
	.w4(32'hbb5d807e),
	.w5(32'hbb1dfb73),
	.w6(32'h3c123066),
	.w7(32'h3c1161c0),
	.w8(32'h3b6347ed),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef31b),
	.w1(32'h3a8a480d),
	.w2(32'hbceac5b9),
	.w3(32'hb99804fa),
	.w4(32'h3ab51500),
	.w5(32'hbce1e566),
	.w6(32'h3b3d6ee5),
	.w7(32'h3baf97c8),
	.w8(32'hbbe6b69d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba83e5),
	.w1(32'hbcb7bb74),
	.w2(32'hbc94a744),
	.w3(32'hbd28d238),
	.w4(32'hbd1eb4dc),
	.w5(32'hbcf10355),
	.w6(32'hbcc6002f),
	.w7(32'hbceff813),
	.w8(32'hbc22c38c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e70da),
	.w1(32'hbb4e1277),
	.w2(32'hbbd0095b),
	.w3(32'hbd3acd42),
	.w4(32'hbcf269ea),
	.w5(32'hbc40d9e6),
	.w6(32'hbcf78745),
	.w7(32'hbcc1db36),
	.w8(32'hbc7ec422),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf086b),
	.w1(32'hbc3a7e7d),
	.w2(32'h3ae2fe0c),
	.w3(32'hbc8a4bfe),
	.w4(32'hbc3007a4),
	.w5(32'h3a9dbd9d),
	.w6(32'hbc951ef5),
	.w7(32'hbccee687),
	.w8(32'h3ba49891),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d8de9),
	.w1(32'h3b04943c),
	.w2(32'hba7f277d),
	.w3(32'h39ae1775),
	.w4(32'hba85bee5),
	.w5(32'h3ac1beec),
	.w6(32'h3b3be983),
	.w7(32'h3b4e655c),
	.w8(32'h3b58850c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bfba3),
	.w1(32'h3b18b3d9),
	.w2(32'hb9ef8d5e),
	.w3(32'h38a8a4dd),
	.w4(32'h3a84679b),
	.w5(32'h3b700728),
	.w6(32'h3b871ce3),
	.w7(32'h3acf86c0),
	.w8(32'h3be3f458),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2eebb),
	.w1(32'hbb655e9c),
	.w2(32'h39f1ea61),
	.w3(32'hbc170b4c),
	.w4(32'hbc3f7528),
	.w5(32'hba2955a6),
	.w6(32'hbb366a63),
	.w7(32'hbc1552a6),
	.w8(32'h3b8a1a6a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880a428),
	.w1(32'h3b86f0b7),
	.w2(32'hbcd18ef3),
	.w3(32'hbb0d99fc),
	.w4(32'h3b8258f1),
	.w5(32'hbce5433a),
	.w6(32'h3a13ac81),
	.w7(32'h3b850f5d),
	.w8(32'hbc24c16a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfabb8c),
	.w1(32'hbc824f17),
	.w2(32'hbc8deea6),
	.w3(32'hbd4c23e4),
	.w4(32'hbd16b393),
	.w5(32'hbc0385fa),
	.w6(32'hbd19b302),
	.w7(32'hbd080997),
	.w8(32'hbabbd900),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93cd7e),
	.w1(32'h39cad9de),
	.w2(32'hbc10900e),
	.w3(32'hbccd1cf5),
	.w4(32'hbc71fb82),
	.w5(32'h3a05bf08),
	.w6(32'hbc3afd8d),
	.w7(32'hbcb86579),
	.w8(32'h3c1f0078),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a3d4),
	.w1(32'h3c491860),
	.w2(32'h3bd31ca6),
	.w3(32'h3aa06776),
	.w4(32'h3bf4452c),
	.w5(32'h3a0efa4a),
	.w6(32'h3c076370),
	.w7(32'h3a6d00cc),
	.w8(32'h3c5ea1b5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule