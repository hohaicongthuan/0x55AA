module layer_10_featuremap_488(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e1683),
	.w1(32'h3aca4026),
	.w2(32'h3acc16f4),
	.w3(32'h3a095adb),
	.w4(32'h3a954ce0),
	.w5(32'hb9a794b4),
	.w6(32'h3abc9576),
	.w7(32'h3ab2da7b),
	.w8(32'h39d7716d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf9252),
	.w1(32'hbae2966f),
	.w2(32'hbb0bcd4b),
	.w3(32'hba2b69b8),
	.w4(32'hbaa110dc),
	.w5(32'hbab55c40),
	.w6(32'h3991296d),
	.w7(32'hbab4be65),
	.w8(32'hbb24af82),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba3a7d),
	.w1(32'hba282278),
	.w2(32'h398440f4),
	.w3(32'hba0aa6f8),
	.w4(32'hbb4c2d00),
	.w5(32'hbb126e5f),
	.w6(32'hbb053afd),
	.w7(32'hbb66d6f4),
	.w8(32'hbb469a21),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddb636),
	.w1(32'hbb283be2),
	.w2(32'h3a38b407),
	.w3(32'h3b182093),
	.w4(32'hbab8ff92),
	.w5(32'h3b31318e),
	.w6(32'h378ddb05),
	.w7(32'hbaec633d),
	.w8(32'hb8e47937),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce6d2),
	.w1(32'h3ac1360a),
	.w2(32'h3a7de978),
	.w3(32'hba52ca0a),
	.w4(32'h384ee56b),
	.w5(32'hb9956bdc),
	.w6(32'hbaba6a7d),
	.w7(32'hb9f091ff),
	.w8(32'hba25c43a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac693e6),
	.w1(32'hba2b50c9),
	.w2(32'hbb191a3a),
	.w3(32'h3aa02119),
	.w4(32'hbaf5d4b1),
	.w5(32'hbb3452fb),
	.w6(32'h3a9a0fd1),
	.w7(32'hba5d487c),
	.w8(32'hb9ef5326),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a803a),
	.w1(32'h3a718138),
	.w2(32'h3ab81754),
	.w3(32'hb97ef336),
	.w4(32'h3a0e33c3),
	.w5(32'h3aae50c2),
	.w6(32'h3ab8b212),
	.w7(32'h3a302f0c),
	.w8(32'hb9e20959),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06ca5b),
	.w1(32'h3a889da9),
	.w2(32'h3b0eebcb),
	.w3(32'h3a8647f1),
	.w4(32'hba26d369),
	.w5(32'h3b07df00),
	.w6(32'h395c856e),
	.w7(32'hbba3bcf1),
	.w8(32'hba89eebc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec29c),
	.w1(32'hbb003d9f),
	.w2(32'hba6a0d37),
	.w3(32'h3aae893c),
	.w4(32'h396c5ac2),
	.w5(32'h3903ebef),
	.w6(32'hb9f12861),
	.w7(32'hb9fabd70),
	.w8(32'hbae79633),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01a64e),
	.w1(32'hba5a0dd5),
	.w2(32'hb890c7e2),
	.w3(32'hbb2122df),
	.w4(32'hbadd5130),
	.w5(32'h38fcbcc4),
	.w6(32'hbb186a7f),
	.w7(32'h39974ee0),
	.w8(32'h3a27d6da),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d13ebf),
	.w1(32'hbaed190f),
	.w2(32'hbac11347),
	.w3(32'hbab67f2d),
	.w4(32'hbab00c6c),
	.w5(32'hbb3088a2),
	.w6(32'hba260a4a),
	.w7(32'h3a09ccc0),
	.w8(32'hbaeaf19d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad6f0),
	.w1(32'h3ac953cd),
	.w2(32'h3ac36a27),
	.w3(32'hba3f2383),
	.w4(32'h3ad02ac6),
	.w5(32'h3b48cd31),
	.w6(32'hbb017700),
	.w7(32'h3a98ea0d),
	.w8(32'h3af997ee),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd00fe),
	.w1(32'hbb0698d6),
	.w2(32'hba9fddaf),
	.w3(32'h3a39fa9f),
	.w4(32'hbaca0056),
	.w5(32'h3a4203d0),
	.w6(32'h3b30f747),
	.w7(32'hbb211c13),
	.w8(32'hbb08886e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125190),
	.w1(32'hba2c784c),
	.w2(32'hba6f84bb),
	.w3(32'hba0786a2),
	.w4(32'hbb45b39d),
	.w5(32'hbbab07c7),
	.w6(32'h39c32422),
	.w7(32'hbafc4f94),
	.w8(32'hbb319081),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57a51a),
	.w1(32'hba14548a),
	.w2(32'hba6368e5),
	.w3(32'hbaa29df9),
	.w4(32'hbb211699),
	.w5(32'hbaf389a1),
	.w6(32'hba74c9b7),
	.w7(32'hbb4b5e4f),
	.w8(32'hbaffae5e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba218748),
	.w1(32'h3a16fc09),
	.w2(32'h3a4753ce),
	.w3(32'hbaabb58c),
	.w4(32'hba9000eb),
	.w5(32'h3adfe915),
	.w6(32'h3945c4c8),
	.w7(32'hbb1bdbb4),
	.w8(32'h3a149123),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69b7a1),
	.w1(32'hb9bf8b3a),
	.w2(32'hb9aabaf0),
	.w3(32'hba973459),
	.w4(32'hb4b3f14c),
	.w5(32'h3ae1f5dd),
	.w6(32'h39c40f7f),
	.w7(32'hba8696a6),
	.w8(32'hb9b3347c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0220ae),
	.w1(32'h3951a1f3),
	.w2(32'hb581174e),
	.w3(32'h3ab8e405),
	.w4(32'h38da8dff),
	.w5(32'hba0f73dd),
	.w6(32'h39c3d56f),
	.w7(32'hb8833676),
	.w8(32'hb9610ad7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab958f2),
	.w1(32'hbb1679d9),
	.w2(32'hba4fb120),
	.w3(32'hba5958c5),
	.w4(32'hbb372b20),
	.w5(32'h3995feba),
	.w6(32'h38f7723e),
	.w7(32'hbaa98691),
	.w8(32'hb846cf30),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f97ac1),
	.w1(32'hbb7551dc),
	.w2(32'hbb762f48),
	.w3(32'h3a0a7c76),
	.w4(32'hbb2de1f1),
	.w5(32'hbb4bbf06),
	.w6(32'h3b051016),
	.w7(32'hbaeb3e2a),
	.w8(32'hbb15be7a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aa922),
	.w1(32'hb9b74c86),
	.w2(32'h39e3ad44),
	.w3(32'hbbc40844),
	.w4(32'h3a416a95),
	.w5(32'h3aeb3dc7),
	.w6(32'hbb52fd7d),
	.w7(32'hb8c74137),
	.w8(32'h3acecf01),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5dd46),
	.w1(32'h3a6362e7),
	.w2(32'hbb00ce99),
	.w3(32'h3b527bef),
	.w4(32'hba375f0b),
	.w5(32'hb98f89a3),
	.w6(32'h3b84dbd6),
	.w7(32'hbb43f086),
	.w8(32'hbaef55e6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079313),
	.w1(32'h37d8bfa2),
	.w2(32'h3ad732a4),
	.w3(32'hbb17619e),
	.w4(32'hb896520d),
	.w5(32'h3a19bbeb),
	.w6(32'hba973e38),
	.w7(32'h3a343363),
	.w8(32'h3ac6385c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeb497),
	.w1(32'hbaacf421),
	.w2(32'hbac2cc80),
	.w3(32'hb8fd3fb0),
	.w4(32'hbb86ec95),
	.w5(32'hbb6c2af7),
	.w6(32'h3a9593c4),
	.w7(32'hbaba2e83),
	.w8(32'hbaf9d68e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af661),
	.w1(32'hbafe92c5),
	.w2(32'h3a7de55c),
	.w3(32'hbb301117),
	.w4(32'hbaf1d975),
	.w5(32'h39ab2c50),
	.w6(32'hba3a4eba),
	.w7(32'h3a458278),
	.w8(32'h3ad4d2d0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0627ca),
	.w1(32'hba944892),
	.w2(32'hbb69b28a),
	.w3(32'h39e8a4f7),
	.w4(32'h3a8860c8),
	.w5(32'hb98f358c),
	.w6(32'hba2834e4),
	.w7(32'h3adffcd3),
	.w8(32'h3ba094a0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e550c),
	.w1(32'hb8a769f5),
	.w2(32'h3a991d33),
	.w3(32'hbae093ff),
	.w4(32'h39c74ffc),
	.w5(32'h3ad5885e),
	.w6(32'h3b14ec8d),
	.w7(32'hba56be73),
	.w8(32'h39e6c5e2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19dc32),
	.w1(32'h3958d35d),
	.w2(32'h3a29db2f),
	.w3(32'h3a028de5),
	.w4(32'hb928f133),
	.w5(32'h3a27cc08),
	.w6(32'h39c9c814),
	.w7(32'h39c92004),
	.w8(32'h3a3ba4b2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc0e54),
	.w1(32'h3a76e229),
	.w2(32'h38a79547),
	.w3(32'h3924011d),
	.w4(32'hba5ddbe7),
	.w5(32'h393551e4),
	.w6(32'h3a69bc6a),
	.w7(32'hba46f6c4),
	.w8(32'hba9d8f8d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1f78d),
	.w1(32'h3970d9ae),
	.w2(32'h39a78d2d),
	.w3(32'hb96ab437),
	.w4(32'h3a59a1cc),
	.w5(32'h390927ec),
	.w6(32'h38ce3792),
	.w7(32'h3a9578a0),
	.w8(32'h3ac5640e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fdf1c),
	.w1(32'h398bd544),
	.w2(32'hba8bc5f1),
	.w3(32'h3b14dc06),
	.w4(32'h3ad98ff1),
	.w5(32'h392fae27),
	.w6(32'h3b7d99b7),
	.w7(32'hb9bbaee9),
	.w8(32'hba4a0a2f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ac4f1),
	.w1(32'hbb1ff6b9),
	.w2(32'hb915599d),
	.w3(32'h399ec0d9),
	.w4(32'hbb6c3b59),
	.w5(32'hba9ee27c),
	.w6(32'hb9bd41de),
	.w7(32'hbb1ea1e7),
	.w8(32'hbadb23a3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24bc4f),
	.w1(32'hba496df6),
	.w2(32'hbab0b950),
	.w3(32'h3a95b83a),
	.w4(32'hb90ae791),
	.w5(32'hb986e39f),
	.w6(32'h39979f95),
	.w7(32'h3a2f23bd),
	.w8(32'hbabb72fe),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20319a),
	.w1(32'h39964022),
	.w2(32'h3a9f2e16),
	.w3(32'hbabef851),
	.w4(32'h391da06b),
	.w5(32'h3aa1a7c9),
	.w6(32'hb92d58c1),
	.w7(32'h3a59a524),
	.w8(32'h39c91632),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c243b),
	.w1(32'h3b54e4ec),
	.w2(32'h3b486d3e),
	.w3(32'hba181c38),
	.w4(32'hb95c0030),
	.w5(32'h3a101f2c),
	.w6(32'h3a3402af),
	.w7(32'hbb62747f),
	.w8(32'hb9b9213c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b232797),
	.w1(32'hb9f845ee),
	.w2(32'h3a3b6a86),
	.w3(32'hbaad30fa),
	.w4(32'hb9885d78),
	.w5(32'h3a920d08),
	.w6(32'hb99b98c2),
	.w7(32'hba60b8a9),
	.w8(32'hba8c8ea0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390db09f),
	.w1(32'hb9a71ff6),
	.w2(32'hbae9719e),
	.w3(32'hba5ebb7a),
	.w4(32'h3b246380),
	.w5(32'hba982a36),
	.w6(32'hbac1bb3b),
	.w7(32'h3ba3d237),
	.w8(32'hb94f6377),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47b278),
	.w1(32'h3a0ec54a),
	.w2(32'h39f2f380),
	.w3(32'h3984e2e4),
	.w4(32'hba99d606),
	.w5(32'hbae5bc88),
	.w6(32'hba3a528c),
	.w7(32'h3a11b53d),
	.w8(32'hbacaa80d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6ca3),
	.w1(32'h3af20acc),
	.w2(32'hba4ec9b9),
	.w3(32'h39a8056b),
	.w4(32'hb882c1b9),
	.w5(32'hbb7fe13d),
	.w6(32'hba3f41ed),
	.w7(32'h3a06f45f),
	.w8(32'hbaeade67),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93ff27),
	.w1(32'hba1e2c0e),
	.w2(32'h3a3ffcb4),
	.w3(32'hbb4c8012),
	.w4(32'hb9543c5c),
	.w5(32'h3aa61a60),
	.w6(32'hbb275e6e),
	.w7(32'h3a98ebc2),
	.w8(32'h3afdc436),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388bba70),
	.w1(32'hbb38f78d),
	.w2(32'hbb29aaca),
	.w3(32'h39495558),
	.w4(32'hbb708d91),
	.w5(32'hbae03710),
	.w6(32'hba358692),
	.w7(32'hba866fd9),
	.w8(32'hba818095),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc671d),
	.w1(32'hbac2be7a),
	.w2(32'hbada3994),
	.w3(32'hbb391d7c),
	.w4(32'hbaa44035),
	.w5(32'h393e27c1),
	.w6(32'hba8ec3d2),
	.w7(32'hbb061c2f),
	.w8(32'hbac68da2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9affbd7),
	.w1(32'hbb759878),
	.w2(32'hbade38a5),
	.w3(32'hba91280f),
	.w4(32'hbb276b43),
	.w5(32'h3a45f30f),
	.w6(32'hba31497d),
	.w7(32'hbabb4f61),
	.w8(32'hbadacdc3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95b322),
	.w1(32'h3a83b0b9),
	.w2(32'h3a8cc179),
	.w3(32'hbb30fdba),
	.w4(32'h3a48b7ea),
	.w5(32'h3a3852ca),
	.w6(32'hba37590e),
	.w7(32'h3aefc968),
	.w8(32'h3a8a044d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cad91),
	.w1(32'h3a55ef9d),
	.w2(32'h3a5e6290),
	.w3(32'h3ad424fe),
	.w4(32'h3acf2490),
	.w5(32'h3b430750),
	.w6(32'h3a843e05),
	.w7(32'h3a97e9b9),
	.w8(32'h3acaacff),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9e0c),
	.w1(32'hb928af7c),
	.w2(32'hbaaad61d),
	.w3(32'hb9004ffa),
	.w4(32'hb9f29fea),
	.w5(32'hbabdca2b),
	.w6(32'h3a2eae2a),
	.w7(32'hbb367dc9),
	.w8(32'hbb0557aa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2b9f6),
	.w1(32'h3a1d7bd5),
	.w2(32'hba97cade),
	.w3(32'hbb6aa3cc),
	.w4(32'h3a798157),
	.w5(32'h3a8a8c18),
	.w6(32'hbb11950d),
	.w7(32'hb947689a),
	.w8(32'h39aae27d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f8186),
	.w1(32'hba2778d7),
	.w2(32'hba99ea9d),
	.w3(32'hba0dd438),
	.w4(32'h3905aecf),
	.w5(32'hbab71615),
	.w6(32'h38523ecc),
	.w7(32'hba5ac57c),
	.w8(32'hbb0b2078),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba967c2a),
	.w1(32'h3a73ad16),
	.w2(32'h38bd0da6),
	.w3(32'hbb2b4f85),
	.w4(32'h3a9a395a),
	.w5(32'h3a96dd03),
	.w6(32'hbb2c0c8e),
	.w7(32'h390c6ef1),
	.w8(32'h3abf406b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a4825),
	.w1(32'hba23e52a),
	.w2(32'h3a87398d),
	.w3(32'h390d5694),
	.w4(32'hba03ce74),
	.w5(32'h3b0e216c),
	.w6(32'hb9e38de3),
	.w7(32'hba9a9b7e),
	.w8(32'h3b257f1d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b8ef1),
	.w1(32'h3acdccaa),
	.w2(32'h3aa7e3ba),
	.w3(32'h3aad267e),
	.w4(32'hb8883a01),
	.w5(32'hb95640eb),
	.w6(32'h3af0eeea),
	.w7(32'hba7ca4c1),
	.w8(32'hba7f5ed8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c6f9),
	.w1(32'hbad7c774),
	.w2(32'hbb051965),
	.w3(32'h3a6c56ea),
	.w4(32'hbace2409),
	.w5(32'hbb1821fc),
	.w6(32'h3aa9fe7e),
	.w7(32'hbaa2a13d),
	.w8(32'hbb0643ba),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ccce7),
	.w1(32'hb8f3561c),
	.w2(32'hb91bf9fe),
	.w3(32'hbb545bed),
	.w4(32'h39163a74),
	.w5(32'h3a19c517),
	.w6(32'hbb85f284),
	.w7(32'h395544bc),
	.w8(32'h3a867bb4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f2530),
	.w1(32'h3b25e73f),
	.w2(32'h3b447295),
	.w3(32'h3990c408),
	.w4(32'h3a15c50a),
	.w5(32'h3a8ad08f),
	.w6(32'h3ab08602),
	.w7(32'h3a4cb4a3),
	.w8(32'h3a94e48a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa2fb9),
	.w1(32'hba874dd5),
	.w2(32'hbabfac1b),
	.w3(32'h3b26725d),
	.w4(32'hbb34b7f1),
	.w5(32'h3a40294a),
	.w6(32'h3a881cd6),
	.w7(32'hbb23b04b),
	.w8(32'hba405513),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e302),
	.w1(32'hbb10aeca),
	.w2(32'hbace517c),
	.w3(32'hbaca54b9),
	.w4(32'hbb5db0e6),
	.w5(32'hbb153ebb),
	.w6(32'hbb5e56db),
	.w7(32'h3a89bbca),
	.w8(32'hba9b95dc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49976e),
	.w1(32'h3a78ce8c),
	.w2(32'h3acc6683),
	.w3(32'h393433e3),
	.w4(32'h39e89049),
	.w5(32'hba717c9b),
	.w6(32'hba2f3e8f),
	.w7(32'h3a92c3f6),
	.w8(32'h3ab67461),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf857),
	.w1(32'hbb5872fc),
	.w2(32'hbbbd1da2),
	.w3(32'h3b183d65),
	.w4(32'hbb3d6cc5),
	.w5(32'hbbb4be23),
	.w6(32'h3b51f303),
	.w7(32'hbac5f945),
	.w8(32'hbbaf1543),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb689176),
	.w1(32'hb93c0097),
	.w2(32'hba5bad2e),
	.w3(32'hbb966a40),
	.w4(32'hba0df25a),
	.w5(32'h39037511),
	.w6(32'hbb5ccd7b),
	.w7(32'hbadf76b6),
	.w8(32'hb9db5d41),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7ef66),
	.w1(32'hbb7922c6),
	.w2(32'hba86abc9),
	.w3(32'hbab312e3),
	.w4(32'hba614e81),
	.w5(32'hbaf0df92),
	.w6(32'hb99c2b94),
	.w7(32'hba6b8486),
	.w8(32'h3a8f3a59),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8811f1),
	.w1(32'h3a8e260b),
	.w2(32'hba415c15),
	.w3(32'hba2dc8b8),
	.w4(32'h39b1f311),
	.w5(32'h39bc59a0),
	.w6(32'hb8b3e600),
	.w7(32'hba8c8cb2),
	.w8(32'h3aedc827),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab32a40),
	.w1(32'hb885f91c),
	.w2(32'hba442fd4),
	.w3(32'hba8c7e8c),
	.w4(32'hb94c4c20),
	.w5(32'hbad9a4c9),
	.w6(32'h38efc178),
	.w7(32'hba0fc962),
	.w8(32'hbaa2348c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb781bdd4),
	.w1(32'hbb36c461),
	.w2(32'hb99f1735),
	.w3(32'hb93c4128),
	.w4(32'hbaddf370),
	.w5(32'h39848d24),
	.w6(32'hb97a267b),
	.w7(32'hba9f3b50),
	.w8(32'hba9ab32c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9a1c0),
	.w1(32'h3a96c326),
	.w2(32'h3a008810),
	.w3(32'hbb3107c9),
	.w4(32'h3a23df7c),
	.w5(32'h3a41a8da),
	.w6(32'hbb013b94),
	.w7(32'h3ab3ece3),
	.w8(32'h3b06c579),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895bb6a),
	.w1(32'h3b06d4be),
	.w2(32'h3b41309e),
	.w3(32'h3a202c1f),
	.w4(32'h3aa11c3e),
	.w5(32'h3af2d6a8),
	.w6(32'h3b332ca4),
	.w7(32'h3b36aa2a),
	.w8(32'h3b98dec9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a3ae9),
	.w1(32'h3a9cb580),
	.w2(32'hb9d16ff0),
	.w3(32'h3b60c79b),
	.w4(32'h3a8554e3),
	.w5(32'h3a645c1f),
	.w6(32'h3b9e2fef),
	.w7(32'h3a7f9794),
	.w8(32'h3b0b5e72),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f1f28),
	.w1(32'hba81d74a),
	.w2(32'hbaeae7dc),
	.w3(32'hb7cf9904),
	.w4(32'hb9e473f1),
	.w5(32'h397e5d05),
	.w6(32'h3a87a860),
	.w7(32'hbb0cfe2a),
	.w8(32'hba76fc94),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad88ecf),
	.w1(32'hbb2963b0),
	.w2(32'hbb6f9cff),
	.w3(32'hbadc50ba),
	.w4(32'hbb0b1ed9),
	.w5(32'hbb158268),
	.w6(32'hbb280b44),
	.w7(32'hbb7e9f21),
	.w8(32'hbb5fdf8f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0072ac),
	.w1(32'h3b136138),
	.w2(32'h3a2793f1),
	.w3(32'hbacb87a7),
	.w4(32'h3b06c99d),
	.w5(32'h3ab6ecdb),
	.w6(32'hbb0a8b11),
	.w7(32'h39209c1b),
	.w8(32'hbad9ffc9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371651af),
	.w1(32'hbaaa2e2c),
	.w2(32'hba8d7a59),
	.w3(32'hbb1a7dc8),
	.w4(32'hbb09e761),
	.w5(32'hbbb17921),
	.w6(32'hbb3a148a),
	.w7(32'h3a803735),
	.w8(32'hbb326a63),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd7c5),
	.w1(32'hbac377a2),
	.w2(32'hbbc6c707),
	.w3(32'hbab47de8),
	.w4(32'hbb848d87),
	.w5(32'h3a231659),
	.w6(32'h37fca4b2),
	.w7(32'h3b03ca16),
	.w8(32'h39bb9410),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf807e),
	.w1(32'h3a3e8a77),
	.w2(32'hb99bfb93),
	.w3(32'h3a5de96b),
	.w4(32'h3b33140e),
	.w5(32'h3bfe00c3),
	.w6(32'h3b1ea969),
	.w7(32'hbaf11800),
	.w8(32'hbb0c827c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e70bc0),
	.w1(32'hbb837bc9),
	.w2(32'hbba0933e),
	.w3(32'hba5013d2),
	.w4(32'hbb05d343),
	.w5(32'hbb8c2546),
	.w6(32'h3b5f9778),
	.w7(32'hbb27c9b9),
	.w8(32'hbb473ab9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89f28d),
	.w1(32'hbb569c91),
	.w2(32'hbb41668f),
	.w3(32'hbb15bd94),
	.w4(32'hbafa42bb),
	.w5(32'hba6930d3),
	.w6(32'h3b0702d8),
	.w7(32'hbb09870b),
	.w8(32'h3aa68144),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47b31a),
	.w1(32'h3909a1d1),
	.w2(32'h3a5ea2fa),
	.w3(32'h3a9ff46d),
	.w4(32'h3b854dc7),
	.w5(32'h3b7267cc),
	.w6(32'h3a9c4b1a),
	.w7(32'h3bce3414),
	.w8(32'h3bbcee96),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08066),
	.w1(32'hbb9e8e43),
	.w2(32'hbb0331b3),
	.w3(32'h3b9bd6c5),
	.w4(32'hbb3c9a4e),
	.w5(32'h3b219c19),
	.w6(32'h3bee769d),
	.w7(32'h3abbea92),
	.w8(32'hb8ff0523),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885dbd),
	.w1(32'hbb45474a),
	.w2(32'h3a17808a),
	.w3(32'h3af65582),
	.w4(32'hbb256ea3),
	.w5(32'hbb0bdecb),
	.w6(32'hb9caf642),
	.w7(32'hbbafcf77),
	.w8(32'hbb82ee71),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f252d),
	.w1(32'h39f3a705),
	.w2(32'h3ab55943),
	.w3(32'hbb802e52),
	.w4(32'h3b4ee904),
	.w5(32'hb96c438a),
	.w6(32'hbb0afdbe),
	.w7(32'hbaf89e8a),
	.w8(32'h3ac34dd1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebc034),
	.w1(32'hba791f4b),
	.w2(32'hbbc8173c),
	.w3(32'hbacdef81),
	.w4(32'hba422266),
	.w5(32'hbb03c60e),
	.w6(32'hbacedaab),
	.w7(32'h390e65b4),
	.w8(32'hbb9b7735),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51d69b),
	.w1(32'h3a3e76cf),
	.w2(32'h3b435734),
	.w3(32'h3a85dc62),
	.w4(32'h3ac676f9),
	.w5(32'hbbd464c3),
	.w6(32'hbb2f086b),
	.w7(32'hbb75cfee),
	.w8(32'hbbd8b8f7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822dcd),
	.w1(32'h3b0d4a14),
	.w2(32'h3b6711ed),
	.w3(32'hbb48dd9b),
	.w4(32'h3bedb511),
	.w5(32'h3ba81001),
	.w6(32'hbb16e042),
	.w7(32'h3b4bbfb0),
	.w8(32'h3a99c911),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac03357),
	.w1(32'h3ad3390d),
	.w2(32'h3ad881be),
	.w3(32'h3acf451d),
	.w4(32'h3bb70b9a),
	.w5(32'h3af8f1be),
	.w6(32'h3a29b712),
	.w7(32'h3aeb6df4),
	.w8(32'h3b6b7f80),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11421f),
	.w1(32'hba87c6ad),
	.w2(32'hbab42404),
	.w3(32'h3a606986),
	.w4(32'hbb2935bc),
	.w5(32'h3b5b1b89),
	.w6(32'h3b51bea3),
	.w7(32'hbad1dffd),
	.w8(32'h399e2f4c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6a970),
	.w1(32'h3b2b8774),
	.w2(32'h395c56df),
	.w3(32'hbabd5b8e),
	.w4(32'h397ae89c),
	.w5(32'hba4980cf),
	.w6(32'h39d7a764),
	.w7(32'h3b6cce72),
	.w8(32'h3c54809f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17dea2),
	.w1(32'h3a742c2a),
	.w2(32'hbaa22077),
	.w3(32'h3bd8a99b),
	.w4(32'h3b9507d1),
	.w5(32'h3acbf00f),
	.w6(32'h3a3e390e),
	.w7(32'h3ae95086),
	.w8(32'h3b2f8a6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65cc02),
	.w1(32'hbb63923d),
	.w2(32'hbc50ec28),
	.w3(32'h3b06165c),
	.w4(32'hba1b704d),
	.w5(32'h3bdc5604),
	.w6(32'h3bb9535b),
	.w7(32'h3af4f62e),
	.w8(32'h3b13bd0f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b766714),
	.w1(32'hbb9b47fa),
	.w2(32'hbbb27a84),
	.w3(32'hbb262a79),
	.w4(32'hbbedb7da),
	.w5(32'hbb892346),
	.w6(32'hbac9c019),
	.w7(32'h3b41a03a),
	.w8(32'h3aac6111),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa248),
	.w1(32'hbb50b3ac),
	.w2(32'hbbad0f56),
	.w3(32'hbb2bdf4f),
	.w4(32'hbb09f010),
	.w5(32'h3bca079f),
	.w6(32'h3ab14d9d),
	.w7(32'h39b658c4),
	.w8(32'h3b1d16f2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a102bb6),
	.w1(32'h3ba3fba7),
	.w2(32'h3ba786b7),
	.w3(32'h3adaf07e),
	.w4(32'hbb09b251),
	.w5(32'hbafc26ea),
	.w6(32'hba37eb4f),
	.w7(32'h3af5d8d6),
	.w8(32'h3a673f5d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb7d7),
	.w1(32'hbbb25029),
	.w2(32'hbabaac91),
	.w3(32'h3bbb0935),
	.w4(32'hb89aad9f),
	.w5(32'h3b915602),
	.w6(32'h3be78d1b),
	.w7(32'hbb8d2f0d),
	.w8(32'h3b2a8aef),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbdf2a),
	.w1(32'hbb8a7f66),
	.w2(32'hba698183),
	.w3(32'h3bbd159b),
	.w4(32'hba616e65),
	.w5(32'hb99fb69e),
	.w6(32'h3b300462),
	.w7(32'h39bdb9aa),
	.w8(32'h3a538bda),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357471),
	.w1(32'hbb590d39),
	.w2(32'hbc2c7917),
	.w3(32'hb9ce2b9c),
	.w4(32'h3bacea66),
	.w5(32'h3c786fb0),
	.w6(32'h3b8fbb28),
	.w7(32'h3be1103f),
	.w8(32'h39697cad),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70f09),
	.w1(32'hb6cb582a),
	.w2(32'hba85e8f5),
	.w3(32'h3c2ccfda),
	.w4(32'hb9f61d39),
	.w5(32'h3c08290f),
	.w6(32'hba9d7ade),
	.w7(32'hba874111),
	.w8(32'hbb2aedd3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f407e0),
	.w1(32'hba1e7703),
	.w2(32'hba6600df),
	.w3(32'hbb06336c),
	.w4(32'hbb037fbb),
	.w5(32'h3b067f38),
	.w6(32'hba9b0e95),
	.w7(32'hbb68577b),
	.w8(32'hbb8e64db),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80404f),
	.w1(32'h3b890282),
	.w2(32'h3b4d8307),
	.w3(32'h3ae5c8f6),
	.w4(32'hbc0188c9),
	.w5(32'hbbd7da3d),
	.w6(32'hbbba02fa),
	.w7(32'h3be79e2d),
	.w8(32'hbaaa5074),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80af71),
	.w1(32'h3a05953d),
	.w2(32'h3b168d82),
	.w3(32'hbb705c0a),
	.w4(32'h3a981f28),
	.w5(32'hbc369c93),
	.w6(32'h3a5b908b),
	.w7(32'hb91efe9c),
	.w8(32'hbb83f24f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8725b),
	.w1(32'hbb03262a),
	.w2(32'hbb98edb6),
	.w3(32'h3ab83dec),
	.w4(32'h3b83f302),
	.w5(32'hbb148870),
	.w6(32'h3b6eb08d),
	.w7(32'h3b676bd4),
	.w8(32'h3a7298b6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2dcee),
	.w1(32'hbba074e0),
	.w2(32'hba621271),
	.w3(32'h3b8bb2bf),
	.w4(32'hbb426e4f),
	.w5(32'h3ac69885),
	.w6(32'h3ab20e55),
	.w7(32'hbb5c0f85),
	.w8(32'hbb559723),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932771),
	.w1(32'hbbc43320),
	.w2(32'hbb7178b3),
	.w3(32'hbbca33b5),
	.w4(32'h3b156c5e),
	.w5(32'hb7dd1e25),
	.w6(32'hb9e48f94),
	.w7(32'hbbff39f1),
	.w8(32'hbc2a1eea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf49867),
	.w1(32'h3a328751),
	.w2(32'h3a6f6ba7),
	.w3(32'h3806dc68),
	.w4(32'h39f26f8d),
	.w5(32'h3bff8646),
	.w6(32'hbb980a13),
	.w7(32'hbb4c9c50),
	.w8(32'hbb2a5f88),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf08b54),
	.w1(32'h3a5dda57),
	.w2(32'hb9465907),
	.w3(32'h3bfe7866),
	.w4(32'h3931e8a3),
	.w5(32'h37bcb568),
	.w6(32'hba9c536c),
	.w7(32'h39b36a29),
	.w8(32'hba0f4ca9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51e0d4),
	.w1(32'hb87901e0),
	.w2(32'hbba46171),
	.w3(32'h3b274e28),
	.w4(32'hba96a9a0),
	.w5(32'hbb869ee1),
	.w6(32'hba3d26ac),
	.w7(32'h3a22f675),
	.w8(32'hbb6381b2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5993bd),
	.w1(32'h3a015d61),
	.w2(32'h3b5e4655),
	.w3(32'h3aae8ce7),
	.w4(32'h3ae98eff),
	.w5(32'hb9b51889),
	.w6(32'h39340d27),
	.w7(32'hbafec996),
	.w8(32'hbb399d92),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b866),
	.w1(32'h3ad6cfc5),
	.w2(32'hbb7aaa69),
	.w3(32'hbb8babad),
	.w4(32'h3a33b86b),
	.w5(32'hbabed5cf),
	.w6(32'h3b05e3e9),
	.w7(32'h3a5bd8f3),
	.w8(32'h3a976a7f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388deba2),
	.w1(32'hb89d5f79),
	.w2(32'h3a2f181d),
	.w3(32'h3ab2d006),
	.w4(32'hbb918011),
	.w5(32'h3c12b4bb),
	.w6(32'h3a2d9622),
	.w7(32'hbafcb9b2),
	.w8(32'hbbb298c4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add0a20),
	.w1(32'h3abc53b6),
	.w2(32'hbab45dde),
	.w3(32'h3bd5f908),
	.w4(32'hb8b14358),
	.w5(32'hba38e6a2),
	.w6(32'h3a17e8e2),
	.w7(32'h3a5e7c2f),
	.w8(32'h3a043369),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080942),
	.w1(32'hbad7b586),
	.w2(32'hbaa26112),
	.w3(32'h3adba735),
	.w4(32'hba89e5b6),
	.w5(32'hba2eeeac),
	.w6(32'h3b6b18d9),
	.w7(32'hbaf67f75),
	.w8(32'h3bb5a23b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c0f3c),
	.w1(32'hb9cb35f7),
	.w2(32'hb9b72fd3),
	.w3(32'hbafd342f),
	.w4(32'hba723ea5),
	.w5(32'hb9568691),
	.w6(32'h3b28b70b),
	.w7(32'hbb17e5f3),
	.w8(32'hbb9de4e0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717b2e),
	.w1(32'hb959734b),
	.w2(32'h3af8b005),
	.w3(32'h3a499685),
	.w4(32'h3a5beb4f),
	.w5(32'h3c49c00e),
	.w6(32'hbb6b5e77),
	.w7(32'h3a7330a8),
	.w8(32'h39db35ad),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b106dd0),
	.w1(32'hbbad40c7),
	.w2(32'hbc0fb0d0),
	.w3(32'h3b8af3e8),
	.w4(32'hbb928c17),
	.w5(32'hbb363219),
	.w6(32'h3b421865),
	.w7(32'h3ab7318a),
	.w8(32'hbbc6a8bc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5442b6),
	.w1(32'hbb881a2d),
	.w2(32'h3ba5a726),
	.w3(32'hbb363920),
	.w4(32'h3c598dc6),
	.w5(32'h3c032c08),
	.w6(32'hbb354261),
	.w7(32'h3aaabf97),
	.w8(32'h3b2f0b62),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c517760),
	.w1(32'h3b6c7ba1),
	.w2(32'hbbce9c00),
	.w3(32'hb90df942),
	.w4(32'hbab71ee1),
	.w5(32'h3a331c2e),
	.w6(32'hbb04f186),
	.w7(32'hbb208851),
	.w8(32'hbb37d357),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea3766),
	.w1(32'hbb1ca857),
	.w2(32'h39c08a2e),
	.w3(32'h3bd349f1),
	.w4(32'hbb6b409b),
	.w5(32'hbaab62fd),
	.w6(32'h3ab550a4),
	.w7(32'h3a4fec02),
	.w8(32'h3ae3e74e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51cfcf),
	.w1(32'hbae17659),
	.w2(32'hbae210c4),
	.w3(32'hbb0c5010),
	.w4(32'hbb5569ce),
	.w5(32'hbbbaf0da),
	.w6(32'h3a77d9ba),
	.w7(32'h39937f7b),
	.w8(32'h3bc74923),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f73b7),
	.w1(32'h3b42e364),
	.w2(32'hb8839192),
	.w3(32'h3b15fba1),
	.w4(32'hbb3fa8be),
	.w5(32'hba01b838),
	.w6(32'h3ad7229f),
	.w7(32'h3b764c16),
	.w8(32'h392e4ab7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6c848),
	.w1(32'hbb0ff0d2),
	.w2(32'hbac3ef6e),
	.w3(32'hb9aff36f),
	.w4(32'hbac6b960),
	.w5(32'hbb07871e),
	.w6(32'h3aa5bb66),
	.w7(32'hbb2525db),
	.w8(32'hba2a51ca),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ee1bc),
	.w1(32'hbb74446d),
	.w2(32'hba3d73d6),
	.w3(32'hba859fca),
	.w4(32'hbb3b759c),
	.w5(32'hbb251146),
	.w6(32'h3baef9a5),
	.w7(32'h3b4cdcd7),
	.w8(32'h3a595524),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeba79),
	.w1(32'h3a30dc94),
	.w2(32'hbb205ac3),
	.w3(32'hbacb392b),
	.w4(32'hbb2541eb),
	.w5(32'h3aec72d9),
	.w6(32'hb90a5fa0),
	.w7(32'h3a0f82a9),
	.w8(32'hbb966df6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40fd09),
	.w1(32'hbbabf4fc),
	.w2(32'hbaa9d405),
	.w3(32'hbb723b55),
	.w4(32'hbaadb2fa),
	.w5(32'h3aad2536),
	.w6(32'hbbcb7a6d),
	.w7(32'hb9ff75d1),
	.w8(32'h3b3537df),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba017c89),
	.w1(32'hbae0c623),
	.w2(32'h3b8df668),
	.w3(32'hba631c4e),
	.w4(32'hba5e8646),
	.w5(32'hbacc2216),
	.w6(32'h3b68ffd4),
	.w7(32'h3b1a76f2),
	.w8(32'hbb03ecd6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b95f98),
	.w1(32'hbb320ff5),
	.w2(32'hbb28261b),
	.w3(32'hbac4764d),
	.w4(32'hbab12b7f),
	.w5(32'h3a04baaf),
	.w6(32'h3b67d83f),
	.w7(32'hba7aa242),
	.w8(32'h37d5308a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1f02),
	.w1(32'hbbb455d8),
	.w2(32'h3b3eecc4),
	.w3(32'hbaa8112a),
	.w4(32'h3b94b997),
	.w5(32'h3c37f264),
	.w6(32'h3a43b187),
	.w7(32'hbb09f987),
	.w8(32'hbb8b3ee4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b0d5),
	.w1(32'h3a94fa3b),
	.w2(32'hba9ff2b9),
	.w3(32'h3be8e251),
	.w4(32'hbb633b3e),
	.w5(32'h399f72c8),
	.w6(32'hbbf35881),
	.w7(32'h3b2790df),
	.w8(32'h3a27d33a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912aa61),
	.w1(32'h3bab4140),
	.w2(32'h3a2bea55),
	.w3(32'hba3107a6),
	.w4(32'h3bbfc590),
	.w5(32'h3bec2a30),
	.w6(32'hba60a790),
	.w7(32'hba056359),
	.w8(32'hba6297bd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c98b8),
	.w1(32'hbb3a8c61),
	.w2(32'hb6886b6a),
	.w3(32'h3bd438c3),
	.w4(32'hbb82bdb4),
	.w5(32'h3bdb9843),
	.w6(32'hbb9b979f),
	.w7(32'hba8f3a0f),
	.w8(32'hbb4da425),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb420263),
	.w1(32'hbb6f3159),
	.w2(32'hbace2778),
	.w3(32'hbad90f0b),
	.w4(32'hbb215466),
	.w5(32'h3be0692e),
	.w6(32'h3a7ed748),
	.w7(32'hb9fe59a0),
	.w8(32'h3b6914a2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1745b0),
	.w1(32'h3af77e9d),
	.w2(32'h3b6c1406),
	.w3(32'h3b811491),
	.w4(32'hbb9dffe1),
	.w5(32'hbbfc2b5e),
	.w6(32'h3ad6b0af),
	.w7(32'h3b251cbf),
	.w8(32'h3ac6239d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae97aad),
	.w1(32'h3bdf8919),
	.w2(32'h3b2ffb5b),
	.w3(32'hbaf908ae),
	.w4(32'h3ab39c62),
	.w5(32'h3c21fcb9),
	.w6(32'hba5708fa),
	.w7(32'hba918350),
	.w8(32'h3bb83029),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d8522),
	.w1(32'h3aea53c4),
	.w2(32'h3aa38301),
	.w3(32'h3c8c8dd1),
	.w4(32'h3b457ca3),
	.w5(32'h3b85e29e),
	.w6(32'h3bd7019e),
	.w7(32'hbae085e4),
	.w8(32'h39bb2a3f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbcaea),
	.w1(32'hbb5520fc),
	.w2(32'hbb43027c),
	.w3(32'h3ad2f90a),
	.w4(32'hbbeefb0d),
	.w5(32'hbba802de),
	.w6(32'h3afe0ce2),
	.w7(32'hbb833b7b),
	.w8(32'hbabc5b52),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6d1d6),
	.w1(32'hbb16dc5a),
	.w2(32'hbb0ab089),
	.w3(32'hbb1a9ec0),
	.w4(32'hbb52896d),
	.w5(32'h3adaeac8),
	.w6(32'h3a770979),
	.w7(32'h3b4e5b6d),
	.w8(32'h3b6753dd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0027d),
	.w1(32'hbbc5b7a1),
	.w2(32'hb9c3df80),
	.w3(32'h3b796b18),
	.w4(32'hbb59ce9f),
	.w5(32'h3a004234),
	.w6(32'h3bb34142),
	.w7(32'h3abed6fc),
	.w8(32'hbb41af7f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28acd0),
	.w1(32'h3af8f8a8),
	.w2(32'h3b13b969),
	.w3(32'hbae5aaf3),
	.w4(32'h3b5a6d04),
	.w5(32'h3b0c7fc4),
	.w6(32'h38de6028),
	.w7(32'hba21d803),
	.w8(32'hbb0b5d26),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad87003),
	.w1(32'h3b3f83e5),
	.w2(32'h3a875830),
	.w3(32'h3ac2938f),
	.w4(32'hbbd72212),
	.w5(32'h3a905837),
	.w6(32'h3b28bd1f),
	.w7(32'hbb3ed973),
	.w8(32'hba933dbb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c276f),
	.w1(32'hba82590d),
	.w2(32'h3b6de31d),
	.w3(32'h3a9d520a),
	.w4(32'h3b97dbc9),
	.w5(32'h3bd055b5),
	.w6(32'hbbb1cf7e),
	.w7(32'hbb14995f),
	.w8(32'hbb0d672f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa68561),
	.w1(32'hbae7e94d),
	.w2(32'h3b69dbce),
	.w3(32'h3c19a860),
	.w4(32'hbb464ac8),
	.w5(32'hbaba1ebb),
	.w6(32'h39bf23d4),
	.w7(32'hbb2974ce),
	.w8(32'hbb02cb1b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2674a),
	.w1(32'hb9f3b758),
	.w2(32'hbb8acd62),
	.w3(32'hba6a4af7),
	.w4(32'h3aa1eec8),
	.w5(32'hbac180f7),
	.w6(32'hbb4b9985),
	.w7(32'h3b84eb40),
	.w8(32'hbb3d0080),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21b690),
	.w1(32'hb82050d3),
	.w2(32'h3b15011c),
	.w3(32'h3b3d1b10),
	.w4(32'hba3592bf),
	.w5(32'h3b93f25f),
	.w6(32'h3b157bab),
	.w7(32'hb9b98e39),
	.w8(32'hbb481289),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8ab23),
	.w1(32'h3b806d58),
	.w2(32'h3ad76304),
	.w3(32'hba0f56f5),
	.w4(32'h3ae5dc08),
	.w5(32'h3adccab7),
	.w6(32'h3b3b7565),
	.w7(32'hba570220),
	.w8(32'h381f7f88),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b935aa3),
	.w1(32'h3ad7bc33),
	.w2(32'hb7ed4577),
	.w3(32'h39fa9d83),
	.w4(32'h3aabfc3e),
	.w5(32'hba4427b1),
	.w6(32'h3b737f04),
	.w7(32'h3a8d43c9),
	.w8(32'h3b1acdc8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dee2b),
	.w1(32'hbb98c50b),
	.w2(32'hbbaea048),
	.w3(32'hbb3069e1),
	.w4(32'hbb0d79bd),
	.w5(32'hb9929fb5),
	.w6(32'h3a824cd4),
	.w7(32'hbb873e2e),
	.w8(32'h3bbd6c8b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08d2ce),
	.w1(32'h3b345234),
	.w2(32'hbb94ae63),
	.w3(32'h3b1fabd4),
	.w4(32'h39564bff),
	.w5(32'h3b1024e6),
	.w6(32'h3b740d36),
	.w7(32'hba9a1176),
	.w8(32'h3b4dc1f4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea3321),
	.w1(32'hb8e0a0c2),
	.w2(32'hba18d3aa),
	.w3(32'hb8e5f3c1),
	.w4(32'hb911afca),
	.w5(32'hb9936216),
	.w6(32'h3b01ecf4),
	.w7(32'h3abe39f2),
	.w8(32'h3afb84be),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915f0d),
	.w1(32'h3b194d20),
	.w2(32'hba8bf227),
	.w3(32'hbae0c5fa),
	.w4(32'hba98a23e),
	.w5(32'hbb42d51b),
	.w6(32'h3b680c41),
	.w7(32'h3abebf11),
	.w8(32'h3b8150d4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b493bf0),
	.w1(32'h3acddab1),
	.w2(32'h3b7f572d),
	.w3(32'hbb412276),
	.w4(32'hbaa459c6),
	.w5(32'h3a617638),
	.w6(32'h3b2d23c5),
	.w7(32'h39909ada),
	.w8(32'h3b159791),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89eda9),
	.w1(32'hb887355e),
	.w2(32'h3b843822),
	.w3(32'hb8d14e6a),
	.w4(32'hb983f3da),
	.w5(32'hba238777),
	.w6(32'h3b0c0013),
	.w7(32'hba69a93a),
	.w8(32'h3a5966a5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad35f2a),
	.w1(32'h3ac9b7e7),
	.w2(32'h389c9ccb),
	.w3(32'hbb0d9e8f),
	.w4(32'hb9f123f9),
	.w5(32'hbb3b2371),
	.w6(32'h394816e6),
	.w7(32'h3aebceb1),
	.w8(32'h3ae5c763),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e93d2),
	.w1(32'hbaf2374b),
	.w2(32'h3a8e35a5),
	.w3(32'h3b2491dc),
	.w4(32'hba5bc1f9),
	.w5(32'h377738fb),
	.w6(32'h3b25adda),
	.w7(32'h3a38d1f6),
	.w8(32'h3ab6b7d4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30faa6),
	.w1(32'h3a3f3b0d),
	.w2(32'hbb2f0ddf),
	.w3(32'h3a9c83e3),
	.w4(32'hbaa1ff59),
	.w5(32'h3b093100),
	.w6(32'h3aea84b1),
	.w7(32'h39b93488),
	.w8(32'h3a4bc4e5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80bc74),
	.w1(32'hbb30187a),
	.w2(32'hbb3974ce),
	.w3(32'h3b1b5ee6),
	.w4(32'h3b404710),
	.w5(32'hbbd2232a),
	.w6(32'hba8e446e),
	.w7(32'h3a8e56a4),
	.w8(32'hbaf5ae10),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb513406),
	.w1(32'hbb35d436),
	.w2(32'h3bd0cd0b),
	.w3(32'hbbe17fbe),
	.w4(32'h3b08a7ef),
	.w5(32'hbaeaf9d3),
	.w6(32'hbab6468c),
	.w7(32'hbad018c9),
	.w8(32'hbaaf0bdd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a080),
	.w1(32'hba352e1d),
	.w2(32'hb9fd5a8a),
	.w3(32'hba31b9cd),
	.w4(32'hbbb5d5f1),
	.w5(32'hbb8267f6),
	.w6(32'h3a27c78b),
	.w7(32'h3b77abb1),
	.w8(32'h3af4ffcb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57a1a8),
	.w1(32'h3a158470),
	.w2(32'h3c03290c),
	.w3(32'hbb8d2b82),
	.w4(32'hbb294d94),
	.w5(32'hbbab2163),
	.w6(32'h3a542dcb),
	.w7(32'h3b0df70a),
	.w8(32'hb9a82a53),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed1fea),
	.w1(32'hbafb3719),
	.w2(32'hbb5cad64),
	.w3(32'hbaeb65c6),
	.w4(32'hbb6239ab),
	.w5(32'h3b691b57),
	.w6(32'hbaa3a1b7),
	.w7(32'hbb685a09),
	.w8(32'hbb637777),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8e275),
	.w1(32'h3ae05058),
	.w2(32'hbb500aad),
	.w3(32'hb9ad0c47),
	.w4(32'h3c0cc8bb),
	.w5(32'h3bddd5a0),
	.w6(32'hbba60171),
	.w7(32'h3c09d8f8),
	.w8(32'h3bf07172),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b73787),
	.w1(32'hbb7c64e7),
	.w2(32'h3a8fec13),
	.w3(32'h3bbdaccb),
	.w4(32'hbae28908),
	.w5(32'h396479c6),
	.w6(32'h3b8b1ad6),
	.w7(32'hbaf22eb8),
	.w8(32'hba8a8d06),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaaff0),
	.w1(32'h3be27cd7),
	.w2(32'h3c1901e3),
	.w3(32'h399a3751),
	.w4(32'h3c01c1e2),
	.w5(32'hba62c5d1),
	.w6(32'h3a48050c),
	.w7(32'hbae74958),
	.w8(32'hba7fddea),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34f562),
	.w1(32'h3b34bffc),
	.w2(32'h39c26ce4),
	.w3(32'hba9e6c8b),
	.w4(32'h3ace4a3b),
	.w5(32'h3b2bd0d1),
	.w6(32'h3a705fa8),
	.w7(32'hba7e33c7),
	.w8(32'h3babda59),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b95a),
	.w1(32'h3bacfc96),
	.w2(32'h3b8563f3),
	.w3(32'h3b899d8a),
	.w4(32'hbb8ba2c0),
	.w5(32'hbad70cbe),
	.w6(32'hba7b726b),
	.w7(32'hbb708de6),
	.w8(32'hbaa1874a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb813b3),
	.w1(32'hbba1f2a1),
	.w2(32'hbb19f40b),
	.w3(32'hbba530a6),
	.w4(32'h3b10a246),
	.w5(32'h3978ea80),
	.w6(32'hbab94456),
	.w7(32'h3b16d006),
	.w8(32'h3b2e1f26),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33c4a6),
	.w1(32'hbab3a860),
	.w2(32'hbbdd7736),
	.w3(32'h3a1a3c6d),
	.w4(32'hbb178e35),
	.w5(32'h3af2fbbf),
	.w6(32'h3bd24d87),
	.w7(32'h3a9b3c53),
	.w8(32'h3b9833fe),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1a1a8),
	.w1(32'h3aeda996),
	.w2(32'h3b9d61a5),
	.w3(32'h3b0ac3d7),
	.w4(32'hbb2329d0),
	.w5(32'h3ae3ad71),
	.w6(32'h3b6dc1b7),
	.w7(32'hbb4623a5),
	.w8(32'hbb180016),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b664),
	.w1(32'h3ae09956),
	.w2(32'hbb8196eb),
	.w3(32'hba274c62),
	.w4(32'h39c55444),
	.w5(32'h3b3b45f0),
	.w6(32'hba4a296b),
	.w7(32'hbb4cdd09),
	.w8(32'h3b4608e5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58b4c3),
	.w1(32'h3a4fed78),
	.w2(32'hba91e46b),
	.w3(32'hbb914281),
	.w4(32'h390ffbc2),
	.w5(32'hbb0e9c6e),
	.w6(32'hbba34bbf),
	.w7(32'h3a4fcc6e),
	.w8(32'hbb65f329),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e5eb3),
	.w1(32'h3b4a5e88),
	.w2(32'hba3cd415),
	.w3(32'hbaa110c0),
	.w4(32'h3b8b0cd3),
	.w5(32'h3abd3878),
	.w6(32'hbb584680),
	.w7(32'h3a51f3bb),
	.w8(32'hb9afcf13),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9490dcb),
	.w1(32'hbb3c0371),
	.w2(32'hbb2921ff),
	.w3(32'h3afa04c2),
	.w4(32'hba09691d),
	.w5(32'hbb8aabf0),
	.w6(32'h3af33ccb),
	.w7(32'hbb0cb5a1),
	.w8(32'hb9c8f2f6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e62211),
	.w1(32'h3a473e9d),
	.w2(32'h3ade48c8),
	.w3(32'hbb15f5a8),
	.w4(32'hbac60df3),
	.w5(32'hbbcb4f71),
	.w6(32'h3b4baa6a),
	.w7(32'h3b5c6284),
	.w8(32'h3989dbd7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ceda5),
	.w1(32'hbbd2d039),
	.w2(32'hbb6a6ee7),
	.w3(32'hba63077f),
	.w4(32'hba9ae4b2),
	.w5(32'h3b272137),
	.w6(32'h39e08010),
	.w7(32'hba0d3941),
	.w8(32'hbaa2f269),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee094),
	.w1(32'h3a5ad967),
	.w2(32'h3ad2f638),
	.w3(32'hbb075b99),
	.w4(32'hba72e86f),
	.w5(32'h3afc122d),
	.w6(32'hbb577227),
	.w7(32'hbbfd4f55),
	.w8(32'hbb2cdf55),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f1f42),
	.w1(32'h397a6b61),
	.w2(32'hba8945f3),
	.w3(32'hbbe3cd6d),
	.w4(32'hb8c1eed4),
	.w5(32'hbb6704f1),
	.w6(32'hbb3d7dbe),
	.w7(32'h3a30b58e),
	.w8(32'hbb672442),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb019c98),
	.w1(32'hbbbf11e8),
	.w2(32'h3a251efb),
	.w3(32'hbb65ba03),
	.w4(32'hb9d86ddc),
	.w5(32'hbb263ea4),
	.w6(32'hbb08b2e8),
	.w7(32'hbb2cbaa4),
	.w8(32'hb9729278),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cab59),
	.w1(32'h3a8b153c),
	.w2(32'h3b075e88),
	.w3(32'hbb1247e9),
	.w4(32'hbb8b1ee7),
	.w5(32'hbabdf53d),
	.w6(32'h3aea9367),
	.w7(32'hbaa9b56d),
	.w8(32'h39e53077),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade762f),
	.w1(32'hbb409807),
	.w2(32'hbb9d5904),
	.w3(32'hbb268fac),
	.w4(32'hbb9dd32f),
	.w5(32'hbbb08f97),
	.w6(32'hb928b9a4),
	.w7(32'hbb99ae87),
	.w8(32'hbaddc8b6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c6a8),
	.w1(32'h381b1509),
	.w2(32'hbba1a097),
	.w3(32'hbb0880dc),
	.w4(32'hba926f33),
	.w5(32'hbb093f98),
	.w6(32'hba9a428a),
	.w7(32'h3ae04d47),
	.w8(32'h394d6a28),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125c66),
	.w1(32'hbbe38e90),
	.w2(32'hbbcfe909),
	.w3(32'hbb344b10),
	.w4(32'h39dc256f),
	.w5(32'h3c2318d6),
	.w6(32'h3a3349d0),
	.w7(32'h38c996da),
	.w8(32'hbbc8c946),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a3ef7),
	.w1(32'h3b111800),
	.w2(32'h3aa4da24),
	.w3(32'hba833dc8),
	.w4(32'h3b44d7c7),
	.w5(32'hba5944ad),
	.w6(32'hbb00fcd4),
	.w7(32'h3b5ced01),
	.w8(32'h3a975576),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb8146),
	.w1(32'h3b90e958),
	.w2(32'hba40415f),
	.w3(32'hba7035f3),
	.w4(32'h3b7ccc67),
	.w5(32'hb8b3aacb),
	.w6(32'hb9ed1276),
	.w7(32'h3ba0bf74),
	.w8(32'hbb23ca9a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2356f3),
	.w1(32'hbb5988c4),
	.w2(32'hba794c7e),
	.w3(32'hbb5e0092),
	.w4(32'hbb53a951),
	.w5(32'hbb1f3f00),
	.w6(32'hbb49287e),
	.w7(32'hba42dac5),
	.w8(32'hbb973f53),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61696e),
	.w1(32'h3a8ecb43),
	.w2(32'h3a796694),
	.w3(32'hbb9624ea),
	.w4(32'hbb92b6b9),
	.w5(32'hbb0a48f7),
	.w6(32'hbb967203),
	.w7(32'h3a0211cc),
	.w8(32'hbab703b9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff825),
	.w1(32'hbb4659d1),
	.w2(32'hbbcffda3),
	.w3(32'hbb3833f0),
	.w4(32'hbbbb880c),
	.w5(32'hbb9403ee),
	.w6(32'h39524e14),
	.w7(32'hbb0551a3),
	.w8(32'hbba0d39b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d51c6),
	.w1(32'h3aed2912),
	.w2(32'h3a838462),
	.w3(32'hbc022408),
	.w4(32'hba5afca5),
	.w5(32'h3ac88dcd),
	.w6(32'hbb116253),
	.w7(32'hba95380b),
	.w8(32'h3ab2424d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abedf),
	.w1(32'h3adb4ee9),
	.w2(32'h3998a414),
	.w3(32'h3a700fc2),
	.w4(32'hbb683da1),
	.w5(32'hbaac36a0),
	.w6(32'hbac61851),
	.w7(32'hb8a0b66e),
	.w8(32'hba026279),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2292d),
	.w1(32'hbbc392c9),
	.w2(32'hbaf2bac8),
	.w3(32'hbb02adc5),
	.w4(32'hb9d3ef94),
	.w5(32'h389ac1fe),
	.w6(32'hbbaf4d4c),
	.w7(32'h3a8b963e),
	.w8(32'h39b4ad3a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a284),
	.w1(32'hbb4da93b),
	.w2(32'hbb99056e),
	.w3(32'hba3db75f),
	.w4(32'hbb94c2b3),
	.w5(32'hbbcd9bf0),
	.w6(32'h3bb42769),
	.w7(32'h398d3f12),
	.w8(32'h3a4da389),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b074a0f),
	.w1(32'h3bbbe125),
	.w2(32'h3bb9ce3d),
	.w3(32'hba81b48e),
	.w4(32'h3bdad6be),
	.w5(32'h3c536cbd),
	.w6(32'h3710d09b),
	.w7(32'h3b16a639),
	.w8(32'h3b938d54),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ed58),
	.w1(32'hbb8bd2e5),
	.w2(32'hbb820209),
	.w3(32'h3c41bc44),
	.w4(32'hbb71d7a6),
	.w5(32'hbbfe4a16),
	.w6(32'h3b9949bc),
	.w7(32'hbb922914),
	.w8(32'hbaf1262a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb682c75),
	.w1(32'hbaa3ca0c),
	.w2(32'h3b00496c),
	.w3(32'hbb67a33d),
	.w4(32'hba2cca54),
	.w5(32'hbab04cae),
	.w6(32'h39bb43c5),
	.w7(32'hbaa94c4b),
	.w8(32'h3a9d97f0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafca465),
	.w1(32'hbae61c87),
	.w2(32'hbb492009),
	.w3(32'hbb71791c),
	.w4(32'hbb74f047),
	.w5(32'hbb461eaa),
	.w6(32'h39e68787),
	.w7(32'hbaeb1d8a),
	.w8(32'hba85070a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10228c),
	.w1(32'hbc10d1d0),
	.w2(32'hbc206622),
	.w3(32'h3b1c16a5),
	.w4(32'h3bd2e01b),
	.w5(32'h3cad2762),
	.w6(32'hbb520b0f),
	.w7(32'hbb814fbb),
	.w8(32'hbbb1632e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc9d8f),
	.w1(32'hbb0967b7),
	.w2(32'h3b0d895b),
	.w3(32'h3c328c45),
	.w4(32'h3abaf46c),
	.w5(32'h3af38e1a),
	.w6(32'hbb5f4f5c),
	.w7(32'h3b295ebe),
	.w8(32'h3b641d29),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2950ed),
	.w1(32'hbb942aac),
	.w2(32'h3b8a45ad),
	.w3(32'h3adbbf59),
	.w4(32'h3a5fc0aa),
	.w5(32'hbba139f6),
	.w6(32'h3bfdfbeb),
	.w7(32'h3acfa17d),
	.w8(32'hbb038716),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf59f6),
	.w1(32'hb99924d2),
	.w2(32'h3b2f16b5),
	.w3(32'hba404fd5),
	.w4(32'hbada349c),
	.w5(32'hb87a40fb),
	.w6(32'h3b5490aa),
	.w7(32'hba8ab898),
	.w8(32'hba43b5b9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d070af),
	.w1(32'h3b9bea3d),
	.w2(32'h3b6f60c1),
	.w3(32'hbac27f11),
	.w4(32'h3af6932a),
	.w5(32'h3bb0b2ed),
	.w6(32'h3bd77b90),
	.w7(32'h3ba3054e),
	.w8(32'h3b69207a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac750d),
	.w1(32'h3b38e1f6),
	.w2(32'h3aa8fa90),
	.w3(32'h3a95367c),
	.w4(32'h39bf286b),
	.w5(32'hbb8d4240),
	.w6(32'h3abf52f5),
	.w7(32'h3a8d4906),
	.w8(32'h3982daca),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd0523),
	.w1(32'hba29c2ba),
	.w2(32'h398d938f),
	.w3(32'h3b974f6b),
	.w4(32'h39b0b274),
	.w5(32'h3a89c55b),
	.w6(32'h39f0476d),
	.w7(32'h3b3bb795),
	.w8(32'h3b2f7e8d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb528),
	.w1(32'hbb862282),
	.w2(32'hbb7e40bd),
	.w3(32'h3b80fb21),
	.w4(32'hbb9f6f06),
	.w5(32'h3b830a5f),
	.w6(32'h39f0ff10),
	.w7(32'h38f23978),
	.w8(32'h39852d50),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8725db),
	.w1(32'h3b9f49f5),
	.w2(32'hbb374c0d),
	.w3(32'h3a3da02e),
	.w4(32'h3b4f30b4),
	.w5(32'hbb9b2368),
	.w6(32'h3a8ff718),
	.w7(32'h3b8b9234),
	.w8(32'h3a7cf715),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290b3e),
	.w1(32'h3bc09fd9),
	.w2(32'hb99d3b98),
	.w3(32'h3a566a38),
	.w4(32'h37baf97c),
	.w5(32'hbb9bfddb),
	.w6(32'h3ac5c07b),
	.w7(32'hbb27d431),
	.w8(32'hbc09d572),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2345c5),
	.w1(32'h3acf5f44),
	.w2(32'h3b285ffd),
	.w3(32'h3b964610),
	.w4(32'hb98c9338),
	.w5(32'hbb3fff28),
	.w6(32'hb9983572),
	.w7(32'hbbf51cf3),
	.w8(32'hbbcd3a77),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89af2c),
	.w1(32'h3aab491a),
	.w2(32'h3b516ac7),
	.w3(32'hbbbeefcf),
	.w4(32'hbbcbeb49),
	.w5(32'h3ab51553),
	.w6(32'hbc1bab12),
	.w7(32'hba06df67),
	.w8(32'hbbc2d487),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b591c),
	.w1(32'h3b30f00c),
	.w2(32'h3b4f4c87),
	.w3(32'hbc39517e),
	.w4(32'h3b8b7cd0),
	.w5(32'h3c277fd3),
	.w6(32'hbb5dc678),
	.w7(32'hba3e2ce1),
	.w8(32'h3ba0910c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf57a9),
	.w1(32'hbbefb7fe),
	.w2(32'hbc1dcf6b),
	.w3(32'h3b199409),
	.w4(32'hbb913f6f),
	.w5(32'hbc27257e),
	.w6(32'hbb0475a2),
	.w7(32'hbbbe27f1),
	.w8(32'hbc140755),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87611b),
	.w1(32'hbc2c2e94),
	.w2(32'hbb04c286),
	.w3(32'hbb8f446f),
	.w4(32'hbbb7b780),
	.w5(32'hbadcdfd9),
	.w6(32'hbbca2ca3),
	.w7(32'h399990cf),
	.w8(32'h3bb71ad0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dc671),
	.w1(32'hbc0257c2),
	.w2(32'hbb9d756f),
	.w3(32'h3b3001e7),
	.w4(32'hbc0f4d7d),
	.w5(32'hbc1961ba),
	.w6(32'h3b97b43e),
	.w7(32'hbc2708ae),
	.w8(32'hbbefe834),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d64e),
	.w1(32'hbb8bf66d),
	.w2(32'hbbaad682),
	.w3(32'h39f0f9b9),
	.w4(32'hbbb3689f),
	.w5(32'hbbe28cc8),
	.w6(32'h3aa13695),
	.w7(32'hbbbc85ca),
	.w8(32'hbba40fe6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1169bb),
	.w1(32'h3c1322a2),
	.w2(32'h3b4429c5),
	.w3(32'hba5402e6),
	.w4(32'h3c7281f8),
	.w5(32'h3c3966d9),
	.w6(32'h3ae0438e),
	.w7(32'h3b52c168),
	.w8(32'h3c9d324e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01969b),
	.w1(32'h3c1751f2),
	.w2(32'h3c1c0916),
	.w3(32'h3b617979),
	.w4(32'h3c168b75),
	.w5(32'h3c547dc5),
	.w6(32'h398706dc),
	.w7(32'h3c2431ec),
	.w8(32'h3c48a1a3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d5259),
	.w1(32'hbabf43f1),
	.w2(32'hbbb92a20),
	.w3(32'h3c4d2c32),
	.w4(32'h3bbd12ee),
	.w5(32'hbb0bc4a8),
	.w6(32'h3c65e8f5),
	.w7(32'h3b7f4ae7),
	.w8(32'h3b36c87f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88edf0),
	.w1(32'hba69523a),
	.w2(32'h3a689382),
	.w3(32'h3ad03245),
	.w4(32'h3aafc2b9),
	.w5(32'h3bdb8ed1),
	.w6(32'h3a638af3),
	.w7(32'hba18c528),
	.w8(32'h3b399fe9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e6e0),
	.w1(32'h3a27ae0d),
	.w2(32'hbaca36e7),
	.w3(32'hbb4e8381),
	.w4(32'h391ba3ad),
	.w5(32'h3ab0af66),
	.w6(32'hbbb45948),
	.w7(32'hb9c41df3),
	.w8(32'hbb229e45),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e5018),
	.w1(32'hbbb96b03),
	.w2(32'hbb6305e9),
	.w3(32'hba8c29a1),
	.w4(32'hbb9d1f52),
	.w5(32'hba1b1cac),
	.w6(32'hba90c9e9),
	.w7(32'hbb8f498d),
	.w8(32'hbbd58c15),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a797fa0),
	.w1(32'h39bf721f),
	.w2(32'h3a00e8db),
	.w3(32'hba177800),
	.w4(32'h3b4d7e66),
	.w5(32'hbb82ad11),
	.w6(32'hbb5f99e0),
	.w7(32'hbb455176),
	.w8(32'hbbdfcc00),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856519),
	.w1(32'h3a2ba526),
	.w2(32'hba68087c),
	.w3(32'h3b190472),
	.w4(32'h3bcf8afb),
	.w5(32'h3bda35ce),
	.w6(32'hbace67f6),
	.w7(32'h3bafecf7),
	.w8(32'h3b826390),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a692996),
	.w1(32'h3b8d7927),
	.w2(32'hbc214e4f),
	.w3(32'hbb6f98d1),
	.w4(32'hbb53f982),
	.w5(32'h39fb24c1),
	.w6(32'hbb06547d),
	.w7(32'hbc15b1da),
	.w8(32'hbb8c7e3a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0583d7),
	.w1(32'h3bc1d4ed),
	.w2(32'hbb49ac59),
	.w3(32'hbb9931e4),
	.w4(32'h3c2c21d4),
	.w5(32'h3c4015a3),
	.w6(32'h3ba7cb80),
	.w7(32'h3b5a97de),
	.w8(32'h3b251b47),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa041),
	.w1(32'h3c0e98ce),
	.w2(32'hbc1ab0e4),
	.w3(32'h3b63005e),
	.w4(32'h3bf357a4),
	.w5(32'hbab7a0b7),
	.w6(32'h3a806720),
	.w7(32'h3b62f286),
	.w8(32'h3b5c58c9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fe8bb),
	.w1(32'hbacaf5d7),
	.w2(32'hbabd8848),
	.w3(32'h3ab80a8f),
	.w4(32'hba9645d7),
	.w5(32'hbbaf8e08),
	.w6(32'h3bf27845),
	.w7(32'hba52c9a7),
	.w8(32'hba5de1cb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fe1cc),
	.w1(32'hba0f1397),
	.w2(32'h3abf5963),
	.w3(32'h3b9f3ea8),
	.w4(32'hb9c0f977),
	.w5(32'h3be0eb8b),
	.w6(32'h3be0c3d5),
	.w7(32'h3b99014d),
	.w8(32'h3b527f1e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba050c4b),
	.w1(32'h3bcaebfd),
	.w2(32'hbc09ec9a),
	.w3(32'hb949c390),
	.w4(32'h3ba79b57),
	.w5(32'hbbc499bc),
	.w6(32'h3bbb6eab),
	.w7(32'hbadae458),
	.w8(32'hbbf33e07),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9a405),
	.w1(32'h3baa13f3),
	.w2(32'hbb3db576),
	.w3(32'hbb9b63be),
	.w4(32'h39af282c),
	.w5(32'hbb0f9b6d),
	.w6(32'hba84dc72),
	.w7(32'hbb124e3a),
	.w8(32'hbba49706),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789aba),
	.w1(32'h3a84ecb8),
	.w2(32'h3aadc825),
	.w3(32'h380dea43),
	.w4(32'hbb186419),
	.w5(32'h398591de),
	.w6(32'hb96cfca3),
	.w7(32'hbada7457),
	.w8(32'h3b6de159),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26e828),
	.w1(32'h38207800),
	.w2(32'h3b8a92e1),
	.w3(32'hbc118260),
	.w4(32'h3979effc),
	.w5(32'h3b2cc85b),
	.w6(32'hbaae8c77),
	.w7(32'hbb498473),
	.w8(32'h3c09acb6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b89ba),
	.w1(32'hbb86f3ff),
	.w2(32'hb991ca39),
	.w3(32'hbb74c5cc),
	.w4(32'h3bc19f9a),
	.w5(32'h3baa7191),
	.w6(32'h3b2db924),
	.w7(32'h3a8af248),
	.w8(32'h3c0ff371),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac02eba),
	.w1(32'h39779b0d),
	.w2(32'hbbed25f6),
	.w3(32'h3b14e23d),
	.w4(32'hbc1b71f5),
	.w5(32'hbb8e846d),
	.w6(32'h3af6074d),
	.w7(32'hbbbc89b7),
	.w8(32'hbbf20f20),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a26a4),
	.w1(32'hb9d2efc1),
	.w2(32'hbc086276),
	.w3(32'hbba9af0f),
	.w4(32'hb94baf01),
	.w5(32'hbc3c100b),
	.w6(32'hbb4e2913),
	.w7(32'hb9c4be9f),
	.w8(32'hbc29458b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e3b3),
	.w1(32'h3b542aea),
	.w2(32'h3b1b7fc6),
	.w3(32'hbba14ad1),
	.w4(32'h3bbfd80b),
	.w5(32'h3c2b86b3),
	.w6(32'hbbac7471),
	.w7(32'h3bcf6853),
	.w8(32'h3a40fb70),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d6ea),
	.w1(32'hbb47c4ac),
	.w2(32'hbbcf8637),
	.w3(32'h3a955172),
	.w4(32'hbb1e8bbf),
	.w5(32'hbc4c2156),
	.w6(32'h3abd8a20),
	.w7(32'h3ad66bd6),
	.w8(32'hbc030cf0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562a38),
	.w1(32'hbbace34c),
	.w2(32'h3b0f7744),
	.w3(32'h3b4d4f04),
	.w4(32'hbb7d262e),
	.w5(32'hbb97a723),
	.w6(32'h3a9a7311),
	.w7(32'h3acf37bd),
	.w8(32'hba014d0f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd82e),
	.w1(32'h3ad433bb),
	.w2(32'hbb3deb6b),
	.w3(32'hb9a96fe4),
	.w4(32'h3bac7b1f),
	.w5(32'hbaee9615),
	.w6(32'hbb2dba8d),
	.w7(32'h3b81f22d),
	.w8(32'h3aacee17),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006594),
	.w1(32'hbb9c6e02),
	.w2(32'hbc1a7f40),
	.w3(32'h3ab516b3),
	.w4(32'hbb2ca884),
	.w5(32'hbc2affd5),
	.w6(32'h3b5136bb),
	.w7(32'h3b6316ba),
	.w8(32'hbc07bfe4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c38778),
	.w1(32'h3c28d779),
	.w2(32'hbc543e4a),
	.w3(32'hbc1e9adf),
	.w4(32'h3a8218b4),
	.w5(32'hbc087187),
	.w6(32'hbb289cb3),
	.w7(32'hbaaea252),
	.w8(32'hbbf4142c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110aad),
	.w1(32'h3c1b1134),
	.w2(32'h3c61bda2),
	.w3(32'h3b0301d8),
	.w4(32'h3c9bb4f8),
	.w5(32'h3ce9d79f),
	.w6(32'h3b9a0c4e),
	.w7(32'h3c2520b1),
	.w8(32'h3cad890e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879faf0),
	.w1(32'hbbb6f4ee),
	.w2(32'hbac91e35),
	.w3(32'h3c04aff0),
	.w4(32'hbc34fac9),
	.w5(32'hbace80ff),
	.w6(32'h3ba7c907),
	.w7(32'hbc19d5ca),
	.w8(32'hbb87c042),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33feb7),
	.w1(32'hb9882684),
	.w2(32'hbb0eccf9),
	.w3(32'hbb78f6f8),
	.w4(32'hba677f8c),
	.w5(32'hbb517f37),
	.w6(32'h39802892),
	.w7(32'hbaa63fba),
	.w8(32'hbb8766a2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118102),
	.w1(32'hbadb0f14),
	.w2(32'h39bf3347),
	.w3(32'hbb0e543d),
	.w4(32'h39e617ec),
	.w5(32'hb9779b3c),
	.w6(32'hbb740517),
	.w7(32'hba8fbba0),
	.w8(32'hba19afd8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b7be),
	.w1(32'h3a6368ca),
	.w2(32'hbbc87c15),
	.w3(32'hba105ed2),
	.w4(32'h3b7bf610),
	.w5(32'hbb8d6690),
	.w6(32'hbb78a7c2),
	.w7(32'h3ba82cf3),
	.w8(32'hb90c3643),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921f207),
	.w1(32'hbb6aac67),
	.w2(32'h3a8dc799),
	.w3(32'h38ba6366),
	.w4(32'hbc28235d),
	.w5(32'hba42f540),
	.w6(32'hbac270b2),
	.w7(32'hbba5d5a6),
	.w8(32'hbc0fe304),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f41cc),
	.w1(32'h3ad7c505),
	.w2(32'hba89238e),
	.w3(32'hba3fd891),
	.w4(32'hbbd95942),
	.w5(32'hbbc34872),
	.w6(32'h3a2e9f83),
	.w7(32'hbb2be4b3),
	.w8(32'hbac001fc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf89a0),
	.w1(32'hbbc4377a),
	.w2(32'hba802ab3),
	.w3(32'hbc1a97dd),
	.w4(32'hbb957ee9),
	.w5(32'hbb05712d),
	.w6(32'h3b776de1),
	.w7(32'h3c142922),
	.w8(32'h3c1049cf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f1095),
	.w1(32'h3a15de3b),
	.w2(32'hbb1b7c5d),
	.w3(32'hb6fdcaef),
	.w4(32'hbac8cdd3),
	.w5(32'h399d097b),
	.w6(32'h3c1041c9),
	.w7(32'h3a49db33),
	.w8(32'hbc5b1e1b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e74a0),
	.w1(32'h3a90afef),
	.w2(32'hbb822413),
	.w3(32'hbb0d163d),
	.w4(32'h3bc49eb7),
	.w5(32'hba0e38d0),
	.w6(32'hbbd6f59c),
	.w7(32'h3b940bf2),
	.w8(32'hbb311e1a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba653d6),
	.w1(32'hbc1e2c27),
	.w2(32'h3c0c9db1),
	.w3(32'hbbe0c7ed),
	.w4(32'hbc0ac8d5),
	.w5(32'h3bb60458),
	.w6(32'hbb9c94ed),
	.w7(32'hbc1da32c),
	.w8(32'h3b5fb562),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b78e2),
	.w1(32'h3b828737),
	.w2(32'h3ba5e0eb),
	.w3(32'h3c4da390),
	.w4(32'h3b61cc9a),
	.w5(32'h3ba0aa91),
	.w6(32'h3baef653),
	.w7(32'h3bceaf8a),
	.w8(32'h3bdea9d4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f70f7),
	.w1(32'h3a2cdbe8),
	.w2(32'h3a859344),
	.w3(32'hbabaa55a),
	.w4(32'h3b0e9949),
	.w5(32'hb9842c70),
	.w6(32'hbae69806),
	.w7(32'hbaa97f9f),
	.w8(32'hbb0b516b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc688de),
	.w1(32'hbb3da918),
	.w2(32'hbc507c51),
	.w3(32'hbbe5f908),
	.w4(32'hbb84f408),
	.w5(32'hbc4dbf4b),
	.w6(32'hbbc11abf),
	.w7(32'hbb011091),
	.w8(32'hbc231d45),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bcb84),
	.w1(32'h3b97cd4b),
	.w2(32'h3c7e1094),
	.w3(32'hbc8ae6aa),
	.w4(32'h3b099881),
	.w5(32'h3c6cc6f4),
	.w6(32'hbc338ca0),
	.w7(32'h3bc32f74),
	.w8(32'h3ca4edb7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ef36f),
	.w1(32'h3b8ea80f),
	.w2(32'hbc089c1b),
	.w3(32'h3b2c22ae),
	.w4(32'h3b8638b3),
	.w5(32'hb8c3cafb),
	.w6(32'h3c2bfbd5),
	.w7(32'h3b619070),
	.w8(32'hb82c5a8b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a47a),
	.w1(32'h3ad9a863),
	.w2(32'hbbecb430),
	.w3(32'h3a772cad),
	.w4(32'hbbc196c7),
	.w5(32'hbb90bc2e),
	.w6(32'h3929ed5e),
	.w7(32'hbbe7bb69),
	.w8(32'hbc424c31),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2fb5),
	.w1(32'hbb8093dd),
	.w2(32'h3b29bb07),
	.w3(32'hbc26fc7d),
	.w4(32'hbba3a85c),
	.w5(32'hb93e3c9d),
	.w6(32'hbc0ccd9e),
	.w7(32'hbbb8620e),
	.w8(32'h3aded6b3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac22dc2),
	.w1(32'h3b980df2),
	.w2(32'h3b02b812),
	.w3(32'hbb96d344),
	.w4(32'hbb48e94c),
	.w5(32'hbbaeec89),
	.w6(32'hbbb61bd6),
	.w7(32'hbbdde5aa),
	.w8(32'hbbba8a84),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fda9),
	.w1(32'h3b848400),
	.w2(32'hbc0d30b2),
	.w3(32'h3a45be13),
	.w4(32'h3b9a8ba9),
	.w5(32'hbc18b971),
	.w6(32'hb9aad008),
	.w7(32'hbb57b6ca),
	.w8(32'hbc145d00),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db92b),
	.w1(32'hbba5a30c),
	.w2(32'hbc859a1a),
	.w3(32'hbbc44998),
	.w4(32'hbc09503f),
	.w5(32'hbc45d0b2),
	.w6(32'hbbf91c15),
	.w7(32'hbbcc1fda),
	.w8(32'hbc7ff48c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a0bd4),
	.w1(32'h3b2e8847),
	.w2(32'h3b4fe16c),
	.w3(32'hbca50613),
	.w4(32'hbb08088e),
	.w5(32'hbb3b1470),
	.w6(32'hbc95d742),
	.w7(32'h3c0a22d4),
	.w8(32'hb903258b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc21dc),
	.w1(32'h3c146ebd),
	.w2(32'h3cbc18ee),
	.w3(32'hbc19fb69),
	.w4(32'h3bccebfb),
	.w5(32'h3cb0dbde),
	.w6(32'h3a748b49),
	.w7(32'h3c5857d8),
	.w8(32'h3cd79659),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be543),
	.w1(32'h3bc9cf17),
	.w2(32'h3bc52657),
	.w3(32'h39e3b530),
	.w4(32'h3bd883b6),
	.w5(32'hbbde1132),
	.w6(32'h3c41cdf9),
	.w7(32'h3bed9e10),
	.w8(32'h3b2c7b38),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae42fe8),
	.w1(32'hbad79fc3),
	.w2(32'hbb8a5008),
	.w3(32'hbb3c8296),
	.w4(32'hbc0129f3),
	.w5(32'hbbee4b4d),
	.w6(32'hbb114ef8),
	.w7(32'hbbead870),
	.w8(32'hbc075db2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule