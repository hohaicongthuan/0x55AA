module layer_10_featuremap_380(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b870fe),
	.w1(32'hb3d0c46e),
	.w2(32'h352ddb6f),
	.w3(32'hb3494e7f),
	.w4(32'hb5b95b2c),
	.w5(32'hb559617e),
	.w6(32'h35dee964),
	.w7(32'hb58a7fab),
	.w8(32'hb50d8852),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8922da4),
	.w1(32'hb835731d),
	.w2(32'hb897119a),
	.w3(32'h380c8957),
	.w4(32'h3813495c),
	.w5(32'h374294cd),
	.w6(32'h3815f994),
	.w7(32'h38d6b17f),
	.w8(32'h3872f7ff),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c9aaa3),
	.w1(32'hb3d7c393),
	.w2(32'h348a0093),
	.w3(32'h35348e37),
	.w4(32'hb556a565),
	.w5(32'hb4dd4150),
	.w6(32'h34eefc0b),
	.w7(32'h3607c204),
	.w8(32'h36117248),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b667cf),
	.w1(32'h37fad4ca),
	.w2(32'hb553a277),
	.w3(32'h3775f17f),
	.w4(32'h380826a3),
	.w5(32'h381572a6),
	.w6(32'h34d37b66),
	.w7(32'hb793699f),
	.w8(32'hb7186745),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e21d2e),
	.w1(32'h3630a1c4),
	.w2(32'h36062362),
	.w3(32'h364e3c99),
	.w4(32'h3645a755),
	.w5(32'h35be5c7e),
	.w6(32'h360c8dee),
	.w7(32'h36a7f9be),
	.w8(32'h3669e56e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3308ff1a),
	.w1(32'h35526913),
	.w2(32'hb459e7d9),
	.w3(32'hb5d97f22),
	.w4(32'h34f2b6f4),
	.w5(32'hb585d74f),
	.w6(32'hb5770aaf),
	.w7(32'hb52e6dc7),
	.w8(32'hb5775ae3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8281c26),
	.w1(32'hb8ad5919),
	.w2(32'hb8a39a40),
	.w3(32'hb80c9387),
	.w4(32'hb8285cf4),
	.w5(32'hb8155df3),
	.w6(32'hb88cd324),
	.w7(32'hb8afb7aa),
	.w8(32'hb82f1ee5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e87d3),
	.w1(32'h392aa174),
	.w2(32'h38a9e9da),
	.w3(32'h38b24fdf),
	.w4(32'h390343a7),
	.w5(32'h38e837f8),
	.w6(32'hb9969d1f),
	.w7(32'hb8bc9476),
	.w8(32'hb9dd25f5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a38e7f),
	.w1(32'h3741e152),
	.w2(32'h381a0607),
	.w3(32'h379ad6b7),
	.w4(32'h37a44852),
	.w5(32'h377dccdb),
	.w6(32'h37c149f1),
	.w7(32'h381792dd),
	.w8(32'h37bc36e6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf65e0),
	.w1(32'hb9c5b3c5),
	.w2(32'hb99c6a67),
	.w3(32'hb91b261d),
	.w4(32'hb91ae9fa),
	.w5(32'hb8a66b42),
	.w6(32'hb9039b53),
	.w7(32'hb92aa40a),
	.w8(32'hb8847f09),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c50dc3),
	.w1(32'hb6c5c759),
	.w2(32'h37a1a067),
	.w3(32'h37f7462b),
	.w4(32'hb67524f3),
	.w5(32'h3767f4e1),
	.w6(32'h37f38ebd),
	.w7(32'hb6ab22dd),
	.w8(32'h37a4c33e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f3d9f1),
	.w1(32'hb63eb96e),
	.w2(32'hb8aae908),
	.w3(32'hb83b8aa1),
	.w4(32'h38b49cf4),
	.w5(32'hb75ca78f),
	.w6(32'hb8d9df94),
	.w7(32'hb85769f1),
	.w8(32'hb893811a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f76dc),
	.w1(32'hb9cb7703),
	.w2(32'hb96e5779),
	.w3(32'hb8eae0e7),
	.w4(32'hb941d28a),
	.w5(32'hb81d2e18),
	.w6(32'hb915b805),
	.w7(32'hb9160630),
	.w8(32'hb8943334),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc9a20),
	.w1(32'h368902e0),
	.w2(32'h36cccad9),
	.w3(32'h34ef434d),
	.w4(32'h364df431),
	.w5(32'h3588b9e0),
	.w6(32'h3715cd0f),
	.w7(32'h357748ab),
	.w8(32'h36d26e2a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b07924),
	.w1(32'hb8ac5076),
	.w2(32'hb90d8ce4),
	.w3(32'h38928c52),
	.w4(32'hb7486b18),
	.w5(32'hb6a6cc37),
	.w6(32'hb8dbbc90),
	.w7(32'hb7f05d58),
	.w8(32'h37ecf22f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b4bb5),
	.w1(32'hb946b72b),
	.w2(32'hb8a1268f),
	.w3(32'h36a96a55),
	.w4(32'h37416c29),
	.w5(32'h38971806),
	.w6(32'hb8ede97f),
	.w7(32'hb8d83316),
	.w8(32'hb8dd94fd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37096d85),
	.w1(32'hb79e7e4c),
	.w2(32'h37078373),
	.w3(32'hb59b8090),
	.w4(32'hb7a7f5f8),
	.w5(32'hb53456de),
	.w6(32'h370bd409),
	.w7(32'hb79fb415),
	.w8(32'h372436e3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376ce01c),
	.w1(32'hb8ff8056),
	.w2(32'h37abc026),
	.w3(32'h38814df0),
	.w4(32'h38d4cd18),
	.w5(32'h394aa58f),
	.w6(32'hb9d4a75c),
	.w7(32'hb9c5616f),
	.w8(32'hb95145d7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f076c0),
	.w1(32'hb9128300),
	.w2(32'hb8830374),
	.w3(32'hb8d516d5),
	.w4(32'hb8ab53fc),
	.w5(32'h37d1636d),
	.w6(32'hb93c1a93),
	.w7(32'hb91281b9),
	.w8(32'hb8455f5c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ad305a),
	.w1(32'hb611291f),
	.w2(32'h3601b307),
	.w3(32'h34358397),
	.w4(32'h34fe3bfe),
	.w5(32'h35a1786a),
	.w6(32'hb44906c3),
	.w7(32'hb50ad543),
	.w8(32'h35b40422),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364d2414),
	.w1(32'h36458cb0),
	.w2(32'hb4cc9a47),
	.w3(32'h359a92f3),
	.w4(32'h36185f73),
	.w5(32'hb6292dfb),
	.w6(32'hb415ef71),
	.w7(32'h3520e7ef),
	.w8(32'hb61e494c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e9f6f7),
	.w1(32'h372d369c),
	.w2(32'hb7defd8c),
	.w3(32'h3624544c),
	.w4(32'h37936d2e),
	.w5(32'hb7f69146),
	.w6(32'hb68181f0),
	.w7(32'hb725a681),
	.w8(32'hb8493fc6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a0b099),
	.w1(32'hb8b6ef99),
	.w2(32'hb9e895d1),
	.w3(32'hb911ae5c),
	.w4(32'h39ebff11),
	.w5(32'hb80516ee),
	.w6(32'hb9a7349c),
	.w7(32'h38c632b2),
	.w8(32'hba06b55d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acc154),
	.w1(32'hb99a467e),
	.w2(32'hb9635f89),
	.w3(32'hb92d127b),
	.w4(32'hb8f5f1fd),
	.w5(32'hb8e253d3),
	.w6(32'hb8ddcd26),
	.w7(32'hb91c1efb),
	.w8(32'hb8d46b46),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6f715),
	.w1(32'hb99cb2c1),
	.w2(32'hb9b6ef84),
	.w3(32'hb8aa9437),
	.w4(32'hb39ee11f),
	.w5(32'hb91912e0),
	.w6(32'h381bde36),
	.w7(32'hb81c7677),
	.w8(32'hb7e44a40),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ff3c3d),
	.w1(32'hb708f367),
	.w2(32'hb6b2ab22),
	.w3(32'hb6e199e4),
	.w4(32'hb77573eb),
	.w5(32'hb75fdd28),
	.w6(32'hb7005ecd),
	.w7(32'hb7838b52),
	.w8(32'hb6e6ddff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366cef77),
	.w1(32'h369c7c4d),
	.w2(32'hb5c6c4e6),
	.w3(32'h358ad99d),
	.w4(32'h35d135ec),
	.w5(32'hb634444d),
	.w6(32'h3657e3f1),
	.w7(32'h3546de14),
	.w8(32'h34f6574f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b9267),
	.w1(32'hb8cf9496),
	.w2(32'hb903863d),
	.w3(32'h38962b6a),
	.w4(32'h373614d0),
	.w5(32'hb7fbe34e),
	.w6(32'h390b2cc3),
	.w7(32'h378b5600),
	.w8(32'hb80f476c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38544fba),
	.w1(32'h3704a0c7),
	.w2(32'h3838d63f),
	.w3(32'h3840e7dc),
	.w4(32'h37acba30),
	.w5(32'h37c9baa6),
	.w6(32'h37b79745),
	.w7(32'hb5fa58ac),
	.w8(32'hb72bdf3e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991a41d),
	.w1(32'hb98636f2),
	.w2(32'hb9584379),
	.w3(32'hb8af5f9f),
	.w4(32'hb870ed2b),
	.w5(32'hb90b4e1b),
	.w6(32'hb7ef15d4),
	.w7(32'hb7a5adcc),
	.w8(32'hb875a665),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362cab4a),
	.w1(32'hb6951b1d),
	.w2(32'hb662e023),
	.w3(32'hb488e1aa),
	.w4(32'hb6b4a6ff),
	.w5(32'hb63103a2),
	.w6(32'h34a773b1),
	.w7(32'hb5dd9341),
	.w8(32'hb5aa513b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fa026f),
	.w1(32'hb692745a),
	.w2(32'h3660e59b),
	.w3(32'h36ac3d59),
	.w4(32'hb7224967),
	.w5(32'h36be5e90),
	.w6(32'h369b8ef7),
	.w7(32'hb7009f58),
	.w8(32'h36b957b1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fcf8c4),
	.w1(32'hb8fd30e1),
	.w2(32'hb8b9608c),
	.w3(32'hb877ee6c),
	.w4(32'hb81bb144),
	.w5(32'h35b888c2),
	.w6(32'hb8b8ddab),
	.w7(32'hb88fbefd),
	.w8(32'hb8387f59),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2e96f),
	.w1(32'hb84d6ad2),
	.w2(32'hb8269f08),
	.w3(32'h358d1f72),
	.w4(32'h37f3330e),
	.w5(32'h32725d13),
	.w6(32'h37672826),
	.w7(32'h3810046d),
	.w8(32'h37a2800b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69277f6),
	.w1(32'hb608e7bd),
	.w2(32'h3591a745),
	.w3(32'hb5e4b06c),
	.w4(32'h35dc3b76),
	.w5(32'h3685117e),
	.w6(32'hb6c7343c),
	.w7(32'hb6fe7d1b),
	.w8(32'h3669bf31),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8884bd7),
	.w1(32'hb864a811),
	.w2(32'hb7fa137c),
	.w3(32'hb8431509),
	.w4(32'hb7677b39),
	.w5(32'h3683cda1),
	.w6(32'hb8c54d48),
	.w7(32'hb86be1e7),
	.w8(32'hb803a017),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba1aa9),
	.w1(32'hb7a56feb),
	.w2(32'hb94c0ab5),
	.w3(32'h3829dbb8),
	.w4(32'h388f8356),
	.w5(32'hb8bf1915),
	.w6(32'hb925c0f7),
	.w7(32'hb926eb63),
	.w8(32'hb981e18d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998e1ea),
	.w1(32'hb8b3bf1e),
	.w2(32'hb9c10876),
	.w3(32'h3802ac25),
	.w4(32'h393940a4),
	.w5(32'hb9501efb),
	.w6(32'h38f4ee3a),
	.w7(32'h39b6df75),
	.w8(32'hb85591a0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef013a),
	.w1(32'hb7cdbc5b),
	.w2(32'hb958c339),
	.w3(32'h3933f690),
	.w4(32'h39670e11),
	.w5(32'h37c4a36f),
	.w6(32'h3958a97a),
	.w7(32'h39876772),
	.w8(32'h38d4ac61),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c4493),
	.w1(32'hb752bb45),
	.w2(32'hb875955e),
	.w3(32'h37b6e9c0),
	.w4(32'h38345e01),
	.w5(32'hb808dcc1),
	.w6(32'h38044249),
	.w7(32'h381de680),
	.w8(32'hb6c6876a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3739c6b9),
	.w1(32'h377e9351),
	.w2(32'h35a91242),
	.w3(32'h36c41095),
	.w4(32'h370e2682),
	.w5(32'hb6973ba4),
	.w6(32'h36f25a93),
	.w7(32'h36b5a912),
	.w8(32'h35f76132),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f0465),
	.w1(32'hb6eeeaa1),
	.w2(32'hb6d76de2),
	.w3(32'hb791c71f),
	.w4(32'hb73ed2f1),
	.w5(32'hb7c9b35a),
	.w6(32'hb74cfa10),
	.w7(32'hb759236c),
	.w8(32'hb82269ae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c758a9),
	.w1(32'hb815a04b),
	.w2(32'hb77c3c59),
	.w3(32'hb7a88795),
	.w4(32'hb81ba207),
	.w5(32'hb8089065),
	.w6(32'hb752cffd),
	.w7(32'hb77c0f05),
	.w8(32'hb73ecede),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fee47),
	.w1(32'hb9a26f97),
	.w2(32'hb93e6ecd),
	.w3(32'hb93892a6),
	.w4(32'hb90bd921),
	.w5(32'h37924670),
	.w6(32'hb972aece),
	.w7(32'hb9321933),
	.w8(32'hb872d333),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9945eb2),
	.w1(32'hb99fb241),
	.w2(32'hb944c49f),
	.w3(32'hb89720c1),
	.w4(32'hb906061c),
	.w5(32'hb8426336),
	.w6(32'hb87a659d),
	.w7(32'hb892affe),
	.w8(32'hb804fd16),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d81896),
	.w1(32'hb9b92b97),
	.w2(32'hb999a5ab),
	.w3(32'hb97341ed),
	.w4(32'hb914201d),
	.w5(32'hb8d2d292),
	.w6(32'hb92792b9),
	.w7(32'hb8fbffbd),
	.w8(32'hb9205846),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d4a62),
	.w1(32'hb91cf594),
	.w2(32'hb939ea5c),
	.w3(32'hb907cfd2),
	.w4(32'h3803d5c0),
	.w5(32'hb8a79e32),
	.w6(32'hb8ca8841),
	.w7(32'hb942f214),
	.w8(32'hb97fa2a1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87230ab),
	.w1(32'hb810612c),
	.w2(32'hb96a7491),
	.w3(32'hb8a85b27),
	.w4(32'h37825a93),
	.w5(32'hb7e30787),
	.w6(32'hb9fb1c85),
	.w7(32'hb9ec4c48),
	.w8(32'hb98552c9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3574d2c2),
	.w1(32'h36ac50fc),
	.w2(32'h373b5d71),
	.w3(32'hb766e0d1),
	.w4(32'hb7acc4fc),
	.w5(32'h355af978),
	.w6(32'hb709fdd3),
	.w7(32'hb7b299ed),
	.w8(32'h36c0bb06),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb699e628),
	.w1(32'h35f7aea3),
	.w2(32'h37927d44),
	.w3(32'hb7528230),
	.w4(32'h37bab065),
	.w5(32'h375eec5c),
	.w6(32'hb6618a56),
	.w7(32'h37c7c16f),
	.w8(32'h37faca79),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a382ef),
	.w1(32'hb656860d),
	.w2(32'h37ab4d42),
	.w3(32'hb78bbb84),
	.w4(32'hb6aea48f),
	.w5(32'h37ac0cf3),
	.w6(32'h37522eeb),
	.w7(32'hb61e2465),
	.w8(32'h377dead4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef578),
	.w1(32'hb918220b),
	.w2(32'hb91edd2b),
	.w3(32'hb800513f),
	.w4(32'hb719ad93),
	.w5(32'hb7fb4861),
	.w6(32'hb88bad9d),
	.w7(32'hb896369a),
	.w8(32'hb89e313b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8249433),
	.w1(32'hb79bca35),
	.w2(32'hb83d2408),
	.w3(32'hb79eb833),
	.w4(32'h379e81cc),
	.w5(32'hb7b3bcd9),
	.w6(32'hb8084400),
	.w7(32'hb83621c7),
	.w8(32'hb88fc966),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938ada2),
	.w1(32'hb92f5ec6),
	.w2(32'hb98932de),
	.w3(32'hb9234524),
	.w4(32'hb7eb5042),
	.w5(32'h32a513f9),
	.w6(32'hb9c3d96a),
	.w7(32'hb9a103e1),
	.w8(32'hb9912ca7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37690245),
	.w1(32'h366ddd64),
	.w2(32'h367b47d3),
	.w3(32'h381c8c13),
	.w4(32'h381daebd),
	.w5(32'hb7b6a8ef),
	.w6(32'hb83eb046),
	.w7(32'hb822710f),
	.w8(32'hb8d5c6b5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ab0394),
	.w1(32'hb588796c),
	.w2(32'hb662b1c9),
	.w3(32'hb6745ae9),
	.w4(32'hb5e5df01),
	.w5(32'hb6b6d65f),
	.w6(32'hb6580b7a),
	.w7(32'h32e80425),
	.w8(32'hb63a7f52),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fb4b05),
	.w1(32'hb412e5b9),
	.w2(32'hb44dc4c9),
	.w3(32'hb595dfca),
	.w4(32'hb52dc268),
	.w5(32'hb5b77f3e),
	.w6(32'h33c6b783),
	.w7(32'hb4e96097),
	.w8(32'hb578e5af),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4c435ff),
	.w1(32'hb68c12a2),
	.w2(32'hb636c85d),
	.w3(32'hb566a4ad),
	.w4(32'hb6608fa8),
	.w5(32'h352800aa),
	.w6(32'hb465ffe4),
	.w7(32'hb6a0c904),
	.w8(32'hb493e5d0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3c293),
	.w1(32'hb73099b7),
	.w2(32'h36b2b36a),
	.w3(32'h3702009e),
	.w4(32'hb6763a11),
	.w5(32'h36adb441),
	.w6(32'h370c0daf),
	.w7(32'h3694bc0b),
	.w8(32'h3704d64f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5c8af),
	.w1(32'hb67f868d),
	.w2(32'hb689396e),
	.w3(32'hb69c8fea),
	.w4(32'hb75919a6),
	.w5(32'hb701b667),
	.w6(32'hb6e74be0),
	.w7(32'hb7696a46),
	.w8(32'hb68b3dfc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8442a5a),
	.w1(32'hb853747f),
	.w2(32'hb84058cf),
	.w3(32'hb8556d64),
	.w4(32'h37da8d84),
	.w5(32'h37f27b2c),
	.w6(32'hb8c60ceb),
	.w7(32'hb905b3d7),
	.w8(32'hb830d9a9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386098ef),
	.w1(32'hb7ee0cbe),
	.w2(32'h381e3dc1),
	.w3(32'h38272c9b),
	.w4(32'h38d846c1),
	.w5(32'h386be6a4),
	.w6(32'h366128c2),
	.w7(32'hb80ba0a5),
	.w8(32'hb870e810),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57ac844),
	.w1(32'h363d4244),
	.w2(32'h3676a179),
	.w3(32'hb6b67440),
	.w4(32'h359924f0),
	.w5(32'h36998f4f),
	.w6(32'hb7112745),
	.w7(32'hb614fa65),
	.w8(32'h3681b783),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350e42f7),
	.w1(32'h352794ab),
	.w2(32'h34252b65),
	.w3(32'h357cd65d),
	.w4(32'hb5d4e0f5),
	.w5(32'hb6032360),
	.w6(32'hb453b6ca),
	.w7(32'hb4feb710),
	.w8(32'hb602446e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3680732c),
	.w1(32'hb6eeee2b),
	.w2(32'hb5daeb4f),
	.w3(32'h35ccc962),
	.w4(32'hb6d4c8c0),
	.w5(32'hb573e18d),
	.w6(32'h350568a7),
	.w7(32'hb6b9e9b9),
	.w8(32'h3586b368),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b02100),
	.w1(32'h366b049e),
	.w2(32'h35a44d6d),
	.w3(32'h361d773b),
	.w4(32'h3668658d),
	.w5(32'h34e73d94),
	.w6(32'h3674276e),
	.w7(32'h353cb507),
	.w8(32'hb56d9eb5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb864b0cf),
	.w1(32'hb780a150),
	.w2(32'hb76d56d0),
	.w3(32'h378fe467),
	.w4(32'h3846ff37),
	.w5(32'h38f3d434),
	.w6(32'hb9163360),
	.w7(32'hb8c1f6e2),
	.w8(32'hb884ea4b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998273b),
	.w1(32'hb9a4a53a),
	.w2(32'hb83bb2b0),
	.w3(32'hb8a172a4),
	.w4(32'hb911be15),
	.w5(32'hb73c4736),
	.w6(32'hb8bd74c1),
	.w7(32'hb9654bd8),
	.w8(32'hb89a50e5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882bac7),
	.w1(32'hb96e263f),
	.w2(32'hb8c9dbf5),
	.w3(32'hb82710c5),
	.w4(32'h37f4a367),
	.w5(32'h376d47e3),
	.w6(32'hb9b0d8c2),
	.w7(32'hb9e063c4),
	.w8(32'hb9f7d8d5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e2a8d),
	.w1(32'hb995da1e),
	.w2(32'hba72b0f9),
	.w3(32'hb8a35e78),
	.w4(32'hba4a31ab),
	.w5(32'hbb26f9b6),
	.w6(32'hb84ceeaa),
	.w7(32'hbb072d9b),
	.w8(32'hbb9472d1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04d557),
	.w1(32'hbaa44367),
	.w2(32'hb9e50bc4),
	.w3(32'hbaf6f1f8),
	.w4(32'hba8a8da9),
	.w5(32'hb9b85a03),
	.w6(32'hbaf19c49),
	.w7(32'hba638a90),
	.w8(32'hba8df324),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0fcf),
	.w1(32'hb9fad152),
	.w2(32'hb918a69b),
	.w3(32'hbad824cc),
	.w4(32'hbb022c67),
	.w5(32'hba32d8fa),
	.w6(32'hba0e2790),
	.w7(32'hb961e658),
	.w8(32'hb998e73b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1b105),
	.w1(32'h3a675ac3),
	.w2(32'h3920a284),
	.w3(32'h3823acaa),
	.w4(32'h3a858813),
	.w5(32'h3a23a19a),
	.w6(32'h3a825665),
	.w7(32'h3ad2364e),
	.w8(32'hb968782c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bacc7f),
	.w1(32'h3a85c7e9),
	.w2(32'h3915140a),
	.w3(32'h3820ced0),
	.w4(32'h38d2f10c),
	.w5(32'hba23e1af),
	.w6(32'h3a80978d),
	.w7(32'hb957acd8),
	.w8(32'hba020627),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927377d),
	.w1(32'hbb3a72ac),
	.w2(32'hba95f95c),
	.w3(32'h393c34e3),
	.w4(32'hbb459bcb),
	.w5(32'hbaa40366),
	.w6(32'hba8e6394),
	.w7(32'hba95bf7c),
	.w8(32'hba323d2b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac36cf1),
	.w1(32'h3aa9fb7e),
	.w2(32'h38f6d6a1),
	.w3(32'hbac7b0c6),
	.w4(32'hba105fdc),
	.w5(32'hb9a732f1),
	.w6(32'hbb0896ac),
	.w7(32'hba362a22),
	.w8(32'hba9e2d83),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e8a5c),
	.w1(32'h3a72b4bd),
	.w2(32'hba160b02),
	.w3(32'hb7e1068d),
	.w4(32'h3a557ba0),
	.w5(32'hba0552ea),
	.w6(32'hba5a39d5),
	.w7(32'hba9c1258),
	.w8(32'hbb100c68),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18848b),
	.w1(32'hb96e03e5),
	.w2(32'hb9c0ffda),
	.w3(32'h38dc126d),
	.w4(32'hb995b749),
	.w5(32'hba7631b3),
	.w6(32'hbb1c5256),
	.w7(32'h384a246b),
	.w8(32'hb818c8c1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f73b),
	.w1(32'hb9201351),
	.w2(32'hba120cf8),
	.w3(32'hba8bcac6),
	.w4(32'hba33831a),
	.w5(32'h399f4d45),
	.w6(32'h3950cdd9),
	.w7(32'hb9275c7f),
	.w8(32'h3ae7e6bf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030ef1),
	.w1(32'hb983534b),
	.w2(32'hbabac94f),
	.w3(32'hb9ff6b19),
	.w4(32'hba88704a),
	.w5(32'hbb1d215b),
	.w6(32'h3abe29db),
	.w7(32'h39c4de2f),
	.w8(32'hba9da1e3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94703c),
	.w1(32'h3aa48cd9),
	.w2(32'h3afb4c04),
	.w3(32'hba55c4d3),
	.w4(32'h3b281514),
	.w5(32'h3b8a539f),
	.w6(32'hbaad9190),
	.w7(32'h3a9f2aca),
	.w8(32'h3b4d8507),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a73a0),
	.w1(32'h3a5f3a23),
	.w2(32'hb8fcf03f),
	.w3(32'h3b4a09ff),
	.w4(32'h3a481cd1),
	.w5(32'hb903ef1e),
	.w6(32'h3b11643b),
	.w7(32'h3ae15f12),
	.w8(32'h39ac56d2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39738684),
	.w1(32'h3a4307ef),
	.w2(32'h387ad8a6),
	.w3(32'h394ef5a3),
	.w4(32'h39fc3649),
	.w5(32'hb9e7a666),
	.w6(32'hb91bb2ff),
	.w7(32'h3b4a94a1),
	.w8(32'h3ac4a610),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8003452),
	.w1(32'h3b2b2ff3),
	.w2(32'h3b33783b),
	.w3(32'h3aac7dff),
	.w4(32'h3af4fdaa),
	.w5(32'h3b38f551),
	.w6(32'h3a9c83bd),
	.w7(32'h3a948e2c),
	.w8(32'h3abb1dc3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa4f5),
	.w1(32'hba0109d4),
	.w2(32'hba273a58),
	.w3(32'h3b23df14),
	.w4(32'h3a91e364),
	.w5(32'h399acfeb),
	.w6(32'h3b0f916d),
	.w7(32'h3ac66bfd),
	.w8(32'h390b6267),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4dd6),
	.w1(32'hbacb208f),
	.w2(32'hbb2880d1),
	.w3(32'hb9cab943),
	.w4(32'hbb2370f3),
	.w5(32'hbb143554),
	.w6(32'h3a256726),
	.w7(32'hba9d0dfa),
	.w8(32'hbaafce4b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e42847),
	.w1(32'hb98f1ba5),
	.w2(32'hba5aef4a),
	.w3(32'hba0c2c1b),
	.w4(32'hb926cc35),
	.w5(32'hba67a496),
	.w6(32'hba333961),
	.w7(32'hba45aa02),
	.w8(32'hba7dd0dc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9932f5),
	.w1(32'h39c47f48),
	.w2(32'hb9d7d708),
	.w3(32'hba9d5099),
	.w4(32'hbaaa907a),
	.w5(32'hbb6a3de2),
	.w6(32'hba9551d7),
	.w7(32'h39b48475),
	.w8(32'h3a51da25),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbb9df),
	.w1(32'hbaf99f63),
	.w2(32'h38db2e03),
	.w3(32'hba8cbe40),
	.w4(32'h39bb28ce),
	.w5(32'h39d46764),
	.w6(32'hb9ccb6b4),
	.w7(32'hbb44ac00),
	.w8(32'hb9de9c92),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8afd86),
	.w1(32'h3ab620f5),
	.w2(32'hb9fe3101),
	.w3(32'hb98d636d),
	.w4(32'h3b261693),
	.w5(32'h39faba18),
	.w6(32'hbb3e7ef7),
	.w7(32'hba8aa130),
	.w8(32'hb991c7c6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f0150),
	.w1(32'hba8b0ed4),
	.w2(32'hb953243f),
	.w3(32'hbaf023ae),
	.w4(32'hb979b52e),
	.w5(32'hba86d73a),
	.w6(32'hba3536da),
	.w7(32'hb9ca7d07),
	.w8(32'hbab94d0e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9908959),
	.w1(32'hba6df781),
	.w2(32'hb97f3ea3),
	.w3(32'hbab12a12),
	.w4(32'hbab0e43a),
	.w5(32'h3a4d937b),
	.w6(32'hbaab9f3b),
	.w7(32'hbb58b5f6),
	.w8(32'hb97ef795),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab550f),
	.w1(32'h3a4ed42c),
	.w2(32'h3aaf601d),
	.w3(32'hba1d9126),
	.w4(32'h3a43a281),
	.w5(32'h38233cbf),
	.w6(32'hbaf22cb3),
	.w7(32'h3ac555e3),
	.w8(32'h3ab0db5d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e54237),
	.w1(32'h3a725676),
	.w2(32'h3a191697),
	.w3(32'h3ae2f48a),
	.w4(32'h3941c7c9),
	.w5(32'h39b21e1b),
	.w6(32'h3abfe7ea),
	.w7(32'hbaab78fc),
	.w8(32'hba8b0c76),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f75ff8),
	.w1(32'hbaf39c50),
	.w2(32'hba55d0b2),
	.w3(32'h3abd1832),
	.w4(32'hba68e68c),
	.w5(32'h3aa1f71f),
	.w6(32'hba1ab79b),
	.w7(32'hbab202b4),
	.w8(32'h3927bcb9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb214b),
	.w1(32'hbaa916d2),
	.w2(32'hba87a002),
	.w3(32'h3a4b11e9),
	.w4(32'h3a653e25),
	.w5(32'hb986fd3a),
	.w6(32'hbb1880ef),
	.w7(32'h3a3c7b59),
	.w8(32'hbb06d2c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5338fa),
	.w1(32'hb9452d4a),
	.w2(32'hb905b15f),
	.w3(32'h39f6c060),
	.w4(32'hba8c8510),
	.w5(32'hba807bfd),
	.w6(32'h385b47d2),
	.w7(32'hb967183a),
	.w8(32'h3a1968b0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899b74b),
	.w1(32'h3a916b63),
	.w2(32'h3a3a43b8),
	.w3(32'hba32590d),
	.w4(32'h3a326403),
	.w5(32'hb9314236),
	.w6(32'hb6c0eb2e),
	.w7(32'h3aa80d33),
	.w8(32'h38929e7a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad22a9a),
	.w1(32'hb9a23f37),
	.w2(32'hba62c8eb),
	.w3(32'h3a0856d2),
	.w4(32'hba0454e7),
	.w5(32'hbac4b29d),
	.w6(32'h3a684e04),
	.w7(32'hbae2f311),
	.w8(32'hbada910f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13cc6f),
	.w1(32'hba6d3467),
	.w2(32'hbac54b1a),
	.w3(32'hbb1f1c2c),
	.w4(32'hba08654e),
	.w5(32'h3967d320),
	.w6(32'hbb28868d),
	.w7(32'hbac139b7),
	.w8(32'h3a118b11),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad2936),
	.w1(32'h39ce1b4f),
	.w2(32'h3a066706),
	.w3(32'hbac5c39d),
	.w4(32'hb91f447e),
	.w5(32'hb96f9178),
	.w6(32'hba884fbf),
	.w7(32'hba94bdc9),
	.w8(32'hb96eb3ac),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b32970),
	.w1(32'hbaa96413),
	.w2(32'hba4e8e0b),
	.w3(32'h39b3f17e),
	.w4(32'h3a42227c),
	.w5(32'hba4d477f),
	.w6(32'hbab75b8f),
	.w7(32'h3912a652),
	.w8(32'hbb027870),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba510491),
	.w1(32'h3aa2662d),
	.w2(32'h39f1b5e6),
	.w3(32'hb8944b7e),
	.w4(32'hba419490),
	.w5(32'hbb4b1273),
	.w6(32'h38e8febc),
	.w7(32'hba23f5bc),
	.w8(32'h391e72f5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb4650),
	.w1(32'hba13d9c0),
	.w2(32'hbacde68b),
	.w3(32'hbad93244),
	.w4(32'hb9d1742c),
	.w5(32'hb9e36796),
	.w6(32'h3999bc97),
	.w7(32'h39506f16),
	.w8(32'h3aa91b12),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00910e),
	.w1(32'h3a4a34b1),
	.w2(32'h3a79e269),
	.w3(32'hbae22fa0),
	.w4(32'h3af7209b),
	.w5(32'h3ae1cbc6),
	.w6(32'h36a945b1),
	.w7(32'h3a5343ea),
	.w8(32'h3ad35b04),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b9d3f),
	.w1(32'hb9dfbd47),
	.w2(32'hba6e0d9f),
	.w3(32'h3b095233),
	.w4(32'h3934eaf4),
	.w5(32'hba3983c9),
	.w6(32'h3a89defa),
	.w7(32'h3ae6e0bb),
	.w8(32'h3a537716),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9b500),
	.w1(32'h38809ff1),
	.w2(32'hba908bd6),
	.w3(32'h395f7e71),
	.w4(32'h3a10e2b8),
	.w5(32'hb8ec3967),
	.w6(32'h3a811467),
	.w7(32'h398ebda1),
	.w8(32'hba330f88),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed9bd2),
	.w1(32'hbac32d4a),
	.w2(32'hb928b448),
	.w3(32'h3a6e4709),
	.w4(32'hb9b2bf8d),
	.w5(32'hb9ad93d1),
	.w6(32'hb9cbe11c),
	.w7(32'hb9949adc),
	.w8(32'hbabaff35),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382e9e89),
	.w1(32'hb89528fe),
	.w2(32'h39847129),
	.w3(32'hbae88274),
	.w4(32'hb96e6510),
	.w5(32'hbaa28256),
	.w6(32'hbaa73934),
	.w7(32'hba906e47),
	.w8(32'hb9b0d5ef),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eadc50),
	.w1(32'hb9eccc6f),
	.w2(32'h3ab9619d),
	.w3(32'h39236b39),
	.w4(32'h39496558),
	.w5(32'hba0d875c),
	.w6(32'h391573ad),
	.w7(32'hb9f54618),
	.w8(32'hba99b02a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0812ca),
	.w1(32'hb9ca981b),
	.w2(32'hba9c0964),
	.w3(32'h3b00960b),
	.w4(32'hba98d38a),
	.w5(32'h3a2fcf11),
	.w6(32'h39f3dcf3),
	.w7(32'hba96f6e2),
	.w8(32'hba289bbc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ec9d3),
	.w1(32'hb81b7837),
	.w2(32'h3884c192),
	.w3(32'hb9b08b0c),
	.w4(32'hba66e2b7),
	.w5(32'hb9a02c72),
	.w6(32'h39d44fb5),
	.w7(32'hba70253f),
	.w8(32'hb98a4a7b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d51de),
	.w1(32'hba8b6ada),
	.w2(32'hbb0e3f50),
	.w3(32'hb9352d39),
	.w4(32'hb60c7b1b),
	.w5(32'hb9a3f4c9),
	.w6(32'hb85f977f),
	.w7(32'hb97036e0),
	.w8(32'hb9618d25),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9720c),
	.w1(32'hb9dad02e),
	.w2(32'hb9cd680a),
	.w3(32'hbb01e676),
	.w4(32'hba54a2dc),
	.w5(32'hbb269d9d),
	.w6(32'hbac514b8),
	.w7(32'hba8cbb49),
	.w8(32'hbb4752c5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab1111),
	.w1(32'h39874d21),
	.w2(32'hb9a7e9e8),
	.w3(32'h3a87115b),
	.w4(32'hb8db451d),
	.w5(32'h381461f8),
	.w6(32'hbadc1301),
	.w7(32'hb9a5ffa3),
	.w8(32'hb9b3160b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f00f0),
	.w1(32'hbab2f277),
	.w2(32'hb9e48fdf),
	.w3(32'hb8dc1cfb),
	.w4(32'hba5ddaed),
	.w5(32'hb9bea641),
	.w6(32'hb991b72e),
	.w7(32'h3a31333c),
	.w8(32'hba673542),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1a477),
	.w1(32'h3a59199d),
	.w2(32'h3a743b1a),
	.w3(32'h3a187e45),
	.w4(32'h3a1d597c),
	.w5(32'h3adb7112),
	.w6(32'h3a3a5453),
	.w7(32'h3af0698f),
	.w8(32'h3a0fe938),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a5ba),
	.w1(32'h3aec9431),
	.w2(32'hb9bc255c),
	.w3(32'hb9c15b42),
	.w4(32'h3a61be1a),
	.w5(32'hb9073aae),
	.w6(32'h387ae373),
	.w7(32'hbac214fb),
	.w8(32'hba87ab8f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3c469),
	.w1(32'h3ae3dc57),
	.w2(32'h3a53d552),
	.w3(32'h3af044ad),
	.w4(32'h3a519c0e),
	.w5(32'hbaf02213),
	.w6(32'hba513cb6),
	.w7(32'hb945e5cf),
	.w8(32'h3a1f6a40),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56bb0e),
	.w1(32'hba637a08),
	.w2(32'hba702e6e),
	.w3(32'h39e0e4be),
	.w4(32'hbad8cff7),
	.w5(32'h3ad02a16),
	.w6(32'h396319e7),
	.w7(32'hba7206a3),
	.w8(32'h3a11f17d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a6b2),
	.w1(32'hba332dcc),
	.w2(32'h39257444),
	.w3(32'hb8c2eaab),
	.w4(32'hba4f70de),
	.w5(32'hb9c5051c),
	.w6(32'h398ed695),
	.w7(32'hb9e44a62),
	.w8(32'hba1c9db4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcd445),
	.w1(32'h3908cb0a),
	.w2(32'h3a84a9ad),
	.w3(32'h3a6b189f),
	.w4(32'hba4e9999),
	.w5(32'hb9b6e74c),
	.w6(32'hbad14357),
	.w7(32'hbb4b8f9e),
	.w8(32'hbb0e2465),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d7143),
	.w1(32'hbaa7179c),
	.w2(32'hbabcd2af),
	.w3(32'hbab1dceb),
	.w4(32'hbaa343e0),
	.w5(32'hba09d8f8),
	.w6(32'hbb121857),
	.w7(32'hb95668e7),
	.w8(32'h3a4bd6b8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba374d32),
	.w1(32'hbb13220c),
	.w2(32'hba379087),
	.w3(32'hbad9746d),
	.w4(32'hb9967847),
	.w5(32'h3b02d038),
	.w6(32'hb9605dfc),
	.w7(32'hb8f32a46),
	.w8(32'h3a6d5824),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67fa91),
	.w1(32'hb921fcd4),
	.w2(32'h375277b7),
	.w3(32'h3a1aaa8d),
	.w4(32'hba9945f6),
	.w5(32'hbad2b8bb),
	.w6(32'hb96d13c0),
	.w7(32'hbaf7d682),
	.w8(32'hbb1c9ee4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa54b68),
	.w1(32'h39e414b6),
	.w2(32'hba487e9a),
	.w3(32'hba496c97),
	.w4(32'hbac5fa5e),
	.w5(32'hbb3cbbe1),
	.w6(32'hbb09753f),
	.w7(32'hbb1847c2),
	.w8(32'hbb1cc348),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9f173),
	.w1(32'h39cb2fb3),
	.w2(32'hbadb01ff),
	.w3(32'hba55ffb3),
	.w4(32'hba68e5f5),
	.w5(32'hbb55a4a5),
	.w6(32'hbaa1483a),
	.w7(32'hbb053219),
	.w8(32'hbb14c3d0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15a5c6),
	.w1(32'h3a137d27),
	.w2(32'hba024954),
	.w3(32'hbb93e0a1),
	.w4(32'h392ef6b5),
	.w5(32'h39ff3ff5),
	.w6(32'hbb37a6f7),
	.w7(32'hb951bc31),
	.w8(32'hba4c0cf9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884f235),
	.w1(32'hbb01dc75),
	.w2(32'hbabc4a36),
	.w3(32'h3ac84881),
	.w4(32'hba7484e3),
	.w5(32'hba1d2a98),
	.w6(32'h399dd03b),
	.w7(32'hbb039772),
	.w8(32'hba6320ed),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7f4be),
	.w1(32'hb7d804bd),
	.w2(32'hba2fd990),
	.w3(32'hba8400b8),
	.w4(32'hba9e2b72),
	.w5(32'h3a169d74),
	.w6(32'hb9f29f06),
	.w7(32'hba40ce3f),
	.w8(32'hb9c83786),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fd0ab),
	.w1(32'h3b33dabf),
	.w2(32'h3a9a2b63),
	.w3(32'hba3eb3c8),
	.w4(32'h3a98794c),
	.w5(32'hba2ba18e),
	.w6(32'h388ca423),
	.w7(32'hb9e63241),
	.w8(32'h35cae32a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8076f6d),
	.w1(32'hb9a5f4ac),
	.w2(32'hbab0c40e),
	.w3(32'h39a7973a),
	.w4(32'hbae178e7),
	.w5(32'hbad76386),
	.w6(32'h3823673b),
	.w7(32'hbab2c411),
	.w8(32'hbb0419fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002094),
	.w1(32'hbaadd50d),
	.w2(32'hba543368),
	.w3(32'hba991fe7),
	.w4(32'hb9687db3),
	.w5(32'hb8f72805),
	.w6(32'hbaa948db),
	.w7(32'hba49987c),
	.w8(32'hba0f7b83),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e698d),
	.w1(32'h39e09cc4),
	.w2(32'h3985eb66),
	.w3(32'hb93904b1),
	.w4(32'h3a96fc0e),
	.w5(32'h3b20834c),
	.w6(32'hb9a02631),
	.w7(32'h398117ee),
	.w8(32'hb9ac741f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41ce8a),
	.w1(32'h3a741270),
	.w2(32'hba009b0b),
	.w3(32'h39b5d43d),
	.w4(32'h39b64e5d),
	.w5(32'hb9201113),
	.w6(32'hba80c907),
	.w7(32'hb9e77e6b),
	.w8(32'h3a8f54d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4f3c7),
	.w1(32'h3b37c086),
	.w2(32'h3ad306e7),
	.w3(32'hb8102366),
	.w4(32'h3a8f908e),
	.w5(32'h39c57f80),
	.w6(32'h3abbc769),
	.w7(32'hba0fd44e),
	.w8(32'hba0ef855),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ffdd5),
	.w1(32'hba49855e),
	.w2(32'hbaff3f86),
	.w3(32'h396803f1),
	.w4(32'hbaa6a22b),
	.w5(32'hb9e27d51),
	.w6(32'hba81addc),
	.w7(32'hba3dccca),
	.w8(32'h39783cc4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77c5b5),
	.w1(32'h3aab3b79),
	.w2(32'h3a2c91c7),
	.w3(32'hba97830e),
	.w4(32'h399cf34a),
	.w5(32'hba0a8a86),
	.w6(32'hba28d82f),
	.w7(32'hbaa7ace0),
	.w8(32'hba5aecb9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935d630),
	.w1(32'hb9d140e9),
	.w2(32'h39168980),
	.w3(32'hba89a94f),
	.w4(32'h3a417036),
	.w5(32'h3a8caf9f),
	.w6(32'hba71429b),
	.w7(32'h3b330f93),
	.w8(32'h3b01e282),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935a83c),
	.w1(32'hb9bb5542),
	.w2(32'hb9efe287),
	.w3(32'h391da268),
	.w4(32'h39e2080e),
	.w5(32'h3745bef8),
	.w6(32'h3abd6fed),
	.w7(32'h39ff6b85),
	.w8(32'hb928ad35),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8b04c),
	.w1(32'hb99bb76c),
	.w2(32'hba2c2339),
	.w3(32'hb84d7bcc),
	.w4(32'h37c2ba3a),
	.w5(32'hba3c266e),
	.w6(32'hba172213),
	.w7(32'h3a82d27e),
	.w8(32'hbab9e757),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977b3fc),
	.w1(32'hba2ea3f9),
	.w2(32'h3a29f103),
	.w3(32'h3a3acbf6),
	.w4(32'hb9e6e787),
	.w5(32'hba2381f4),
	.w6(32'hba36a89e),
	.w7(32'h39b41a3d),
	.w8(32'h3a4d8c36),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a554aa5),
	.w1(32'hb9ef5a8a),
	.w2(32'hb9b53e6e),
	.w3(32'h3a8596d3),
	.w4(32'hb9c1069f),
	.w5(32'hba0bdef3),
	.w6(32'h3ad7a4ec),
	.w7(32'hba1a3eea),
	.w8(32'hbb1a5388),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67da4),
	.w1(32'hb739d771),
	.w2(32'h39d00942),
	.w3(32'hba541b2a),
	.w4(32'hba5442e5),
	.w5(32'hb9ba0ef9),
	.w6(32'hba70a998),
	.w7(32'hba863eee),
	.w8(32'hbb0b19fe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3bb8f),
	.w1(32'hba0c8aac),
	.w2(32'hba4fb6b8),
	.w3(32'h3a30926d),
	.w4(32'hbab354f6),
	.w5(32'hbb073cec),
	.w6(32'h3a1658c3),
	.w7(32'hba799c2c),
	.w8(32'hbaa552dd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d2780),
	.w1(32'h3921a95f),
	.w2(32'h3a6bc186),
	.w3(32'hbb44c408),
	.w4(32'h3ae71f11),
	.w5(32'h3b0bcec0),
	.w6(32'hba91f21f),
	.w7(32'h393312a6),
	.w8(32'h3928b54a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa86830),
	.w1(32'h39ef9bcc),
	.w2(32'h3a8338ea),
	.w3(32'h3a86abcb),
	.w4(32'h3aa6142c),
	.w5(32'h3b08dab4),
	.w6(32'hb8acadb9),
	.w7(32'h3a117981),
	.w8(32'h3a909b10),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88da09b),
	.w1(32'hba6396b1),
	.w2(32'hbb030e66),
	.w3(32'h3a18554b),
	.w4(32'hba84653d),
	.w5(32'hbb15299f),
	.w6(32'h39f0d1a8),
	.w7(32'h3aba3e70),
	.w8(32'hb6b03bc2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d121),
	.w1(32'hb91dbf37),
	.w2(32'hb9fdaec2),
	.w3(32'hba778c1f),
	.w4(32'h39526982),
	.w5(32'hb928f259),
	.w6(32'hba83d898),
	.w7(32'h3999439d),
	.w8(32'h3a334a6e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5959e1),
	.w1(32'h3958ccb1),
	.w2(32'hb9ff1a70),
	.w3(32'h39db01a8),
	.w4(32'h39ad5ef1),
	.w5(32'hba859c75),
	.w6(32'hba6d34be),
	.w7(32'h3a48a039),
	.w8(32'hbaa24c9a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8648a4),
	.w1(32'hb98963e4),
	.w2(32'hb9f0374f),
	.w3(32'h3a194921),
	.w4(32'hba64d61d),
	.w5(32'h3ab5563b),
	.w6(32'hb984a06e),
	.w7(32'hbaa9e6fa),
	.w8(32'hbac43389),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fc3a2),
	.w1(32'hba93132e),
	.w2(32'hbb1c6d70),
	.w3(32'hba8e4841),
	.w4(32'hb92290e5),
	.w5(32'hbaf06db4),
	.w6(32'hb9a2d298),
	.w7(32'hbb1aa79e),
	.w8(32'hbb5bbca6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e22b3),
	.w1(32'h3aa545d9),
	.w2(32'h3a9ab01b),
	.w3(32'h3a8c69e5),
	.w4(32'h3ad52779),
	.w5(32'h3a753af1),
	.w6(32'hba95b6bd),
	.w7(32'h3a1c5bd3),
	.w8(32'hbabfdb99),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca0128),
	.w1(32'hba1146da),
	.w2(32'h3a3e1c81),
	.w3(32'hbaafdbf5),
	.w4(32'hb63d3a6c),
	.w5(32'h39e7ad99),
	.w6(32'hb8b898c4),
	.w7(32'hbb3468a2),
	.w8(32'hbb47a4e3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de0031),
	.w1(32'h3a6edccb),
	.w2(32'hba723f2e),
	.w3(32'hba2e5cf5),
	.w4(32'hba1de179),
	.w5(32'h393c6a61),
	.w6(32'hbb8c9445),
	.w7(32'hb952b257),
	.w8(32'hba87760b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b4e243),
	.w1(32'h39971b73),
	.w2(32'h3a336694),
	.w3(32'hb915b5b5),
	.w4(32'h3a062484),
	.w5(32'h3988ba7b),
	.w6(32'hba38a1f5),
	.w7(32'h3a62cbc0),
	.w8(32'h395abb78),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a42f7a),
	.w1(32'hba34f803),
	.w2(32'hb9f7c867),
	.w3(32'hba0a9dd2),
	.w4(32'hbb0cbab2),
	.w5(32'h3a1a49be),
	.w6(32'h39e3f434),
	.w7(32'hbb1d5709),
	.w8(32'hba5b5bfe),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab07405),
	.w1(32'h3891f4a6),
	.w2(32'hba710924),
	.w3(32'hba93357a),
	.w4(32'h39eae0ad),
	.w5(32'hba2aa9d7),
	.w6(32'h3a932a17),
	.w7(32'h3a70aee4),
	.w8(32'h3a68a361),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a64ea0),
	.w1(32'hb9ca2413),
	.w2(32'h3a80b0c7),
	.w3(32'h39db480a),
	.w4(32'hb9bcf7ae),
	.w5(32'h3abf379a),
	.w6(32'h3a3b9c39),
	.w7(32'hbacce823),
	.w8(32'h39f02d07),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997641f),
	.w1(32'h3a076d4b),
	.w2(32'h3a180dfe),
	.w3(32'h3a364367),
	.w4(32'hb91ab61c),
	.w5(32'h3b0868f0),
	.w6(32'h3831e262),
	.w7(32'h3910dc19),
	.w8(32'h39ab234c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202ded),
	.w1(32'h3b1bc7ac),
	.w2(32'h3b49604f),
	.w3(32'h398f8037),
	.w4(32'h3a97c30d),
	.w5(32'hbaab8177),
	.w6(32'h3887b11a),
	.w7(32'h39928d73),
	.w8(32'h3b014a79),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e82c9),
	.w1(32'h3a38225c),
	.w2(32'hba3dab96),
	.w3(32'hba12236c),
	.w4(32'hb9922c12),
	.w5(32'hbb25c200),
	.w6(32'h3aa62917),
	.w7(32'h39e26661),
	.w8(32'h3a9149b0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85698a),
	.w1(32'h39ef1080),
	.w2(32'hba8824b5),
	.w3(32'hbab791d0),
	.w4(32'h3a86c8ba),
	.w5(32'hba9ca4dc),
	.w6(32'hb9705a29),
	.w7(32'h3b06e381),
	.w8(32'h3acdbd60),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc25de),
	.w1(32'h39316d1a),
	.w2(32'hba58c6a1),
	.w3(32'h3a87470e),
	.w4(32'hb9b312cb),
	.w5(32'hb92909b2),
	.w6(32'h3b562e20),
	.w7(32'hba1780ef),
	.w8(32'hb95e1d70),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb4ce4),
	.w1(32'h394bed7d),
	.w2(32'h3ab43f09),
	.w3(32'hba6d9122),
	.w4(32'hbac5b99a),
	.w5(32'h394522f2),
	.w6(32'hba57d8ea),
	.w7(32'h3a34e2f2),
	.w8(32'hb85a2e5f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac91906),
	.w1(32'h393f38f6),
	.w2(32'h39db26da),
	.w3(32'h3a8bf93a),
	.w4(32'h3a2342a3),
	.w5(32'h3b142db9),
	.w6(32'h390d80a8),
	.w7(32'h398d93ce),
	.w8(32'h3a0f923d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e12b1d),
	.w1(32'hbacac7b8),
	.w2(32'hb8ae1786),
	.w3(32'h3a40c53c),
	.w4(32'h3afedf05),
	.w5(32'h3affe98d),
	.w6(32'h3a705c9b),
	.w7(32'h3a1954f5),
	.w8(32'hba048a23),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b0a90),
	.w1(32'h38a0775c),
	.w2(32'h3a562fd8),
	.w3(32'h397da33f),
	.w4(32'hb61ee209),
	.w5(32'h3b12fa2e),
	.w6(32'h396ff183),
	.w7(32'hba272b15),
	.w8(32'hba07cb35),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acbe55),
	.w1(32'hbae15c49),
	.w2(32'h3a5892ab),
	.w3(32'hb9949df2),
	.w4(32'hbaba51d1),
	.w5(32'hba5b2a3d),
	.w6(32'hba72c1c4),
	.w7(32'hb9ca018c),
	.w8(32'hb93973dc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36ebae),
	.w1(32'h38b6ee86),
	.w2(32'hba519cf9),
	.w3(32'hba154db0),
	.w4(32'h39eac093),
	.w5(32'hba897519),
	.w6(32'hbae6b4f3),
	.w7(32'h3996479c),
	.w8(32'hba3673c3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6be210),
	.w1(32'hb9d0c456),
	.w2(32'hba899b68),
	.w3(32'hb9a98c6c),
	.w4(32'hb9ad38f9),
	.w5(32'h39b57366),
	.w6(32'h3a23e804),
	.w7(32'hba1cbe4f),
	.w8(32'hbadcbcdc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06cdf3),
	.w1(32'hb9c4a80c),
	.w2(32'h3a570c6a),
	.w3(32'hba8b7611),
	.w4(32'h38db642c),
	.w5(32'h39a71e3f),
	.w6(32'hb99ef39c),
	.w7(32'h37dd9088),
	.w8(32'hb9efdf2d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d76cc),
	.w1(32'hb97023ba),
	.w2(32'hb923a83d),
	.w3(32'hba03f110),
	.w4(32'h386cc1dd),
	.w5(32'h39dfa6d5),
	.w6(32'h39cca274),
	.w7(32'h39d853ae),
	.w8(32'h3a371f31),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380bd8b1),
	.w1(32'hba5826bd),
	.w2(32'hb7fe5e20),
	.w3(32'h398dc3fc),
	.w4(32'hbb1e6032),
	.w5(32'hb9abd8bb),
	.w6(32'h3971dfcc),
	.w7(32'hbb098590),
	.w8(32'hba3c8b9c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2326f2),
	.w1(32'hba9bfb76),
	.w2(32'hbaeb3ffd),
	.w3(32'hba838719),
	.w4(32'hba87766b),
	.w5(32'hba90e61b),
	.w6(32'h3a60b9fc),
	.w7(32'h3a441dc3),
	.w8(32'h3a9d4f54),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12d54),
	.w1(32'h3a1f41ae),
	.w2(32'hb96392f4),
	.w3(32'h3a7eeb13),
	.w4(32'hba86d6e4),
	.w5(32'h38e00f2a),
	.w6(32'h3aac7ad0),
	.w7(32'hb9fc739a),
	.w8(32'h39d46810),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86cd81c),
	.w1(32'hba9803e3),
	.w2(32'hb9d8026e),
	.w3(32'hba4edbc6),
	.w4(32'hb9c777c7),
	.w5(32'h3a89f800),
	.w6(32'h38853305),
	.w7(32'h3aa14676),
	.w8(32'h3b46b61c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b570c),
	.w1(32'hba24f5b7),
	.w2(32'hbaa93298),
	.w3(32'h3aa8c02c),
	.w4(32'hbad77b96),
	.w5(32'h3a4aba59),
	.w6(32'h3b17ba4b),
	.w7(32'h3a4249bb),
	.w8(32'h3ac5f63f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91431d2),
	.w1(32'hb9d98845),
	.w2(32'hba4bd2e1),
	.w3(32'h3ad4a312),
	.w4(32'hba498d20),
	.w5(32'h39d48b5e),
	.w6(32'h3a87d602),
	.w7(32'hba89b050),
	.w8(32'h3a1904fa),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca0245),
	.w1(32'h3aedee9e),
	.w2(32'hb91b0502),
	.w3(32'hba062b74),
	.w4(32'hba9eb16d),
	.w5(32'hbae7d818),
	.w6(32'hba58841c),
	.w7(32'h3a8784d5),
	.w8(32'hb911f34d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae67d81),
	.w1(32'h391e5f6b),
	.w2(32'h3a92ce92),
	.w3(32'h3a19c6b4),
	.w4(32'hb905664e),
	.w5(32'h3aa6e63b),
	.w6(32'h3a8cb7cc),
	.w7(32'hba281d86),
	.w8(32'h3af65370),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7b501),
	.w1(32'h39aedcf8),
	.w2(32'h38c9d9f8),
	.w3(32'h3a218246),
	.w4(32'h3a5105f2),
	.w5(32'h3a067fa1),
	.w6(32'h3a64c801),
	.w7(32'h39d9cc76),
	.w8(32'h3aef781d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e1578d),
	.w1(32'h3a94f4ba),
	.w2(32'h3967e37d),
	.w3(32'hb9f2c1bb),
	.w4(32'h39c6973c),
	.w5(32'hb95a378f),
	.w6(32'h3ae8739e),
	.w7(32'h3a67a4cd),
	.w8(32'hba2cb951),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996dda9),
	.w1(32'hbacf0f15),
	.w2(32'h388f925f),
	.w3(32'hb9fde779),
	.w4(32'h3852309b),
	.w5(32'h3b1be089),
	.w6(32'h3a922f9e),
	.w7(32'hbb14af13),
	.w8(32'h39cf1a68),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ecea2),
	.w1(32'h3a14b3e4),
	.w2(32'h3a53f47c),
	.w3(32'h381a2d7c),
	.w4(32'h3ad670e2),
	.w5(32'h3ad77569),
	.w6(32'h3a994c2e),
	.w7(32'h39b15acd),
	.w8(32'h3aae2fc2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7da43),
	.w1(32'h3a8fd99c),
	.w2(32'hb9034659),
	.w3(32'hba2a3b52),
	.w4(32'h3a1d6a4a),
	.w5(32'hbb051401),
	.w6(32'h37fa59de),
	.w7(32'h3ad8d549),
	.w8(32'hbaf6a9b1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5075ee),
	.w1(32'h3a5b16ed),
	.w2(32'h3a8a7dd5),
	.w3(32'hba7ee07e),
	.w4(32'h3aa0fafb),
	.w5(32'hb9d1416b),
	.w6(32'hbb066c4e),
	.w7(32'h399ccdc2),
	.w8(32'hbaaeadc6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a5144),
	.w1(32'hbb04d986),
	.w2(32'hbad7b2a7),
	.w3(32'hb8f99639),
	.w4(32'hbae12b38),
	.w5(32'hba995726),
	.w6(32'hb97c826b),
	.w7(32'hba726be2),
	.w8(32'hbaeeef3a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75a3e),
	.w1(32'hba5bdcf5),
	.w2(32'hbb0ca46d),
	.w3(32'hbae35c28),
	.w4(32'hba3360d2),
	.w5(32'hbaf0f6e1),
	.w6(32'hbac7a804),
	.w7(32'hba1ee59c),
	.w8(32'hbac1f0c6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba317e63),
	.w1(32'hb9dc3713),
	.w2(32'h3a05c2c1),
	.w3(32'hbb09642c),
	.w4(32'h3a68e2b3),
	.w5(32'h3b2c8239),
	.w6(32'hba71f3da),
	.w7(32'h3a70c4db),
	.w8(32'h39f4851f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e456),
	.w1(32'h3ac579dc),
	.w2(32'h393b9fac),
	.w3(32'hb9e9727f),
	.w4(32'h3ace27db),
	.w5(32'h3a9bdc91),
	.w6(32'hba34ed8c),
	.w7(32'h3a49b963),
	.w8(32'hbac6c005),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28a060),
	.w1(32'hbaa123a4),
	.w2(32'hb9ea5273),
	.w3(32'h3a90acda),
	.w4(32'h39fcd83f),
	.w5(32'h3a6360ec),
	.w6(32'h3a2ddcbf),
	.w7(32'h38f9326d),
	.w8(32'h3a925705),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32c11b),
	.w1(32'h3a1f48b4),
	.w2(32'h3a14af65),
	.w3(32'hb9c19334),
	.w4(32'h3b03804f),
	.w5(32'h3b2e20d2),
	.w6(32'hb9c1cfb1),
	.w7(32'h3b071ecc),
	.w8(32'h3b2a8827),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22a548),
	.w1(32'hbaff9cfc),
	.w2(32'hb997f3e7),
	.w3(32'h3b2c762f),
	.w4(32'h389f8c4c),
	.w5(32'h3aa07d6a),
	.w6(32'h3b0ad833),
	.w7(32'hb92cc7ed),
	.w8(32'hb8dc28cb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae94cc1),
	.w1(32'hb99e2dc7),
	.w2(32'hb9ccdbf2),
	.w3(32'h3b4b34a1),
	.w4(32'hba84e6cb),
	.w5(32'hba2f7556),
	.w6(32'h3b2cf244),
	.w7(32'h39d7a117),
	.w8(32'h3b1c4c60),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5a6ed),
	.w1(32'hb9eec866),
	.w2(32'hba282d01),
	.w3(32'hb9f312f9),
	.w4(32'hb9b67275),
	.w5(32'hba8f6e70),
	.w6(32'h3aefa5e3),
	.w7(32'hba8c4613),
	.w8(32'hba8a23f3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0ee81),
	.w1(32'h39a7af50),
	.w2(32'hba4f1df6),
	.w3(32'hb8b9f3db),
	.w4(32'hbb12ee41),
	.w5(32'hba845eeb),
	.w6(32'hb97b0230),
	.w7(32'hba1b41c8),
	.w8(32'hb9fa4ae7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d36b4),
	.w1(32'hbc76f9ee),
	.w2(32'hbc811b5d),
	.w3(32'hb9e6b54b),
	.w4(32'hbbf7cfc9),
	.w5(32'hbc1bf694),
	.w6(32'h376b0d26),
	.w7(32'hbc94a753),
	.w8(32'hbc8565fd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71855),
	.w1(32'hbca3c127),
	.w2(32'hbc27f6e7),
	.w3(32'h3c192b8f),
	.w4(32'hbcbb6f75),
	.w5(32'hbc03aeb4),
	.w6(32'h3963a96d),
	.w7(32'hbc0092aa),
	.w8(32'h3c20dd5e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bc5ad),
	.w1(32'hbae0a484),
	.w2(32'hb9dd3627),
	.w3(32'h3c8782a4),
	.w4(32'hbbef5a55),
	.w5(32'h3b2785e3),
	.w6(32'h3cac2420),
	.w7(32'hbb2a97ca),
	.w8(32'h3aa6de85),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3916bc),
	.w1(32'hbca78d96),
	.w2(32'hbc13d127),
	.w3(32'h3bf46dea),
	.w4(32'hbcc9c4c1),
	.w5(32'hbc646f57),
	.w6(32'h3bbe96ac),
	.w7(32'hbc8c6f56),
	.w8(32'hbca7b394),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254128),
	.w1(32'h3b17db87),
	.w2(32'h3b9e1262),
	.w3(32'h3b98de3c),
	.w4(32'hba6be98a),
	.w5(32'hbbfe91b5),
	.w6(32'h39a665db),
	.w7(32'hbbb4b503),
	.w8(32'hbb927f61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cefb7),
	.w1(32'h3c257ae1),
	.w2(32'h3b317c0c),
	.w3(32'hbb15de5a),
	.w4(32'h3c036023),
	.w5(32'h3c800c70),
	.w6(32'h3ab43c3c),
	.w7(32'h3bb28a70),
	.w8(32'h3b19cdec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f3050),
	.w1(32'h39b15034),
	.w2(32'h3c09375d),
	.w3(32'h3b5321ad),
	.w4(32'h39f47c17),
	.w5(32'h3c120976),
	.w6(32'h3b932450),
	.w7(32'h3b112f18),
	.w8(32'h3b9adbc4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a042c),
	.w1(32'h3c0ad2f5),
	.w2(32'h3c208051),
	.w3(32'h3c0472db),
	.w4(32'h3c407d42),
	.w5(32'hbae2a1c8),
	.w6(32'h3aac6808),
	.w7(32'hb9befd14),
	.w8(32'h3b575c58),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3145f1),
	.w1(32'hbc321d1a),
	.w2(32'h3b43b5a3),
	.w3(32'hbbda3e4e),
	.w4(32'hbca8cbb8),
	.w5(32'hbc3a4785),
	.w6(32'h396e4019),
	.w7(32'hbc95d3c8),
	.w8(32'hbcb26b25),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c901693),
	.w1(32'h3c147024),
	.w2(32'hba8f83a5),
	.w3(32'h3cadf05a),
	.w4(32'h3d132785),
	.w5(32'h3c23d004),
	.w6(32'h3c243c7e),
	.w7(32'h3caacdc1),
	.w8(32'h3ba52957),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5255a1),
	.w1(32'h3bacaf6a),
	.w2(32'h3b3367e8),
	.w3(32'hbc65f4f0),
	.w4(32'hbaa99949),
	.w5(32'hbbee0c08),
	.w6(32'hbc293d56),
	.w7(32'hbbc38bd4),
	.w8(32'hbb16e6cf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb637955),
	.w1(32'h3d420034),
	.w2(32'h3b40d5f9),
	.w3(32'hbadd2afe),
	.w4(32'h3da35db3),
	.w5(32'h3c01a662),
	.w6(32'hbb987901),
	.w7(32'h3d68b0d9),
	.w8(32'h3bc1b520),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5813de),
	.w1(32'h3baff517),
	.w2(32'hbaf09f70),
	.w3(32'hbda3bb3d),
	.w4(32'hbaccfd8e),
	.w5(32'hbbbf266d),
	.w6(32'hbd7018f5),
	.w7(32'h3a5644b0),
	.w8(32'hbbecb1c1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6848a),
	.w1(32'hb9475a5c),
	.w2(32'hbc07191c),
	.w3(32'hbb9b20f4),
	.w4(32'h3b23991c),
	.w5(32'hbbb9be22),
	.w6(32'hbbd557e1),
	.w7(32'hb97b8778),
	.w8(32'hbb4aa6fe),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc39d04),
	.w1(32'h3b9d667d),
	.w2(32'hbc431c06),
	.w3(32'hb9977259),
	.w4(32'hbbcda2be),
	.w5(32'hbb21598e),
	.w6(32'h3ba1a9c8),
	.w7(32'h3a989d5d),
	.w8(32'hbb4e38c1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ca04),
	.w1(32'hbbb82637),
	.w2(32'h3bd38399),
	.w3(32'h3b1ab52e),
	.w4(32'hbc19df7c),
	.w5(32'hbc15560c),
	.w6(32'h3ac24f0b),
	.w7(32'hbc2295fd),
	.w8(32'hbc4dba44),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a231d),
	.w1(32'hbc0aa4c2),
	.w2(32'hbbaf8bdd),
	.w3(32'h3c48b023),
	.w4(32'hbc8f7acb),
	.w5(32'h3b8193ce),
	.w6(32'h3b91fb15),
	.w7(32'hbbacbb7b),
	.w8(32'h3c55561e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd9e5d),
	.w1(32'hbc626b2c),
	.w2(32'h3c37ff37),
	.w3(32'hbb389e87),
	.w4(32'hbc638312),
	.w5(32'hbc03d896),
	.w6(32'h3c1870f2),
	.w7(32'hbc7f6a06),
	.w8(32'hba1580cd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdd8f3),
	.w1(32'h3adc2837),
	.w2(32'h3ba6ccd7),
	.w3(32'h3cbdbddc),
	.w4(32'hb980bd8b),
	.w5(32'hba0d8f51),
	.w6(32'h3bf4f159),
	.w7(32'hbb96483a),
	.w8(32'hbbe911a6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f37e5),
	.w1(32'hb95321c2),
	.w2(32'h3af308fd),
	.w3(32'h3ac4efc4),
	.w4(32'hbbb74a01),
	.w5(32'h3c1a0b95),
	.w6(32'h3b058a87),
	.w7(32'hbaa00512),
	.w8(32'hbb44a29b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443561),
	.w1(32'hbb9797ec),
	.w2(32'hbad1a64d),
	.w3(32'h3b687dd7),
	.w4(32'hbc881e7e),
	.w5(32'h3c27b055),
	.w6(32'h3bffc971),
	.w7(32'hbc6ea6b7),
	.w8(32'hbb25f99c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb479fd),
	.w1(32'hbca57669),
	.w2(32'hbbb799dd),
	.w3(32'h3b9c461d),
	.w4(32'hbce9ab06),
	.w5(32'hbba3644e),
	.w6(32'hb9ab957e),
	.w7(32'hbcb0f5a7),
	.w8(32'hbc0d5e5a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c4ea),
	.w1(32'h3a1edf89),
	.w2(32'h3b74350f),
	.w3(32'h3c30c4b7),
	.w4(32'hbc1d2d51),
	.w5(32'h3c11e7c2),
	.w6(32'h3b3db719),
	.w7(32'hbb4daf02),
	.w8(32'hbbcbeddb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2707),
	.w1(32'h3c024dc3),
	.w2(32'h3ad70e5d),
	.w3(32'h3b4b349f),
	.w4(32'h3cbc0d4b),
	.w5(32'h3bbc8962),
	.w6(32'hbc1596f7),
	.w7(32'h3c9603d3),
	.w8(32'h3ad9caa3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ac3a3),
	.w1(32'h3c201197),
	.w2(32'h3b2fc317),
	.w3(32'hbcd75b94),
	.w4(32'h3c17ec4d),
	.w5(32'hbae1c608),
	.w6(32'hbc87d8e0),
	.w7(32'h3c4886b9),
	.w8(32'h3b743b43),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73a7ae),
	.w1(32'h3b3aa570),
	.w2(32'hbac8d7de),
	.w3(32'hbc917c1e),
	.w4(32'hbc42f683),
	.w5(32'h3b6c5991),
	.w6(32'hbb80668c),
	.w7(32'hbccecd9b),
	.w8(32'hbcae8b3a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298f96),
	.w1(32'hbc2189ab),
	.w2(32'h3aeca187),
	.w3(32'h3b8a7edc),
	.w4(32'hbc15b25c),
	.w5(32'hbcc972d6),
	.w6(32'hbbfa4d55),
	.w7(32'hbbcc2e49),
	.w8(32'h3b20f768),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28c3dc),
	.w1(32'hba58638b),
	.w2(32'hbc1bba2e),
	.w3(32'h3cd94e62),
	.w4(32'hbc422b7d),
	.w5(32'hbc78cec4),
	.w6(32'h3caa6125),
	.w7(32'hbc4abdaa),
	.w8(32'hbc03e0f6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909ed2),
	.w1(32'hbbbfacfc),
	.w2(32'h3b954a99),
	.w3(32'h3cde8d18),
	.w4(32'hbc031540),
	.w5(32'h3af0bc33),
	.w6(32'h3cb8f63d),
	.w7(32'hbc7bc6b9),
	.w8(32'h3b491d22),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96866a),
	.w1(32'h3af4e9fb),
	.w2(32'h3bbb1f73),
	.w3(32'hbbc5b1f6),
	.w4(32'hbb381365),
	.w5(32'h3b02867b),
	.w6(32'h39af7633),
	.w7(32'hbab23c05),
	.w8(32'hbb0b1ae7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0226c9),
	.w1(32'hbbf50b7c),
	.w2(32'hbac1dd0f),
	.w3(32'hba962b8f),
	.w4(32'hbc889b53),
	.w5(32'h3bf9fbcf),
	.w6(32'hbb7bf98d),
	.w7(32'hbc254d80),
	.w8(32'hbca2d7e6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c500b),
	.w1(32'hbafcbd2b),
	.w2(32'hbac90b7e),
	.w3(32'h3b864170),
	.w4(32'hbb8e86eb),
	.w5(32'hbbabf9ac),
	.w6(32'hbacb314a),
	.w7(32'hbc0d4d74),
	.w8(32'hbbb489f6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b455529),
	.w1(32'hbbeaaac2),
	.w2(32'hba66eaae),
	.w3(32'h3b400b63),
	.w4(32'hbc7edfdc),
	.w5(32'hb90c0c0a),
	.w6(32'h3c29b6ad),
	.w7(32'hbc2503b3),
	.w8(32'hbbcfb243),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b629c74),
	.w1(32'hbadc7e62),
	.w2(32'hbc6fd1e5),
	.w3(32'h3c614aad),
	.w4(32'hbaa9bf6e),
	.w5(32'hbc95cd92),
	.w6(32'h3b311caa),
	.w7(32'hbbf1aa55),
	.w8(32'hbba0668b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65538),
	.w1(32'hbc737090),
	.w2(32'h3acba803),
	.w3(32'h3ca54fea),
	.w4(32'hbd04fc33),
	.w5(32'hbb8d0814),
	.w6(32'h3c69882e),
	.w7(32'hbc9122f2),
	.w8(32'hbc7d0f13),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f941e),
	.w1(32'h3affff1e),
	.w2(32'hb9d01e11),
	.w3(32'h3c3ab0c0),
	.w4(32'hba212c07),
	.w5(32'h38ac7ff7),
	.w6(32'h3b06b7fe),
	.w7(32'h3b20dd8f),
	.w8(32'h3c1a4b58),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b0c7d),
	.w1(32'h3b860acc),
	.w2(32'h3b5494ee),
	.w3(32'h3a28d4d3),
	.w4(32'h3c013253),
	.w5(32'h3b666ff8),
	.w6(32'h3c426595),
	.w7(32'h39ca0697),
	.w8(32'hb9715a84),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3023),
	.w1(32'h3a0f1097),
	.w2(32'hb9f06ba1),
	.w3(32'h3acebba6),
	.w4(32'h39e3ac10),
	.w5(32'h3b95a326),
	.w6(32'h3b269d51),
	.w7(32'hba91df8a),
	.w8(32'h3a038db1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae0592),
	.w1(32'hbc5f07dc),
	.w2(32'h3b08d248),
	.w3(32'h3a9a91e3),
	.w4(32'hbca614f9),
	.w5(32'hbc2b9788),
	.w6(32'hbb292226),
	.w7(32'hbccb2e1a),
	.w8(32'hbbead72b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15174b),
	.w1(32'hbacce90c),
	.w2(32'h3bc716f7),
	.w3(32'h3af8f327),
	.w4(32'hbba19601),
	.w5(32'hbbc1dcf0),
	.w6(32'hbc5fecae),
	.w7(32'h3b0ef5d6),
	.w8(32'h3b8877fa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b555b03),
	.w1(32'hbbddaa82),
	.w2(32'hbae0585c),
	.w3(32'hbaebc8ee),
	.w4(32'hbbed6a14),
	.w5(32'hbbec3548),
	.w6(32'h3bf76e87),
	.w7(32'hbc0be114),
	.w8(32'hbb8810b6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d6d96),
	.w1(32'hbc87de8d),
	.w2(32'hbb960459),
	.w3(32'h3cafedbe),
	.w4(32'hbcbe63cc),
	.w5(32'h3aff67f3),
	.w6(32'h3c196d80),
	.w7(32'hbb5f5d80),
	.w8(32'h3bef1c9f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b8492),
	.w1(32'hbc1f7d0a),
	.w2(32'hbb972d1d),
	.w3(32'h3bca8ca8),
	.w4(32'hbc88c9b1),
	.w5(32'h39536a67),
	.w6(32'h3b34e5aa),
	.w7(32'hbcad0bde),
	.w8(32'hbba27605),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab94d5),
	.w1(32'h3adf944c),
	.w2(32'h3a9ab446),
	.w3(32'h3cb4819d),
	.w4(32'h3b799f74),
	.w5(32'hbb8f4668),
	.w6(32'h3ca5605f),
	.w7(32'hbbaefd4d),
	.w8(32'hbb87eda4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87766f),
	.w1(32'h3a992690),
	.w2(32'h3c26d3f8),
	.w3(32'hbb8b6b99),
	.w4(32'h3ca28c9b),
	.w5(32'hbb1b3995),
	.w6(32'hbbb7a291),
	.w7(32'h3b7a10c3),
	.w8(32'h3b709cd7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822e38),
	.w1(32'h3b979425),
	.w2(32'h3c2e4c55),
	.w3(32'hbb5b6bdf),
	.w4(32'h3b58b7fe),
	.w5(32'h3c946ead),
	.w6(32'hbabf1cf5),
	.w7(32'hbaf5a449),
	.w8(32'hba3c9051),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92405a),
	.w1(32'hbc3dafb7),
	.w2(32'hbc11ca2b),
	.w3(32'hbbd316b7),
	.w4(32'hbc7bd496),
	.w5(32'hbc2cf0da),
	.w6(32'hbc5e579f),
	.w7(32'hbc03551c),
	.w8(32'h3a71234a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ae4e5),
	.w1(32'hbb981b29),
	.w2(32'h3bac7e20),
	.w3(32'h3cbd70fc),
	.w4(32'h3990e0d3),
	.w5(32'h3c94e43c),
	.w6(32'h3c9051cd),
	.w7(32'hb8d87ee6),
	.w8(32'hbb864ed9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0a49),
	.w1(32'h3a0b6cc4),
	.w2(32'hb8984551),
	.w3(32'h3afe7ae9),
	.w4(32'hbc056f55),
	.w5(32'hbc927082),
	.w6(32'hbc19669b),
	.w7(32'h3b5861b8),
	.w8(32'hbbd9eb1e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62ef55),
	.w1(32'hbb2f91ac),
	.w2(32'h3b85e315),
	.w3(32'hbbb92fd1),
	.w4(32'hbaa5e0f8),
	.w5(32'h3b55371f),
	.w6(32'h3beb48c2),
	.w7(32'hbacccef7),
	.w8(32'h3c1e7226),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c359090),
	.w1(32'hbc6bc0cd),
	.w2(32'hbbf66423),
	.w3(32'h35b7b56e),
	.w4(32'hbd018b7c),
	.w5(32'hbcf053e3),
	.w6(32'h3c2df12d),
	.w7(32'hbca0516d),
	.w8(32'hbc0e174f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c617658),
	.w1(32'h3c0bbb44),
	.w2(32'hbba7ad1a),
	.w3(32'h3ca25420),
	.w4(32'h3c18595f),
	.w5(32'hbc1e64b0),
	.w6(32'h3c2bfde9),
	.w7(32'h3c20fd2f),
	.w8(32'hbbbcaff4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7b5a),
	.w1(32'hbc972342),
	.w2(32'hbc0558b1),
	.w3(32'hbc608d6f),
	.w4(32'hbc3fedab),
	.w5(32'hbc5965a4),
	.w6(32'hbc2f3943),
	.w7(32'hbc6b92a8),
	.w8(32'h3c06077c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba597b),
	.w1(32'h3a10282c),
	.w2(32'h38da7896),
	.w3(32'h3bb5644f),
	.w4(32'hbbf93906),
	.w5(32'hbb53e125),
	.w6(32'h3c9ae82e),
	.w7(32'h3a6d753d),
	.w8(32'h3c64c60a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adec9d5),
	.w1(32'h3b788e23),
	.w2(32'h3c22dc0b),
	.w3(32'h3c8a5d37),
	.w4(32'h3c8311a8),
	.w5(32'h3cb4db7d),
	.w6(32'h3c9a8f22),
	.w7(32'h3aafb2cb),
	.w8(32'h3c14e7c3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3110e5),
	.w1(32'hbb280f13),
	.w2(32'h3c57e674),
	.w3(32'hbbc21cbb),
	.w4(32'hbc6378cc),
	.w5(32'hbbeebc5f),
	.w6(32'hbc43cd53),
	.w7(32'hbbcacd2b),
	.w8(32'hbbfabad8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5eeacf),
	.w1(32'hbc01636a),
	.w2(32'hba120958),
	.w3(32'h3bcc6261),
	.w4(32'hbc2d2180),
	.w5(32'hbb3a0730),
	.w6(32'h3bb01750),
	.w7(32'hbbba243b),
	.w8(32'h3bc4d638),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b471b18),
	.w1(32'hbc7c4730),
	.w2(32'hbb4c527b),
	.w3(32'h3b7205b7),
	.w4(32'hbcba0119),
	.w5(32'hbb4b084b),
	.w6(32'h3bb13cfa),
	.w7(32'hbc77a79c),
	.w8(32'hbc268dfa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9de547),
	.w1(32'hbb4223bc),
	.w2(32'hbc5ddb18),
	.w3(32'h3d15110d),
	.w4(32'hbc4320b0),
	.w5(32'hbbcf355b),
	.w6(32'h3c8d9b87),
	.w7(32'hbbfa9f98),
	.w8(32'h3b523f28),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule