module layer_8_featuremap_39(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897bc3),
	.w1(32'hbab4e5fe),
	.w2(32'h3a0e7239),
	.w3(32'hbb1e1a92),
	.w4(32'hba6f0a43),
	.w5(32'h3843f6a6),
	.w6(32'hbaae67ed),
	.w7(32'hba478afe),
	.w8(32'hb892f5fe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501149),
	.w1(32'h3b420350),
	.w2(32'h3b2d34fa),
	.w3(32'h3b4f5712),
	.w4(32'h3b159c3f),
	.w5(32'h3a99f5dc),
	.w6(32'h3b402122),
	.w7(32'h3b0b52f9),
	.w8(32'h3af1539b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18fc8d),
	.w1(32'h3ad650ac),
	.w2(32'h3a91f6b7),
	.w3(32'h3b6c0f78),
	.w4(32'h3adcfaa9),
	.w5(32'h3a7bb002),
	.w6(32'h3b8cd67d),
	.w7(32'h3b380e7c),
	.w8(32'h3ab6803d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa748b8),
	.w1(32'hbb2039d2),
	.w2(32'hba31fb1e),
	.w3(32'h39b0c871),
	.w4(32'hba9f3420),
	.w5(32'hba896c23),
	.w6(32'h3a169842),
	.w7(32'h3997fd77),
	.w8(32'h39c1beb8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1b7d3),
	.w1(32'h3af1b5d0),
	.w2(32'h3b552b2f),
	.w3(32'hb8776b38),
	.w4(32'h3a2ea1bf),
	.w5(32'h3b1c87a6),
	.w6(32'h39b5fd7c),
	.w7(32'h3a38896f),
	.w8(32'h3b690811),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8558),
	.w1(32'h3b46c324),
	.w2(32'h3bb7031d),
	.w3(32'h3ace5c93),
	.w4(32'h3b21dfd1),
	.w5(32'h3b774215),
	.w6(32'h3aeaa27b),
	.w7(32'h3b0e8ef3),
	.w8(32'h3b9a5a16),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a257e34),
	.w1(32'h3a4e88fe),
	.w2(32'h3a214542),
	.w3(32'h39e65a48),
	.w4(32'h3a37b14f),
	.w5(32'h3a2a07f2),
	.w6(32'h3a324ebb),
	.w7(32'h39bacba0),
	.w8(32'hb7d35b02),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db24b7),
	.w1(32'h3a87b972),
	.w2(32'h3b4c7a3d),
	.w3(32'h3a85ab04),
	.w4(32'h39e7c776),
	.w5(32'h3ad48954),
	.w6(32'hba4abf5f),
	.w7(32'hba89a0cb),
	.w8(32'h3ad33c30),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab1979),
	.w1(32'h3b3d3bf9),
	.w2(32'h3b6abda7),
	.w3(32'h3b0092aa),
	.w4(32'h3b2a565c),
	.w5(32'h3b819a5c),
	.w6(32'h3b0aa799),
	.w7(32'h3b2c5338),
	.w8(32'h3b23cd11),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb505e02),
	.w1(32'hbaaecea6),
	.w2(32'hbb07eca4),
	.w3(32'h3a73fc8e),
	.w4(32'hbb14d129),
	.w5(32'hbb0eac32),
	.w6(32'hba21f956),
	.w7(32'hbad68007),
	.w8(32'hba9eb1f2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e49e6),
	.w1(32'hbaa8300e),
	.w2(32'h39fed121),
	.w3(32'hbb46b9a1),
	.w4(32'hbad4fe85),
	.w5(32'hb989f1e0),
	.w6(32'hbb252ced),
	.w7(32'hba967025),
	.w8(32'h39d88f5c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba314245),
	.w1(32'h3a620f62),
	.w2(32'h3b088398),
	.w3(32'hb9fca9d4),
	.w4(32'h3a9ccc14),
	.w5(32'h3adde5b5),
	.w6(32'h3a9379d2),
	.w7(32'h3acaef55),
	.w8(32'h3b047aac),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09f394),
	.w1(32'h3abd486e),
	.w2(32'h3ad3e141),
	.w3(32'h3b2a1c63),
	.w4(32'h3b0da10b),
	.w5(32'h3b35f4bd),
	.w6(32'h3b0ac908),
	.w7(32'h3b2a70ac),
	.w8(32'h3b9a9b65),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c680),
	.w1(32'h3a9f95b8),
	.w2(32'h3a67b1a5),
	.w3(32'h3b1a4ae3),
	.w4(32'h3abae4b2),
	.w5(32'h3a16902c),
	.w6(32'h3a79f64a),
	.w7(32'h3a4020b0),
	.w8(32'h3a2f0b31),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a882eef),
	.w1(32'h3a2fa3e1),
	.w2(32'h39ea227b),
	.w3(32'h3a906307),
	.w4(32'h3a6dff98),
	.w5(32'h3994a6b1),
	.w6(32'h3a0925c9),
	.w7(32'h399e0415),
	.w8(32'hb999a94b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbde3e),
	.w1(32'hb9d8b34d),
	.w2(32'hb9aa82c5),
	.w3(32'hb9221890),
	.w4(32'hb9101c50),
	.w5(32'hb946a277),
	.w6(32'hb8ec75fa),
	.w7(32'h392ea39b),
	.w8(32'h3a18b99c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba746f11),
	.w1(32'hbab2eb52),
	.w2(32'hbae7c78c),
	.w3(32'hb900d1af),
	.w4(32'hb9c1fe19),
	.w5(32'hba5e4ff5),
	.w6(32'h39b03b3d),
	.w7(32'h3a30d609),
	.w8(32'hb9a0a8ac),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39141967),
	.w1(32'hb9f08a14),
	.w2(32'h3942c5f1),
	.w3(32'h3a269ad6),
	.w4(32'hb88ae3e4),
	.w5(32'hb9b99017),
	.w6(32'h3ac45305),
	.w7(32'hba052ca1),
	.w8(32'h3a0abf65),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb950235),
	.w1(32'hba8dd860),
	.w2(32'h3b01d420),
	.w3(32'hbb474fcc),
	.w4(32'h3a2a30c2),
	.w5(32'h3a98d533),
	.w6(32'hba2c4282),
	.w7(32'hb916250e),
	.w8(32'h3a124b9e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c31f),
	.w1(32'hbadec851),
	.w2(32'h3bb61646),
	.w3(32'hbc051905),
	.w4(32'hbb9d460a),
	.w5(32'h3b555060),
	.w6(32'hbb7ea564),
	.w7(32'h392248b6),
	.w8(32'h3c0c9d07),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393cda2f),
	.w1(32'h3a93e8d4),
	.w2(32'h3b045f93),
	.w3(32'h3a14deeb),
	.w4(32'h3b23a1f4),
	.w5(32'h3b64ec6a),
	.w6(32'h3af6a27c),
	.w7(32'h3b0a317f),
	.w8(32'h3b7838aa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6837),
	.w1(32'h3b1ecd6f),
	.w2(32'h3b440c24),
	.w3(32'h3b9aa2d1),
	.w4(32'h3b476b36),
	.w5(32'h3b34832f),
	.w6(32'h3b868582),
	.w7(32'h3b17028e),
	.w8(32'h3b35c965),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa867e9),
	.w1(32'h38ed3e1c),
	.w2(32'h3b0455d2),
	.w3(32'hbad0f2a8),
	.w4(32'hbb4d5535),
	.w5(32'hbb5f16ed),
	.w6(32'hbb0d80e9),
	.w7(32'hbafd5736),
	.w8(32'hbb30fd09),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204f79),
	.w1(32'hba88d08a),
	.w2(32'h3b3e929e),
	.w3(32'hbb3fb8b1),
	.w4(32'hbb1968aa),
	.w5(32'h3a6ecd1a),
	.w6(32'hbadb2681),
	.w7(32'h3a6ffc58),
	.w8(32'h3b353dc5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09c9eb),
	.w1(32'h3a08f03a),
	.w2(32'h3a7101b3),
	.w3(32'h3a0fc281),
	.w4(32'hb7738ed7),
	.w5(32'h3a08ecaa),
	.w6(32'h3a5b8da6),
	.w7(32'h3aa3fe56),
	.w8(32'h3a606082),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb382e20),
	.w1(32'h3a6a01d6),
	.w2(32'h3baa28ca),
	.w3(32'hbb4f14a2),
	.w4(32'hba56ac28),
	.w5(32'h3af5bf3c),
	.w6(32'hbaf05b58),
	.w7(32'h39f7407e),
	.w8(32'h3b4d1e51),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940a07f),
	.w1(32'hba247b8f),
	.w2(32'hb9b3269b),
	.w3(32'hb9562415),
	.w4(32'hba6d0a9e),
	.w5(32'hb9fb959d),
	.w6(32'hb90ea229),
	.w7(32'hb91df934),
	.w8(32'h3a5a537f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ebfb),
	.w1(32'h3c284c0b),
	.w2(32'h3c4dbef4),
	.w3(32'h3b22d56f),
	.w4(32'h3c0edce1),
	.w5(32'h3c8b9bf9),
	.w6(32'h3bf0cbaa),
	.w7(32'h3c08d419),
	.w8(32'h3b9eaae8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8829e),
	.w1(32'h3aa9ebca),
	.w2(32'h3b10f744),
	.w3(32'hb8b30f8b),
	.w4(32'h3aadf8f3),
	.w5(32'h3a8aa429),
	.w6(32'hba31200d),
	.w7(32'h3acf1caf),
	.w8(32'h3b1fad3b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbd6a4),
	.w1(32'h3a2c468e),
	.w2(32'h3a357a4a),
	.w3(32'h39c9a1c2),
	.w4(32'h39f814f8),
	.w5(32'h3a023aa4),
	.w6(32'h39e9b046),
	.w7(32'h3a022d59),
	.w8(32'h3adebab3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b6608),
	.w1(32'hbab7e97a),
	.w2(32'hba19cce2),
	.w3(32'h3b0fa48e),
	.w4(32'h3a76dd0d),
	.w5(32'h39fe580a),
	.w6(32'h39ceee62),
	.w7(32'h3a8b8c5a),
	.w8(32'h3a31b892),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f7f84),
	.w1(32'h3a191de9),
	.w2(32'h3b2bade5),
	.w3(32'hba39bada),
	.w4(32'h39b390d3),
	.w5(32'h3b6255c4),
	.w6(32'hb6e80994),
	.w7(32'h3a521688),
	.w8(32'h3b8b9901),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2202b9),
	.w1(32'hba3916c0),
	.w2(32'hb9d7dea3),
	.w3(32'h3abd9b39),
	.w4(32'h39106296),
	.w5(32'hba985d90),
	.w6(32'h3ad4df72),
	.w7(32'h3aee863d),
	.w8(32'h3a57ddaf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e6ca),
	.w1(32'hba06b1e0),
	.w2(32'hba2fc8c5),
	.w3(32'h39956f01),
	.w4(32'hb9be0ad9),
	.w5(32'hba402fd6),
	.w6(32'h3ac8af75),
	.w7(32'h3ab2aea6),
	.w8(32'h3ac2fc73),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af63eac),
	.w1(32'hb8e6c3e9),
	.w2(32'h39d78f7c),
	.w3(32'h3a91c454),
	.w4(32'hba91def8),
	.w5(32'h3a2ed91f),
	.w6(32'h3ad8f837),
	.w7(32'h398c1dde),
	.w8(32'h3a97bf10),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe034),
	.w1(32'hba591cc8),
	.w2(32'h3a331c24),
	.w3(32'hbac5b8c3),
	.w4(32'h39a28e23),
	.w5(32'h3a75dcf7),
	.w6(32'hba303691),
	.w7(32'h3977af08),
	.w8(32'h3a505086),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1acdb4),
	.w1(32'hba7a5f82),
	.w2(32'hb98e5be8),
	.w3(32'hb9cfc731),
	.w4(32'hbab18a23),
	.w5(32'hba257730),
	.w6(32'hb9584121),
	.w7(32'h39469edf),
	.w8(32'hb919fb68),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5089dd),
	.w1(32'h3b42857b),
	.w2(32'h3b340185),
	.w3(32'h3b58a728),
	.w4(32'h3b2a89c5),
	.w5(32'h3b16f21f),
	.w6(32'h3b25e475),
	.w7(32'h3ade179e),
	.w8(32'h3b3576cf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed01c9),
	.w1(32'h3aa0aa77),
	.w2(32'h3a619b87),
	.w3(32'h3b02cf6d),
	.w4(32'h3ae26109),
	.w5(32'h39d41a1e),
	.w6(32'h3a7937be),
	.w7(32'h3a1b6a95),
	.w8(32'h3a67bd90),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f370b),
	.w1(32'h38073ba0),
	.w2(32'h396ddb3f),
	.w3(32'h39727d25),
	.w4(32'h38d3fd86),
	.w5(32'h399e4fb4),
	.w6(32'h39bd89f5),
	.w7(32'h39aaffb8),
	.w8(32'h39016604),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2701fb),
	.w1(32'h3a8ace99),
	.w2(32'h3bc934f0),
	.w3(32'hba7b63ae),
	.w4(32'h3aac5be0),
	.w5(32'h3ba3f593),
	.w6(32'h3a3c5900),
	.w7(32'h3b4df0bf),
	.w8(32'h3c1e3054),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb443f),
	.w1(32'h3a021877),
	.w2(32'h39f1ad3c),
	.w3(32'h3ad61fb6),
	.w4(32'h3a71f636),
	.w5(32'h3a926554),
	.w6(32'h3b39fc07),
	.w7(32'h3abf2a5b),
	.w8(32'hbb213740),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e2a3),
	.w1(32'hbb55eb9e),
	.w2(32'hbaf297d1),
	.w3(32'hbb4024ef),
	.w4(32'hbb63a173),
	.w5(32'hbabd5534),
	.w6(32'hbbae8f43),
	.w7(32'hba90605b),
	.w8(32'h3a5a5fe0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a741),
	.w1(32'h3a2aefb0),
	.w2(32'h3ae708ad),
	.w3(32'hbb1ed040),
	.w4(32'hba62b439),
	.w5(32'h3a57d959),
	.w6(32'h3a9e0e15),
	.w7(32'h3a63b209),
	.w8(32'h3b1297fd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9b5bc),
	.w1(32'h3b3c9fbb),
	.w2(32'h3b89de55),
	.w3(32'h3a2622c8),
	.w4(32'h3aaf714d),
	.w5(32'h3a782ace),
	.w6(32'h3aabac41),
	.w7(32'h3a5e9e20),
	.w8(32'h3b877242),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e2abe),
	.w1(32'h3b431c38),
	.w2(32'h3ae43b18),
	.w3(32'h3b33d3db),
	.w4(32'h3afa9f83),
	.w5(32'h3aa61e41),
	.w6(32'h3bae423a),
	.w7(32'h3b4497fe),
	.w8(32'h3afc9131),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba331581),
	.w1(32'h3aa3f568),
	.w2(32'h3ab225ac),
	.w3(32'hba708856),
	.w4(32'hb9a995ed),
	.w5(32'h3956567e),
	.w6(32'hba0ffc23),
	.w7(32'hbacd27ed),
	.w8(32'h3b4b871f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a430ff0),
	.w1(32'h3b63e6f8),
	.w2(32'h3b497314),
	.w3(32'hbaa720be),
	.w4(32'hb8623fe1),
	.w5(32'h3ac65c28),
	.w6(32'h3aaef4c5),
	.w7(32'h39ee975c),
	.w8(32'h3b036b60),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0bdad),
	.w1(32'hbab48370),
	.w2(32'h398cae06),
	.w3(32'hb9dfa56c),
	.w4(32'hbaa3f91e),
	.w5(32'hba119198),
	.w6(32'h3ada4cc7),
	.w7(32'h3b557148),
	.w8(32'h3b5414c4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae28005),
	.w1(32'h3a5f6dcc),
	.w2(32'h3a86e50a),
	.w3(32'h3aa73e9b),
	.w4(32'h3a1c19ef),
	.w5(32'hb9653fc4),
	.w6(32'h3af6b531),
	.w7(32'h39dab10c),
	.w8(32'h3a75dcac),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c291daf),
	.w1(32'h3c242f63),
	.w2(32'h3c2f6202),
	.w3(32'h3c20e3b2),
	.w4(32'h3c05c075),
	.w5(32'h3c23a818),
	.w6(32'h3c0cdcda),
	.w7(32'h3c01d9b7),
	.w8(32'h3c2f5fbb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa645b4),
	.w1(32'h3bc0e95e),
	.w2(32'h3c470855),
	.w3(32'hba524b13),
	.w4(32'h3b51554b),
	.w5(32'h3bc7c668),
	.w6(32'h38b0c0aa),
	.w7(32'h3aebd776),
	.w8(32'h3a96344d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26129a),
	.w1(32'h3a851f1e),
	.w2(32'h3bb01a08),
	.w3(32'hbb1f85e3),
	.w4(32'hb99e354a),
	.w5(32'h3b71a71d),
	.w6(32'hbb892ad3),
	.w7(32'hba165304),
	.w8(32'h3b8b3317),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0a74),
	.w1(32'hba8e9e97),
	.w2(32'hb97287ee),
	.w3(32'hb9282543),
	.w4(32'hba0dd821),
	.w5(32'hbacaabe2),
	.w6(32'h39822c88),
	.w7(32'h3a6e4a83),
	.w8(32'hbae682f5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c068a),
	.w1(32'h39e7fb9f),
	.w2(32'h38daafc8),
	.w3(32'h3a22dfa0),
	.w4(32'hba7e4b0e),
	.w5(32'hba924212),
	.w6(32'hbad18086),
	.w7(32'hba15b5ea),
	.w8(32'hbb76f9ad),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1f32f),
	.w1(32'hbac77cc1),
	.w2(32'hbb19005e),
	.w3(32'hbb328ed4),
	.w4(32'h38f40c5f),
	.w5(32'hba76b6de),
	.w6(32'hb8c8210a),
	.w7(32'hbabaf103),
	.w8(32'h3a8c4ec9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432705),
	.w1(32'hba47cfd1),
	.w2(32'hba1b2c57),
	.w3(32'hba667ef4),
	.w4(32'hba94067f),
	.w5(32'h3922760d),
	.w6(32'h37e0302d),
	.w7(32'hba26e008),
	.w8(32'hbb5709c9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd1a6),
	.w1(32'hbac7e6ed),
	.w2(32'hba918671),
	.w3(32'hbb4adc7b),
	.w4(32'hbad1dde8),
	.w5(32'hba90e7c6),
	.w6(32'hbb2dda99),
	.w7(32'hbb316009),
	.w8(32'h3b949a8a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95344a0),
	.w1(32'hb93e3b32),
	.w2(32'h3a15bc3b),
	.w3(32'hb910ff31),
	.w4(32'hba044667),
	.w5(32'h3a23bca9),
	.w6(32'h3b01c811),
	.w7(32'h3b6f8fd8),
	.w8(32'hb9d37a62),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2020d2),
	.w1(32'h39cf06c0),
	.w2(32'h3a5f66c4),
	.w3(32'h39f84646),
	.w4(32'hb8a68e1f),
	.w5(32'hba17f328),
	.w6(32'h39ad2c8f),
	.w7(32'h3aa51d4f),
	.w8(32'h3b45fa2e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f7786),
	.w1(32'h3a8b9279),
	.w2(32'h39fdd071),
	.w3(32'h3823208b),
	.w4(32'h399152db),
	.w5(32'h3a8d1576),
	.w6(32'h3a6c834b),
	.w7(32'h38af298e),
	.w8(32'h3b7e25e5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fbe99),
	.w1(32'h3b5928c8),
	.w2(32'h3b26de6b),
	.w3(32'h3ad1e596),
	.w4(32'h3ab72afa),
	.w5(32'h3aee136c),
	.w6(32'h3b8e789c),
	.w7(32'h3b2847d5),
	.w8(32'hb98e8c2e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8a696),
	.w1(32'h3af6c636),
	.w2(32'h3be3acba),
	.w3(32'h3a2d6aea),
	.w4(32'h3ac03b90),
	.w5(32'h3bd5fdb6),
	.w6(32'h3a9ee017),
	.w7(32'h3b39a2d5),
	.w8(32'h3b3409b1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1f749),
	.w1(32'hb9d5c2d0),
	.w2(32'hbafe0363),
	.w3(32'hb9dbeac3),
	.w4(32'hba2ddbea),
	.w5(32'hba401bcc),
	.w6(32'hbae5e6ed),
	.w7(32'hbb3a59b7),
	.w8(32'h3ab03c82),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7aac8),
	.w1(32'h3a7a83dd),
	.w2(32'h39fc0585),
	.w3(32'h3a8fea4e),
	.w4(32'hb9bfabf4),
	.w5(32'h39734f7b),
	.w6(32'h3ab0c5b8),
	.w7(32'h39e0b7bb),
	.w8(32'hba88f63a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b06868),
	.w1(32'h395c6fe5),
	.w2(32'h3a77fc72),
	.w3(32'hba308dcb),
	.w4(32'hba3d9250),
	.w5(32'hb9392b48),
	.w6(32'hba663d8e),
	.w7(32'hba5ae7aa),
	.w8(32'h3a84a449),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065592),
	.w1(32'h3b1d1df1),
	.w2(32'h3b84d4d4),
	.w3(32'h3ac0ebbc),
	.w4(32'h3aa8f6f8),
	.w5(32'h3b21597a),
	.w6(32'h3b52119e),
	.w7(32'h3b446696),
	.w8(32'h3b5718f5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71838c),
	.w1(32'h3aad4841),
	.w2(32'h3b1bc5d7),
	.w3(32'hba991702),
	.w4(32'hba2ada77),
	.w5(32'h3a99e1f2),
	.w6(32'h3acc34d3),
	.w7(32'h3abaff73),
	.w8(32'h3b35452f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cee0),
	.w1(32'h3a890f23),
	.w2(32'h3a589864),
	.w3(32'h3aa23fb9),
	.w4(32'h3a3507de),
	.w5(32'h3a7cc996),
	.w6(32'h3aae5907),
	.w7(32'h3a0ab96a),
	.w8(32'h3b7a66b4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d0349),
	.w1(32'h3991e4a4),
	.w2(32'h3bb16e5e),
	.w3(32'hbbad699d),
	.w4(32'hba06dc2d),
	.w5(32'h3b8a6f6c),
	.w6(32'hba0f9977),
	.w7(32'h3b2a4753),
	.w8(32'h3a8e995a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85712b),
	.w1(32'h3a5fd9a8),
	.w2(32'h3a2f39fc),
	.w3(32'h3a940545),
	.w4(32'h3a09ee03),
	.w5(32'h3a7844c8),
	.w6(32'h3ab1a242),
	.w7(32'h3a5a05fe),
	.w8(32'h3abaa822),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e8b57),
	.w1(32'h3aaae4e8),
	.w2(32'h3b3f0633),
	.w3(32'hba7b457c),
	.w4(32'h3a24214d),
	.w5(32'h3b5f0731),
	.w6(32'h3aa541b4),
	.w7(32'h3afc3e9a),
	.w8(32'h3b868c69),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad11d69),
	.w1(32'h3ac03496),
	.w2(32'h3a411b46),
	.w3(32'h3abb48a7),
	.w4(32'h3a739652),
	.w5(32'h3a11fb37),
	.w6(32'h3af770ae),
	.w7(32'h3a76a358),
	.w8(32'hbafe3172),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15a968),
	.w1(32'h396f6fa1),
	.w2(32'hba8cd121),
	.w3(32'h3a453d2e),
	.w4(32'hba00c91d),
	.w5(32'hbaa90be6),
	.w6(32'h39aab7aa),
	.w7(32'h38977328),
	.w8(32'h3b940b0b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64be95),
	.w1(32'h3b6722ca),
	.w2(32'h3b1bc02f),
	.w3(32'h3b1164fa),
	.w4(32'h3b00c498),
	.w5(32'h3b120825),
	.w6(32'h3b754214),
	.w7(32'h3b353e07),
	.w8(32'h3a8e6fe4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b65691),
	.w1(32'h3af39b00),
	.w2(32'h3b327aa6),
	.w3(32'hba347ec0),
	.w4(32'h3a4edaa6),
	.w5(32'h3b171c7e),
	.w6(32'h3952f66e),
	.w7(32'h3ab4033f),
	.w8(32'h3b84b5c5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad85886),
	.w1(32'h3ae9b300),
	.w2(32'h3ab2907a),
	.w3(32'h3a9d3d63),
	.w4(32'h3a45c730),
	.w5(32'h3a93e076),
	.w6(32'h3b10a13a),
	.w7(32'h3ac6d885),
	.w8(32'h3ba718cb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ef6f),
	.w1(32'h3aff8c63),
	.w2(32'h3bc394bd),
	.w3(32'h399ea53a),
	.w4(32'h3a8270fc),
	.w5(32'h3bd56bfd),
	.w6(32'h3b97a587),
	.w7(32'h3bc05ce2),
	.w8(32'h3b890bd3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914277c),
	.w1(32'h399e6e6a),
	.w2(32'h38f35e1b),
	.w3(32'h3a438c3d),
	.w4(32'hb8bb6f8f),
	.w5(32'h399dce6e),
	.w6(32'h3b234247),
	.w7(32'h3a5398ba),
	.w8(32'hbb0480de),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba029e73),
	.w1(32'hb9e6aa82),
	.w2(32'hb7ef27ed),
	.w3(32'hba54587a),
	.w4(32'hba4c16a7),
	.w5(32'hb902194c),
	.w6(32'hb9f685f5),
	.w7(32'hba0de185),
	.w8(32'h3a70cfbd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb4a8b),
	.w1(32'hbb0d4228),
	.w2(32'hbb0018fe),
	.w3(32'h3a732fa5),
	.w4(32'h3a96e065),
	.w5(32'h3abc4291),
	.w6(32'h39132025),
	.w7(32'h3a078884),
	.w8(32'h3b50f4de),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b765d1a),
	.w1(32'h3b923155),
	.w2(32'h3ba1a87d),
	.w3(32'h3adaa72c),
	.w4(32'h3b11e683),
	.w5(32'h3b1e9baf),
	.w6(32'h3b6efe37),
	.w7(32'h3b72e696),
	.w8(32'h3b987ee3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b070c52),
	.w1(32'h3ba40be5),
	.w2(32'h3bd0b3fc),
	.w3(32'h3aae89b2),
	.w4(32'h3b263d63),
	.w5(32'h3babc18a),
	.w6(32'h3b27bc34),
	.w7(32'h3b20fded),
	.w8(32'h3bfd8375),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef1b71),
	.w1(32'h3ba2535c),
	.w2(32'h3c1d09dd),
	.w3(32'h3ba42f61),
	.w4(32'h3bceaf65),
	.w5(32'h3c1ab7db),
	.w6(32'h3bc454bd),
	.w7(32'h3b84a76d),
	.w8(32'h3c2f83f9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76897e),
	.w1(32'h3b6606e5),
	.w2(32'h3be99e50),
	.w3(32'hbb0104b1),
	.w4(32'h3aca01ed),
	.w5(32'h3b508d17),
	.w6(32'hb930de41),
	.w7(32'h3b44af27),
	.w8(32'h3bd70610),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980b41e),
	.w1(32'h3b532273),
	.w2(32'h3bc02303),
	.w3(32'hba11734d),
	.w4(32'h38dcfc19),
	.w5(32'h3b5c14e2),
	.w6(32'hba94a0fe),
	.w7(32'h39bc5fbe),
	.w8(32'h3bd5beb8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a97ca2),
	.w1(32'hbae1bd20),
	.w2(32'hbadf2891),
	.w3(32'hb8618b54),
	.w4(32'hbae9ed4b),
	.w5(32'hbb455057),
	.w6(32'h3adbe3df),
	.w7(32'h3b624c2a),
	.w8(32'h3b3dba1a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3441de),
	.w1(32'h3b05e738),
	.w2(32'h3ad4514c),
	.w3(32'h3b1ab6eb),
	.w4(32'h39e99c72),
	.w5(32'h3ac0f154),
	.w6(32'h3b5af77d),
	.w7(32'h3ad4db6a),
	.w8(32'h3a8cf25d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38018cbf),
	.w1(32'hbaae1475),
	.w2(32'hbaa0013b),
	.w3(32'h3723af35),
	.w4(32'hba837e9a),
	.w5(32'hbabce2ec),
	.w6(32'hb742cb2a),
	.w7(32'h3a83ca3e),
	.w8(32'h3b8b2f36),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992a7c4),
	.w1(32'hbac51592),
	.w2(32'hba3beffb),
	.w3(32'h393ca24c),
	.w4(32'hbadcc786),
	.w5(32'hbb316e38),
	.w6(32'h3b0567a0),
	.w7(32'h3b6cf16d),
	.w8(32'h3b9437d8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f920fc),
	.w1(32'hba27f5b6),
	.w2(32'hb93dd66d),
	.w3(32'h38c1cc54),
	.w4(32'hb9e43041),
	.w5(32'hba9ff8ee),
	.w6(32'h3af870ac),
	.w7(32'h3b68756e),
	.w8(32'h3b46d1ef),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f90d),
	.w1(32'h391c9507),
	.w2(32'h37a70d9a),
	.w3(32'h3a207fda),
	.w4(32'hb7a851b8),
	.w5(32'hba48b8aa),
	.w6(32'h3a8c2440),
	.w7(32'h3abf9667),
	.w8(32'h3a8622c6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d578a5),
	.w1(32'hbab26bd9),
	.w2(32'h3abe1c15),
	.w3(32'hbaff1168),
	.w4(32'hbb650657),
	.w5(32'h3b178a9d),
	.w6(32'hbb245a85),
	.w7(32'hbb0bf7a6),
	.w8(32'h3b26f50e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eceaf),
	.w1(32'h3b0db3dd),
	.w2(32'h3b6a89cb),
	.w3(32'h3a281866),
	.w4(32'h3a959b82),
	.w5(32'h3b28282c),
	.w6(32'h3aef9e08),
	.w7(32'h3ae45c72),
	.w8(32'h3b411c85),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3bc15),
	.w1(32'hba5077be),
	.w2(32'hba6aaa19),
	.w3(32'hb9cc3028),
	.w4(32'hb73c75c0),
	.w5(32'h39e0a55a),
	.w6(32'h3b5ad041),
	.w7(32'h3b2b9064),
	.w8(32'h3b0e3044),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f854),
	.w1(32'hbb579e63),
	.w2(32'hbade4e1b),
	.w3(32'hbb31483d),
	.w4(32'hbb48a8e0),
	.w5(32'hbb5ebe93),
	.w6(32'hba819c0f),
	.w7(32'h3a0e25dd),
	.w8(32'h3ad3f39c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f58b4),
	.w1(32'h3b8fe232),
	.w2(32'h3bec95ea),
	.w3(32'h39d6b0d1),
	.w4(32'h3b2597c2),
	.w5(32'h3be29af1),
	.w6(32'h3b4f4b69),
	.w7(32'h3ba756dc),
	.w8(32'h3bed2991),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387cffd6),
	.w1(32'h3ab00d57),
	.w2(32'h3ab0e99d),
	.w3(32'h396a36c3),
	.w4(32'h3ab7197c),
	.w5(32'h3b1a5fab),
	.w6(32'h3a12a31a),
	.w7(32'h39eb28a1),
	.w8(32'h3b9074ed),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfc1ed),
	.w1(32'h3a9b2560),
	.w2(32'h3b098235),
	.w3(32'h3b108d33),
	.w4(32'h3a61d356),
	.w5(32'h3b55377d),
	.w6(32'h3b9f35b7),
	.w7(32'h3b8eb70a),
	.w8(32'h3b1a16d3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06426b),
	.w1(32'h3ab6f0a9),
	.w2(32'h3a6a5f54),
	.w3(32'h3ad30769),
	.w4(32'h37f55df2),
	.w5(32'h3a1952c4),
	.w6(32'h3b219fc4),
	.w7(32'h3a78d00a),
	.w8(32'h3aba3a68),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a045985),
	.w1(32'hb9f6bc75),
	.w2(32'hb9e47f3a),
	.w3(32'hb8108e19),
	.w4(32'hba040453),
	.w5(32'hba8126df),
	.w6(32'h3a0fe6b8),
	.w7(32'h3acdfef3),
	.w8(32'h3b2cf825),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874be1),
	.w1(32'h3b8244cb),
	.w2(32'h3b5a2c2a),
	.w3(32'h3b5ca84f),
	.w4(32'h3b20ceac),
	.w5(32'h3b175148),
	.w6(32'h3b97c03b),
	.w7(32'h3b6fc902),
	.w8(32'h3b4f6ae7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed619),
	.w1(32'h3ae396f0),
	.w2(32'h3b190181),
	.w3(32'h3af869eb),
	.w4(32'h3a123f4e),
	.w5(32'h3b56e0a7),
	.w6(32'h3b98d946),
	.w7(32'h3b4909a7),
	.w8(32'h3a11c7be),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9673c),
	.w1(32'hbaabc5a1),
	.w2(32'hb87952ba),
	.w3(32'hbb2f903a),
	.w4(32'hbb76959d),
	.w5(32'hbb049336),
	.w6(32'hb955d529),
	.w7(32'h39fc50f4),
	.w8(32'h3b51b6db),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76233),
	.w1(32'hbac9d69b),
	.w2(32'hba864a88),
	.w3(32'hba3a7c1e),
	.w4(32'hbac1423b),
	.w5(32'hbaa5078f),
	.w6(32'h3981bc36),
	.w7(32'h3a292951),
	.w8(32'hb926407a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225ea1),
	.w1(32'h3a2cfa8b),
	.w2(32'h3b4687ed),
	.w3(32'hbb86d1c3),
	.w4(32'hb9b5cd64),
	.w5(32'h3a07aff2),
	.w6(32'hbb34f40d),
	.w7(32'hb8fdf160),
	.w8(32'hbb284a4e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c6b2a),
	.w1(32'hb81ccfdb),
	.w2(32'h3b3a8557),
	.w3(32'hbb7f855f),
	.w4(32'hb980368c),
	.w5(32'h3a456981),
	.w6(32'h380a7d40),
	.w7(32'h393776dd),
	.w8(32'h3a7b5843),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa09a04),
	.w1(32'hbaa71e36),
	.w2(32'hb8c6db74),
	.w3(32'hba46dd8d),
	.w4(32'hba683f80),
	.w5(32'h39c1f1e4),
	.w6(32'hba66ada5),
	.w7(32'hba340caa),
	.w8(32'h3a9422cc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f06a63),
	.w1(32'hbaabdda0),
	.w2(32'hba5515f5),
	.w3(32'h394ad987),
	.w4(32'hba942a91),
	.w5(32'hba57724d),
	.w6(32'h38dcb412),
	.w7(32'hba1e93f9),
	.w8(32'h39f80a6d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fd3b5),
	.w1(32'h3b26a4ab),
	.w2(32'h3af9fcb9),
	.w3(32'h3b9f7bff),
	.w4(32'h3b2de26d),
	.w5(32'h3b00d086),
	.w6(32'h3b497e29),
	.w7(32'h3b428fd8),
	.w8(32'h3ad798b8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003a0d),
	.w1(32'hba08b826),
	.w2(32'hbb31b95d),
	.w3(32'hbabc40c2),
	.w4(32'h3937064f),
	.w5(32'h3a626507),
	.w6(32'hbb098f39),
	.w7(32'hbb1102c0),
	.w8(32'h3b289527),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba746a1a),
	.w1(32'hbb01584f),
	.w2(32'h3a8f8153),
	.w3(32'hba23e66f),
	.w4(32'hbacc32ff),
	.w5(32'h3a789379),
	.w6(32'hbaa9e2f8),
	.w7(32'hba84e583),
	.w8(32'h3b124ada),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0101da),
	.w1(32'hbb7d29ef),
	.w2(32'hbb33a042),
	.w3(32'hbb1efe4d),
	.w4(32'hbb7a474b),
	.w5(32'hbb247162),
	.w6(32'hb9f77ea6),
	.w7(32'hbacb336a),
	.w8(32'hbaa8a563),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc7792),
	.w1(32'hb8bc189f),
	.w2(32'h3826da71),
	.w3(32'h3a0eb3a0),
	.w4(32'h3919d8f7),
	.w5(32'h384e7dab),
	.w6(32'hb8bf8126),
	.w7(32'h3a0953cb),
	.w8(32'hb9fe4195),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce86c8),
	.w1(32'hb9a9e583),
	.w2(32'hb9767f8b),
	.w3(32'h396a5224),
	.w4(32'h3966b6da),
	.w5(32'hb9af5a78),
	.w6(32'hb97d6192),
	.w7(32'h3932cb0e),
	.w8(32'hba1d23a1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb9ddf),
	.w1(32'h3a8976ca),
	.w2(32'h3a01bc57),
	.w3(32'h3ae3486e),
	.w4(32'h3a6c8837),
	.w5(32'h39baabdd),
	.w6(32'h38d6689c),
	.w7(32'h39e6f7b4),
	.w8(32'h3a86c251),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58295f),
	.w1(32'hbb225031),
	.w2(32'hbb0c1ab2),
	.w3(32'h3615ee41),
	.w4(32'hba19234f),
	.w5(32'hb954826b),
	.w6(32'hb9b59a82),
	.w7(32'hbafe4bf6),
	.w8(32'h3ac599f0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82da99c),
	.w1(32'h39c6d032),
	.w2(32'h3af73289),
	.w3(32'h39659336),
	.w4(32'h3a888662),
	.w5(32'h3b11b733),
	.w6(32'h3a06620b),
	.w7(32'h3abf51ed),
	.w8(32'h3b37dee6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed5b52),
	.w1(32'hba9b9843),
	.w2(32'hbb5cf1ca),
	.w3(32'h38da656f),
	.w4(32'hb9a4b49d),
	.w5(32'hbb1a0372),
	.w6(32'hba5f52a2),
	.w7(32'hbb56e684),
	.w8(32'hba8120e6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42fc52),
	.w1(32'hbab1af60),
	.w2(32'hbb252817),
	.w3(32'hba4d1fda),
	.w4(32'hb942bc96),
	.w5(32'hba80fa1b),
	.w6(32'hbadec67f),
	.w7(32'hbaaba19b),
	.w8(32'hb98906f2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0988cc),
	.w1(32'hb7e430b0),
	.w2(32'hba9f1bc7),
	.w3(32'h3a88e5cf),
	.w4(32'hba790fce),
	.w5(32'h3a1f7ca5),
	.w6(32'h3a06a9d7),
	.w7(32'h3a380fd3),
	.w8(32'h3a6f1217),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dab79c),
	.w1(32'hbb40a4a4),
	.w2(32'hbb0d92a8),
	.w3(32'h399bd5fc),
	.w4(32'hba31eb53),
	.w5(32'hbab6aadd),
	.w6(32'hbab6ebec),
	.w7(32'hbb14ba6a),
	.w8(32'h3a270c10),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af7ee4),
	.w1(32'hb9e11701),
	.w2(32'hb8939bd3),
	.w3(32'hb9c6f3fd),
	.w4(32'hb997bc86),
	.w5(32'h392d3682),
	.w6(32'h3aebdc0f),
	.w7(32'h3b096efb),
	.w8(32'hbad6da87),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadde6ff),
	.w1(32'hbb286d3d),
	.w2(32'hbb36b35e),
	.w3(32'hbae06794),
	.w4(32'hbb1df8ee),
	.w5(32'hbae46b15),
	.w6(32'hbb0b6848),
	.w7(32'hbb56a01f),
	.w8(32'hb81eba87),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8ba73),
	.w1(32'h3ad7e08d),
	.w2(32'hb82a1817),
	.w3(32'h3b754914),
	.w4(32'h3b714a47),
	.w5(32'h3b35287e),
	.w6(32'h3b0ca1e9),
	.w7(32'hb92e1e4d),
	.w8(32'h3b0a422d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab61ae0),
	.w1(32'h3af7723e),
	.w2(32'h3a8cd1d8),
	.w3(32'h3b204512),
	.w4(32'h3ade8c13),
	.w5(32'h3ad4dea2),
	.w6(32'h388a5fe3),
	.w7(32'h394e524e),
	.w8(32'hb8451058),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c90a7),
	.w1(32'hba26be6a),
	.w2(32'hba29958d),
	.w3(32'hba20b07b),
	.w4(32'hba9048b1),
	.w5(32'hba182853),
	.w6(32'hb9d3e1e8),
	.w7(32'hb7ae2817),
	.w8(32'h3957779c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d72ea),
	.w1(32'hbb8a0303),
	.w2(32'hba929ec9),
	.w3(32'hbae65e44),
	.w4(32'hbb15f05b),
	.w5(32'hbb1eb459),
	.w6(32'hb9ba6200),
	.w7(32'h3945d924),
	.w8(32'hb9c92bf1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule