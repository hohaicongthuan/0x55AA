module layer_10_featuremap_454(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f781d),
	.w1(32'h3bb17120),
	.w2(32'h3a19cda6),
	.w3(32'hba358df3),
	.w4(32'h3b83913b),
	.w5(32'hb9deec92),
	.w6(32'h39975126),
	.w7(32'h3baa493b),
	.w8(32'h3bdf45f7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821f04),
	.w1(32'hb9924393),
	.w2(32'hb7eb50f2),
	.w3(32'h39a1ecfa),
	.w4(32'hbc04ae6b),
	.w5(32'hbc204420),
	.w6(32'h3c7899f7),
	.w7(32'h3b8b2534),
	.w8(32'h3b1e4e68),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93441d),
	.w1(32'hbbb8e31a),
	.w2(32'h3bdfcb1b),
	.w3(32'h3c8beb4b),
	.w4(32'hbada8cad),
	.w5(32'h3c98b11e),
	.w6(32'h3baf5466),
	.w7(32'h3b6c30e6),
	.w8(32'hbb28ec6b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7cb3),
	.w1(32'hb8c4f1d6),
	.w2(32'hbb875e42),
	.w3(32'h3c420c5a),
	.w4(32'hbc2f7aae),
	.w5(32'hbc050473),
	.w6(32'hbbd8b0a9),
	.w7(32'h3c119dc0),
	.w8(32'h3c21d965),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b434),
	.w1(32'hbbaa3918),
	.w2(32'hbb97c3b6),
	.w3(32'h3c251ab7),
	.w4(32'hba785f8d),
	.w5(32'h3af69e10),
	.w6(32'h3c08509a),
	.w7(32'hbbb2e9f4),
	.w8(32'h3b833097),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb336bdb),
	.w1(32'h3be5e4f0),
	.w2(32'h3c1517d8),
	.w3(32'h3b94f7af),
	.w4(32'h3c065cf8),
	.w5(32'hbab2f2be),
	.w6(32'h3bedce96),
	.w7(32'h3b2cb8ca),
	.w8(32'h3b0b1894),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c2e5),
	.w1(32'hbbcdb499),
	.w2(32'h3ba89888),
	.w3(32'h3bb5dbc5),
	.w4(32'h3be8fa97),
	.w5(32'h3ca21cdc),
	.w6(32'hbc20b2a2),
	.w7(32'hbca960e6),
	.w8(32'hbc1c0ae8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12d2df),
	.w1(32'h3c9f03bd),
	.w2(32'h3cc0a103),
	.w3(32'h3c06ad7a),
	.w4(32'hbbc2333a),
	.w5(32'hbc00fd73),
	.w6(32'hbd091b28),
	.w7(32'hbd2d60f0),
	.w8(32'hbd898ae3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd6f5b7),
	.w1(32'hbabe361b),
	.w2(32'hbb5cc57b),
	.w3(32'hbbd8eabe),
	.w4(32'h3c2db6cc),
	.w5(32'h3af18abd),
	.w6(32'hbd1b551a),
	.w7(32'hbba3dc43),
	.w8(32'hbc344c1b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44463d),
	.w1(32'hbb00ff52),
	.w2(32'hbb1577cf),
	.w3(32'hbc6e489b),
	.w4(32'h3ba262c6),
	.w5(32'h3b5306f8),
	.w6(32'hbc88feaf),
	.w7(32'hba8bcd47),
	.w8(32'h3bb6ff39),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a30b),
	.w1(32'hbc01137d),
	.w2(32'h3ae652b1),
	.w3(32'h3c45f1bf),
	.w4(32'hbc56cbd9),
	.w5(32'h3b5284b4),
	.w6(32'hbb88d89a),
	.w7(32'hbc9b6522),
	.w8(32'hbb892749),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896ab9),
	.w1(32'h3c1da823),
	.w2(32'h3c12f8c3),
	.w3(32'hbbb00f1d),
	.w4(32'h3c45a7c3),
	.w5(32'h3c7f0d33),
	.w6(32'hbc7b20cc),
	.w7(32'hbb78b611),
	.w8(32'h3c301e4c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5636e),
	.w1(32'hba879dc6),
	.w2(32'hbb8ac191),
	.w3(32'h3bfd59dc),
	.w4(32'hbb85777d),
	.w5(32'hbc43bc24),
	.w6(32'hbb4b3139),
	.w7(32'h3b748b95),
	.w8(32'h3ad06da6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bccac),
	.w1(32'hbc240479),
	.w2(32'hbcad8c25),
	.w3(32'h3c9a48b8),
	.w4(32'hbb024d5f),
	.w5(32'hbc29f360),
	.w6(32'h3aa50aea),
	.w7(32'h3b1541c9),
	.w8(32'h3c9d4209),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a0612),
	.w1(32'hbc031884),
	.w2(32'hbc15a35b),
	.w3(32'hbc3c5546),
	.w4(32'hba69627e),
	.w5(32'h3a5a181b),
	.w6(32'h3c37dc30),
	.w7(32'h3ab5512c),
	.w8(32'h3bf8604e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801868),
	.w1(32'h3c473e7e),
	.w2(32'hb93eebad),
	.w3(32'hbb840c6b),
	.w4(32'h3bc630b0),
	.w5(32'h3acb144b),
	.w6(32'h3bbd9d9e),
	.w7(32'h3b6a1545),
	.w8(32'hbbb87cfa),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cb87f),
	.w1(32'hb9a1f54c),
	.w2(32'h3a3bcb60),
	.w3(32'hbbf95770),
	.w4(32'h3b43686c),
	.w5(32'h3acfcd4e),
	.w6(32'hbb091a95),
	.w7(32'hbb946da0),
	.w8(32'hbb25508f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86ccf),
	.w1(32'h3bd4af7f),
	.w2(32'hbb0fb2d1),
	.w3(32'h3bde3d69),
	.w4(32'h3bee3cec),
	.w5(32'hba54b542),
	.w6(32'hbc80cc9f),
	.w7(32'hbbe09598),
	.w8(32'hbc07bc44),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a484ef8),
	.w1(32'hbba60f5b),
	.w2(32'hb930c2d4),
	.w3(32'hb8b99b2b),
	.w4(32'h3c0c83c2),
	.w5(32'h3c875b73),
	.w6(32'hbc1461bc),
	.w7(32'hbc455c3d),
	.w8(32'hbbed0144),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f7e3),
	.w1(32'hbb8e928a),
	.w2(32'h3b44ab08),
	.w3(32'hba5d8c2a),
	.w4(32'h3976a455),
	.w5(32'h3a693fcf),
	.w6(32'hbb2fc09c),
	.w7(32'hbc161c35),
	.w8(32'h3befa184),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05dae1),
	.w1(32'h3c1a219b),
	.w2(32'h3c66752a),
	.w3(32'hbb27f542),
	.w4(32'h3c85ff25),
	.w5(32'h3c8e9299),
	.w6(32'h39506b6a),
	.w7(32'h3b3a3d19),
	.w8(32'h3b917fab),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474390),
	.w1(32'hbbc1030c),
	.w2(32'h3b2ad2be),
	.w3(32'hbab49ecf),
	.w4(32'h3a89a33f),
	.w5(32'h397022ac),
	.w6(32'hb9da6429),
	.w7(32'h3b4ee2ea),
	.w8(32'h3bf85338),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77dd67),
	.w1(32'h3b012f7c),
	.w2(32'h3a147b8e),
	.w3(32'h3bcb419c),
	.w4(32'h3baefb50),
	.w5(32'hba1dded3),
	.w6(32'hbb270d89),
	.w7(32'hbb905258),
	.w8(32'hbae31363),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec29c4),
	.w1(32'h3ba1f791),
	.w2(32'hbb969981),
	.w3(32'h3c0bb235),
	.w4(32'h3c474fea),
	.w5(32'h3bf48952),
	.w6(32'h3ab1bfad),
	.w7(32'hbb12916d),
	.w8(32'hbc2cd859),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd9419),
	.w1(32'hbc3fa443),
	.w2(32'h3b59c4f1),
	.w3(32'h3cb63f9a),
	.w4(32'hbc159545),
	.w5(32'hbb6abac0),
	.w6(32'h3c726787),
	.w7(32'hbbe9a60d),
	.w8(32'h3a97f8f2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587803),
	.w1(32'h3c54b375),
	.w2(32'h3c204fc6),
	.w3(32'hbc068cd4),
	.w4(32'h3b9f816c),
	.w5(32'h3aec00bc),
	.w6(32'hbb777121),
	.w7(32'h3c095926),
	.w8(32'h3bb6ac8b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b86e),
	.w1(32'hbc286a10),
	.w2(32'hbb1f0f35),
	.w3(32'hbb09269c),
	.w4(32'hbb2c5839),
	.w5(32'h3b96fc7a),
	.w6(32'h3baa04cb),
	.w7(32'hbb51a146),
	.w8(32'h3b6d08b3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20d9d9),
	.w1(32'hbc18a97f),
	.w2(32'hb8e760f0),
	.w3(32'h3b8decc5),
	.w4(32'hbbb7c91b),
	.w5(32'hbc0dbeb2),
	.w6(32'h3c8850bd),
	.w7(32'h3c1c6f5a),
	.w8(32'h3ba2b38b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3bdf8),
	.w1(32'h3aa163de),
	.w2(32'h3b5aa088),
	.w3(32'h3a87ba30),
	.w4(32'h3b70182a),
	.w5(32'hbbba5e4b),
	.w6(32'hba1ae7e1),
	.w7(32'h3bb8d260),
	.w8(32'hbb7f351d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01c34d),
	.w1(32'hbb939629),
	.w2(32'hbb846f87),
	.w3(32'h3bf38dda),
	.w4(32'h3aa097ae),
	.w5(32'h3a6cea10),
	.w6(32'h3c463673),
	.w7(32'h3c300641),
	.w8(32'h3c18334c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb633d27),
	.w1(32'h3b88ab97),
	.w2(32'hbae18cbe),
	.w3(32'hbbc474db),
	.w4(32'hba50a288),
	.w5(32'hbc2a08c1),
	.w6(32'hbade008e),
	.w7(32'hbb08b16d),
	.w8(32'h3b0e7a81),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad85da4),
	.w1(32'hbbd0087b),
	.w2(32'hbc5609a3),
	.w3(32'hba318405),
	.w4(32'hbc2c441b),
	.w5(32'hbca0d401),
	.w6(32'hbb41ce50),
	.w7(32'hbc2a4cc3),
	.w8(32'hbc9e7d30),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ce957),
	.w1(32'hbc1ca8fe),
	.w2(32'hbbc8314e),
	.w3(32'hb9719a9e),
	.w4(32'hbc0f3739),
	.w5(32'hbaea7b16),
	.w6(32'hbca9d21c),
	.w7(32'hbc01e5a7),
	.w8(32'hbba3867f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19a087),
	.w1(32'h3b28be5b),
	.w2(32'h3c0146fa),
	.w3(32'hba6082de),
	.w4(32'h3b9d32bf),
	.w5(32'h3aa58e44),
	.w6(32'hba29d7ce),
	.w7(32'h3b487261),
	.w8(32'hbbffd8e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf68fe7),
	.w1(32'hbc57bef8),
	.w2(32'hbc8e0fcd),
	.w3(32'hbbed5f9d),
	.w4(32'hbc1745b3),
	.w5(32'hbae3dfb3),
	.w6(32'hbb8dd94e),
	.w7(32'h3ca14e72),
	.w8(32'h3d00ebc9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c73b2),
	.w1(32'hbb3439bd),
	.w2(32'hbb9a4ede),
	.w3(32'hbc12bd54),
	.w4(32'hbb5c7a9b),
	.w5(32'hbb829642),
	.w6(32'h3c22bfb3),
	.w7(32'hbb347bab),
	.w8(32'hb98baab0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11b411),
	.w1(32'hbb70a6d8),
	.w2(32'h3c938177),
	.w3(32'hba25d05a),
	.w4(32'h3c81450e),
	.w5(32'h3c5ad523),
	.w6(32'h3bc52d4e),
	.w7(32'hbc2351b7),
	.w8(32'h3c74e438),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f7204),
	.w1(32'hbc65b8a6),
	.w2(32'hbb996d4e),
	.w3(32'h3b350753),
	.w4(32'hbc751331),
	.w5(32'hbc50271e),
	.w6(32'h3c8bb88e),
	.w7(32'hba937fcc),
	.w8(32'hbc2a77ff),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a137b),
	.w1(32'hbc4918ce),
	.w2(32'hba1e1fe8),
	.w3(32'h3cbee6d7),
	.w4(32'hbbb4f1e8),
	.w5(32'h3c047fd6),
	.w6(32'h3c554120),
	.w7(32'hba9d6eee),
	.w8(32'h3bdb0ae7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bb19c),
	.w1(32'h3af8ad63),
	.w2(32'h3c040bc3),
	.w3(32'hbc308a66),
	.w4(32'hbb888a1b),
	.w5(32'h3a7d7590),
	.w6(32'h3bab7d41),
	.w7(32'h39bc7317),
	.w8(32'h3b12ad68),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b36a39),
	.w1(32'h3baf5e70),
	.w2(32'h3b21af33),
	.w3(32'h3bedbf33),
	.w4(32'hbb33646c),
	.w5(32'hbbfc9a3f),
	.w6(32'h3a215976),
	.w7(32'hbafb54de),
	.w8(32'h3ab4111d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f22d),
	.w1(32'hbc49594d),
	.w2(32'h3b02f533),
	.w3(32'hbc64802e),
	.w4(32'hbbdafa72),
	.w5(32'h3bfb0ec9),
	.w6(32'hbc1d3f54),
	.w7(32'hbc29752a),
	.w8(32'h3bd2c6d6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f853),
	.w1(32'hba874b1f),
	.w2(32'hbc00f5ec),
	.w3(32'h3b0f256d),
	.w4(32'hbbd1dd46),
	.w5(32'hbca37ce5),
	.w6(32'h3b3652fa),
	.w7(32'h398c54bf),
	.w8(32'hbbfd85e2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62815f),
	.w1(32'h3c20cd73),
	.w2(32'h3b7ef109),
	.w3(32'h3c4be44d),
	.w4(32'hbb18136a),
	.w5(32'h3b915524),
	.w6(32'hbc00ac86),
	.w7(32'h3b5a2f1d),
	.w8(32'h3bdc1bfc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c03a1),
	.w1(32'hbb705e00),
	.w2(32'hb983cd34),
	.w3(32'hbb36f1dd),
	.w4(32'h3bbdb363),
	.w5(32'hb9f95c60),
	.w6(32'h3bf07b25),
	.w7(32'hbb08af3c),
	.w8(32'hbbf21755),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c379ddf),
	.w1(32'h3c03f5ca),
	.w2(32'h3b588550),
	.w3(32'hbb586688),
	.w4(32'h3a95d5ca),
	.w5(32'h3b9501d6),
	.w6(32'h3b2d1903),
	.w7(32'hbb3650a4),
	.w8(32'hbbf5995f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc944f9),
	.w1(32'hbbee8ae3),
	.w2(32'hbbbae8df),
	.w3(32'h3b95d42d),
	.w4(32'hbb3d0dc0),
	.w5(32'hba28f557),
	.w6(32'h3b5418d2),
	.w7(32'h3b0a7cf5),
	.w8(32'h3c2375ed),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7715),
	.w1(32'h3a7fdd2b),
	.w2(32'h39cfb1df),
	.w3(32'hbbacf6be),
	.w4(32'h3bfbb97c),
	.w5(32'hb92f0595),
	.w6(32'hbc97c2ab),
	.w7(32'hbbafbb8f),
	.w8(32'hbbfc1d63),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee94ef),
	.w1(32'h3ba72b88),
	.w2(32'h3b802c00),
	.w3(32'hbc4639df),
	.w4(32'h3c4e834c),
	.w5(32'h3c9bb949),
	.w6(32'hbc282036),
	.w7(32'hbb26ad7f),
	.w8(32'h3b41c1bc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15103a),
	.w1(32'h3adee467),
	.w2(32'hbb8c8345),
	.w3(32'hbc3b811c),
	.w4(32'hbc2c8aa1),
	.w5(32'hbb2e3bce),
	.w6(32'hbc119e8f),
	.w7(32'hbbbb6d3e),
	.w8(32'hbb919c85),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8f43b),
	.w1(32'hbb05165c),
	.w2(32'hbbeacb38),
	.w3(32'h3c2cfd15),
	.w4(32'h3b2bad90),
	.w5(32'hbc08579f),
	.w6(32'h398bdb43),
	.w7(32'hbb217119),
	.w8(32'hbc067728),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375b1a),
	.w1(32'h39c2cdf3),
	.w2(32'hba592220),
	.w3(32'h3bcad6ce),
	.w4(32'hbbdd6ad4),
	.w5(32'hbbf684d2),
	.w6(32'hba226f6c),
	.w7(32'hbb8b2ab9),
	.w8(32'hbc6727fc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827f207),
	.w1(32'h3c7a737f),
	.w2(32'h3c363279),
	.w3(32'hbbd6c73b),
	.w4(32'h3c3f471d),
	.w5(32'h3b9f10f7),
	.w6(32'hbc02e513),
	.w7(32'hbc27bb22),
	.w8(32'hbc84f606),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c204b62),
	.w1(32'h3c938a24),
	.w2(32'h3c4b6e63),
	.w3(32'h3b17c3f8),
	.w4(32'h3c100dca),
	.w5(32'h3c07f2b1),
	.w6(32'hbcf18db5),
	.w7(32'hbc9a6305),
	.w8(32'hbcae5977),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c346809),
	.w1(32'hbb7ebe53),
	.w2(32'hbaf4a80a),
	.w3(32'h3b9a3edb),
	.w4(32'hbb11a158),
	.w5(32'h3b8cb31e),
	.w6(32'hbcab504c),
	.w7(32'hbbaab4dc),
	.w8(32'h3bbccb68),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d64f8),
	.w1(32'h3ae0bd3c),
	.w2(32'h3b2f1e62),
	.w3(32'h3c07875e),
	.w4(32'hbba728c2),
	.w5(32'hbbdbbed1),
	.w6(32'h3b014189),
	.w7(32'hbb617c12),
	.w8(32'hbba6938f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be01910),
	.w1(32'hbba1d6c7),
	.w2(32'hbb901fa8),
	.w3(32'h3c8650ce),
	.w4(32'hbc0edf50),
	.w5(32'hbc1d16a5),
	.w6(32'hbbb97346),
	.w7(32'hbb4b2847),
	.w8(32'hbba5138f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb455839),
	.w1(32'h3b75728b),
	.w2(32'h3b81b426),
	.w3(32'hbb4bd4e2),
	.w4(32'hbaa0df57),
	.w5(32'hbabb2d57),
	.w6(32'hbb85d8e2),
	.w7(32'h3aa43d65),
	.w8(32'h3ad48020),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae79169),
	.w1(32'hbbde1657),
	.w2(32'h3a0226ed),
	.w3(32'hbba31673),
	.w4(32'hbb96c936),
	.w5(32'h3b4c2841),
	.w6(32'hb9f40833),
	.w7(32'hbb682d53),
	.w8(32'h3b70fb8a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14ed75),
	.w1(32'h3be56504),
	.w2(32'h3c08cdb0),
	.w3(32'h3c0e7c72),
	.w4(32'h3c31f9cc),
	.w5(32'h3a6e1d42),
	.w6(32'h3a9a9c43),
	.w7(32'hbae3ac3c),
	.w8(32'h3b959c01),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b1556),
	.w1(32'hba618f6a),
	.w2(32'h3c4aaa99),
	.w3(32'hb92703ca),
	.w4(32'h39f165b0),
	.w5(32'h3c01fb45),
	.w6(32'hbb1b7c22),
	.w7(32'hbb8176a2),
	.w8(32'hbb581dbf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47a56d),
	.w1(32'hbc16e373),
	.w2(32'hbc4db598),
	.w3(32'hbad8a232),
	.w4(32'hbb4c1ade),
	.w5(32'h3a6266df),
	.w6(32'hbbca6c89),
	.w7(32'hbbff67f0),
	.w8(32'h3b148557),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23a7a0),
	.w1(32'hbbd78010),
	.w2(32'hbb7edc6e),
	.w3(32'hbc2e5400),
	.w4(32'hbc2c2006),
	.w5(32'hbbb3b02c),
	.w6(32'h3a7d35f0),
	.w7(32'hbb35cea1),
	.w8(32'hb982a6a4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3b5f),
	.w1(32'h3a2dfca2),
	.w2(32'hbaf9330e),
	.w3(32'h3c922f92),
	.w4(32'hba935c1f),
	.w5(32'hbb9307fc),
	.w6(32'h3c075e16),
	.w7(32'h3bcafbb9),
	.w8(32'h3b9f1f1f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57bfc7),
	.w1(32'h3bc91c9b),
	.w2(32'h3af5ad41),
	.w3(32'h3b3886d3),
	.w4(32'h3b9e4d90),
	.w5(32'hbaed5cc9),
	.w6(32'h3b015aa1),
	.w7(32'h3b49f192),
	.w8(32'hbb85c002),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb9a0),
	.w1(32'hbb70def3),
	.w2(32'hba61ae92),
	.w3(32'h3a1bfab4),
	.w4(32'h39cbd394),
	.w5(32'h3c785c51),
	.w6(32'hbb926729),
	.w7(32'hbc064f13),
	.w8(32'hb9357707),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891b43),
	.w1(32'h3a47d93b),
	.w2(32'hbbf48b7c),
	.w3(32'h3bc86a8e),
	.w4(32'h3b70c53c),
	.w5(32'hbcc56cb9),
	.w6(32'hbbfac3c7),
	.w7(32'h3bf40553),
	.w8(32'h3c106dc2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049596),
	.w1(32'hbabc4e6b),
	.w2(32'hbadf76d8),
	.w3(32'hbcaa3296),
	.w4(32'h3abea13c),
	.w5(32'hbbfb9fa5),
	.w6(32'hbc656b41),
	.w7(32'hbc17d958),
	.w8(32'h3bace847),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e92c),
	.w1(32'h3bf391b0),
	.w2(32'hba871b6d),
	.w3(32'hbc5dfb75),
	.w4(32'hbac98d00),
	.w5(32'hbbb74be0),
	.w6(32'hbba60af3),
	.w7(32'h3a8d198b),
	.w8(32'hbb8d1695),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139eb9),
	.w1(32'hbc16ee56),
	.w2(32'hbb1032c5),
	.w3(32'h3c96748c),
	.w4(32'hbbc485f7),
	.w5(32'h3b27f0d6),
	.w6(32'h3cc15a46),
	.w7(32'h39f019a9),
	.w8(32'h3bbe0043),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3f44a),
	.w1(32'h3b78e6eb),
	.w2(32'h3b8b8734),
	.w3(32'hbb8fdea1),
	.w4(32'h3bcb87ef),
	.w5(32'h375704e8),
	.w6(32'hb84ac69a),
	.w7(32'h39147e31),
	.w8(32'h3aa3adf8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86b2f51),
	.w1(32'h3b8167ad),
	.w2(32'h39e5f327),
	.w3(32'hbb8c03f2),
	.w4(32'h3bc3ba2d),
	.w5(32'hbb4cff7f),
	.w6(32'hbb8d9f17),
	.w7(32'h3b708ab4),
	.w8(32'h3b1e4957),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a9c06),
	.w1(32'hbba24a22),
	.w2(32'h3bb82155),
	.w3(32'hb95e2665),
	.w4(32'hbabf1f06),
	.w5(32'h3be1f34b),
	.w6(32'h3bdfcedf),
	.w7(32'hbb6cd0a9),
	.w8(32'h3b9b69b7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac64469),
	.w1(32'h3a627b93),
	.w2(32'hbae86f4a),
	.w3(32'hba845326),
	.w4(32'hba32b346),
	.w5(32'hbadb3796),
	.w6(32'h3a7b5187),
	.w7(32'hbaf3fbd1),
	.w8(32'hbb965343),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160bf2),
	.w1(32'hbae4d00e),
	.w2(32'h3af14152),
	.w3(32'h3b05de01),
	.w4(32'h3b8cd7a4),
	.w5(32'h3afe6389),
	.w6(32'hb903d6c0),
	.w7(32'h390cf8cd),
	.w8(32'h3b3572a4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037e4e),
	.w1(32'h3a0dfe2c),
	.w2(32'h3a711c7e),
	.w3(32'h3a487461),
	.w4(32'h3bb923c6),
	.w5(32'hbb06afed),
	.w6(32'hbb04ed31),
	.w7(32'hbae7f56a),
	.w8(32'h392aedc9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cb0a4),
	.w1(32'h3be94696),
	.w2(32'hbac0c829),
	.w3(32'h3b03c41d),
	.w4(32'h3bed39f6),
	.w5(32'hbb3af304),
	.w6(32'hbc6972e7),
	.w7(32'hbbe43bda),
	.w8(32'hbc199823),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa57564),
	.w1(32'h3a43404d),
	.w2(32'h3bb2cb21),
	.w3(32'h3ac0d2fc),
	.w4(32'h3b8c02ea),
	.w5(32'h3b9c325c),
	.w6(32'h3c13fa7a),
	.w7(32'h3bcaa3bd),
	.w8(32'h3b13920f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39caa5),
	.w1(32'h3ac1bc66),
	.w2(32'h370e10a0),
	.w3(32'hba8c3b74),
	.w4(32'h3b8ddb2e),
	.w5(32'hba49a466),
	.w6(32'hbbfae09f),
	.w7(32'h3b6e5398),
	.w8(32'hbb41023c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca931a),
	.w1(32'h398f04db),
	.w2(32'hbb6c034d),
	.w3(32'h3bac210a),
	.w4(32'h3aba9872),
	.w5(32'hbbd2f47d),
	.w6(32'h3b234386),
	.w7(32'h3b2bded5),
	.w8(32'h3a9afc7d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5cb1c),
	.w1(32'h3bb0c924),
	.w2(32'h3abdafa3),
	.w3(32'h3b9093fb),
	.w4(32'h3bb0f568),
	.w5(32'h3a3de625),
	.w6(32'h3bc28612),
	.w7(32'h3bf1b536),
	.w8(32'h3b3f053a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2b7a4),
	.w1(32'h3bb1d8e9),
	.w2(32'h3b58f381),
	.w3(32'h3c05cf47),
	.w4(32'h3b80a1f8),
	.w5(32'h3bbccfd3),
	.w6(32'h3b1f093c),
	.w7(32'h3968e037),
	.w8(32'h3b826c48),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1904c3),
	.w1(32'hbaf98bcf),
	.w2(32'hbab0b8fa),
	.w3(32'hba227b78),
	.w4(32'hbb30bcda),
	.w5(32'h3ae04240),
	.w6(32'hbb01b319),
	.w7(32'hba14dd7e),
	.w8(32'h3b492b8e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b635e),
	.w1(32'h3bb111dc),
	.w2(32'h3807d744),
	.w3(32'hbb1f9ac0),
	.w4(32'h3c46f343),
	.w5(32'h3be019e4),
	.w6(32'h3a0de150),
	.w7(32'h3be1d91f),
	.w8(32'h3c081f96),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943cfe),
	.w1(32'h3b2a95b4),
	.w2(32'h3a2b6e94),
	.w3(32'hbc202d65),
	.w4(32'h3b97109b),
	.w5(32'h3bb11c91),
	.w6(32'hbbb5ad0b),
	.w7(32'h3b003b9f),
	.w8(32'h3b042411),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12ef4d),
	.w1(32'h3a3b1c3f),
	.w2(32'h3c32ff80),
	.w3(32'hbaa39aee),
	.w4(32'hbb449205),
	.w5(32'h3cd0a642),
	.w6(32'h3b59902f),
	.w7(32'h3bb1dd93),
	.w8(32'h3ba651f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989dcfd),
	.w1(32'hbbfb34d1),
	.w2(32'hba9f0392),
	.w3(32'h3acc6c35),
	.w4(32'hbb3e5043),
	.w5(32'hbb3d54f0),
	.w6(32'h3b2a8ef1),
	.w7(32'h3ab8a6f2),
	.w8(32'hbb98e070),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399683c6),
	.w1(32'hbb094f4a),
	.w2(32'hbba94228),
	.w3(32'hba0f6c29),
	.w4(32'h39cbd7e1),
	.w5(32'hbbe13a12),
	.w6(32'h3bbf1fab),
	.w7(32'hba33d0e7),
	.w8(32'hbb835dba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b422c7c),
	.w1(32'h3a4af7a7),
	.w2(32'hbbb397e4),
	.w3(32'hbbf98e38),
	.w4(32'h3a86c1fd),
	.w5(32'hbbb0cf85),
	.w6(32'hbbcbe863),
	.w7(32'hba9b3a06),
	.w8(32'hbb0c7b56),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3fe12),
	.w1(32'h3bad266d),
	.w2(32'hbad99fc4),
	.w3(32'hb98e5122),
	.w4(32'hbba230bd),
	.w5(32'h39f3a9e3),
	.w6(32'hbc8b6766),
	.w7(32'hbc0402cd),
	.w8(32'hbc1acc31),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0645a4),
	.w1(32'h39eb84e3),
	.w2(32'h3b2e5306),
	.w3(32'h3bb743ec),
	.w4(32'h3afba6a4),
	.w5(32'h3ba30477),
	.w6(32'h3c07e0e2),
	.w7(32'h3b8fcda6),
	.w8(32'h3c07ce5f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0235d2),
	.w1(32'h3ab84e21),
	.w2(32'h3be42dde),
	.w3(32'hbb073ab3),
	.w4(32'h3b22fdc4),
	.w5(32'h3aefdf04),
	.w6(32'hbc762546),
	.w7(32'h3b839fbf),
	.w8(32'h3c02e429),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0878),
	.w1(32'hbaff2e02),
	.w2(32'h3a42d26c),
	.w3(32'h3bf3aaff),
	.w4(32'h39d0b68b),
	.w5(32'hba16a06d),
	.w6(32'h3c0153d1),
	.w7(32'h3b86ebb6),
	.w8(32'h3b280e20),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb9148),
	.w1(32'h3a666e0f),
	.w2(32'hbaab0b26),
	.w3(32'h3b4209ca),
	.w4(32'hb9ad356f),
	.w5(32'h3aa764bc),
	.w6(32'hbba493c6),
	.w7(32'hbb17195c),
	.w8(32'hbb013ff9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcba5fa),
	.w1(32'h3b6f6077),
	.w2(32'h3b8ac037),
	.w3(32'h3c06e444),
	.w4(32'h3bd22d14),
	.w5(32'h3a93df8f),
	.w6(32'h3bacc7a3),
	.w7(32'h3bef0ba4),
	.w8(32'h3b725bba),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6460e7),
	.w1(32'hbc5c9884),
	.w2(32'hbc708a83),
	.w3(32'h3bed01e7),
	.w4(32'hbbeb856f),
	.w5(32'hbbf362e3),
	.w6(32'h3c1a5f01),
	.w7(32'h3b55e4fa),
	.w8(32'hbb175461),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4c96c),
	.w1(32'h3a4c7c3b),
	.w2(32'hbab0721f),
	.w3(32'h3bdaa5c3),
	.w4(32'h3a316442),
	.w5(32'h3bbcc78b),
	.w6(32'h3be73cb0),
	.w7(32'h3b3cd721),
	.w8(32'h3bb294e7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae37083),
	.w1(32'h3ad58943),
	.w2(32'hba3ba853),
	.w3(32'hbaef5ab2),
	.w4(32'hbb5900e7),
	.w5(32'h3b12060f),
	.w6(32'hbc8517f3),
	.w7(32'hbb1caa85),
	.w8(32'hbb09bc2b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92365b),
	.w1(32'h39c1128e),
	.w2(32'h3aea95d9),
	.w3(32'h3b61b99b),
	.w4(32'hbb72d2c7),
	.w5(32'hbb9c3d0a),
	.w6(32'hbb0f94af),
	.w7(32'hbc26173c),
	.w8(32'h3b232c45),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4133ce),
	.w1(32'h3c4d2f76),
	.w2(32'h3c241c3d),
	.w3(32'hbc4b63c0),
	.w4(32'h3bae8689),
	.w5(32'h3c0da9e7),
	.w6(32'hbc2f6d44),
	.w7(32'hbc11fde7),
	.w8(32'h3af6ecc2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046e30),
	.w1(32'hbbdbf4e9),
	.w2(32'hbbabc1c9),
	.w3(32'h3c155a4e),
	.w4(32'hbaba1436),
	.w5(32'hbc159bb8),
	.w6(32'h3ca37a48),
	.w7(32'hba9b3747),
	.w8(32'hbb73ae6e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0afaea),
	.w1(32'hbb02439f),
	.w2(32'hbb658bd1),
	.w3(32'h3b61688b),
	.w4(32'hba58ac6c),
	.w5(32'h39c460ad),
	.w6(32'h3bb8300b),
	.w7(32'h3ae2f42f),
	.w8(32'hbad0933e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c875),
	.w1(32'hb9c14a4a),
	.w2(32'hbb917b35),
	.w3(32'hbb300591),
	.w4(32'h3bb2acce),
	.w5(32'h3a63c30f),
	.w6(32'hbc4aa6c2),
	.w7(32'hbb3e840a),
	.w8(32'h3c1927de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66ab9b),
	.w1(32'hba619fb2),
	.w2(32'hba8d5960),
	.w3(32'hbba4a6f8),
	.w4(32'hbb0250e1),
	.w5(32'hba779d10),
	.w6(32'hbb11f383),
	.w7(32'hbaf2906d),
	.w8(32'hbb92814e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fe2a9),
	.w1(32'hba9f06c8),
	.w2(32'hbbfb4eb1),
	.w3(32'hbbff59bb),
	.w4(32'h3c185e1c),
	.w5(32'h3ad735b7),
	.w6(32'hbc02334d),
	.w7(32'hbb156531),
	.w8(32'hbb0a9795),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404dd0),
	.w1(32'hbba5d0db),
	.w2(32'h3c18d064),
	.w3(32'hba45571a),
	.w4(32'hbb22d3b0),
	.w5(32'h3c524224),
	.w6(32'hbb71652d),
	.w7(32'hb93bbfb2),
	.w8(32'h3c29691f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace8d3),
	.w1(32'h37610f77),
	.w2(32'h3b3f2c47),
	.w3(32'h3a3d4bb1),
	.w4(32'hba9e98af),
	.w5(32'hb8bd9ced),
	.w6(32'hba9a7fee),
	.w7(32'hbaf3bdad),
	.w8(32'hba682192),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b701671),
	.w1(32'h3b03de6b),
	.w2(32'hbae0591d),
	.w3(32'hba5d3d90),
	.w4(32'h3ab104ea),
	.w5(32'hbb57d3dd),
	.w6(32'h39e66484),
	.w7(32'hbab7e10c),
	.w8(32'hbbc61ac8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23549f),
	.w1(32'h3b1a7b37),
	.w2(32'hba67bb5c),
	.w3(32'h3c5b9afa),
	.w4(32'h3b990ac9),
	.w5(32'hba73a5fe),
	.w6(32'h3b883991),
	.w7(32'hbb65cd42),
	.w8(32'hba62fd21),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ad9ac),
	.w1(32'hbb1120fd),
	.w2(32'hbb34dc41),
	.w3(32'h3b6a12c3),
	.w4(32'h3ada71e6),
	.w5(32'hbb4fa293),
	.w6(32'h3c1229c2),
	.w7(32'hba18f448),
	.w8(32'h3ad72f87),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384aa2),
	.w1(32'hbc0b7fa4),
	.w2(32'hbb228ff5),
	.w3(32'h3b983d8a),
	.w4(32'hbc22b972),
	.w5(32'h393244d3),
	.w6(32'h3c15c5c8),
	.w7(32'h3b09551c),
	.w8(32'h3a53abd1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e06c),
	.w1(32'hbba29912),
	.w2(32'h3bae4b2f),
	.w3(32'h3adbd811),
	.w4(32'hbc62fc45),
	.w5(32'h3c33d85f),
	.w6(32'h3bab365b),
	.w7(32'hbb16ddd4),
	.w8(32'h3b8a4c12),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcfc73),
	.w1(32'h3a63012a),
	.w2(32'h3b8c4375),
	.w3(32'hbc26c1bf),
	.w4(32'hbb453184),
	.w5(32'h3bf6bff6),
	.w6(32'hbcab7c7d),
	.w7(32'hbc832702),
	.w8(32'hbb96770a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ee69),
	.w1(32'h3c55ab80),
	.w2(32'h3b727964),
	.w3(32'h3c11ede7),
	.w4(32'h3c3fddff),
	.w5(32'hbb75f9a8),
	.w6(32'h3bdae055),
	.w7(32'h3badf88b),
	.w8(32'hbabd8496),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba802940),
	.w1(32'hbb919765),
	.w2(32'h3b921b78),
	.w3(32'h3ac7bb90),
	.w4(32'hbb911973),
	.w5(32'h3b54563f),
	.w6(32'hba528fa7),
	.w7(32'hbb08764f),
	.w8(32'h3bdda191),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b358b),
	.w1(32'h3a8a46f1),
	.w2(32'hba0886e4),
	.w3(32'hbbbf54d4),
	.w4(32'hba3a601d),
	.w5(32'hbb3bb691),
	.w6(32'h3b0f8f95),
	.w7(32'hb9f5d8f3),
	.w8(32'h397dc44e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a660281),
	.w1(32'hb9bf1f02),
	.w2(32'h3ad9dc59),
	.w3(32'h39383837),
	.w4(32'hba8b6198),
	.w5(32'hba36ff4f),
	.w6(32'h39d5f1c4),
	.w7(32'h3a06c0ba),
	.w8(32'h3bbb025e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21fc26),
	.w1(32'h39be0475),
	.w2(32'h3ba55eae),
	.w3(32'hbb8e8475),
	.w4(32'hbbbdecc6),
	.w5(32'hba9c0c9a),
	.w6(32'hbac370a2),
	.w7(32'h388357c5),
	.w8(32'h3a7aeba4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a4ec1),
	.w1(32'h3ba47a88),
	.w2(32'h39111a82),
	.w3(32'h3ba0358b),
	.w4(32'h3bf765b9),
	.w5(32'hba1e5430),
	.w6(32'h3bd43c91),
	.w7(32'h3ba7edde),
	.w8(32'h38d264f5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eeb4c),
	.w1(32'hbbf2ac4a),
	.w2(32'h3aeb328b),
	.w3(32'h39f72e77),
	.w4(32'hbbe89836),
	.w5(32'h3b9f29c3),
	.w6(32'hba9c311b),
	.w7(32'hbb66b256),
	.w8(32'h3b4aee48),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb821b29),
	.w1(32'h3c1080fc),
	.w2(32'hbb35978e),
	.w3(32'hbbbcdcba),
	.w4(32'h3c3d75d1),
	.w5(32'hbb95c6c0),
	.w6(32'hbb6e1e3e),
	.w7(32'h3c1c600c),
	.w8(32'hbb326a9a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc3709),
	.w1(32'hbb996d46),
	.w2(32'hbbbb1e69),
	.w3(32'h3ad7fd50),
	.w4(32'h3ba04612),
	.w5(32'hbb3c37ba),
	.w6(32'hbb4c671a),
	.w7(32'hbb5cce82),
	.w8(32'hbadfaa5b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2014f6),
	.w1(32'hbb86850b),
	.w2(32'hbbd760f9),
	.w3(32'h3c60b1d9),
	.w4(32'hb8f9be32),
	.w5(32'hb9fbf7d3),
	.w6(32'h3c570dac),
	.w7(32'h3baf71ac),
	.w8(32'h3b9edd8e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032dfa),
	.w1(32'hbaee8249),
	.w2(32'hbba2e01c),
	.w3(32'hbbaf99c2),
	.w4(32'hbbab63b2),
	.w5(32'hbba18222),
	.w6(32'hbbdcad29),
	.w7(32'hbb513c75),
	.w8(32'hbbb00051),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec9ef),
	.w1(32'h3b6c3890),
	.w2(32'hbb778e59),
	.w3(32'hbb8c83e4),
	.w4(32'h3ba49aa9),
	.w5(32'hbc17aa46),
	.w6(32'hbb774840),
	.w7(32'h3ae656bc),
	.w8(32'hbb320e34),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff643e),
	.w1(32'h3b33879d),
	.w2(32'h3a293339),
	.w3(32'hbac195c9),
	.w4(32'h3bc5a2a7),
	.w5(32'hbb38af3b),
	.w6(32'hb992e941),
	.w7(32'h3b48aaad),
	.w8(32'hba21eead),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d1b1),
	.w1(32'hbc0096bc),
	.w2(32'h3c4c8c27),
	.w3(32'hbb53ff7a),
	.w4(32'hbc0aa340),
	.w5(32'h3c56a96d),
	.w6(32'h3ae4a94d),
	.w7(32'hbb735344),
	.w8(32'h3c51c600),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb71614),
	.w1(32'h3c5fedc4),
	.w2(32'h3c269c10),
	.w3(32'hbb6e8af0),
	.w4(32'h3c13c72c),
	.w5(32'h3c406f4e),
	.w6(32'hbcdd4ca3),
	.w7(32'hbc9a000b),
	.w8(32'hbc535e23),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b097b37),
	.w1(32'h3b881a62),
	.w2(32'hbb6a31d8),
	.w3(32'h3b3d8c5d),
	.w4(32'h3ba7c1b2),
	.w5(32'h3b1a08be),
	.w6(32'hbc512712),
	.w7(32'hbb8e535c),
	.w8(32'hbb2557ed),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a806a25),
	.w1(32'hb7a41b6d),
	.w2(32'h3a478a1f),
	.w3(32'h3b993934),
	.w4(32'h38eaf220),
	.w5(32'h3a925bbe),
	.w6(32'h3b90e353),
	.w7(32'h3863873a),
	.w8(32'hba11360a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fc36b),
	.w1(32'h3b094015),
	.w2(32'h3a5b613c),
	.w3(32'hbb79e0f2),
	.w4(32'hbb3df53c),
	.w5(32'hbb5be70c),
	.w6(32'hbac75af8),
	.w7(32'hbb532b07),
	.w8(32'hbbc96671),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba536fb2),
	.w1(32'hbb9e7bfd),
	.w2(32'hbafa05ae),
	.w3(32'hbb390cb8),
	.w4(32'h3a255081),
	.w5(32'hbb78dc68),
	.w6(32'hbb90a61a),
	.w7(32'h399308e4),
	.w8(32'h39f07e98),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b506663),
	.w1(32'hba15998c),
	.w2(32'hbb971f4c),
	.w3(32'h3b4faf9a),
	.w4(32'hba8f6fa6),
	.w5(32'hbb8b565f),
	.w6(32'h3b4b97ec),
	.w7(32'hbb592fc5),
	.w8(32'hbbb1143b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb189b7),
	.w1(32'hbba4eef4),
	.w2(32'h3b513d0e),
	.w3(32'h3bfef9eb),
	.w4(32'hbbfaf0cd),
	.w5(32'h3b4caf10),
	.w6(32'h3bf3909c),
	.w7(32'hbab05c3b),
	.w8(32'h3bbbe47d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc16b9),
	.w1(32'h3a4b56db),
	.w2(32'hbbd52f5a),
	.w3(32'hba693d2b),
	.w4(32'h3c18179b),
	.w5(32'h3ad940f0),
	.w6(32'hbc78ef11),
	.w7(32'hbaeba88c),
	.w8(32'hbad1e1fd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaa26f),
	.w1(32'hbb92e768),
	.w2(32'h383beb46),
	.w3(32'h3b52928a),
	.w4(32'hbb9688a3),
	.w5(32'hba7dfe2f),
	.w6(32'h3b90e57d),
	.w7(32'h3a09a898),
	.w8(32'h394e7b26),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231233),
	.w1(32'h398b4da6),
	.w2(32'h3bc7b252),
	.w3(32'h3b817da5),
	.w4(32'hba8c8b77),
	.w5(32'h3ac032ad),
	.w6(32'hbb8cfa90),
	.w7(32'hbb85b0e7),
	.w8(32'h3b398888),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8c6e2),
	.w1(32'hbad6243a),
	.w2(32'hbba8b25e),
	.w3(32'h3bcfa0cd),
	.w4(32'hba5612fb),
	.w5(32'hbb239c3e),
	.w6(32'hbbc63eef),
	.w7(32'hbbf42796),
	.w8(32'hb9ddfd46),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7225e),
	.w1(32'h3b635709),
	.w2(32'h39d3e61b),
	.w3(32'hbbe4b778),
	.w4(32'hbaca4d71),
	.w5(32'hbb35493e),
	.w6(32'h3b9fc134),
	.w7(32'hbb64b385),
	.w8(32'hbb9b77d5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53982c),
	.w1(32'h3bde2e11),
	.w2(32'h3b780a48),
	.w3(32'h3a4de6b8),
	.w4(32'h3bb0f150),
	.w5(32'h3b7b6bd6),
	.w6(32'hbb84b039),
	.w7(32'h3aea8668),
	.w8(32'h3b6235c5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466c3f),
	.w1(32'hba1bbb5a),
	.w2(32'h3b53c3d0),
	.w3(32'hbb2d18e9),
	.w4(32'hbb13b083),
	.w5(32'h3b5ffeb0),
	.w6(32'hbb26e040),
	.w7(32'hba2ca820),
	.w8(32'hbaa9bddf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3afa50),
	.w1(32'hbc274a6b),
	.w2(32'hbc21648e),
	.w3(32'h3b8947ae),
	.w4(32'hbbb1c680),
	.w5(32'hbb6efdf4),
	.w6(32'h3c402b28),
	.w7(32'h3ba48e57),
	.w8(32'h3b9df24b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba71cc),
	.w1(32'h3bff395c),
	.w2(32'h3ba23d67),
	.w3(32'hb8d5c716),
	.w4(32'h3b8f67a2),
	.w5(32'h3c003c19),
	.w6(32'h3be137ae),
	.w7(32'h3b5daa09),
	.w8(32'h3bcedf87),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd11af5),
	.w1(32'h3ad6dce2),
	.w2(32'hb98f8c20),
	.w3(32'hbbc2e3f2),
	.w4(32'h3b03d1f2),
	.w5(32'h3a1a6cc1),
	.w6(32'hbbadcdcf),
	.w7(32'h3a341cb8),
	.w8(32'h3b21f41e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f4b9a),
	.w1(32'h3a2db8ea),
	.w2(32'hba7021f2),
	.w3(32'hbb428eb8),
	.w4(32'h3b08498b),
	.w5(32'h38102def),
	.w6(32'hbb04b375),
	.w7(32'hb85308dd),
	.w8(32'h398bc061),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0759d),
	.w1(32'hba105f61),
	.w2(32'hbae2c9b4),
	.w3(32'hbb54b4c9),
	.w4(32'h3aea67d6),
	.w5(32'hbadae8be),
	.w6(32'hbb210aee),
	.w7(32'h3a45bb64),
	.w8(32'hba73bb2b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f87b4),
	.w1(32'hbbac4046),
	.w2(32'hbb960ad7),
	.w3(32'h3bc65346),
	.w4(32'hbbaabc19),
	.w5(32'hbb8f4d31),
	.w6(32'h3c3273ce),
	.w7(32'hbac728cf),
	.w8(32'hbae3603e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db846),
	.w1(32'h3b8f90b9),
	.w2(32'h3b997273),
	.w3(32'hbb0f07a9),
	.w4(32'h3c3d5716),
	.w5(32'h3bb890b3),
	.w6(32'hbbe09378),
	.w7(32'h3b34672b),
	.w8(32'h3ad71947),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe03a1),
	.w1(32'h3ac1aae5),
	.w2(32'h39e224d6),
	.w3(32'hbbd47cfa),
	.w4(32'hb9fd786c),
	.w5(32'hbaa0a5da),
	.w6(32'hbb809a2d),
	.w7(32'hb9c0a333),
	.w8(32'h3b6475d1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166232),
	.w1(32'h3b5cb862),
	.w2(32'h3c511387),
	.w3(32'h3b856220),
	.w4(32'h3c1ced75),
	.w5(32'h3cc1086b),
	.w6(32'hbb52dcea),
	.w7(32'h3b04ea5c),
	.w8(32'h3c8a2e46),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc779),
	.w1(32'h3b41c77b),
	.w2(32'hbb9f1aef),
	.w3(32'hbb3d855d),
	.w4(32'hb9e93fb5),
	.w5(32'hbbd8cfa5),
	.w6(32'hbc01f4c4),
	.w7(32'hbbafde67),
	.w8(32'h3a903873),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3ec3),
	.w1(32'h3894a2a8),
	.w2(32'hba99b2c2),
	.w3(32'hbacfe9ae),
	.w4(32'h3ba61d8b),
	.w5(32'hbb9f7c10),
	.w6(32'hbb4cdd3f),
	.w7(32'hbb441043),
	.w8(32'hbb015878),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054e94),
	.w1(32'hbc4aa75b),
	.w2(32'hbb26ea00),
	.w3(32'h3b72dd4e),
	.w4(32'hbc07b2f8),
	.w5(32'hbb26f271),
	.w6(32'h3c279f77),
	.w7(32'hba0a3899),
	.w8(32'h3bd287a0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763e29),
	.w1(32'hbbd73964),
	.w2(32'hb9630355),
	.w3(32'hbc1232cc),
	.w4(32'hbc34ab7f),
	.w5(32'h3b766097),
	.w6(32'hb9a70bb4),
	.w7(32'hbba2c326),
	.w8(32'h3ae1dd11),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64e5d8),
	.w1(32'h3b1e344b),
	.w2(32'hbbb9909e),
	.w3(32'h3aadc091),
	.w4(32'h3b096ac7),
	.w5(32'h3a354fcb),
	.w6(32'h3b3daf09),
	.w7(32'h3b41b960),
	.w8(32'h3b7a8c5a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980d225),
	.w1(32'hbc032209),
	.w2(32'hbb9af52a),
	.w3(32'hb86c2de1),
	.w4(32'hbb6a7d95),
	.w5(32'hba3573b0),
	.w6(32'hba739fd3),
	.w7(32'hbb1af42d),
	.w8(32'h3985a1ca),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a229464),
	.w1(32'h3b982b3c),
	.w2(32'hbaa1f27a),
	.w3(32'h3b52d775),
	.w4(32'h3a850d8b),
	.w5(32'hbb0cbb2e),
	.w6(32'h3beb5c97),
	.w7(32'h3b674fc2),
	.w8(32'hb7941e16),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef249d),
	.w1(32'h3b98f552),
	.w2(32'h3bd36aad),
	.w3(32'h3bbce64e),
	.w4(32'h3aebee23),
	.w5(32'h3b9299f9),
	.w6(32'h3c7ab3f7),
	.w7(32'h3ba7e37c),
	.w8(32'h3bc6f171),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a7489),
	.w1(32'h3ae8ef9b),
	.w2(32'hbb773dcd),
	.w3(32'hb79ae64c),
	.w4(32'h3bf95acc),
	.w5(32'hbb5ba845),
	.w6(32'hbb6ca98f),
	.w7(32'h39a0aacb),
	.w8(32'hbbe8c6af),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f4198),
	.w1(32'hbb088db3),
	.w2(32'h3b92dd7e),
	.w3(32'hbb57e34d),
	.w4(32'hbb60ec8c),
	.w5(32'h3b9d5e2a),
	.w6(32'h3b1c68aa),
	.w7(32'hbb29f8e2),
	.w8(32'h3b2a29d5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f287),
	.w1(32'h3bb1ee93),
	.w2(32'h3b925a00),
	.w3(32'hbb9bc760),
	.w4(32'h3ae95f3d),
	.w5(32'h3b5223ec),
	.w6(32'hbc60f262),
	.w7(32'hbb517db1),
	.w8(32'hba70fe12),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82d873),
	.w1(32'hbbab137e),
	.w2(32'hbb03f14e),
	.w3(32'hbb25ce3b),
	.w4(32'hbb98b5f5),
	.w5(32'hba455c1f),
	.w6(32'hb96974b2),
	.w7(32'hbb0ac95b),
	.w8(32'hb9a88a3f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde51e),
	.w1(32'hbb785250),
	.w2(32'hbbc54adc),
	.w3(32'h3b0d5bd4),
	.w4(32'hbc1bb7be),
	.w5(32'hbae61340),
	.w6(32'h3ae30a1a),
	.w7(32'hb92d6689),
	.w8(32'h3a16c214),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908eac),
	.w1(32'h3a9da16b),
	.w2(32'h3990c6d4),
	.w3(32'h3b549c54),
	.w4(32'h3b2bb116),
	.w5(32'hbb937681),
	.w6(32'h3be0b966),
	.w7(32'h3b1f38e9),
	.w8(32'hbb223f52),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18b13),
	.w1(32'h3b9bacff),
	.w2(32'hbb18a4e4),
	.w3(32'h3b87b7f8),
	.w4(32'h3c1ef7e2),
	.w5(32'hba6c140f),
	.w6(32'h3a38fa47),
	.w7(32'h3b0ca9de),
	.w8(32'hbbd82c12),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e9512),
	.w1(32'hbafbff6c),
	.w2(32'h3b43431f),
	.w3(32'hbbb11049),
	.w4(32'hba4f2a02),
	.w5(32'h39ff6272),
	.w6(32'hbba153ca),
	.w7(32'hbb0cf9af),
	.w8(32'hbbba9ea9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edf9c),
	.w1(32'hbab65515),
	.w2(32'hbb7af007),
	.w3(32'hbac797f8),
	.w4(32'hba107c8d),
	.w5(32'hbb84b1ca),
	.w6(32'hbb51c3d6),
	.w7(32'hbb0ac58a),
	.w8(32'hba8c1054),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a7f8),
	.w1(32'hbbb98647),
	.w2(32'hbb9942a9),
	.w3(32'h3b3b9a4b),
	.w4(32'hbabafe81),
	.w5(32'hbba3b770),
	.w6(32'h3c3177c6),
	.w7(32'h3a96ebba),
	.w8(32'hbb3ccc9f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1ef80),
	.w1(32'h3b41cb46),
	.w2(32'h3b8e6bab),
	.w3(32'hbb8bc862),
	.w4(32'h3c00dc42),
	.w5(32'h3ba3a7b9),
	.w6(32'hbc7633e3),
	.w7(32'hbbfbbfdc),
	.w8(32'hbb981495),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b468e2c),
	.w1(32'h3b05d5d0),
	.w2(32'hba8ff747),
	.w3(32'hba99566e),
	.w4(32'h3b3d3b8a),
	.w5(32'h3be9b004),
	.w6(32'h3ac246d7),
	.w7(32'h3b430ec4),
	.w8(32'h3bda0385),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba391ae),
	.w1(32'hbb61833b),
	.w2(32'hbbaf453a),
	.w3(32'hbb1f9598),
	.w4(32'hbb09fc9d),
	.w5(32'hbb7b7377),
	.w6(32'hbaccd298),
	.w7(32'h3a82ddf7),
	.w8(32'hbb37649f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cd5ca),
	.w1(32'hbc2acc4f),
	.w2(32'hbb94877a),
	.w3(32'hba355b33),
	.w4(32'hbc0fa445),
	.w5(32'hbad3c6df),
	.w6(32'h3a4c0340),
	.w7(32'hbbb451f0),
	.w8(32'hbb2e876c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6aad2a),
	.w1(32'h3b1b7c49),
	.w2(32'hbbb60207),
	.w3(32'h3be39432),
	.w4(32'h3b92720c),
	.w5(32'hbbaaa86c),
	.w6(32'h3bc1c250),
	.w7(32'h3b64666f),
	.w8(32'hbae3d5a7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939b121),
	.w1(32'h3c03c46b),
	.w2(32'h3b8d7281),
	.w3(32'h3a2538c4),
	.w4(32'h3bc9fb77),
	.w5(32'h39600493),
	.w6(32'hbaa2040a),
	.w7(32'h3ba13f70),
	.w8(32'h3b798d65),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1d271),
	.w1(32'h3bcd2a21),
	.w2(32'h3a47c77d),
	.w3(32'hbad79c05),
	.w4(32'h3bec712b),
	.w5(32'h3b889fe9),
	.w6(32'hbc218167),
	.w7(32'hbb9f1db6),
	.w8(32'h3a926abb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48a9be),
	.w1(32'h35bb3a53),
	.w2(32'h3b9f4a4b),
	.w3(32'h3af4a1e2),
	.w4(32'hbac431fa),
	.w5(32'h3bcc29e5),
	.w6(32'h3ad585db),
	.w7(32'hbb070600),
	.w8(32'h3bd63b83),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9f93d),
	.w1(32'h3b38c4c6),
	.w2(32'h3b5f3673),
	.w3(32'h3c111327),
	.w4(32'h3b5bd6a1),
	.w5(32'h3b290519),
	.w6(32'h3c10d25a),
	.w7(32'h3ae4364d),
	.w8(32'h3be80bdc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a99df),
	.w1(32'h3bcd17e0),
	.w2(32'h3bb58bb7),
	.w3(32'h3ae62fda),
	.w4(32'h3b8e790e),
	.w5(32'h3b155ca9),
	.w6(32'h3b35dc86),
	.w7(32'h3b9054e9),
	.w8(32'h3c06e260),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf61f73),
	.w1(32'h3a58c71b),
	.w2(32'hbc1c589b),
	.w3(32'hbba401e4),
	.w4(32'hba845c4c),
	.w5(32'hbc472578),
	.w6(32'hbb8579b9),
	.w7(32'hba00d7b1),
	.w8(32'hbc052995),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc2f45),
	.w1(32'hbb056d62),
	.w2(32'hbad35d30),
	.w3(32'hbad18403),
	.w4(32'hb9b6e833),
	.w5(32'hbb1d7450),
	.w6(32'h3b47f483),
	.w7(32'h3b223239),
	.w8(32'h3abc43a0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac16c0a),
	.w1(32'h3b99d4d4),
	.w2(32'h3b44c321),
	.w3(32'h3c0d9cf8),
	.w4(32'h3b23146b),
	.w5(32'h3a87926f),
	.w6(32'h3bae0563),
	.w7(32'h3baa3277),
	.w8(32'h3b9f9ca0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dccb3),
	.w1(32'hbb65c364),
	.w2(32'hbad8f1e8),
	.w3(32'h3aaffba8),
	.w4(32'hb87c3145),
	.w5(32'hbb7ebbb2),
	.w6(32'h3a29df0b),
	.w7(32'h3b71c399),
	.w8(32'h3ab9af05),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d10c),
	.w1(32'hbb2d29ad),
	.w2(32'hbb05189f),
	.w3(32'h3b745296),
	.w4(32'h3b2897f4),
	.w5(32'h3a9d6f94),
	.w6(32'h3bc3b693),
	.w7(32'h3aacaff4),
	.w8(32'hbaf77ff3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3e4d2),
	.w1(32'hb90f04fe),
	.w2(32'h3ad807c8),
	.w3(32'hbb08f7e2),
	.w4(32'h3aafcac4),
	.w5(32'h3adadad5),
	.w6(32'hba064649),
	.w7(32'h3a396a9d),
	.w8(32'hbae951af),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e7249),
	.w1(32'h3bb41e4d),
	.w2(32'hba0498d0),
	.w3(32'h3b901346),
	.w4(32'h3bbc1cf6),
	.w5(32'hbb9fce43),
	.w6(32'h3bc013e3),
	.w7(32'h3b636126),
	.w8(32'h3ae546f0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b171f83),
	.w1(32'h38afc18f),
	.w2(32'h3c1af5b2),
	.w3(32'hbad55f56),
	.w4(32'h3b47432b),
	.w5(32'h3c5c7579),
	.w6(32'hbb37d147),
	.w7(32'h3abe41db),
	.w8(32'h3be243af),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39819e29),
	.w1(32'h3ad48949),
	.w2(32'hbb6de2a6),
	.w3(32'h3a37c664),
	.w4(32'h3bc39256),
	.w5(32'hbb76828e),
	.w6(32'h3a798e9e),
	.w7(32'h3ba8fbeb),
	.w8(32'hbb9436bd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1da62),
	.w1(32'h3aa04e51),
	.w2(32'hbac75ed7),
	.w3(32'hbb30ab40),
	.w4(32'h3bbc5126),
	.w5(32'hba8c8862),
	.w6(32'hbc6bf9fe),
	.w7(32'hbb2bf4e9),
	.w8(32'hbc1ebf76),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f84ede),
	.w1(32'h3af420e5),
	.w2(32'h3b6f8c17),
	.w3(32'h3c10ebdd),
	.w4(32'hbc32f8a1),
	.w5(32'h3ac1d229),
	.w6(32'h3c7fd3fe),
	.w7(32'h3b98f736),
	.w8(32'h3bc29843),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75b992),
	.w1(32'hba8cd1c8),
	.w2(32'hbab1a2fc),
	.w3(32'h3b828b41),
	.w4(32'h3b9224bc),
	.w5(32'hba0e1be0),
	.w6(32'hbb7b7203),
	.w7(32'hba4f0ded),
	.w8(32'hba2402d6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922cf1f),
	.w1(32'hbbb29b61),
	.w2(32'hbbb486ee),
	.w3(32'hbb08f18a),
	.w4(32'hbb53500e),
	.w5(32'hbb73303f),
	.w6(32'hbb35ea10),
	.w7(32'hbb86646a),
	.w8(32'hbb87b26e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530ca0),
	.w1(32'h3b129a08),
	.w2(32'hbafe533b),
	.w3(32'h3b955469),
	.w4(32'h3b156906),
	.w5(32'hbbd86668),
	.w6(32'h3ba69d48),
	.w7(32'h3a405859),
	.w8(32'hbb10f256),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba717143),
	.w1(32'hb9c0d522),
	.w2(32'h399850af),
	.w3(32'hbb040562),
	.w4(32'h3abbe4ec),
	.w5(32'hbb33096c),
	.w6(32'hbb2dc05b),
	.w7(32'h39cf7a49),
	.w8(32'hbaa0f899),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbaca5),
	.w1(32'h3b837da1),
	.w2(32'hbaba1bd5),
	.w3(32'h3c031de7),
	.w4(32'h3bed80d4),
	.w5(32'h3a00d077),
	.w6(32'h3b0dd481),
	.w7(32'hbba5c416),
	.w8(32'hba33ed9b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b56aa),
	.w1(32'hbc05d064),
	.w2(32'h3adfc525),
	.w3(32'hbb7cb94e),
	.w4(32'hbc03a5a3),
	.w5(32'h3ba0375a),
	.w6(32'hba92b910),
	.w7(32'hbc08fc2c),
	.w8(32'hba032317),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba715636),
	.w1(32'h39eb7528),
	.w2(32'h3aaa0f84),
	.w3(32'hb986d078),
	.w4(32'hbbdac51d),
	.w5(32'h3a90a3d1),
	.w6(32'h3bc37cb3),
	.w7(32'h3b482b65),
	.w8(32'h3b9020e5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c628ada),
	.w1(32'hba5c59b2),
	.w2(32'h3a665b4c),
	.w3(32'h3c30a343),
	.w4(32'hbae7aad3),
	.w5(32'h3b383e94),
	.w6(32'h3ba44f9c),
	.w7(32'h3a845df5),
	.w8(32'hbb372bbb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc855f),
	.w1(32'h3a2a6dc7),
	.w2(32'hbb8da7fa),
	.w3(32'hba83c571),
	.w4(32'h3bb58c43),
	.w5(32'hbb269133),
	.w6(32'hba68ed9e),
	.w7(32'hb98880ad),
	.w8(32'hbb1c2c99),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0c224),
	.w1(32'hbbf65ed0),
	.w2(32'h3a9ab16d),
	.w3(32'hbace2dc3),
	.w4(32'h3b7196e0),
	.w5(32'hbb7a7af5),
	.w6(32'hbc1d6c5c),
	.w7(32'h3b1cef14),
	.w8(32'hbc2e70c2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb459f07),
	.w1(32'hbb473d00),
	.w2(32'hbc863ffe),
	.w3(32'hbc0a1420),
	.w4(32'hbbfe6dfa),
	.w5(32'hbc97696c),
	.w6(32'h3917784c),
	.w7(32'hbc43600a),
	.w8(32'hba6c0e0f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee02dc),
	.w1(32'h3c06dc27),
	.w2(32'hbb1fa6f3),
	.w3(32'h39c9cc45),
	.w4(32'h3c4bbd15),
	.w5(32'hbc39d6d0),
	.w6(32'hbc7f0526),
	.w7(32'h3bc5fbc7),
	.w8(32'h3b8f4c2d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b153a),
	.w1(32'h3aec3e99),
	.w2(32'hbb7e8841),
	.w3(32'hbae87118),
	.w4(32'hbb507f8d),
	.w5(32'hbc364769),
	.w6(32'h3a9d4f7b),
	.w7(32'hbc168aa2),
	.w8(32'h3bdc89f7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37493f),
	.w1(32'h3bdf781b),
	.w2(32'h3be5fb50),
	.w3(32'hbae5f18f),
	.w4(32'h3b8ea4a3),
	.w5(32'h3bc052ab),
	.w6(32'hbaaff12d),
	.w7(32'h3c331206),
	.w8(32'h3be18203),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22f9b4),
	.w1(32'hbb3667a2),
	.w2(32'hbbe0f54e),
	.w3(32'hbb4faf77),
	.w4(32'h3be87782),
	.w5(32'hbb7ff899),
	.w6(32'h3b61a184),
	.w7(32'h3b6e99a4),
	.w8(32'h3d3814a2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaf932),
	.w1(32'h3bca5342),
	.w2(32'hbb17f493),
	.w3(32'h3b9793a4),
	.w4(32'hbba5c062),
	.w5(32'h3c8fb0ce),
	.w6(32'h3c4d52f0),
	.w7(32'h3b35ea52),
	.w8(32'h39245323),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae01d9f),
	.w1(32'hbb9ff21c),
	.w2(32'hbc6789bd),
	.w3(32'h3bf53a15),
	.w4(32'hbbb3b901),
	.w5(32'hbcf88439),
	.w6(32'hb920e40f),
	.w7(32'hbad1a541),
	.w8(32'hbaad31fc),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ed1b),
	.w1(32'hbc258557),
	.w2(32'h3ad5b666),
	.w3(32'hbcb834b3),
	.w4(32'hbcabb581),
	.w5(32'h3b5a2fa4),
	.w6(32'hbb96021f),
	.w7(32'hbc35e4fe),
	.w8(32'hbbe3e216),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2f42),
	.w1(32'hba1eaf65),
	.w2(32'hbbb9ce28),
	.w3(32'h3bf792e3),
	.w4(32'h3b5616c5),
	.w5(32'h3aa956f8),
	.w6(32'hba4b5a4d),
	.w7(32'h3bd3c3a9),
	.w8(32'hbba39878),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0070b2),
	.w1(32'h3b2940de),
	.w2(32'h3b5c4edd),
	.w3(32'hbbf6476b),
	.w4(32'h3bcabd89),
	.w5(32'h3be06036),
	.w6(32'hbb68941a),
	.w7(32'h3bb077c9),
	.w8(32'h3b7dd40a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c144),
	.w1(32'h3b29989a),
	.w2(32'h3b78756b),
	.w3(32'h3b340dcb),
	.w4(32'h3c32f6b4),
	.w5(32'h3bfc99a0),
	.w6(32'h3bce1450),
	.w7(32'hb8da2335),
	.w8(32'h3c104ba7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1b35b),
	.w1(32'h3c544864),
	.w2(32'h3c9bbdec),
	.w3(32'hbc6de96e),
	.w4(32'h3bdb1e48),
	.w5(32'h3b89a879),
	.w6(32'hbb485c1c),
	.w7(32'h3bd02c8a),
	.w8(32'hbc37e8cd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928b40),
	.w1(32'h3ad161c7),
	.w2(32'h3b8047f1),
	.w3(32'hbccf28b5),
	.w4(32'hbbb87454),
	.w5(32'h3a4fc2a0),
	.w6(32'hbca70d2c),
	.w7(32'hbc9b0697),
	.w8(32'h3889d1ee),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebdf37),
	.w1(32'hbc997cda),
	.w2(32'hbc1d6f05),
	.w3(32'hbbaa01b6),
	.w4(32'hbcb948bd),
	.w5(32'hbc83bd3e),
	.w6(32'hbb1befd4),
	.w7(32'hbcd00b8c),
	.w8(32'hbca0d2c6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934a60),
	.w1(32'hbb8845bf),
	.w2(32'h3af0bccf),
	.w3(32'hbcce8b8c),
	.w4(32'hba532efc),
	.w5(32'hbc365e05),
	.w6(32'hbbfb7d42),
	.w7(32'hbbd25a16),
	.w8(32'hbb899599),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c162f),
	.w1(32'hbb41bcbd),
	.w2(32'h3c1234f1),
	.w3(32'h3b08f343),
	.w4(32'h3bb83c77),
	.w5(32'h3ca138ee),
	.w6(32'h3bb9169e),
	.w7(32'h3c316921),
	.w8(32'h3b851928),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba930b1),
	.w1(32'hbba6ffb4),
	.w2(32'h3c37cb24),
	.w3(32'h3c914002),
	.w4(32'h3b25b7ef),
	.w5(32'h3ce421a4),
	.w6(32'h39eafec2),
	.w7(32'h3bc6d734),
	.w8(32'hbb461603),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1379d0),
	.w1(32'h3b0a76c7),
	.w2(32'hb9c1a5a9),
	.w3(32'h3c199ee3),
	.w4(32'h3accc2eb),
	.w5(32'h3ced7ec9),
	.w6(32'hba112ca3),
	.w7(32'hb9567908),
	.w8(32'hbbe9b5bc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded3ca),
	.w1(32'h3aba0268),
	.w2(32'h3c801b22),
	.w3(32'hb8d13532),
	.w4(32'h3c021dfd),
	.w5(32'h3c11b3c1),
	.w6(32'hbca82f82),
	.w7(32'hbc21b51a),
	.w8(32'h3bf881ba),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e416d5),
	.w1(32'h3c0534f5),
	.w2(32'hba84e590),
	.w3(32'hbb741c9a),
	.w4(32'h3be9f292),
	.w5(32'hbc50c02b),
	.w6(32'hbca4d107),
	.w7(32'hbc3fa1e5),
	.w8(32'hbcaf2bfd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f62b2),
	.w1(32'hba3de969),
	.w2(32'h3ab5dcb9),
	.w3(32'hbc902c39),
	.w4(32'h3c020cdc),
	.w5(32'h3b220dc6),
	.w6(32'hbca926ff),
	.w7(32'hba64dac3),
	.w8(32'h3b2812ff),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24457),
	.w1(32'h3a122e9d),
	.w2(32'hb9be8428),
	.w3(32'h3c3a4fd7),
	.w4(32'hb877a7d1),
	.w5(32'h3b92c156),
	.w6(32'h3c5d6885),
	.w7(32'h3b10ff2d),
	.w8(32'h3a02ed8c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad496a5),
	.w1(32'h3acd134a),
	.w2(32'hbbf14cf2),
	.w3(32'h3b2b094a),
	.w4(32'h3c3d08d5),
	.w5(32'h3bf98ec9),
	.w6(32'h3c75b0df),
	.w7(32'h3c3424bc),
	.w8(32'h3c4645dd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19d7e2),
	.w1(32'hbc27c1e7),
	.w2(32'h3b0a22f4),
	.w3(32'hbb0ffadf),
	.w4(32'hbb326241),
	.w5(32'hb90edb53),
	.w6(32'hba8f30cc),
	.w7(32'h3bf800b7),
	.w8(32'h39942406),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2dab),
	.w1(32'hbbdc6076),
	.w2(32'hbc81f5ea),
	.w3(32'hbb0f27d9),
	.w4(32'hbc07aba7),
	.w5(32'hbcc94a4c),
	.w6(32'h3c1f39fe),
	.w7(32'hbbddd4ce),
	.w8(32'hbc8446e0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4de976),
	.w1(32'hbcd2ae95),
	.w2(32'hbcd4bc55),
	.w3(32'hbb3413a0),
	.w4(32'hbc99a3a7),
	.w5(32'hbca76657),
	.w6(32'hbc43fc8d),
	.w7(32'hbca200b0),
	.w8(32'hbc5016dc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7783),
	.w1(32'hbbda55d3),
	.w2(32'hba4e130b),
	.w3(32'hbc2031c6),
	.w4(32'hbad2dfda),
	.w5(32'hbac9aac9),
	.w6(32'hbc115ec8),
	.w7(32'hbbbad2c5),
	.w8(32'h3bf1dbe4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c3c75),
	.w1(32'hbb8c7a1e),
	.w2(32'hbb645fc7),
	.w3(32'h3b06a47a),
	.w4(32'hbae5ef99),
	.w5(32'hbad253e3),
	.w6(32'hba9e7d81),
	.w7(32'h39fbd3b8),
	.w8(32'h3bb5e74b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5d87),
	.w1(32'h3c3bff33),
	.w2(32'hba79f172),
	.w3(32'hbc1ee23b),
	.w4(32'h3b0a7d00),
	.w5(32'hbbdc8938),
	.w6(32'hbc244113),
	.w7(32'hbb671cdb),
	.w8(32'h3ac634ad),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c588a91),
	.w1(32'hbcdc8ce2),
	.w2(32'hbcd02a68),
	.w3(32'h3ac8aac5),
	.w4(32'hbc98ef81),
	.w5(32'hbcd465ed),
	.w6(32'hbbadf77c),
	.w7(32'hbc9362c0),
	.w8(32'hbca17423),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc18bb),
	.w1(32'h3b26af97),
	.w2(32'hbaa766d7),
	.w3(32'hbc512276),
	.w4(32'hba984f3a),
	.w5(32'h3b400003),
	.w6(32'hbc997a51),
	.w7(32'h3b0aaed2),
	.w8(32'hbc00d6e4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66a5e2),
	.w1(32'hbae5cc57),
	.w2(32'h3cc8c522),
	.w3(32'hbbb2f459),
	.w4(32'h3c836244),
	.w5(32'h3d00e105),
	.w6(32'hbca03477),
	.w7(32'hbcb5f2d6),
	.w8(32'hbc167748),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd05a08),
	.w1(32'hbc975bb0),
	.w2(32'hbc0e00c0),
	.w3(32'hbc8f0413),
	.w4(32'hbbe5b064),
	.w5(32'h3b11c1de),
	.w6(32'hbbf87d1f),
	.w7(32'hbc0b79a6),
	.w8(32'hbcd7a8a5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca282b1),
	.w1(32'h3a1afa5d),
	.w2(32'h3bd80e2c),
	.w3(32'h3c233fa5),
	.w4(32'hbba73c1c),
	.w5(32'h3ae12d1e),
	.w6(32'hbca1e91f),
	.w7(32'hbbdec2ff),
	.w8(32'hbc9ee315),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d18cd),
	.w1(32'hbc51e2d6),
	.w2(32'hbc1fb159),
	.w3(32'hbb62d393),
	.w4(32'hbc603b18),
	.w5(32'hbbeb04b7),
	.w6(32'hbc9a92b5),
	.w7(32'hbba317c8),
	.w8(32'hba118831),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9cb5a),
	.w1(32'h3b825758),
	.w2(32'h3b33acb8),
	.w3(32'hbad77221),
	.w4(32'h3cacf1f0),
	.w5(32'hbbbcb252),
	.w6(32'h3b0149b7),
	.w7(32'hba9c5ba5),
	.w8(32'h3a9554ed),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ccb34),
	.w1(32'hbb6a49ed),
	.w2(32'hba7723d1),
	.w3(32'hbc58dff5),
	.w4(32'hbc449885),
	.w5(32'hbc2d1655),
	.w6(32'hbab7208c),
	.w7(32'hbc11ffe1),
	.w8(32'hb9bcc8f2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b383dc2),
	.w1(32'hb9cc354c),
	.w2(32'hba0aa785),
	.w3(32'h3bb13e39),
	.w4(32'h3b943e42),
	.w5(32'hbc0fb9fa),
	.w6(32'hbc17dc82),
	.w7(32'h39f7255a),
	.w8(32'h3c28787e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b2216),
	.w1(32'hbb09bc3b),
	.w2(32'hbbaa5339),
	.w3(32'hbbbd479a),
	.w4(32'hbc0a6ad4),
	.w5(32'hbc1d4e1d),
	.w6(32'h3b9579ce),
	.w7(32'hbc4c6ea8),
	.w8(32'hbc048aae),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace07b5),
	.w1(32'hbba423ac),
	.w2(32'h3c17a289),
	.w3(32'hbc12627d),
	.w4(32'h3983c7e9),
	.w5(32'hbc8c0fbd),
	.w6(32'hbc3b56cb),
	.w7(32'h3a81b2ec),
	.w8(32'hbb7395bc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3cd91),
	.w1(32'h3b54122f),
	.w2(32'h3907384b),
	.w3(32'h3b659ae5),
	.w4(32'hbb34578d),
	.w5(32'hbbdd49d4),
	.w6(32'h3b08bc12),
	.w7(32'hbb94a5f6),
	.w8(32'h3b5213ff),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7fe36),
	.w1(32'h3c5c85a9),
	.w2(32'h3c831841),
	.w3(32'h3be0cf74),
	.w4(32'h3c749374),
	.w5(32'h3ca5a4e3),
	.w6(32'hbbea3e84),
	.w7(32'h3b2d19bf),
	.w8(32'h3aac3434),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82f76d),
	.w1(32'h3c54314c),
	.w2(32'hbbb8a73f),
	.w3(32'hbc57395d),
	.w4(32'h3cab46e2),
	.w5(32'hbca1b1a0),
	.w6(32'hbc1e4899),
	.w7(32'h3b0e3364),
	.w8(32'h3cc433e2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20a5c1),
	.w1(32'hbc08ef02),
	.w2(32'hbae9b6cf),
	.w3(32'h3cd3178e),
	.w4(32'hbc8b6e71),
	.w5(32'hbbb57ac0),
	.w6(32'hbb0bd5d0),
	.w7(32'hbb3e0ae2),
	.w8(32'hba595bc9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ea4a3),
	.w1(32'h3ba3e18a),
	.w2(32'h3b660e84),
	.w3(32'h3c87a5fd),
	.w4(32'h3b1d0918),
	.w5(32'hba832b93),
	.w6(32'h3b66f39c),
	.w7(32'h3bb2b047),
	.w8(32'h3abc00c4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35d80),
	.w1(32'h3ba163d2),
	.w2(32'hbbcb0d96),
	.w3(32'h3a3629b0),
	.w4(32'h3c7cab88),
	.w5(32'hbb99ac20),
	.w6(32'h3ba6ac34),
	.w7(32'h3c26f7bf),
	.w8(32'h3b4403e1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0d29),
	.w1(32'hbc614108),
	.w2(32'hbcbd8f38),
	.w3(32'hbc9a7de1),
	.w4(32'hbb302c0e),
	.w5(32'h3c55cb1d),
	.w6(32'hbbcd7912),
	.w7(32'h3b0a0455),
	.w8(32'h3ca886ed),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee3cb9),
	.w1(32'hba4361b3),
	.w2(32'hbc123ad8),
	.w3(32'h3bf18012),
	.w4(32'hbb581073),
	.w5(32'hbc13d770),
	.w6(32'h3abe1586),
	.w7(32'hba6db4ed),
	.w8(32'h3c205299),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cbb41),
	.w1(32'hbbd3d9dc),
	.w2(32'hbbefbc74),
	.w3(32'hbc428b95),
	.w4(32'h3bf59be2),
	.w5(32'hbb08e805),
	.w6(32'h3b237ce2),
	.w7(32'hbc8e7926),
	.w8(32'hbc13c238),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca294d8),
	.w1(32'h3b8044f0),
	.w2(32'h3b60b2c9),
	.w3(32'hbcdb49fb),
	.w4(32'hbbab8fe1),
	.w5(32'h3ce6f63e),
	.w6(32'hbc8a51f1),
	.w7(32'hbbce14b7),
	.w8(32'hbb8a3f22),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a960abc),
	.w1(32'h3b17b228),
	.w2(32'hbb32c10c),
	.w3(32'hbb1cc525),
	.w4(32'hbba09f60),
	.w5(32'hbc0562db),
	.w6(32'hbab22593),
	.w7(32'hbc0f4699),
	.w8(32'h3b9ebe84),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b085),
	.w1(32'h3be5c64f),
	.w2(32'h3cf79bb2),
	.w3(32'h3ad9062b),
	.w4(32'h3cf1bc2e),
	.w5(32'h3d6cbff0),
	.w6(32'h3b83990b),
	.w7(32'h3bfe927d),
	.w8(32'h3a8f7b69),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd58d59),
	.w1(32'h3bad90d4),
	.w2(32'hbb42af32),
	.w3(32'h3c5a4af3),
	.w4(32'h3bf920e4),
	.w5(32'h3c92ce1f),
	.w6(32'h3c372782),
	.w7(32'h3a00aa18),
	.w8(32'h3be3e428),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833a3a),
	.w1(32'h3b651e88),
	.w2(32'hbbb7da46),
	.w3(32'hbc71d6e2),
	.w4(32'h3c713b1d),
	.w5(32'h3c62ef5f),
	.w6(32'hbbe6f371),
	.w7(32'hbad23877),
	.w8(32'h3cf33772),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5a3e7),
	.w1(32'h3c4f262b),
	.w2(32'hbbe5752f),
	.w3(32'h3c7afc27),
	.w4(32'h3b5bc474),
	.w5(32'hbc1f496f),
	.w6(32'h3c5491f3),
	.w7(32'h3b25ca2d),
	.w8(32'h3c3bfafc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25d364),
	.w1(32'hb9bc9011),
	.w2(32'hbaa8ce85),
	.w3(32'hbb2e881f),
	.w4(32'hba62f3ab),
	.w5(32'hbbfa4fd9),
	.w6(32'h395aed55),
	.w7(32'h3b0495ee),
	.w8(32'hbbbb60ac),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9c05),
	.w1(32'hba1866da),
	.w2(32'h3b783d1a),
	.w3(32'hbbf482ee),
	.w4(32'hbbba7a2b),
	.w5(32'h3b8ae04e),
	.w6(32'hbc4b9210),
	.w7(32'hbc8512c3),
	.w8(32'h3a5371f6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule