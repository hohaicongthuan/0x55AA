module layer_8_featuremap_202(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc934db5),
	.w1(32'h3b5c20fe),
	.w2(32'hbae1acb1),
	.w3(32'hbc617878),
	.w4(32'hba59265b),
	.w5(32'h3b95c6af),
	.w6(32'hbba5b2e9),
	.w7(32'hbb9944d8),
	.w8(32'h3baa8da0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb388c14),
	.w1(32'h3b52eeec),
	.w2(32'h3b0a899d),
	.w3(32'hbafc25af),
	.w4(32'hbb4f4150),
	.w5(32'hba9c5580),
	.w6(32'hbbaac6a2),
	.w7(32'hbbd39723),
	.w8(32'h3b280c5a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22c76d),
	.w1(32'hbbd59b6a),
	.w2(32'hbbd661c0),
	.w3(32'h3ba54ff2),
	.w4(32'hbbcc71a9),
	.w5(32'hbab7a970),
	.w6(32'hbbaa0bcc),
	.w7(32'hbc849686),
	.w8(32'hbc2efabb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24dc74),
	.w1(32'hbba0f7dc),
	.w2(32'hbb7b2813),
	.w3(32'hbbd1361d),
	.w4(32'hb9fadb0e),
	.w5(32'h3b374924),
	.w6(32'hbb8e8fe6),
	.w7(32'hbc20ca14),
	.w8(32'hbb3fb6bb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f173b),
	.w1(32'h3ba5116e),
	.w2(32'h399ef345),
	.w3(32'hbb973fff),
	.w4(32'h3c826719),
	.w5(32'h3c92ca90),
	.w6(32'hbc3030b2),
	.w7(32'hbc873d25),
	.w8(32'hbbd3454c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a1d9),
	.w1(32'hbb33d013),
	.w2(32'hbb9f9d7b),
	.w3(32'h3c80f876),
	.w4(32'hbb9240e0),
	.w5(32'hba97e081),
	.w6(32'h3bb54fad),
	.w7(32'h3b00e55e),
	.w8(32'hbc21ff58),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968204a),
	.w1(32'hbb4715b6),
	.w2(32'hbb760af9),
	.w3(32'h3bffb3b7),
	.w4(32'h3b6dd119),
	.w5(32'h3b04a77a),
	.w6(32'hbb5b7d3a),
	.w7(32'hbc1b2d5d),
	.w8(32'hbbe260cd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6600ea),
	.w1(32'hbaa8561b),
	.w2(32'hbbfe42a4),
	.w3(32'h3acbdc30),
	.w4(32'h3ad9845c),
	.w5(32'h3bf6e8ed),
	.w6(32'hbbd7c684),
	.w7(32'hbbe487f6),
	.w8(32'hbbe037d5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08862f),
	.w1(32'h3c31935b),
	.w2(32'h39899553),
	.w3(32'h3b074db7),
	.w4(32'h3ce7715f),
	.w5(32'h3d055179),
	.w6(32'hbd1cb87e),
	.w7(32'hbd540c7e),
	.w8(32'hbd0fb9d6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ed74b),
	.w1(32'hbba3719c),
	.w2(32'hbc4fda01),
	.w3(32'h3cbb6085),
	.w4(32'hbc9ad7cc),
	.w5(32'hbca8b49b),
	.w6(32'h3c1fd9eb),
	.w7(32'hbbabb097),
	.w8(32'h3bbb514b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8c3e),
	.w1(32'hbb39ed71),
	.w2(32'hba971ff1),
	.w3(32'hbc90d546),
	.w4(32'h3c1ab11d),
	.w5(32'h3c082f9d),
	.w6(32'hbc19ba56),
	.w7(32'hbc2180d6),
	.w8(32'hbc21301e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67cf5a),
	.w1(32'h3b035f90),
	.w2(32'hbbdc586d),
	.w3(32'h3aa36dde),
	.w4(32'hba7b76a7),
	.w5(32'hbc6e9e82),
	.w6(32'h3ba02784),
	.w7(32'hba0cc16e),
	.w8(32'h3c53406f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22b80a),
	.w1(32'h3c1ea354),
	.w2(32'h3b841976),
	.w3(32'hbbcc87c1),
	.w4(32'h3bb6fb06),
	.w5(32'h3c08ddcf),
	.w6(32'h3aa055ec),
	.w7(32'hbb4a0a78),
	.w8(32'hbb25be73),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b7217),
	.w1(32'hba804d9b),
	.w2(32'h3acf6c4a),
	.w3(32'h3c1f85d7),
	.w4(32'hbb0ec1f7),
	.w5(32'hbae47854),
	.w6(32'hbb461ecd),
	.w7(32'hbbc76026),
	.w8(32'hbb8af557),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb704c094),
	.w1(32'hbbb41bd9),
	.w2(32'hbb55ee51),
	.w3(32'hbb2a07e0),
	.w4(32'h3c67326a),
	.w5(32'h3c95adda),
	.w6(32'hbcc47c10),
	.w7(32'hbce694e2),
	.w8(32'hbce0d7c5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba646fd),
	.w1(32'h3c4c1cce),
	.w2(32'h3c15cc31),
	.w3(32'h3c574cc2),
	.w4(32'h3ad8e7e3),
	.w5(32'hbbaff7b4),
	.w6(32'hbb67bbb4),
	.w7(32'h3b050949),
	.w8(32'h3b0f05f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c4260),
	.w1(32'h3b313155),
	.w2(32'hbad6f5bc),
	.w3(32'hbb244d80),
	.w4(32'hbb7bdf31),
	.w5(32'hbc36ef42),
	.w6(32'hba8adc58),
	.w7(32'hba546dcc),
	.w8(32'hbbe59d30),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82b392),
	.w1(32'hb91b1580),
	.w2(32'h3b6d6530),
	.w3(32'hbb95b1fb),
	.w4(32'hba04a917),
	.w5(32'h3b89b541),
	.w6(32'h3b0cfe77),
	.w7(32'h3b192856),
	.w8(32'h3c02cf2e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96d87),
	.w1(32'h3c649ac0),
	.w2(32'h3c778780),
	.w3(32'h3c48d1f7),
	.w4(32'h3c3f03bf),
	.w5(32'h3c653a70),
	.w6(32'h3c8d54d4),
	.w7(32'h3bd7a2b0),
	.w8(32'h3beb5991),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088c8b),
	.w1(32'h3c1464de),
	.w2(32'h3c167056),
	.w3(32'h3c0ce944),
	.w4(32'h3cdb70fe),
	.w5(32'h3ce321ee),
	.w6(32'h3b416471),
	.w7(32'hbbc0df6d),
	.w8(32'hbc2079a1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3303a0),
	.w1(32'h3ba546d4),
	.w2(32'h3c849f1a),
	.w3(32'h3c5366f7),
	.w4(32'h3be59521),
	.w5(32'h3c1b04ae),
	.w6(32'h3c3ca375),
	.w7(32'h3c11ed23),
	.w8(32'h3c638b4e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c570c9e),
	.w1(32'hbb1b780c),
	.w2(32'hbb59f15e),
	.w3(32'h3b49c7cf),
	.w4(32'h3b975b61),
	.w5(32'h3bc36123),
	.w6(32'hbc7d4fc8),
	.w7(32'hbb9d52eb),
	.w8(32'hbb70adec),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01818d),
	.w1(32'h3c4888af),
	.w2(32'h3c5f40c9),
	.w3(32'h3c2ae431),
	.w4(32'h3c3fb5c1),
	.w5(32'h3c7813e6),
	.w6(32'hbc0bf1af),
	.w7(32'hbc35c836),
	.w8(32'h3bfbe74f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef4554),
	.w1(32'h3b468994),
	.w2(32'hb987df59),
	.w3(32'hb9b7b79d),
	.w4(32'hbb0fb797),
	.w5(32'h3bbbcb8c),
	.w6(32'h382c7038),
	.w7(32'h3ad60c34),
	.w8(32'hbb32731a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a5a7),
	.w1(32'h3c9e19d3),
	.w2(32'h3d1952b6),
	.w3(32'h3ba73fa3),
	.w4(32'h3cad452f),
	.w5(32'h3d09aac1),
	.w6(32'h3c65fbb6),
	.w7(32'h3cd4780a),
	.w8(32'h3c9547da),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cef3fc2),
	.w1(32'h3bf776ca),
	.w2(32'h3c90514d),
	.w3(32'h3cce1daa),
	.w4(32'h3c8e04fe),
	.w5(32'h3ce02f9f),
	.w6(32'h3bb8bb7a),
	.w7(32'h3bd16eda),
	.w8(32'h3bd19096),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7e06),
	.w1(32'hbb84fc5c),
	.w2(32'hbc78d889),
	.w3(32'h3c0a2efc),
	.w4(32'hbbd444a2),
	.w5(32'hbc446505),
	.w6(32'h3a0e79fb),
	.w7(32'h3bfbbefa),
	.w8(32'h3b130d5d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd840049),
	.w1(32'h3c26db8c),
	.w2(32'h3d4779f3),
	.w3(32'hbc4ec9e4),
	.w4(32'h3da2625d),
	.w5(32'h3d62b5de),
	.w6(32'h3d82b893),
	.w7(32'h3db9fea7),
	.w8(32'h3d1aeaa7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d4e7d),
	.w1(32'h3a56afd2),
	.w2(32'hbc326762),
	.w3(32'h3bd5b5ea),
	.w4(32'hbc522cb8),
	.w5(32'hbca96cf6),
	.w6(32'hbc2a776a),
	.w7(32'hbcb5d4a7),
	.w8(32'hbcc3e3a9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1477b),
	.w1(32'h3ac44b15),
	.w2(32'h3b470144),
	.w3(32'h3b456b51),
	.w4(32'h3cb103ef),
	.w5(32'h3ccff81b),
	.w6(32'h3a86916c),
	.w7(32'hbb07593c),
	.w8(32'h3bdf1c40),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aec1e),
	.w1(32'hbcec0741),
	.w2(32'hbd31ab49),
	.w3(32'h3cc5c2f1),
	.w4(32'hbcd7a53c),
	.w5(32'hbd255fd2),
	.w6(32'hbcab657f),
	.w7(32'hbd08a2ef),
	.w8(32'hbcf67813),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc79e7),
	.w1(32'h3c11fafe),
	.w2(32'h3c299f50),
	.w3(32'hbcfcd678),
	.w4(32'h3c3b8d29),
	.w5(32'h3c129862),
	.w6(32'hbbd3f927),
	.w7(32'hbc50971e),
	.w8(32'hbc58a009),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3160),
	.w1(32'h3bb23ac9),
	.w2(32'h3c271087),
	.w3(32'h3bf8db34),
	.w4(32'h3bc4b1c7),
	.w5(32'h3bc30233),
	.w6(32'h3b84a46f),
	.w7(32'h3c2ba9b9),
	.w8(32'h390f8728),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed67a),
	.w1(32'hb81af092),
	.w2(32'hbb46ca35),
	.w3(32'hbb415997),
	.w4(32'hbbb25cd7),
	.w5(32'hbb407742),
	.w6(32'h39817907),
	.w7(32'h39c8feda),
	.w8(32'h3a168050),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb671fad),
	.w1(32'hbc3fb127),
	.w2(32'hbc6597fa),
	.w3(32'h3c07a55f),
	.w4(32'hba8430ac),
	.w5(32'hbb89f761),
	.w6(32'h392ed5fb),
	.w7(32'h3a4db6e2),
	.w8(32'h3b39e196),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80e5fb),
	.w1(32'h3acb5d2c),
	.w2(32'h3bb07fea),
	.w3(32'hbbedf7c3),
	.w4(32'h3b582d73),
	.w5(32'hba2c5923),
	.w6(32'h3c096e07),
	.w7(32'h3bbd6fa3),
	.w8(32'h3a5efcd7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb1aab),
	.w1(32'h3c910b8c),
	.w2(32'h3cb219e5),
	.w3(32'hbc0ac9f8),
	.w4(32'h3cb99f70),
	.w5(32'h3ce1b954),
	.w6(32'h3c99addf),
	.w7(32'h3cc7eaf2),
	.w8(32'h3c9bc336),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91012a),
	.w1(32'hbbf092f0),
	.w2(32'hbb9b75dc),
	.w3(32'h3cbb72ee),
	.w4(32'h3c1b757c),
	.w5(32'h3c6e5166),
	.w6(32'hbcd8a6cd),
	.w7(32'hbcf9ca46),
	.w8(32'hbcb78ad4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47514),
	.w1(32'hb993e8ef),
	.w2(32'h3b60794a),
	.w3(32'h3c1fc1d0),
	.w4(32'h3b3b0f33),
	.w5(32'h3b200c6a),
	.w6(32'hb9b4e23b),
	.w7(32'hbb3a7b6b),
	.w8(32'hbb412da3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7620),
	.w1(32'h3aa1958f),
	.w2(32'h3a0d1107),
	.w3(32'h3aa0993f),
	.w4(32'hbb38d22a),
	.w5(32'hbbc7b79a),
	.w6(32'h3b7ec94b),
	.w7(32'hba5d7aa9),
	.w8(32'h3b2bd9d8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff727),
	.w1(32'h3b22be64),
	.w2(32'hbab09e7a),
	.w3(32'hbbc8b5aa),
	.w4(32'hbb35dbdf),
	.w5(32'hbc04dd62),
	.w6(32'h3bba48da),
	.w7(32'h3ae3cb34),
	.w8(32'h3bbd0cb4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aea8b),
	.w1(32'h39d9ef31),
	.w2(32'h39acbefd),
	.w3(32'h3a20ea4a),
	.w4(32'h3bdee260),
	.w5(32'hbbc9bace),
	.w6(32'hbc60da7d),
	.w7(32'hbc2c334b),
	.w8(32'hbb91cb2e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a336a4f),
	.w1(32'h3c574131),
	.w2(32'h3c7d526c),
	.w3(32'hbc8a20ea),
	.w4(32'h3c13c034),
	.w5(32'h3c25cd4d),
	.w6(32'h3c20b65a),
	.w7(32'h3c130e40),
	.w8(32'h3c28f7a8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b8296),
	.w1(32'h3bc024cf),
	.w2(32'h3aa2a885),
	.w3(32'h3c5a347c),
	.w4(32'h3bd068c9),
	.w5(32'hbb30b82d),
	.w6(32'h3ba54c4b),
	.w7(32'h39e1e66f),
	.w8(32'h3ad5a1a7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c168),
	.w1(32'h3c53f5da),
	.w2(32'h3c6a11c7),
	.w3(32'h3c002ba1),
	.w4(32'h3c3d7ad5),
	.w5(32'h3c69c5f7),
	.w6(32'h3bee66f6),
	.w7(32'h3bf38eb9),
	.w8(32'h3bd86cd2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318637),
	.w1(32'h3bc7d3cd),
	.w2(32'h3b87223d),
	.w3(32'hbb1404c9),
	.w4(32'h3bc7aa6a),
	.w5(32'h3b321b39),
	.w6(32'h3b7c8807),
	.w7(32'hba780a1e),
	.w8(32'hb998bdcb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278bdb),
	.w1(32'hbadf54bf),
	.w2(32'hbb0a8bb3),
	.w3(32'h3b52b86b),
	.w4(32'hbbb250c1),
	.w5(32'hbb4b7eaf),
	.w6(32'hbc072a7e),
	.w7(32'hbbd57a83),
	.w8(32'hbc09f2f7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55a55),
	.w1(32'h3c0ee244),
	.w2(32'h3c637baa),
	.w3(32'h3ae0ef8f),
	.w4(32'h3c857a6c),
	.w5(32'h3c74590a),
	.w6(32'h3c1167a6),
	.w7(32'h3c5f6c87),
	.w8(32'h3c4d1af6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b0b2d),
	.w1(32'hbbbad053),
	.w2(32'hbc01d135),
	.w3(32'hbaead703),
	.w4(32'hbbd6bd6a),
	.w5(32'hbba0cf24),
	.w6(32'hbbc37a86),
	.w7(32'hbb9ddfda),
	.w8(32'hbb0293bb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07702b),
	.w1(32'h3c1189ce),
	.w2(32'h3af6d0a0),
	.w3(32'h3acf4fe6),
	.w4(32'h3b92c3d4),
	.w5(32'hba635ebb),
	.w6(32'hbb0f9ce9),
	.w7(32'hba752e59),
	.w8(32'h3b4ea69b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5cf23),
	.w1(32'h3b96a398),
	.w2(32'h3a99aae2),
	.w3(32'h3a859e8b),
	.w4(32'hba733755),
	.w5(32'hbc222044),
	.w6(32'hbbf6b73d),
	.w7(32'hbbe32e92),
	.w8(32'h3b06d6a6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c837056),
	.w1(32'h3cd0d0ca),
	.w2(32'h3c6e6d74),
	.w3(32'h3c382171),
	.w4(32'h3cdd1ae7),
	.w5(32'h3cc18567),
	.w6(32'h3c4dee2a),
	.w7(32'h3c121dac),
	.w8(32'h3cba13f3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50978f),
	.w1(32'h3c063e4e),
	.w2(32'h3c077927),
	.w3(32'h3be4870c),
	.w4(32'h3c6abcd3),
	.w5(32'h3c941b0e),
	.w6(32'hbba03189),
	.w7(32'hbc3c40d3),
	.w8(32'hb98e6b91),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3b6c8),
	.w1(32'h3befe878),
	.w2(32'h3bf84e48),
	.w3(32'h3c3ca99d),
	.w4(32'hba693a74),
	.w5(32'h3b889592),
	.w6(32'h3c07c4a1),
	.w7(32'h3c4050e8),
	.w8(32'h3b38820b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd51f5),
	.w1(32'h3b9bbf3a),
	.w2(32'hbb2dfdc9),
	.w3(32'h39dd0b7a),
	.w4(32'h3b9fd382),
	.w5(32'hbba487ab),
	.w6(32'h3a28b170),
	.w7(32'h3b16ccf1),
	.w8(32'h3af64743),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac94457),
	.w1(32'h3c59ff28),
	.w2(32'h3c331f5a),
	.w3(32'hbb57f0fc),
	.w4(32'h3bafc4db),
	.w5(32'h3c585ae7),
	.w6(32'hbb4152e7),
	.w7(32'hbb98d522),
	.w8(32'h3c2bdb50),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd388),
	.w1(32'hba8ccf13),
	.w2(32'hbb90667b),
	.w3(32'h3c2e52ac),
	.w4(32'hbb393f5a),
	.w5(32'hbb9a638a),
	.w6(32'hbbb7b9ba),
	.w7(32'hbb3b9afe),
	.w8(32'h3acdb83d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3de4c),
	.w1(32'hbb483845),
	.w2(32'hbc107d4c),
	.w3(32'hbc300eda),
	.w4(32'hb9c7fe92),
	.w5(32'h3bcf309b),
	.w6(32'hbbb333ac),
	.w7(32'hbc981387),
	.w8(32'h39f8f2de),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc253b0),
	.w1(32'hbb65964b),
	.w2(32'hbb0e06b0),
	.w3(32'h3bb8f058),
	.w4(32'hbc0d156b),
	.w5(32'hbc10f006),
	.w6(32'hb9db2201),
	.w7(32'h3a7bb0a7),
	.w8(32'hb758b235),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9daaec),
	.w1(32'hbae5e4f3),
	.w2(32'hb9bf217a),
	.w3(32'hbc09642a),
	.w4(32'hbb374c07),
	.w5(32'h39c472fb),
	.w6(32'hbaa608b8),
	.w7(32'hbb79623e),
	.w8(32'hbc276227),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87ec6),
	.w1(32'h3bb18d7c),
	.w2(32'h3c574452),
	.w3(32'hbb3e0bd3),
	.w4(32'h3b829b66),
	.w5(32'h3c437184),
	.w6(32'hbaf60423),
	.w7(32'hbbf504b6),
	.w8(32'hbba33b84),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2c2fc),
	.w1(32'h3d07de47),
	.w2(32'h3d48688a),
	.w3(32'h3c6cc19f),
	.w4(32'h3d19fd5c),
	.w5(32'h3d68fd2e),
	.w6(32'h3c92d1d9),
	.w7(32'h3cc1f77b),
	.w8(32'h3c79c553),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10f546),
	.w1(32'h3b833f94),
	.w2(32'h38c147dc),
	.w3(32'h3d45ad70),
	.w4(32'hbb5ee491),
	.w5(32'hbbc25754),
	.w6(32'hbb0a72bb),
	.w7(32'hbc319145),
	.w8(32'hbc4c91d0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c4ac2),
	.w1(32'hbc5599a3),
	.w2(32'hbcac70c2),
	.w3(32'hbc07e043),
	.w4(32'hbc2ff71e),
	.w5(32'hbc8fde90),
	.w6(32'h39059c5a),
	.w7(32'hbb9ce5b7),
	.w8(32'hba1c7ccc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a8715),
	.w1(32'h3b394fe7),
	.w2(32'h3bbba6c1),
	.w3(32'hbc331ceb),
	.w4(32'hbb9e82e3),
	.w5(32'hbbaf9970),
	.w6(32'h3a483add),
	.w7(32'h3bb472f8),
	.w8(32'hba92cf59),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2368e2),
	.w1(32'hbb2638d2),
	.w2(32'hbb274c29),
	.w3(32'hbbafe276),
	.w4(32'hbad203db),
	.w5(32'hbb4632f7),
	.w6(32'hbae91e8d),
	.w7(32'hbb8a53ca),
	.w8(32'h3a11248f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2cf80),
	.w1(32'hba965791),
	.w2(32'hba4cd651),
	.w3(32'hbb8939e4),
	.w4(32'h3bb54beb),
	.w5(32'h3aa55eb1),
	.w6(32'h3a14b26a),
	.w7(32'hbbd0dfd1),
	.w8(32'hbb179912),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499a0a),
	.w1(32'h3bfc82f1),
	.w2(32'h3bfe01d7),
	.w3(32'h3c5fc378),
	.w4(32'h3c401343),
	.w5(32'h3c1cf767),
	.w6(32'h3c29d304),
	.w7(32'h3b3f2c2c),
	.w8(32'hbadbce2c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad31a3),
	.w1(32'h3b8ab5da),
	.w2(32'h3b677ac0),
	.w3(32'h3bd1f25b),
	.w4(32'hbbccd698),
	.w5(32'h3a17187e),
	.w6(32'h383becd5),
	.w7(32'hbba4cf6b),
	.w8(32'hb9a4d5cc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ca5ba),
	.w1(32'h3ba523b9),
	.w2(32'h3c34049e),
	.w3(32'h3adbad44),
	.w4(32'h3c517c73),
	.w5(32'h3c88d881),
	.w6(32'h3a8255cf),
	.w7(32'hbc4816c3),
	.w8(32'hbbfa8052),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec73f),
	.w1(32'hbc0085a2),
	.w2(32'hbc329579),
	.w3(32'h3b25cbe7),
	.w4(32'h3b9e830f),
	.w5(32'hbb3de9c0),
	.w6(32'hbcc73299),
	.w7(32'hbcc771cf),
	.w8(32'hbbb8fc40),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a268528),
	.w1(32'h3be100d0),
	.w2(32'h3afa5e8e),
	.w3(32'hbc0a67b9),
	.w4(32'h3babcca5),
	.w5(32'h3bac0cd3),
	.w6(32'h3ad7e42a),
	.w7(32'hb94aa8eb),
	.w8(32'h3b95fa89),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf696),
	.w1(32'hbb931d80),
	.w2(32'hbb644ca7),
	.w3(32'hbb53886a),
	.w4(32'h3b9002b9),
	.w5(32'h3b5af45a),
	.w6(32'hbadfe383),
	.w7(32'hbc1df633),
	.w8(32'hbbe07fd2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33a877),
	.w1(32'hbc511bc2),
	.w2(32'hbca99c1c),
	.w3(32'hbb5fa92c),
	.w4(32'hbba04c82),
	.w5(32'hbbce6cb6),
	.w6(32'hbc653fb2),
	.w7(32'hbcddb161),
	.w8(32'hbc217599),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb685),
	.w1(32'h3c9fb2f1),
	.w2(32'h3d0ce8f9),
	.w3(32'hbbdbe647),
	.w4(32'h3ca13fe3),
	.w5(32'h3d0efd98),
	.w6(32'h3c90d5a1),
	.w7(32'h3cdb2660),
	.w8(32'h3cd4280a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1115ae),
	.w1(32'h3c2cb35b),
	.w2(32'h3c3ac325),
	.w3(32'h3cb198e0),
	.w4(32'h3c31f057),
	.w5(32'h3c1f4ddd),
	.w6(32'h3b866753),
	.w7(32'hbb446023),
	.w8(32'h3bc79952),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd277ae),
	.w1(32'hbaeaad5b),
	.w2(32'hbbc673ed),
	.w3(32'h3b91d815),
	.w4(32'hbaed4691),
	.w5(32'hbbdb139f),
	.w6(32'h3b2a6470),
	.w7(32'hbbfca1d4),
	.w8(32'hba662886),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93b55b),
	.w1(32'h3c120797),
	.w2(32'hbb273368),
	.w3(32'hb927d3df),
	.w4(32'h3bc11856),
	.w5(32'hbb8b63aa),
	.w6(32'h3bd60ee7),
	.w7(32'hbbc01ab8),
	.w8(32'h3acf6d6a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdda9a5),
	.w1(32'hbc1f3d6b),
	.w2(32'hbccf3abe),
	.w3(32'h3a8b6f41),
	.w4(32'h3b17a9ac),
	.w5(32'hbc791c98),
	.w6(32'hbc54a8e4),
	.w7(32'hbc9a72d2),
	.w8(32'hb7a660dc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b234),
	.w1(32'h3bbe0dbe),
	.w2(32'hbbaf0840),
	.w3(32'hbc87c5d2),
	.w4(32'h3b8d9f4a),
	.w5(32'h3ae5dc36),
	.w6(32'h3b558e19),
	.w7(32'hbb234d34),
	.w8(32'hbc02b633),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff7f2d),
	.w1(32'h391095b5),
	.w2(32'hbb0889b8),
	.w3(32'hbb8136f5),
	.w4(32'h3b9f76ac),
	.w5(32'h3a7fbff6),
	.w6(32'hbbfd20c0),
	.w7(32'hbc0e3b6b),
	.w8(32'hbb62adfb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74a9a9),
	.w1(32'hbb6a1936),
	.w2(32'h3a8c170a),
	.w3(32'h3a7303a2),
	.w4(32'hbb4b14eb),
	.w5(32'hbb70d339),
	.w6(32'h3b167649),
	.w7(32'h3b2984a2),
	.w8(32'hbab58cd4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85a7e7),
	.w1(32'h3c473a5a),
	.w2(32'h3c6441f8),
	.w3(32'h3b7f48bd),
	.w4(32'h3b86e986),
	.w5(32'h3c656c94),
	.w6(32'h3bc56304),
	.w7(32'h3b84abff),
	.w8(32'h3b808111),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2952),
	.w1(32'hb92cfe6c),
	.w2(32'h3b4b09eb),
	.w3(32'h3c0c21bd),
	.w4(32'h3b96ef22),
	.w5(32'h3b917c33),
	.w6(32'h3b7221e8),
	.w7(32'h3c2fb557),
	.w8(32'h3bc16f52),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f3c0),
	.w1(32'h3c79208f),
	.w2(32'h3c7ff5f7),
	.w3(32'h3b9e9bb7),
	.w4(32'h3c904cd2),
	.w5(32'h3cbc84a4),
	.w6(32'h3b2ae6db),
	.w7(32'hbc1d718f),
	.w8(32'h3bb2195f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42a930),
	.w1(32'h3c2af8f2),
	.w2(32'h3c0f2aad),
	.w3(32'h3ab111b9),
	.w4(32'h3c98fee7),
	.w5(32'h3c8a486b),
	.w6(32'hbc3462a5),
	.w7(32'hbb800fce),
	.w8(32'hbc12b24f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef841c),
	.w1(32'hbceb67bf),
	.w2(32'hbd37240e),
	.w3(32'h3c6ccbf3),
	.w4(32'hbd13ff89),
	.w5(32'hbd4e41f1),
	.w6(32'hbcd3caa5),
	.w7(32'hbd0fa079),
	.w8(32'hbcfc13a7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20c80d),
	.w1(32'h3d42dbcb),
	.w2(32'h3d8a9fa5),
	.w3(32'hbd40defa),
	.w4(32'h3d19ed4a),
	.w5(32'h3d5fc557),
	.w6(32'h3d1c8f40),
	.w7(32'h3d578f26),
	.w8(32'h3d1e6902),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d60115f),
	.w1(32'hbd4429f4),
	.w2(32'hbd816a13),
	.w3(32'h3d32fb7f),
	.w4(32'hbd2035ad),
	.w5(32'hbd57edd6),
	.w6(32'hbcefd9d2),
	.w7(32'hbd1c0c70),
	.w8(32'hbd0a9968),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd68a97b),
	.w1(32'h3b13996f),
	.w2(32'hbb94a77c),
	.w3(32'hbd5328da),
	.w4(32'hbc27bf1e),
	.w5(32'hbc454969),
	.w6(32'hbc13015b),
	.w7(32'hbba430f8),
	.w8(32'hbc123820),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47fc6a),
	.w1(32'hbb6ec260),
	.w2(32'hbbb9daa5),
	.w3(32'hbc6551c2),
	.w4(32'h3929529d),
	.w5(32'hba6bbefa),
	.w6(32'hbb9f72fa),
	.w7(32'h3a345c96),
	.w8(32'h3b936607),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb564ac5),
	.w1(32'h39b0eeb9),
	.w2(32'hba744874),
	.w3(32'h38825009),
	.w4(32'h3b4d92be),
	.w5(32'hbc2a0f18),
	.w6(32'h3ade1e91),
	.w7(32'hbaabae3a),
	.w8(32'h3b7472d4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced5ce),
	.w1(32'h37d9a511),
	.w2(32'hbb6cd356),
	.w3(32'hba58cf53),
	.w4(32'hbaca83cc),
	.w5(32'hbaa81e3a),
	.w6(32'h3c2ae4ce),
	.w7(32'h3c079c5c),
	.w8(32'h3c1965a9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c5a53),
	.w1(32'h3b3d85ba),
	.w2(32'h3b391f62),
	.w3(32'hbaf536eb),
	.w4(32'hbbc87ccf),
	.w5(32'hbc0470fc),
	.w6(32'h3bdc683d),
	.w7(32'h3bf0b358),
	.w8(32'h3c11f095),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b745403),
	.w1(32'h3c0c56f2),
	.w2(32'hbb7ffa95),
	.w3(32'hbbf3831d),
	.w4(32'h3ca54798),
	.w5(32'h3c4ec041),
	.w6(32'hb909f8d2),
	.w7(32'hbc55c27b),
	.w8(32'hb9480724),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1a878),
	.w1(32'hbc7fe80d),
	.w2(32'hbcd8e22e),
	.w3(32'h3c1c1e2d),
	.w4(32'hbc852c2c),
	.w5(32'hbcd654fd),
	.w6(32'hbc6cbdd6),
	.w7(32'hbcc2ab9d),
	.w8(32'hbcb18ddc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc518f1d),
	.w1(32'h3c9e5b74),
	.w2(32'h3c954b4e),
	.w3(32'hbc69ea00),
	.w4(32'h3c6a252c),
	.w5(32'h3c648542),
	.w6(32'h3c64e1dd),
	.w7(32'h3c5a118c),
	.w8(32'h3c964fc7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdadb31),
	.w1(32'h3ba7c648),
	.w2(32'h3c166631),
	.w3(32'hbb95e2e7),
	.w4(32'hb98b9759),
	.w5(32'h3b92c153),
	.w6(32'h3a450e93),
	.w7(32'hbb09acb9),
	.w8(32'hbaad4299),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6c50a),
	.w1(32'h3bb1c387),
	.w2(32'hbb1c8e84),
	.w3(32'hbb15a41f),
	.w4(32'h3b50bfb7),
	.w5(32'h3acda31a),
	.w6(32'h3b764794),
	.w7(32'h3b3bc986),
	.w8(32'h3bf3f4b2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2e88c),
	.w1(32'hbc0fba69),
	.w2(32'hbc3be3a3),
	.w3(32'h3b835ed6),
	.w4(32'hbbbcce39),
	.w5(32'hbc55bdd5),
	.w6(32'hbc829b88),
	.w7(32'hbc201f37),
	.w8(32'h3b621776),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d298b),
	.w1(32'hbad28bdf),
	.w2(32'h3c054203),
	.w3(32'hbb90c6e0),
	.w4(32'h3aa8bbee),
	.w5(32'hb9d62053),
	.w6(32'h3b97f9a2),
	.w7(32'h3bfb1e32),
	.w8(32'h3b873763),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67612),
	.w1(32'hba556f9a),
	.w2(32'h3c3993e0),
	.w3(32'h3b82df24),
	.w4(32'h3b8c7a8b),
	.w5(32'h3b677c43),
	.w6(32'hba220a37),
	.w7(32'h3bb60796),
	.w8(32'h3c3de3de),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42d528),
	.w1(32'h3b002ce4),
	.w2(32'h3c3a8459),
	.w3(32'h3c5423c4),
	.w4(32'h3baf7950),
	.w5(32'hbb40b6d8),
	.w6(32'h3be407ae),
	.w7(32'h3bc88b0f),
	.w8(32'h3b9c3f12),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5958a),
	.w1(32'hbc29c3ca),
	.w2(32'hbbf2b71d),
	.w3(32'h3ba89486),
	.w4(32'hbc833cea),
	.w5(32'hbc80e49e),
	.w6(32'h3bce4354),
	.w7(32'hbaecc227),
	.w8(32'hbb93a1a5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe522c3),
	.w1(32'h3b640991),
	.w2(32'h3bde93a6),
	.w3(32'hbc0952f9),
	.w4(32'h3b885e07),
	.w5(32'hba96ffef),
	.w6(32'h3b07b929),
	.w7(32'h3b3c7b15),
	.w8(32'hbab0d142),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39daee6c),
	.w1(32'h3c49903a),
	.w2(32'h3c3f1eae),
	.w3(32'h3a79f634),
	.w4(32'h3c31517e),
	.w5(32'h3c3234d1),
	.w6(32'h3bd1f687),
	.w7(32'hba68b162),
	.w8(32'h3a92fd8a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c194069),
	.w1(32'hbcc2c834),
	.w2(32'hbd13f2d7),
	.w3(32'h3ba34b12),
	.w4(32'hbb5b593c),
	.w5(32'hbc4d1ca0),
	.w6(32'hbc5bd810),
	.w7(32'hbcca52b6),
	.w8(32'hbcb39405),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdec622),
	.w1(32'h3c893ca9),
	.w2(32'h3c6f7e04),
	.w3(32'hbc5a7c1d),
	.w4(32'h3c8ec2b5),
	.w5(32'h3caf0110),
	.w6(32'h3c2bd75f),
	.w7(32'h3beede3b),
	.w8(32'h3c190e98),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7e9e),
	.w1(32'h39a8c953),
	.w2(32'hbb408c92),
	.w3(32'h3cb8aad3),
	.w4(32'hbba8eeb8),
	.w5(32'hbc1f2387),
	.w6(32'h3afc887b),
	.w7(32'h3ac07baf),
	.w8(32'h3aa38be0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baddf65),
	.w1(32'h3babdf7d),
	.w2(32'h3bb9e581),
	.w3(32'hbbeb0fb0),
	.w4(32'hbbbf2c3b),
	.w5(32'hbb65f0bf),
	.w6(32'hbab35868),
	.w7(32'h3af97236),
	.w8(32'h3c08b159),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3476eb),
	.w1(32'h3b2998ee),
	.w2(32'h3c0369dc),
	.w3(32'hbbd6977c),
	.w4(32'h39792bc3),
	.w5(32'h3be2263b),
	.w6(32'h3c6eaf2e),
	.w7(32'h3b000530),
	.w8(32'h3b876963),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a344e),
	.w1(32'h3b869ddb),
	.w2(32'h3b5a5050),
	.w3(32'h3bbea67e),
	.w4(32'hbbd4d7c1),
	.w5(32'hbc5eef33),
	.w6(32'h3c492773),
	.w7(32'h3bfd3836),
	.w8(32'h3b7b6d10),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93437b),
	.w1(32'hbc0fec9d),
	.w2(32'hbb931d56),
	.w3(32'hbc0894da),
	.w4(32'hbbab68fd),
	.w5(32'hbc29d9b8),
	.w6(32'hbb65d1d6),
	.w7(32'hbc2f2495),
	.w8(32'hbbb4c63a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eafb6),
	.w1(32'h39d85700),
	.w2(32'hbb01dd2a),
	.w3(32'h3bc7c63a),
	.w4(32'h3c85a17d),
	.w5(32'h3c7145d1),
	.w6(32'hbc04959f),
	.w7(32'hbc345a14),
	.w8(32'hbc2dd305),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba642e48),
	.w1(32'hbccd3ea5),
	.w2(32'hbd16efc9),
	.w3(32'h3c2f0932),
	.w4(32'hbc8f117d),
	.w5(32'hbcf6690b),
	.w6(32'hbcbb5772),
	.w7(32'hbccb3a41),
	.w8(32'hbc8ccead),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf06e6f),
	.w1(32'h3b067ce2),
	.w2(32'h3b8ecadf),
	.w3(32'hbce9f4bd),
	.w4(32'hbba9b1cd),
	.w5(32'hbbc31ced),
	.w6(32'h3b42ab72),
	.w7(32'h3b93b5c3),
	.w8(32'h3b6e5206),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8853fa),
	.w1(32'hbb099adc),
	.w2(32'h3ac7e828),
	.w3(32'hbb3799b1),
	.w4(32'h3bbda1bc),
	.w5(32'h3cb22929),
	.w6(32'h3c0795bc),
	.w7(32'h3b145337),
	.w8(32'hbc86d83d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853716f),
	.w1(32'hba762012),
	.w2(32'h3b1c3958),
	.w3(32'h3ce13ce2),
	.w4(32'h3bc897dc),
	.w5(32'h3a94bdd3),
	.w6(32'h3aa24aa8),
	.w7(32'hbba414ba),
	.w8(32'h388c323b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b46a5),
	.w1(32'hbafe3b9f),
	.w2(32'hbbca844b),
	.w3(32'h3af80b99),
	.w4(32'h3b9eb7c1),
	.w5(32'h3bbdc3ed),
	.w6(32'hbbee49be),
	.w7(32'hbc2ab1db),
	.w8(32'hbc251b2a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae48a),
	.w1(32'h3ba51b98),
	.w2(32'h3c1f8484),
	.w3(32'hbb058329),
	.w4(32'h3bc16f4c),
	.w5(32'h3c29a6f5),
	.w6(32'h3b9bfacc),
	.w7(32'h3c03e80d),
	.w8(32'h3c1e7c96),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0edfe4),
	.w1(32'hba06b98e),
	.w2(32'h3bbe293c),
	.w3(32'h3b16ba8b),
	.w4(32'hbaa42095),
	.w5(32'hba5419ce),
	.w6(32'hb98c8289),
	.w7(32'h3968c3cd),
	.w8(32'h3a165e6f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbbf9d),
	.w1(32'h3a91b18f),
	.w2(32'h3c118bd3),
	.w3(32'h3b8d124b),
	.w4(32'h3beeba9b),
	.w5(32'h3bf50bc4),
	.w6(32'hbbc374de),
	.w7(32'hbc11e200),
	.w8(32'hba84e3a7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8debf4),
	.w1(32'h3b48a3fa),
	.w2(32'hb9ca242a),
	.w3(32'hbb347e8a),
	.w4(32'hbb18d10c),
	.w5(32'hbb80aedc),
	.w6(32'hba0daf9e),
	.w7(32'hba67fec2),
	.w8(32'h3b8ba493),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f0a87),
	.w1(32'hbb1573d4),
	.w2(32'hba0b6f54),
	.w3(32'hba5e2411),
	.w4(32'hbb3a7ce9),
	.w5(32'hbb5a1f5e),
	.w6(32'hbb1a1f65),
	.w7(32'hbbe64481),
	.w8(32'hbb989efd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dc67c),
	.w1(32'hbb9a6de8),
	.w2(32'hbc2433dc),
	.w3(32'hbaaa1ab8),
	.w4(32'h3bbcbc96),
	.w5(32'h3bd065ad),
	.w6(32'hbc270c9e),
	.w7(32'hbc355d06),
	.w8(32'hbc44e2a1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39bcee),
	.w1(32'h3bc191b0),
	.w2(32'h3bfb8df4),
	.w3(32'hbbf6dfaf),
	.w4(32'hba8c796d),
	.w5(32'hba215668),
	.w6(32'h39d7a27e),
	.w7(32'hb91f502b),
	.w8(32'h3bce3f16),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ce442),
	.w1(32'hbad45b87),
	.w2(32'hbadb9445),
	.w3(32'hb9cc6b04),
	.w4(32'h3acd1ee3),
	.w5(32'h3b0bcb93),
	.w6(32'h38642008),
	.w7(32'hbb152c47),
	.w8(32'h3a380282),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6673de),
	.w1(32'hbc18af80),
	.w2(32'h3a373b9e),
	.w3(32'h3a47e543),
	.w4(32'h3a72de82),
	.w5(32'h3aad1be2),
	.w6(32'hbc38303f),
	.w7(32'hbbef3eb4),
	.w8(32'hbb400a07),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule