module layer_10_featuremap_510(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ce5e2),
	.w1(32'h3bf95c3f),
	.w2(32'hbbe63ff7),
	.w3(32'hbc642bad),
	.w4(32'hbabe9c9c),
	.w5(32'h3d158f2e),
	.w6(32'hbb8533e3),
	.w7(32'h39d37626),
	.w8(32'h3bd816f8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e428),
	.w1(32'h3c757701),
	.w2(32'hbcaef2ae),
	.w3(32'hba8b7d27),
	.w4(32'h3c0ab047),
	.w5(32'h3c2948f4),
	.w6(32'h3be30b70),
	.w7(32'h3c80514c),
	.w8(32'h3ca17a69),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f1299),
	.w1(32'h3badc475),
	.w2(32'hbc9034a7),
	.w3(32'hbc4a7f59),
	.w4(32'h3c3688b2),
	.w5(32'h3a2ca0d0),
	.w6(32'h395eb4c7),
	.w7(32'hbb957e20),
	.w8(32'h3b1033c8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a22ce),
	.w1(32'hbc2f60a5),
	.w2(32'h3ae5216f),
	.w3(32'h3af0fa09),
	.w4(32'hbc0254f7),
	.w5(32'hbbf63cce),
	.w6(32'h3bce6fe7),
	.w7(32'h3bb0033b),
	.w8(32'h3c02b27c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60a395),
	.w1(32'hbbcc366c),
	.w2(32'hbaff6159),
	.w3(32'hbc794af4),
	.w4(32'hbc9543e8),
	.w5(32'h3bc06eb1),
	.w6(32'h3c3a18fa),
	.w7(32'h3afa5749),
	.w8(32'hbbe92b39),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99f60f),
	.w1(32'hbc072321),
	.w2(32'h3c0d1842),
	.w3(32'h3b27ca52),
	.w4(32'hbc702593),
	.w5(32'h3cfd4033),
	.w6(32'h3c5117b0),
	.w7(32'h3bd27d8d),
	.w8(32'hbba480ef),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fec7d4),
	.w1(32'hbcef20bb),
	.w2(32'hbb8a08f9),
	.w3(32'h3be8b274),
	.w4(32'h3aad5937),
	.w5(32'hba80e40e),
	.w6(32'h3a626d9e),
	.w7(32'hbbf19fe0),
	.w8(32'hbc0c46eb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd1d14),
	.w1(32'h3c0403e6),
	.w2(32'h3c78b50a),
	.w3(32'hbc9c42ef),
	.w4(32'hbc9ff85a),
	.w5(32'hbb469df1),
	.w6(32'hbd291ad9),
	.w7(32'h3c0d3db2),
	.w8(32'hbc2862ed),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05973b),
	.w1(32'hbc426f36),
	.w2(32'h3bfd1383),
	.w3(32'h3cc3fb75),
	.w4(32'h3cb8c9d0),
	.w5(32'hbc0e5d4d),
	.w6(32'h3c4e8522),
	.w7(32'hbaefa5d9),
	.w8(32'hba25dbb7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8439e),
	.w1(32'hbc061071),
	.w2(32'hbc1450ee),
	.w3(32'hbb93a16b),
	.w4(32'h39b67197),
	.w5(32'hbbb3d966),
	.w6(32'hbc14a133),
	.w7(32'h3ae3aba3),
	.w8(32'h3ca3ba1f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6f4d),
	.w1(32'h3a619da9),
	.w2(32'hbb20df4c),
	.w3(32'h3c339d05),
	.w4(32'hbb836610),
	.w5(32'h3b28e3a6),
	.w6(32'hbb5f104a),
	.w7(32'h3b3f1909),
	.w8(32'h3aed4df3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc746279),
	.w1(32'h3c3e9896),
	.w2(32'hbc0cc46a),
	.w3(32'h3b80fbe8),
	.w4(32'hbb88819d),
	.w5(32'hbbb6e7f4),
	.w6(32'h3bd45d22),
	.w7(32'h3b6094b4),
	.w8(32'h3ba3e412),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4516),
	.w1(32'h3c53894d),
	.w2(32'hbc6df3e6),
	.w3(32'h3c161bb9),
	.w4(32'h3aa15df1),
	.w5(32'hbc8faa60),
	.w6(32'h3bb813da),
	.w7(32'hbb2b4512),
	.w8(32'hbcc6a466),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fde4a),
	.w1(32'hbb9579b9),
	.w2(32'h3aa70a5a),
	.w3(32'h3c1dd303),
	.w4(32'hbc13f649),
	.w5(32'h3a60f36d),
	.w6(32'hbb804477),
	.w7(32'hbc0c5a9a),
	.w8(32'hbab2bd34),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18bc7d),
	.w1(32'hbc88c121),
	.w2(32'h3b95fa11),
	.w3(32'hbc012e40),
	.w4(32'hb96dc95d),
	.w5(32'hbc622494),
	.w6(32'hbc34f8eb),
	.w7(32'h3c84111b),
	.w8(32'hbbb822fa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b65c0),
	.w1(32'h3c5fa4b6),
	.w2(32'hba99c031),
	.w3(32'hbc19b867),
	.w4(32'h3acf698f),
	.w5(32'h3b1a129b),
	.w6(32'h3afbc806),
	.w7(32'hbc0b65f5),
	.w8(32'hb87b8c79),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032f96),
	.w1(32'hbc15cb7e),
	.w2(32'hba9fef70),
	.w3(32'h3bdf95df),
	.w4(32'hb9edafa1),
	.w5(32'hba8e2a60),
	.w6(32'h3c4080e8),
	.w7(32'h3b970ab8),
	.w8(32'hbb16b4b4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d277c),
	.w1(32'hbd0941cb),
	.w2(32'hbc8360f5),
	.w3(32'hbbbd8aaf),
	.w4(32'hbd0428f9),
	.w5(32'hbc4c26ee),
	.w6(32'hbcb2c4f4),
	.w7(32'hbca92bb6),
	.w8(32'hbc949103),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c795f49),
	.w1(32'h3ae295fd),
	.w2(32'hbb1cc316),
	.w3(32'hbbef2276),
	.w4(32'hbbe3c04d),
	.w5(32'hbba5c1b9),
	.w6(32'hbb9f899a),
	.w7(32'hbbb3078b),
	.w8(32'hbace0c17),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb16c83),
	.w1(32'hbbffabf3),
	.w2(32'h3c093980),
	.w3(32'hbb52e9fc),
	.w4(32'h3aa6eba2),
	.w5(32'hbb840702),
	.w6(32'hbb1a5a1c),
	.w7(32'hbc1c7a40),
	.w8(32'hbc13ac4e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3f34),
	.w1(32'hb64d0472),
	.w2(32'h3ba00f40),
	.w3(32'hbc1153bb),
	.w4(32'hbbc4c6ba),
	.w5(32'hbd0e4c8a),
	.w6(32'h3c6e267a),
	.w7(32'hbbb36783),
	.w8(32'hbb7b4b95),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaa9ed),
	.w1(32'h3b05de13),
	.w2(32'hba0f10a7),
	.w3(32'h3c50c242),
	.w4(32'h3c07da38),
	.w5(32'h3ca4edbb),
	.w6(32'hbc4fa898),
	.w7(32'h3b4e1403),
	.w8(32'hbabbabd0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36d195),
	.w1(32'hbbe7081d),
	.w2(32'hbcc34176),
	.w3(32'hbb572b2f),
	.w4(32'hba90e7d2),
	.w5(32'hbcfec696),
	.w6(32'hbc897deb),
	.w7(32'hbd0dfa9b),
	.w8(32'hbc9782f8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc718372),
	.w1(32'h3bf83248),
	.w2(32'h3c31c255),
	.w3(32'h3b0d60ba),
	.w4(32'hbc9e82c6),
	.w5(32'h3d028f13),
	.w6(32'hbbc9c26e),
	.w7(32'hbc441eca),
	.w8(32'h3b3d284f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a9c43),
	.w1(32'h3b031128),
	.w2(32'h3ce3f82b),
	.w3(32'h3c85807b),
	.w4(32'hbabc20cf),
	.w5(32'h3c4472de),
	.w6(32'h3baf340b),
	.w7(32'h3c1751dd),
	.w8(32'hba706431),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c418b3b),
	.w1(32'h3a3e3b62),
	.w2(32'h3d339259),
	.w3(32'hbbb3618a),
	.w4(32'h3c173589),
	.w5(32'hbaafed4c),
	.w6(32'hbb39f856),
	.w7(32'hba2f2692),
	.w8(32'h3a690008),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa688e),
	.w1(32'hbcb37935),
	.w2(32'h3b0ac416),
	.w3(32'hbb8276ff),
	.w4(32'h3be9c577),
	.w5(32'h3b971009),
	.w6(32'h3bbb4937),
	.w7(32'h3c3510f8),
	.w8(32'hbc5f12f2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45e505),
	.w1(32'hbbe41d18),
	.w2(32'hbc177ef8),
	.w3(32'h3bd0dd51),
	.w4(32'hbd57213a),
	.w5(32'h3aec9fdf),
	.w6(32'h3c57562f),
	.w7(32'h3aee437c),
	.w8(32'h3cb2076d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f06f),
	.w1(32'hbab71cb2),
	.w2(32'h3bc36cca),
	.w3(32'hbb40e154),
	.w4(32'hbc179883),
	.w5(32'hbd4d0e20),
	.w6(32'h3b49a3ca),
	.w7(32'hbb513b41),
	.w8(32'hbc44b9e7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe28859),
	.w1(32'h3cc97d63),
	.w2(32'h3c5e9b52),
	.w3(32'h3be42fcc),
	.w4(32'h3bfffb94),
	.w5(32'h3c8c8709),
	.w6(32'h3cfa4565),
	.w7(32'h3a6b2dcf),
	.w8(32'h3cf7a7d5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c625357),
	.w1(32'h39c5b11e),
	.w2(32'h3c6f95e0),
	.w3(32'h3aeb8ff2),
	.w4(32'hbc0da92e),
	.w5(32'h3be53c5a),
	.w6(32'hbbcc04d0),
	.w7(32'h3b495058),
	.w8(32'h3c11f0d4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953af3f),
	.w1(32'hbc0c01f0),
	.w2(32'hbb9b9228),
	.w3(32'hbc12ce25),
	.w4(32'h3ac28545),
	.w5(32'hbc24c2b0),
	.w6(32'h3d8a0cd3),
	.w7(32'hbb266819),
	.w8(32'hbbb7beeb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d4c8e),
	.w1(32'hbc11ce27),
	.w2(32'h3bfa09ac),
	.w3(32'h39654cdc),
	.w4(32'h3c861ebf),
	.w5(32'h3a29cf52),
	.w6(32'hbc3cb4da),
	.w7(32'hbbe92637),
	.w8(32'hbb26ad72),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee29e7),
	.w1(32'hb9c3f98d),
	.w2(32'h3b12d35e),
	.w3(32'hbc0bf81e),
	.w4(32'hbc74b0bd),
	.w5(32'hbc310f44),
	.w6(32'h3b0c692e),
	.w7(32'hbc258abb),
	.w8(32'h391a1f49),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010aff),
	.w1(32'hbb776600),
	.w2(32'hbc1f2441),
	.w3(32'h3c14a0d9),
	.w4(32'hbba49346),
	.w5(32'hb7fab7af),
	.w6(32'hbb3b8558),
	.w7(32'h3b487984),
	.w8(32'h3babdfa6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30d574),
	.w1(32'h3ba9fa71),
	.w2(32'hbbf05cfd),
	.w3(32'h39494e5e),
	.w4(32'hbb4ec772),
	.w5(32'hbab56e21),
	.w6(32'h3a1fd47e),
	.w7(32'hba69cc5c),
	.w8(32'hbb5c57d2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa5c7),
	.w1(32'h3cb49ba6),
	.w2(32'h3a9500e7),
	.w3(32'h3bd86568),
	.w4(32'h3c1fdf3f),
	.w5(32'hb9c85efc),
	.w6(32'h3b14fd99),
	.w7(32'hbac2c893),
	.w8(32'hbc69c1d3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc380cde),
	.w1(32'h3ccf13ce),
	.w2(32'h3cc86ca5),
	.w3(32'hbae8125d),
	.w4(32'h3c763e13),
	.w5(32'h3c9b679f),
	.w6(32'h3c97b5e0),
	.w7(32'h3ccf0b9c),
	.w8(32'h3cb1219e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd002a1),
	.w1(32'hbc56bb05),
	.w2(32'h3cc0a748),
	.w3(32'h3bc209d0),
	.w4(32'h3aa09269),
	.w5(32'h3c3fdaca),
	.w6(32'h3c936702),
	.w7(32'h3ccb42a2),
	.w8(32'h3c811bd5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0627c),
	.w1(32'h3bdbd3e9),
	.w2(32'h3c220ec6),
	.w3(32'hbc2a5c2e),
	.w4(32'h3abd5dfa),
	.w5(32'h3b834c59),
	.w6(32'h3ba9a17b),
	.w7(32'h3c726d5b),
	.w8(32'h3c510669),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e0efc),
	.w1(32'h3b501fe6),
	.w2(32'hb9a6fca4),
	.w3(32'hbc057226),
	.w4(32'h3c27b72e),
	.w5(32'h3cb12b2c),
	.w6(32'h3b785283),
	.w7(32'h3c387e78),
	.w8(32'h3c2d562c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0325),
	.w1(32'h3c1ba9dd),
	.w2(32'h3c19ccb2),
	.w3(32'hbc507f9c),
	.w4(32'h3a635f61),
	.w5(32'h3c04d9e3),
	.w6(32'h3a5dc10d),
	.w7(32'hbc02b1c0),
	.w8(32'h3a964537),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fbd34),
	.w1(32'h39ed761d),
	.w2(32'hbae90f34),
	.w3(32'hbc609fc9),
	.w4(32'hba436457),
	.w5(32'h3c855358),
	.w6(32'hbc57fa94),
	.w7(32'h3b53fad1),
	.w8(32'h3b67c2ff),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0edbaf),
	.w1(32'hbbf16fe2),
	.w2(32'hbbc79992),
	.w3(32'h3c38e8e9),
	.w4(32'hbba75fdb),
	.w5(32'h3a234ea2),
	.w6(32'h3cb96bb7),
	.w7(32'hbc28ae0a),
	.w8(32'h3b98939c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b8fe9),
	.w1(32'hba02087c),
	.w2(32'hbb86852f),
	.w3(32'hbbf21d8a),
	.w4(32'h3b5079d1),
	.w5(32'h3c509cb0),
	.w6(32'h3b6b18a9),
	.w7(32'h3c25c970),
	.w8(32'h3c034b79),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7066e),
	.w1(32'hbbb9598b),
	.w2(32'h3a1220b2),
	.w3(32'hbb36570a),
	.w4(32'h3c55bbe6),
	.w5(32'h3c236b6f),
	.w6(32'hbc285cd6),
	.w7(32'h3c10d61c),
	.w8(32'h3be279f0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6473e),
	.w1(32'hbc4bb5be),
	.w2(32'h3bf28c05),
	.w3(32'hbc1d5f46),
	.w4(32'h3b9cf6a8),
	.w5(32'h3bcece86),
	.w6(32'hbb50645d),
	.w7(32'h3bd926b7),
	.w8(32'hbc4326a7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b7d0a),
	.w1(32'hbcb12eec),
	.w2(32'hbd19c522),
	.w3(32'hbc836c0d),
	.w4(32'hbc9e8d4b),
	.w5(32'hbcb88186),
	.w6(32'hbcbfa28b),
	.w7(32'hbcc84140),
	.w8(32'hbcc30a74),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dedc8),
	.w1(32'hbc1af9bf),
	.w2(32'h3b919edc),
	.w3(32'h3c8bfdcb),
	.w4(32'hbd1878f3),
	.w5(32'hbbce7b3b),
	.w6(32'hbc16d5cd),
	.w7(32'hbc18da47),
	.w8(32'h3bd16456),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0a999),
	.w1(32'hbad24399),
	.w2(32'hbb63072d),
	.w3(32'hbb0491a1),
	.w4(32'hbb8e4a71),
	.w5(32'hbadb661c),
	.w6(32'hbbf4ca5f),
	.w7(32'h3bfd811a),
	.w8(32'h3c9af362),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3a8c),
	.w1(32'h3bbf7c1d),
	.w2(32'h3bcd1791),
	.w3(32'h3b51d605),
	.w4(32'h3c00eb7d),
	.w5(32'hbab100b6),
	.w6(32'hbc3a7ceb),
	.w7(32'h3ab07c31),
	.w8(32'hbbb05c57),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe614bd),
	.w1(32'h3bc8470a),
	.w2(32'h3c51fd3e),
	.w3(32'hbc31fab3),
	.w4(32'h3be39e30),
	.w5(32'h3beceac1),
	.w6(32'hbae5c019),
	.w7(32'h3c2a2edd),
	.w8(32'hbc90fca7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29272a),
	.w1(32'hbc9e8329),
	.w2(32'hbbd15548),
	.w3(32'h3b97b222),
	.w4(32'hbc1e3ddb),
	.w5(32'h3b974fb1),
	.w6(32'hbd02ba6f),
	.w7(32'hbc8ab705),
	.w8(32'h3902887f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b961b20),
	.w1(32'hbc8afa4d),
	.w2(32'hbc28867d),
	.w3(32'h3b97d56e),
	.w4(32'hbc18e3d8),
	.w5(32'hbc920913),
	.w6(32'hbc71322d),
	.w7(32'hbb033820),
	.w8(32'hbc91e18e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d4755),
	.w1(32'hbcb3410f),
	.w2(32'hbb7134af),
	.w3(32'h3a13ce24),
	.w4(32'hbcb3072f),
	.w5(32'hbb2733ad),
	.w6(32'hbd04c057),
	.w7(32'h3c79f8c0),
	.w8(32'h3d35a072),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11cf4a),
	.w1(32'hbc93798a),
	.w2(32'h383742ba),
	.w3(32'hbbf0db34),
	.w4(32'h3d262657),
	.w5(32'h3bc9e0ba),
	.w6(32'hbc007f73),
	.w7(32'hbac2ef17),
	.w8(32'h3d43f415),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c433),
	.w1(32'h3cb38101),
	.w2(32'hbbc172e8),
	.w3(32'hbb4fd78a),
	.w4(32'h3d0588f8),
	.w5(32'h3b40fb50),
	.w6(32'h3a4c5ab4),
	.w7(32'h39e679cb),
	.w8(32'hbca686e9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12e884),
	.w1(32'h3b5a63dc),
	.w2(32'h3bbf6d74),
	.w3(32'hba12741c),
	.w4(32'hbc27e318),
	.w5(32'hbb894392),
	.w6(32'hbd10a630),
	.w7(32'hbb3ee8f9),
	.w8(32'hbb805d06),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf9da88),
	.w1(32'hbba40278),
	.w2(32'h3c9d2e05),
	.w3(32'hbb68f809),
	.w4(32'hba5c1784),
	.w5(32'hbb019511),
	.w6(32'hbad30d80),
	.w7(32'hbc314d2c),
	.w8(32'hbbe80a93),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109e97),
	.w1(32'hbc2e0e30),
	.w2(32'h3d0190dc),
	.w3(32'h3c1ee474),
	.w4(32'hbc03b1a6),
	.w5(32'h3b112c96),
	.w6(32'hbb13f0e0),
	.w7(32'hbc834d5e),
	.w8(32'hbce53518),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bae02),
	.w1(32'hbca84928),
	.w2(32'hbb460045),
	.w3(32'hbc94b65c),
	.w4(32'h3a0dc5c9),
	.w5(32'hbc58570f),
	.w6(32'hbb90880f),
	.w7(32'hbc56dd7a),
	.w8(32'h3b54ec5d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a85a5),
	.w1(32'hbbe07d90),
	.w2(32'hbbb9d08b),
	.w3(32'hbc2ac772),
	.w4(32'hbc10e00d),
	.w5(32'hbaa20103),
	.w6(32'hbc0fe444),
	.w7(32'hbc834bfe),
	.w8(32'h3a297ade),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd21ed09),
	.w1(32'hb8ac7996),
	.w2(32'hbc44999a),
	.w3(32'hb98a312b),
	.w4(32'hbaf98092),
	.w5(32'hbc6a58fb),
	.w6(32'hbb625c0f),
	.w7(32'h3cb7b619),
	.w8(32'hbaed654b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a3a9a),
	.w1(32'hbb16ffe3),
	.w2(32'h3bb1891e),
	.w3(32'h3a9b8e75),
	.w4(32'hbd246314),
	.w5(32'h394b2168),
	.w6(32'h3c1d0da6),
	.w7(32'h3aaf4349),
	.w8(32'hbb0ebcfe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d1b0f),
	.w1(32'hbca6048c),
	.w2(32'hbb904dd8),
	.w3(32'h3c44edee),
	.w4(32'hbc0808eb),
	.w5(32'hbcd0b11b),
	.w6(32'hba8bce3f),
	.w7(32'h3ab42115),
	.w8(32'hbba3ad12),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb2fd6),
	.w1(32'hbc8448cd),
	.w2(32'hbbc57d50),
	.w3(32'hbc25f286),
	.w4(32'hbbb74ced),
	.w5(32'h3b6f0aa2),
	.w6(32'hbc06a9d8),
	.w7(32'h3aa0762b),
	.w8(32'h3bac049a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93bc4),
	.w1(32'hbbde9728),
	.w2(32'hbc1e91ab),
	.w3(32'h3bb6d453),
	.w4(32'hb9d59927),
	.w5(32'hbbf4731d),
	.w6(32'h3ba6a9b7),
	.w7(32'hbc5485ba),
	.w8(32'hbc956e3b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e6294),
	.w1(32'hbbd776c3),
	.w2(32'h3c307079),
	.w3(32'hba09cffc),
	.w4(32'hbc1bde56),
	.w5(32'h3b321b83),
	.w6(32'hbbc018cd),
	.w7(32'hbc740561),
	.w8(32'h3c129fc8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1006e9),
	.w1(32'hbc02ad1e),
	.w2(32'hbc3a3f5a),
	.w3(32'hbcaf40dc),
	.w4(32'hbbddf96c),
	.w5(32'hbcef9cba),
	.w6(32'h3b9fbb2e),
	.w7(32'hbc8f31f1),
	.w8(32'hbbde6bcc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca790ff),
	.w1(32'h3cd0b3ea),
	.w2(32'h3bb919fa),
	.w3(32'hbbd94eda),
	.w4(32'hbbc976f3),
	.w5(32'h3c2aed86),
	.w6(32'h3cb34180),
	.w7(32'h3cbd7b5e),
	.w8(32'h3cd1392a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd694),
	.w1(32'hbb1e23f4),
	.w2(32'hbb843011),
	.w3(32'hba9574e7),
	.w4(32'hbaa4896f),
	.w5(32'h3b78529e),
	.w6(32'h3b32fe3f),
	.w7(32'hbc6a4caf),
	.w8(32'hbb964b51),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69ee47),
	.w1(32'h3b42812c),
	.w2(32'h3ce6c2cc),
	.w3(32'h3c7019b3),
	.w4(32'h3c3f98c4),
	.w5(32'hbbbf113d),
	.w6(32'hba76fe36),
	.w7(32'hbc0be3a6),
	.w8(32'hbc0f2770),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524b1b),
	.w1(32'h3d01f395),
	.w2(32'hbbac9e22),
	.w3(32'hbc7789c5),
	.w4(32'hbc330db9),
	.w5(32'h3b0637a4),
	.w6(32'h3c784677),
	.w7(32'hbc54dcdd),
	.w8(32'hbca6e462),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bc9b1),
	.w1(32'hbabc55e3),
	.w2(32'hbc83e5e7),
	.w3(32'h3bf75a3f),
	.w4(32'hbb96dbf2),
	.w5(32'hbc22f833),
	.w6(32'hbbcfed83),
	.w7(32'h3a2b0bc0),
	.w8(32'h3bda4a8a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63de07),
	.w1(32'hbbfe7602),
	.w2(32'h3c97e9c6),
	.w3(32'hbc2de975),
	.w4(32'h3b2e1106),
	.w5(32'hbc68ad17),
	.w6(32'hba32a69b),
	.w7(32'h3b8a0915),
	.w8(32'hbb5a651d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc2c42),
	.w1(32'hbc940970),
	.w2(32'hbcd05e54),
	.w3(32'hba335257),
	.w4(32'hbc8c993f),
	.w5(32'hbc275de1),
	.w6(32'hbc7717dd),
	.w7(32'hbc773931),
	.w8(32'hbc999746),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9be640),
	.w1(32'hbb80e9f4),
	.w2(32'h3973cef7),
	.w3(32'hbb7d2b8f),
	.w4(32'hbc989891),
	.w5(32'hbcd27732),
	.w6(32'hbbf8d565),
	.w7(32'hbba6d4e7),
	.w8(32'hbd35cb24),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5f68),
	.w1(32'h3b53d274),
	.w2(32'h3c02d8c5),
	.w3(32'h3c040464),
	.w4(32'h3c7e502b),
	.w5(32'hba1b4c80),
	.w6(32'hbbfa228e),
	.w7(32'hbb931ecf),
	.w8(32'h3b42d876),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68b42a),
	.w1(32'h3c0eca84),
	.w2(32'hbbb56cc6),
	.w3(32'hbc072dbe),
	.w4(32'h3b1c76ac),
	.w5(32'hbb27f2d9),
	.w6(32'hbbc6605a),
	.w7(32'h3cb7dc28),
	.w8(32'h3c15d385),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb180e5a),
	.w1(32'hbbe005b6),
	.w2(32'hbc275f2e),
	.w3(32'hba7cc2d4),
	.w4(32'hbc89bea0),
	.w5(32'h3c08f7b7),
	.w6(32'h3a03430e),
	.w7(32'hbb8abb2f),
	.w8(32'h3c252886),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6e662),
	.w1(32'hbc27fa10),
	.w2(32'hbafd86f4),
	.w3(32'h3cb38451),
	.w4(32'hbac60e6f),
	.w5(32'h3c83e786),
	.w6(32'h3c9956af),
	.w7(32'h3c52b636),
	.w8(32'h3c282211),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f37e1),
	.w1(32'hbc3bcce8),
	.w2(32'hbc50555b),
	.w3(32'hbb1a8a5c),
	.w4(32'hbb3c6321),
	.w5(32'hbc388c35),
	.w6(32'hbb099451),
	.w7(32'hbb871f5b),
	.w8(32'hbcd470e9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79ebbd),
	.w1(32'h3c26a65d),
	.w2(32'hbbe2625f),
	.w3(32'h3b9af41d),
	.w4(32'hbc01bc1b),
	.w5(32'h3cb4cfb7),
	.w6(32'h3c38a911),
	.w7(32'hbc5ceafa),
	.w8(32'hbd92bd79),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0a0fd),
	.w1(32'h3c99b92c),
	.w2(32'h3b41b331),
	.w3(32'h3d042c19),
	.w4(32'hbbda9652),
	.w5(32'h3bdd5d70),
	.w6(32'hbbea6f2a),
	.w7(32'h3b4fa91b),
	.w8(32'hbaebb65d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d1476),
	.w1(32'hbbf3016a),
	.w2(32'h3c17e839),
	.w3(32'hbba3be9e),
	.w4(32'hbb34ed6e),
	.w5(32'hb9bfbd78),
	.w6(32'h3c262943),
	.w7(32'hbb2b06a7),
	.w8(32'h3c015bd3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20a45b),
	.w1(32'h3afd32dc),
	.w2(32'h3ca14fe6),
	.w3(32'hbc2fd530),
	.w4(32'h3c5c2728),
	.w5(32'hbc61960c),
	.w6(32'h3d07882e),
	.w7(32'h3bbed122),
	.w8(32'h3ae2e5bf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c711663),
	.w1(32'h39fb4e0b),
	.w2(32'hb9bb326f),
	.w3(32'h3c32ac8e),
	.w4(32'h3bc51225),
	.w5(32'h3cb0781f),
	.w6(32'h3cf18ca7),
	.w7(32'hbbf5f0b6),
	.w8(32'hbca512e4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5ffb6),
	.w1(32'hb9e71ca6),
	.w2(32'hbc38273e),
	.w3(32'h3cc03e9c),
	.w4(32'h3d0bfafd),
	.w5(32'h3b9ee811),
	.w6(32'hbc31e225),
	.w7(32'hbbd4333b),
	.w8(32'hbc5b4dd8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf10bb),
	.w1(32'hbb98009c),
	.w2(32'hbb7325c5),
	.w3(32'hbc47530b),
	.w4(32'h3c907345),
	.w5(32'hbad432c8),
	.w6(32'hbc2adbe3),
	.w7(32'hba54deff),
	.w8(32'hbc8bebc7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14c14b),
	.w1(32'hbbe5206f),
	.w2(32'hbcc1665f),
	.w3(32'hbd1aa101),
	.w4(32'hbc5e0ed6),
	.w5(32'hbd15d6e1),
	.w6(32'hbcea29a0),
	.w7(32'hbc7dde4a),
	.w8(32'hbc610a9f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cdf9e),
	.w1(32'h3cba6edf),
	.w2(32'h3d3cc8e3),
	.w3(32'h3b037942),
	.w4(32'hbb4a9173),
	.w5(32'hbbbaca2d),
	.w6(32'hbb8497a0),
	.w7(32'h3c46305a),
	.w8(32'h3bf78ffe),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e573f),
	.w1(32'hbaac9714),
	.w2(32'hbb9a5839),
	.w3(32'h3b4c6f43),
	.w4(32'hbc728bd0),
	.w5(32'hba253115),
	.w6(32'hbbf98157),
	.w7(32'hbceb647c),
	.w8(32'hbc96446e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeee19),
	.w1(32'h3b15f29f),
	.w2(32'h3cca2da9),
	.w3(32'h3c41aa81),
	.w4(32'h3b9b7985),
	.w5(32'h3c9d8d15),
	.w6(32'h3bd86a13),
	.w7(32'hbc8f524c),
	.w8(32'h3c3101b0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d8053),
	.w1(32'h3b78417a),
	.w2(32'hbba353ed),
	.w3(32'hbbe4dfef),
	.w4(32'hbc2339c4),
	.w5(32'h3bd58fd4),
	.w6(32'h3a4cdba3),
	.w7(32'hbba03d6f),
	.w8(32'h3c72f2e8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09fc2a),
	.w1(32'hbb8a9412),
	.w2(32'hbc0ce9cc),
	.w3(32'hbc39db90),
	.w4(32'hba08ca93),
	.w5(32'h3c0a28f8),
	.w6(32'hbbaee52d),
	.w7(32'hbbb84397),
	.w8(32'hbbd68b6b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f414),
	.w1(32'hbc4204c7),
	.w2(32'h3aca55aa),
	.w3(32'hbc2617ad),
	.w4(32'h3bf41334),
	.w5(32'h3c39a87f),
	.w6(32'h39f17c50),
	.w7(32'hbaddb10f),
	.w8(32'hbc44868e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c2c16),
	.w1(32'hbb2be7a1),
	.w2(32'h3c8195ca),
	.w3(32'h3b2885e9),
	.w4(32'h3c319f48),
	.w5(32'hba985d10),
	.w6(32'hbbe08d56),
	.w7(32'h3b21136d),
	.w8(32'h3b04f65c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4131f9),
	.w1(32'h3c8e575f),
	.w2(32'hbb0100b6),
	.w3(32'h3b30fd25),
	.w4(32'h3c3f0722),
	.w5(32'h3b4fd670),
	.w6(32'hbca7a30e),
	.w7(32'h3a6ec181),
	.w8(32'hbc6f6ea8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fd71),
	.w1(32'h3b37a5be),
	.w2(32'hbbbd282f),
	.w3(32'hbb6e04a8),
	.w4(32'h3cd2e3d3),
	.w5(32'h3c4a8456),
	.w6(32'hba012eb3),
	.w7(32'h3b3773e7),
	.w8(32'hbbebdb9f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc219485),
	.w1(32'h3a9cf30c),
	.w2(32'hbb750fae),
	.w3(32'hbbc34183),
	.w4(32'h3bb54968),
	.w5(32'hbc3444f4),
	.w6(32'hbcbfafc3),
	.w7(32'hbc927a67),
	.w8(32'hbb3e9187),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc910258),
	.w1(32'h3a714203),
	.w2(32'h3c179c26),
	.w3(32'hbc38df85),
	.w4(32'h3c746b07),
	.w5(32'h3c931e3d),
	.w6(32'hba9879a4),
	.w7(32'h3b26c3ae),
	.w8(32'h3c87dc6e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bc57d),
	.w1(32'hba409bca),
	.w2(32'h3ca119d0),
	.w3(32'hbc86104e),
	.w4(32'h3d2fd464),
	.w5(32'h3c74bda0),
	.w6(32'hb8a28f69),
	.w7(32'hba6d68b3),
	.w8(32'h39070755),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960dcc2),
	.w1(32'h3a90b52f),
	.w2(32'hbc3c81ac),
	.w3(32'hbb2cc901),
	.w4(32'h3c036527),
	.w5(32'hbc987895),
	.w6(32'h3ad649cb),
	.w7(32'h3c763293),
	.w8(32'hbc60291b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf3d92),
	.w1(32'h3c805d17),
	.w2(32'hb99784a5),
	.w3(32'h3c1328b1),
	.w4(32'hbbfc9f41),
	.w5(32'hbc50d207),
	.w6(32'hbc9f4a6d),
	.w7(32'hbbdfbc7a),
	.w8(32'h3bd0352f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88cf60),
	.w1(32'hbc49301d),
	.w2(32'hbcc398a3),
	.w3(32'hbc6c6690),
	.w4(32'hbbe29831),
	.w5(32'hbd03f8df),
	.w6(32'hbad4ceda),
	.w7(32'hbc3703e2),
	.w8(32'hbbbf76e2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9848868),
	.w1(32'h3c731335),
	.w2(32'hbc1c6a6e),
	.w3(32'h3bb18e79),
	.w4(32'h3b3c9a6a),
	.w5(32'hba9cecee),
	.w6(32'h3ca5b8b1),
	.w7(32'h3bb269dd),
	.w8(32'hbc54fff9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ffe07),
	.w1(32'hbba21ee2),
	.w2(32'hbbdd88e1),
	.w3(32'h3bf77795),
	.w4(32'h3c27a1b9),
	.w5(32'hba95fdfa),
	.w6(32'h3cfbd71c),
	.w7(32'hbb38d196),
	.w8(32'h3b92c75f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bc3c1),
	.w1(32'h3a81d820),
	.w2(32'hbb930502),
	.w3(32'hbc8f40d1),
	.w4(32'hbc0c0472),
	.w5(32'h3c082edc),
	.w6(32'hbb0a80be),
	.w7(32'h3c45bc9f),
	.w8(32'hbb8f1fe7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c8c0f),
	.w1(32'hbb2cba20),
	.w2(32'h3cf14a36),
	.w3(32'h3c18de92),
	.w4(32'hbbbe8952),
	.w5(32'h3c877d94),
	.w6(32'h3c66808d),
	.w7(32'h3b88118b),
	.w8(32'h3c0a820d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d2427),
	.w1(32'hbc1bf52d),
	.w2(32'h3c0998b6),
	.w3(32'h3be14a28),
	.w4(32'hbb8b3d95),
	.w5(32'h3bfa73c5),
	.w6(32'h3bdbd31c),
	.w7(32'h3c554880),
	.w8(32'h3c0be372),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e58ff),
	.w1(32'h3b02981d),
	.w2(32'hbc90b47b),
	.w3(32'hbaa5859a),
	.w4(32'hbab2384d),
	.w5(32'hbc39f521),
	.w6(32'h3bb40433),
	.w7(32'hbbec2a3f),
	.w8(32'hbbffe7b4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbe543),
	.w1(32'hbc0cb784),
	.w2(32'h3ca73735),
	.w3(32'h3c95048f),
	.w4(32'hbbb28a3e),
	.w5(32'hba90f362),
	.w6(32'h3a6d367e),
	.w7(32'h3c474f52),
	.w8(32'h3c5addc0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd398564),
	.w1(32'h3c2cdec3),
	.w2(32'h3b9edaf0),
	.w3(32'h3b8c5d67),
	.w4(32'hbb863935),
	.w5(32'h3bb7ae67),
	.w6(32'h3bde4995),
	.w7(32'hbab35bee),
	.w8(32'hbb2e83ca),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3e355),
	.w1(32'hbbe9e171),
	.w2(32'hbc190937),
	.w3(32'hbb620ab8),
	.w4(32'hbb553f55),
	.w5(32'hba358c61),
	.w6(32'hbb88fd4f),
	.w7(32'hb89b6f2a),
	.w8(32'h3a8e7b85),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dfa88),
	.w1(32'h3cd3f0da),
	.w2(32'h3c29220c),
	.w3(32'hbbc79c87),
	.w4(32'h3d02b499),
	.w5(32'h3b69066a),
	.w6(32'hbb439cda),
	.w7(32'h3a638de5),
	.w8(32'hbcf3e609),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcef5f6),
	.w1(32'h3b8f0830),
	.w2(32'h3c253d30),
	.w3(32'h3b5b7287),
	.w4(32'hba0f138a),
	.w5(32'hbc2d689b),
	.w6(32'hbc10db58),
	.w7(32'h3c2cb550),
	.w8(32'hbb7e20ad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe20645),
	.w1(32'h3c6c089e),
	.w2(32'h39149152),
	.w3(32'h3c1d5d4d),
	.w4(32'h3b0c5b9e),
	.w5(32'hbad90d96),
	.w6(32'hbaf5f7ef),
	.w7(32'h3cda4eca),
	.w8(32'h3b39505e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4bf3),
	.w1(32'h3c4a654c),
	.w2(32'hbb5850be),
	.w3(32'hbc08466d),
	.w4(32'h3aeb61fd),
	.w5(32'h3cb2346b),
	.w6(32'h3c80030a),
	.w7(32'h3bf03026),
	.w8(32'h3b8e366c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67f031),
	.w1(32'hba4d168f),
	.w2(32'hbaa82ed8),
	.w3(32'hbbbb7cda),
	.w4(32'h3c37e7a7),
	.w5(32'hbadbeb55),
	.w6(32'hb79cb3b6),
	.w7(32'hba4684bc),
	.w8(32'h397be552),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c350f67),
	.w1(32'h3be560ac),
	.w2(32'h3c4838fb),
	.w3(32'h3b79787c),
	.w4(32'hbb082742),
	.w5(32'hbbd89201),
	.w6(32'hbb047209),
	.w7(32'h3cc484ae),
	.w8(32'h3c111fdd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab20b1b),
	.w1(32'hbbbd3a7a),
	.w2(32'hbc28b9bf),
	.w3(32'hbc4f8596),
	.w4(32'h3ba72600),
	.w5(32'h3bdba049),
	.w6(32'h3ba6d6c6),
	.w7(32'h3904b765),
	.w8(32'hbc9b0305),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bd726),
	.w1(32'hbc927305),
	.w2(32'hbbf6a227),
	.w3(32'h3b6c453b),
	.w4(32'hbc25f9c2),
	.w5(32'hbbe57795),
	.w6(32'hbadf8fbf),
	.w7(32'hbbbf35ff),
	.w8(32'h3a441cb3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecff90),
	.w1(32'h3c044608),
	.w2(32'h3ac37bca),
	.w3(32'h3bda35c0),
	.w4(32'h3b1122b8),
	.w5(32'h3bc550a8),
	.w6(32'h3c7ce8b7),
	.w7(32'h3c6a0353),
	.w8(32'hbc8b643a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f0a8),
	.w1(32'h3b7b61fb),
	.w2(32'hbb4d5764),
	.w3(32'hbabba4a5),
	.w4(32'hbc108326),
	.w5(32'hbc874bed),
	.w6(32'h3af5fa53),
	.w7(32'hbc9f0ad2),
	.w8(32'h3c3da24d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babcd90),
	.w1(32'hbb8a28c0),
	.w2(32'h3a46fa83),
	.w3(32'h3bd0e542),
	.w4(32'h3b5c3d74),
	.w5(32'hbba8780e),
	.w6(32'hbb72c2df),
	.w7(32'h3b2dc25f),
	.w8(32'hbb4ac768),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc498158),
	.w1(32'hb8e51be1),
	.w2(32'h3cb05e97),
	.w3(32'hbb4798a0),
	.w4(32'h3b8c6236),
	.w5(32'hbbc7a363),
	.w6(32'h3b6ca507),
	.w7(32'h3b0a9649),
	.w8(32'hbb4859e1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b166),
	.w1(32'hbc9f3c31),
	.w2(32'hbbc091cd),
	.w3(32'h3c320a71),
	.w4(32'hbc51cb30),
	.w5(32'h3c36e389),
	.w6(32'hbc033c47),
	.w7(32'h3b9182f2),
	.w8(32'h3b572ed6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfdeef),
	.w1(32'h3b915d76),
	.w2(32'h3b8e3cb2),
	.w3(32'h3c806c49),
	.w4(32'hba14e717),
	.w5(32'hbbdeb341),
	.w6(32'hb95ca178),
	.w7(32'hbc8290bd),
	.w8(32'hbc0c313f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d6997),
	.w1(32'h3c8d6b0d),
	.w2(32'h3c8b132f),
	.w3(32'h3c0d4d62),
	.w4(32'hbc50da2e),
	.w5(32'h3c23c309),
	.w6(32'hbc1435b7),
	.w7(32'h3c01e174),
	.w8(32'h3b6a092a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4e2c),
	.w1(32'hbc40702b),
	.w2(32'hbba691b1),
	.w3(32'hbb974b77),
	.w4(32'hba9fc2f8),
	.w5(32'h3b129b18),
	.w6(32'h3aea181b),
	.w7(32'h3c0b9cd5),
	.w8(32'hbc0190c7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2992db),
	.w1(32'h3af154cd),
	.w2(32'h3c0ad81a),
	.w3(32'hba80f314),
	.w4(32'hbc33c533),
	.w5(32'hbb788abb),
	.w6(32'hbb5ed72c),
	.w7(32'h3c2d2175),
	.w8(32'h3caec338),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4acf38),
	.w1(32'h3ba74d74),
	.w2(32'h3c0e4c19),
	.w3(32'hbbb1a1c0),
	.w4(32'h3b70102e),
	.w5(32'h3c47208c),
	.w6(32'hbbfb4aca),
	.w7(32'h3b8a2257),
	.w8(32'hb8538634),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cb943),
	.w1(32'h3c9204f2),
	.w2(32'hbb0b590b),
	.w3(32'h3be87178),
	.w4(32'hba01b61f),
	.w5(32'h3a290b4c),
	.w6(32'h3c461b63),
	.w7(32'hbcfb6674),
	.w8(32'hbc1545b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd9b29),
	.w1(32'hb9489700),
	.w2(32'h393949ed),
	.w3(32'h3d00462f),
	.w4(32'h3c80a604),
	.w5(32'h3c581c29),
	.w6(32'h3bf785e8),
	.w7(32'hbc24e009),
	.w8(32'h3c8d1ca0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336930),
	.w1(32'hbc1d281f),
	.w2(32'hbcc94d7c),
	.w3(32'h3b918231),
	.w4(32'hbc67500e),
	.w5(32'hbbcd8147),
	.w6(32'hbc221906),
	.w7(32'hbc15ea83),
	.w8(32'hbbafd701),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051263),
	.w1(32'h3bc9e37c),
	.w2(32'hbbbb187d),
	.w3(32'hb8eeaa54),
	.w4(32'h3c12def9),
	.w5(32'hbc697e20),
	.w6(32'hbb166749),
	.w7(32'h3c03052a),
	.w8(32'h3c396cc3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add78cd),
	.w1(32'hbc7765b7),
	.w2(32'hbb7268f9),
	.w3(32'hbbafd140),
	.w4(32'h3b4e22d1),
	.w5(32'hbbbb477a),
	.w6(32'hb9b2159d),
	.w7(32'h3c2865c4),
	.w8(32'hbb164f74),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05abb9),
	.w1(32'hbc92f47f),
	.w2(32'hbcbbe429),
	.w3(32'hbc272e6d),
	.w4(32'h3bbd00ce),
	.w5(32'hbc4b4a3b),
	.w6(32'hbc282fb1),
	.w7(32'hbbcd3922),
	.w8(32'hbc4a19e3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e110a),
	.w1(32'h3c403f7c),
	.w2(32'h39c2e307),
	.w3(32'hbc44cc01),
	.w4(32'h3b48ff8c),
	.w5(32'h3cb9d829),
	.w6(32'hbcb768a8),
	.w7(32'hbc38e262),
	.w8(32'h3b6568a6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b6043),
	.w1(32'h3bbdc036),
	.w2(32'h3ba72587),
	.w3(32'hba5fba3d),
	.w4(32'hbbf7c114),
	.w5(32'hba99d8b4),
	.w6(32'hbc5103d6),
	.w7(32'h3b917698),
	.w8(32'hbd0f23f5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf75eb),
	.w1(32'hbacd9ddc),
	.w2(32'hbc0ff9c2),
	.w3(32'hbae93f84),
	.w4(32'hbbb7fe14),
	.w5(32'hbc056097),
	.w6(32'h3b8e3a59),
	.w7(32'hbb847384),
	.w8(32'h3ce13882),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1c37),
	.w1(32'h3b8e394c),
	.w2(32'h3bc4fa8a),
	.w3(32'hbb8e7bdd),
	.w4(32'h3cb9d7c2),
	.w5(32'h3c48a8c9),
	.w6(32'h3d0a5fab),
	.w7(32'h3bb766b3),
	.w8(32'h3c539666),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9fc1),
	.w1(32'hbc00279d),
	.w2(32'h3be72371),
	.w3(32'hbc52b6a4),
	.w4(32'hbc0d07cd),
	.w5(32'hbb88cde2),
	.w6(32'hbc07b0a9),
	.w7(32'hbc28e1fc),
	.w8(32'h3c2505a3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a176b),
	.w1(32'h3bf2600c),
	.w2(32'hbc197c24),
	.w3(32'h3ac3b320),
	.w4(32'hbc3642bc),
	.w5(32'h3b860c6c),
	.w6(32'hbb205061),
	.w7(32'hbc6ce777),
	.w8(32'h3ba904f0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947625),
	.w1(32'hbca75e2b),
	.w2(32'h3accf8a9),
	.w3(32'h3c03abe3),
	.w4(32'hba109c81),
	.w5(32'h3c6f7ead),
	.w6(32'h3a8dc1cd),
	.w7(32'h3b9be4c0),
	.w8(32'hbcff4c0b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f46b4),
	.w1(32'h3aacf276),
	.w2(32'hbb6f4372),
	.w3(32'h3b81b9e1),
	.w4(32'h3c2e3f16),
	.w5(32'h3c3c2fe4),
	.w6(32'hbc9a9da9),
	.w7(32'hbb564c33),
	.w8(32'hbbb13faf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc327ddd),
	.w1(32'hbc2d4dd0),
	.w2(32'h3c42584c),
	.w3(32'hbc42b266),
	.w4(32'hbbef7f20),
	.w5(32'h3c259193),
	.w6(32'hbb1b72fe),
	.w7(32'h3a3cfa38),
	.w8(32'h3b59e987),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b412b9b),
	.w1(32'h3b19e962),
	.w2(32'hba8291d2),
	.w3(32'hbb5e330b),
	.w4(32'h3aae41bd),
	.w5(32'hbc45f574),
	.w6(32'hbc3845eb),
	.w7(32'hbc4c4872),
	.w8(32'h3be85431),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c238e63),
	.w1(32'hbc37e061),
	.w2(32'h3a0180f0),
	.w3(32'h3b14915d),
	.w4(32'hbc51b4ed),
	.w5(32'h3b1cc434),
	.w6(32'h3d06a609),
	.w7(32'h3c898709),
	.w8(32'hbc712629),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66e5ce),
	.w1(32'hba9f3fb7),
	.w2(32'h3c149b11),
	.w3(32'hbbd4f4cc),
	.w4(32'h3bb894cc),
	.w5(32'h3b5fb74e),
	.w6(32'hbac6adb7),
	.w7(32'hbc4ae089),
	.w8(32'h3c076e17),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8cdfa),
	.w1(32'h3cb466bb),
	.w2(32'h3cba3d59),
	.w3(32'h3c7da26e),
	.w4(32'hbc0df428),
	.w5(32'h3c2bd2ca),
	.w6(32'h3c05bcb3),
	.w7(32'h3ba395fa),
	.w8(32'h3c66bca0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c86c9),
	.w1(32'h3b0af382),
	.w2(32'hbd0244a4),
	.w3(32'hbbed16cb),
	.w4(32'h3ac2bc3b),
	.w5(32'hbbe2b73a),
	.w6(32'hbc7047b1),
	.w7(32'hbc231796),
	.w8(32'h3b490c93),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4170),
	.w1(32'h3c54418b),
	.w2(32'hbb0fd041),
	.w3(32'hbc35a410),
	.w4(32'h3c9e8d01),
	.w5(32'h3b86498e),
	.w6(32'h3b6fb618),
	.w7(32'h3ab00ccd),
	.w8(32'h3bbf7066),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a55d),
	.w1(32'h3c36d72a),
	.w2(32'h3c5d2e30),
	.w3(32'h3c082014),
	.w4(32'hb9bb16a0),
	.w5(32'h3ade2cb2),
	.w6(32'h3c24047e),
	.w7(32'hbbd9b42e),
	.w8(32'hbbed2e5a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87bf7c),
	.w1(32'hb9f1eb89),
	.w2(32'hbb55428f),
	.w3(32'h3c47aed6),
	.w4(32'h3b32c4ac),
	.w5(32'hbb7da25c),
	.w6(32'hbbf5b656),
	.w7(32'h3c77c3f4),
	.w8(32'h3bd3d471),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb881cd),
	.w1(32'hbac7b96e),
	.w2(32'h3badc27c),
	.w3(32'hbc137bd6),
	.w4(32'h3bcad346),
	.w5(32'h3bcc6bf3),
	.w6(32'hbc1045b2),
	.w7(32'h3bbb4ebe),
	.w8(32'hbcce9ecd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbffee),
	.w1(32'h3b27ec11),
	.w2(32'h38e26e47),
	.w3(32'h3c0275f8),
	.w4(32'hbbc74307),
	.w5(32'h3bd04d87),
	.w6(32'h3c3f0e03),
	.w7(32'h3c8054a2),
	.w8(32'h3b225073),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf377ac),
	.w1(32'h3b2eacaf),
	.w2(32'h3c7e51a9),
	.w3(32'hbadec2b5),
	.w4(32'h3c027572),
	.w5(32'hbc82f1ef),
	.w6(32'h3c39cde0),
	.w7(32'h3bb9b3cd),
	.w8(32'hbb7b71e5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebb9d),
	.w1(32'hbb98fa65),
	.w2(32'hbb9c9362),
	.w3(32'h3b06ef23),
	.w4(32'hbc251b99),
	.w5(32'hbbd38d31),
	.w6(32'hbb734b34),
	.w7(32'hbb0d77b3),
	.w8(32'hbca28ba5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb127d),
	.w1(32'hbc0e3c61),
	.w2(32'hbcd2e4d0),
	.w3(32'hbb8f9e65),
	.w4(32'h3cec3add),
	.w5(32'h3bd8faa6),
	.w6(32'hbb97dbdb),
	.w7(32'hbc3805a6),
	.w8(32'hbb8929bc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddbe0a),
	.w1(32'hbb4ef2f2),
	.w2(32'hbbd5daf3),
	.w3(32'hb990c82d),
	.w4(32'hbc025a77),
	.w5(32'hbbe1b9f6),
	.w6(32'h3a31f384),
	.w7(32'hbaa624ae),
	.w8(32'hbbc05dd4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33ea8a),
	.w1(32'hbc5afe25),
	.w2(32'h3b88b6ef),
	.w3(32'hbba58856),
	.w4(32'hbbf5982f),
	.w5(32'hbbebff13),
	.w6(32'h3a871bb8),
	.w7(32'h3854b855),
	.w8(32'h3bfe4fa2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7f6c),
	.w1(32'hb8324d8f),
	.w2(32'h39d4c340),
	.w3(32'hbc23b4a1),
	.w4(32'h3c0cd839),
	.w5(32'hbbaace2d),
	.w6(32'hbbdadbd8),
	.w7(32'hbac7c683),
	.w8(32'hba9aabe8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71dee3),
	.w1(32'h3b7a374c),
	.w2(32'h3bbbfe15),
	.w3(32'hbc15d198),
	.w4(32'hbb3b0c12),
	.w5(32'h3b7484a5),
	.w6(32'hbc8c6d95),
	.w7(32'hbc6c99c6),
	.w8(32'h3c1c52d3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92dada),
	.w1(32'hbaea9e70),
	.w2(32'h3bb4013d),
	.w3(32'hbb1adc57),
	.w4(32'h3b76bae8),
	.w5(32'hbac2db77),
	.w6(32'h3bd83d11),
	.w7(32'h3bc5ec6e),
	.w8(32'hbbd38c8e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a83cf),
	.w1(32'hbad30553),
	.w2(32'hbc7563e7),
	.w3(32'hbc25fb54),
	.w4(32'h3ba04b8c),
	.w5(32'hbb1c6630),
	.w6(32'hbb43bdd5),
	.w7(32'hbbb77446),
	.w8(32'h39fbb2ce),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c92c3),
	.w1(32'hbbd4e091),
	.w2(32'hbb932118),
	.w3(32'h3b0cac94),
	.w4(32'hba6a5672),
	.w5(32'h39b0c1dc),
	.w6(32'hbba9ef5f),
	.w7(32'h3a6f387c),
	.w8(32'h3c8515bc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94528c),
	.w1(32'h3c053c6e),
	.w2(32'h3ca2ea76),
	.w3(32'hbbcbb7ce),
	.w4(32'h3ac88deb),
	.w5(32'h3b37d5cf),
	.w6(32'h3a9367d1),
	.w7(32'h3b6c9270),
	.w8(32'h3d28c61d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97409b),
	.w1(32'h3bc238f1),
	.w2(32'hbb30ca73),
	.w3(32'hbc08b105),
	.w4(32'h3a8edf1f),
	.w5(32'hbc1948f5),
	.w6(32'hbc749bc9),
	.w7(32'hbc6c50d4),
	.w8(32'hbc919d64),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c666fff),
	.w1(32'hbbed3aaa),
	.w2(32'hbcc3d174),
	.w3(32'hbb78986d),
	.w4(32'h3b9c87d5),
	.w5(32'h3aa42b0d),
	.w6(32'h3bd9082b),
	.w7(32'hbb8c0054),
	.w8(32'h3b3a3836),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae9f5),
	.w1(32'h3ba8fb81),
	.w2(32'h3bcc6e12),
	.w3(32'hbacb5fab),
	.w4(32'h3cb32b81),
	.w5(32'h3cc2d71d),
	.w6(32'h3b95fde5),
	.w7(32'hbc5556cb),
	.w8(32'h3c8b3846),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a706d),
	.w1(32'hbb0c7542),
	.w2(32'h3b6837b1),
	.w3(32'h3a8e9826),
	.w4(32'h3cfabe38),
	.w5(32'hbbdd12d7),
	.w6(32'h3b9affcf),
	.w7(32'hbb9d6865),
	.w8(32'hbad59a63),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587e0a),
	.w1(32'h398f83a0),
	.w2(32'h3a746f84),
	.w3(32'h3be019be),
	.w4(32'hbc85376c),
	.w5(32'hba9042f7),
	.w6(32'hba87747b),
	.w7(32'hbbdbecca),
	.w8(32'hbbf248f5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dcb62),
	.w1(32'hbcfaaa50),
	.w2(32'h3aee52df),
	.w3(32'hbc299bcf),
	.w4(32'h3c9cd4fa),
	.w5(32'hbbdc5522),
	.w6(32'hbabce771),
	.w7(32'hbc69de8c),
	.w8(32'h3c808b2b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a389),
	.w1(32'hbc5ce6c5),
	.w2(32'hbc372268),
	.w3(32'hbc11fe74),
	.w4(32'hbc936324),
	.w5(32'h3c19b578),
	.w6(32'hba636325),
	.w7(32'hbd32f004),
	.w8(32'hbc057154),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e6189),
	.w1(32'hba35dc1b),
	.w2(32'h3bfe7d12),
	.w3(32'h3c5a6d91),
	.w4(32'h3b82979a),
	.w5(32'hbc0e1ee2),
	.w6(32'h3b5b2e51),
	.w7(32'h3bdf8875),
	.w8(32'h3ba7464c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2e9b),
	.w1(32'hbbea4bfc),
	.w2(32'hbbc793be),
	.w3(32'h3c0b8a83),
	.w4(32'hba570560),
	.w5(32'hbbae0405),
	.w6(32'hbc3f2230),
	.w7(32'h3b9333e7),
	.w8(32'hbc00f92d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aa161),
	.w1(32'hbacd6794),
	.w2(32'hbbf179e5),
	.w3(32'h3bcd3d2f),
	.w4(32'h39cea62e),
	.w5(32'hbc16f179),
	.w6(32'h3d0a5ad6),
	.w7(32'hbbd4ff08),
	.w8(32'hbc8b54d4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3f99),
	.w1(32'h3c100f6e),
	.w2(32'hb9acb43a),
	.w3(32'hbba735d4),
	.w4(32'hbb5410c1),
	.w5(32'hbafd7d2f),
	.w6(32'h3a09783a),
	.w7(32'hbc038b1a),
	.w8(32'h3986f14c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08af7),
	.w1(32'h3b67efe7),
	.w2(32'hbb6ca1ca),
	.w3(32'h3b0de4bc),
	.w4(32'hbbb21762),
	.w5(32'hbbfd7df5),
	.w6(32'hbc12f643),
	.w7(32'hbb55c27f),
	.w8(32'h3bf1119a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b1cf),
	.w1(32'h3c00bd4b),
	.w2(32'hbb16ea8e),
	.w3(32'hbc63ebc3),
	.w4(32'hbb92704d),
	.w5(32'hbcb98e8c),
	.w6(32'hbbb16e39),
	.w7(32'hbc738295),
	.w8(32'h3bec5e06),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2147da),
	.w1(32'hb94cbf9e),
	.w2(32'h3c9c3f1a),
	.w3(32'hbaff1d55),
	.w4(32'hbba11311),
	.w5(32'h3c58e586),
	.w6(32'hbc4885b2),
	.w7(32'h3be73ae8),
	.w8(32'hbbaef93c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07bb58),
	.w1(32'h3b167626),
	.w2(32'h3a3767cc),
	.w3(32'h3c0666c4),
	.w4(32'hbae87ef3),
	.w5(32'hba84e4d9),
	.w6(32'h3a423fe3),
	.w7(32'hbb1ddefd),
	.w8(32'h3c42ba84),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8436f6),
	.w1(32'hbbac081e),
	.w2(32'h3c69993b),
	.w3(32'hbc50692a),
	.w4(32'hbc6374ed),
	.w5(32'h3c0f8394),
	.w6(32'hbbff091d),
	.w7(32'h3c1bb957),
	.w8(32'hbb86ba8b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68394),
	.w1(32'hbcf3016a),
	.w2(32'hbc1e0dfe),
	.w3(32'h3c002369),
	.w4(32'hbb5d6c2a),
	.w5(32'hbc05ff6c),
	.w6(32'h3c694e00),
	.w7(32'h3c5acc60),
	.w8(32'hbcd6a82c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65222c),
	.w1(32'h3c559882),
	.w2(32'h3c99d421),
	.w3(32'hbbce122e),
	.w4(32'hbacb4b8c),
	.w5(32'h39487b13),
	.w6(32'hbc97184c),
	.w7(32'h3c47957a),
	.w8(32'hbc65f072),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38bb1b),
	.w1(32'hbbbffd76),
	.w2(32'h3b788d85),
	.w3(32'hbbe9b6a3),
	.w4(32'hbc1012fa),
	.w5(32'h3c253009),
	.w6(32'hbc7e85e6),
	.w7(32'hbbb24ba4),
	.w8(32'hbbad173d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeae99a),
	.w1(32'hbc0bd86c),
	.w2(32'hbce3ef81),
	.w3(32'hbb5868df),
	.w4(32'hbb8733dc),
	.w5(32'hbc1ae710),
	.w6(32'hbbdfaa46),
	.w7(32'hbc820355),
	.w8(32'hbc044f61),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d9e6),
	.w1(32'hbb7e5d2d),
	.w2(32'h3ca4566d),
	.w3(32'h3ae3f561),
	.w4(32'h3c0b9b93),
	.w5(32'h3c975962),
	.w6(32'h3b27a533),
	.w7(32'h3c1f47cf),
	.w8(32'h3caae250),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dba38),
	.w1(32'hba6d4891),
	.w2(32'h3ac6dee7),
	.w3(32'h3986ec8d),
	.w4(32'hbbe4a780),
	.w5(32'hbc33ff87),
	.w6(32'hba73f137),
	.w7(32'hbc32e8bc),
	.w8(32'hbb163730),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d95c0),
	.w1(32'h3c2f4e67),
	.w2(32'hbc77ea32),
	.w3(32'hbc49e6a8),
	.w4(32'hbbb39f78),
	.w5(32'hbb988120),
	.w6(32'hbc0cdb7c),
	.w7(32'h3b469c34),
	.w8(32'hbb8499b6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9421bd),
	.w1(32'h3c1cb6ae),
	.w2(32'hbc529cf1),
	.w3(32'hba170edd),
	.w4(32'hbcdede49),
	.w5(32'h3ba5c846),
	.w6(32'hba114a7d),
	.w7(32'h3c255e08),
	.w8(32'h3b0892f1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0ca7),
	.w1(32'h3ad51c12),
	.w2(32'hbb3b838d),
	.w3(32'hbb73bddb),
	.w4(32'hbb8e49ea),
	.w5(32'hbbb37877),
	.w6(32'h3a08160e),
	.w7(32'hba9ca441),
	.w8(32'h3c093923),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b0d54),
	.w1(32'h3bed6dc0),
	.w2(32'hbaf22c06),
	.w3(32'hbb444416),
	.w4(32'h3c545b0d),
	.w5(32'hbabb735b),
	.w6(32'hbb8e024f),
	.w7(32'h3b76e7a5),
	.w8(32'hbb9c515a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5934ef),
	.w1(32'hbc117a63),
	.w2(32'hbc9f35c0),
	.w3(32'hbc218257),
	.w4(32'hbc8ddf53),
	.w5(32'hbcb30039),
	.w6(32'hbb60f97c),
	.w7(32'h3b69065d),
	.w8(32'hbc14c76f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb047c46),
	.w1(32'h3c38c34e),
	.w2(32'h3c11d4dc),
	.w3(32'hbab72204),
	.w4(32'h3cb4b4d1),
	.w5(32'h3c2891e5),
	.w6(32'h3c181d7d),
	.w7(32'h3b6db7a2),
	.w8(32'h3cb3d53b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfcff21),
	.w1(32'h3cb6fedf),
	.w2(32'hbc0168c9),
	.w3(32'hbc5ab2ae),
	.w4(32'hbcb847e6),
	.w5(32'hbbceb588),
	.w6(32'hbc20c468),
	.w7(32'hbb789125),
	.w8(32'hbbb762e7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f2fd),
	.w1(32'h3bd56514),
	.w2(32'hbae8e0f5),
	.w3(32'hba781958),
	.w4(32'h3bc90383),
	.w5(32'hbc05016e),
	.w6(32'h3b74627d),
	.w7(32'hb9ee8177),
	.w8(32'h39f58424),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31f0d1),
	.w1(32'hbc142068),
	.w2(32'hbc0d7c8d),
	.w3(32'hba99f325),
	.w4(32'h3c13f077),
	.w5(32'h3aafbe1c),
	.w6(32'h3ac3c876),
	.w7(32'h3a5e0aa2),
	.w8(32'h3c5ba461),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d71a),
	.w1(32'hbc160e63),
	.w2(32'hbb8d3514),
	.w3(32'h3af9ed06),
	.w4(32'h3c815257),
	.w5(32'hbbb5d17a),
	.w6(32'hba59cc9b),
	.w7(32'hbbbfa66c),
	.w8(32'h3b4a7fc6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3839e3),
	.w1(32'hbb70aad4),
	.w2(32'h3c0df9fd),
	.w3(32'hbacc0eef),
	.w4(32'h3ae08c96),
	.w5(32'hbb7f51a1),
	.w6(32'hbc310e13),
	.w7(32'h3b247f2d),
	.w8(32'hbc1d9a7d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d014),
	.w1(32'h3ac37ab7),
	.w2(32'hbc2baa7f),
	.w3(32'h3beb789d),
	.w4(32'h3be5d8d8),
	.w5(32'hbcf36849),
	.w6(32'hbb1046da),
	.w7(32'h3c05a757),
	.w8(32'hbaafc918),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07edd4),
	.w1(32'h3c7af624),
	.w2(32'hba81395a),
	.w3(32'hbc8f68fc),
	.w4(32'hbb3eec70),
	.w5(32'h3b2a4fbd),
	.w6(32'hbc8619cf),
	.w7(32'hbbcefd4f),
	.w8(32'hbbb386a9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75bfa),
	.w1(32'h3c05af03),
	.w2(32'h3c372d46),
	.w3(32'h3b48af83),
	.w4(32'h3bd30537),
	.w5(32'h3a54dee1),
	.w6(32'h3baceb90),
	.w7(32'hbbc8165f),
	.w8(32'h3b849753),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb531418),
	.w1(32'h3b96dc4e),
	.w2(32'h3c21850d),
	.w3(32'h3b67d1be),
	.w4(32'h3bf0cce7),
	.w5(32'h3b949175),
	.w6(32'h3ada22aa),
	.w7(32'hbafabd2b),
	.w8(32'h3bac40d8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af0bc),
	.w1(32'hbbae5d1b),
	.w2(32'h3c7af224),
	.w3(32'hbb1da413),
	.w4(32'hbc059ce9),
	.w5(32'h3bcf562e),
	.w6(32'hbb9f8643),
	.w7(32'h3a8b97b8),
	.w8(32'hbbb42b14),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf2f7d),
	.w1(32'hbb32a8f6),
	.w2(32'hbb003cd0),
	.w3(32'h3c36cf90),
	.w4(32'h3c93b91b),
	.w5(32'h3c631a81),
	.w6(32'h3c5605ea),
	.w7(32'h3b68a2a4),
	.w8(32'h3c20260d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54a74f),
	.w1(32'h3b58b96c),
	.w2(32'h3c16bf14),
	.w3(32'hbbe7a5eb),
	.w4(32'hbc1bea41),
	.w5(32'h3a4ec6eb),
	.w6(32'h3aca3ff4),
	.w7(32'h3b4f01dc),
	.w8(32'hba7ed16b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944de7f),
	.w1(32'h3aad90d0),
	.w2(32'h3c0284cc),
	.w3(32'h3b397ba7),
	.w4(32'h3c188f3c),
	.w5(32'h3b44f52f),
	.w6(32'h3bb1e766),
	.w7(32'h3a47f775),
	.w8(32'h3b1040b8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf83518),
	.w1(32'hbbcaa764),
	.w2(32'hbbc19e9d),
	.w3(32'hbc5a8ded),
	.w4(32'h3c700d41),
	.w5(32'hbc23cea6),
	.w6(32'h3b7f4f08),
	.w7(32'h3bd2deab),
	.w8(32'h3a77c309),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4cd70),
	.w1(32'h3b41c779),
	.w2(32'hb8b16db9),
	.w3(32'hbbd97e28),
	.w4(32'hb9f7b1d0),
	.w5(32'h3b525c8b),
	.w6(32'hbb9b5c11),
	.w7(32'h3c4117be),
	.w8(32'h3b31d5ab),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee807c),
	.w1(32'h3b9e1b5b),
	.w2(32'h3c1c3152),
	.w3(32'hbc19cfb7),
	.w4(32'h3c8df890),
	.w5(32'hbc2072b2),
	.w6(32'h3c85aee3),
	.w7(32'h3aaac969),
	.w8(32'hbc440726),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06a994),
	.w1(32'hbc51c3a9),
	.w2(32'hbba34375),
	.w3(32'hbba87585),
	.w4(32'hbbbd0c39),
	.w5(32'hbc9db3fa),
	.w6(32'hbc56f0a1),
	.w7(32'hbb75caba),
	.w8(32'hbc082c48),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc819ed),
	.w1(32'h3b3973fb),
	.w2(32'h3c994957),
	.w3(32'h3bba660b),
	.w4(32'hbaef7560),
	.w5(32'h3c5481c4),
	.w6(32'hbbc3323b),
	.w7(32'h3bff7110),
	.w8(32'hbbf21df1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c873e),
	.w1(32'hbb15cdee),
	.w2(32'h3c87a9e6),
	.w3(32'h3c37483c),
	.w4(32'h3ad4bd8e),
	.w5(32'h3b7770f9),
	.w6(32'hbbfcf29b),
	.w7(32'hbbcc9bd3),
	.w8(32'hbb70d9de),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8df01),
	.w1(32'h3a82e685),
	.w2(32'h3bc4fcc5),
	.w3(32'hbb863e73),
	.w4(32'h37072335),
	.w5(32'h3bc03f8d),
	.w6(32'hb80ae85a),
	.w7(32'hba7a9b50),
	.w8(32'hba138cc5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42054),
	.w1(32'hbbf5c2b0),
	.w2(32'h3a5134a7),
	.w3(32'hba806f3e),
	.w4(32'hbbd118aa),
	.w5(32'hbbad7893),
	.w6(32'hbade36dc),
	.w7(32'hbcabbf71),
	.w8(32'h39b6daf6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965fb4),
	.w1(32'h3be684a7),
	.w2(32'hbb2df014),
	.w3(32'h3c03871a),
	.w4(32'h3c226229),
	.w5(32'hbb2c518c),
	.w6(32'h3c9b0d6f),
	.w7(32'h3b6c2702),
	.w8(32'hbbd5dc86),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b011dad),
	.w1(32'hbb60c9c4),
	.w2(32'hbc543b68),
	.w3(32'hbc6c4e5a),
	.w4(32'hbc5ed281),
	.w5(32'hbc26314d),
	.w6(32'hbc315d47),
	.w7(32'hbc0a3fd5),
	.w8(32'hbc6f5271),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb79bd),
	.w1(32'h3a18b796),
	.w2(32'hbc01aee9),
	.w3(32'hbbcf0483),
	.w4(32'hb9f2ede2),
	.w5(32'hbafcbde3),
	.w6(32'hbbf8720b),
	.w7(32'h3bad4a3f),
	.w8(32'hbca7c916),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17cdf9),
	.w1(32'hbaf834ba),
	.w2(32'h3bb1d86d),
	.w3(32'h3b368040),
	.w4(32'h3b6588ab),
	.w5(32'h3b061bf8),
	.w6(32'h3bbe2b28),
	.w7(32'h3bf0e3fd),
	.w8(32'h3b9dc6f2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f04b),
	.w1(32'h3be634bc),
	.w2(32'hb9b104f1),
	.w3(32'hb955e8c1),
	.w4(32'h3ca96da7),
	.w5(32'h3c0290a0),
	.w6(32'h3c35acee),
	.w7(32'hbb01cb52),
	.w8(32'hbc40a3d2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3caf38),
	.w1(32'hbbf0ffbe),
	.w2(32'hb9a542f7),
	.w3(32'h3b4acde3),
	.w4(32'hbc131093),
	.w5(32'hbb730451),
	.w6(32'h3b416bd6),
	.w7(32'hbc6ff9fc),
	.w8(32'hbc3a21aa),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afb21d),
	.w1(32'hbb864657),
	.w2(32'h3b5e8706),
	.w3(32'hbc3be251),
	.w4(32'hbc2ed38a),
	.w5(32'h3b0f9d94),
	.w6(32'h3ad49110),
	.w7(32'hbbb0db81),
	.w8(32'h3b82c9f7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9efc8),
	.w1(32'hbae87179),
	.w2(32'h3b3aeeda),
	.w3(32'h3be6c1af),
	.w4(32'hbc95d4b8),
	.w5(32'h3bae3f72),
	.w6(32'hbbb6c31e),
	.w7(32'hbc0a7bd2),
	.w8(32'hbb56bb31),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ffb9c),
	.w1(32'hbbb8e7ba),
	.w2(32'h3b61b0c0),
	.w3(32'h3cc53693),
	.w4(32'hbc06e089),
	.w5(32'hbc1433fb),
	.w6(32'h3c3ce4e5),
	.w7(32'h3b045366),
	.w8(32'hbbb10cb7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809e25),
	.w1(32'h3ba33147),
	.w2(32'h39d0ae0d),
	.w3(32'hbd5c1489),
	.w4(32'hbbc0456c),
	.w5(32'h3c896d98),
	.w6(32'hbb455ffc),
	.w7(32'h3cec318c),
	.w8(32'h3ae3f877),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919634a),
	.w1(32'h3b1326e7),
	.w2(32'hbbad4d54),
	.w3(32'h3c27349c),
	.w4(32'hbca52811),
	.w5(32'hbc2bdaa2),
	.w6(32'h3c2d7b50),
	.w7(32'hbc5c0e28),
	.w8(32'hbd1d1084),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a6da9),
	.w1(32'h3bfd327e),
	.w2(32'hbc7e267b),
	.w3(32'hbc319320),
	.w4(32'h3d06a707),
	.w5(32'h3c082888),
	.w6(32'h3b9fa979),
	.w7(32'h3b55a797),
	.w8(32'h3b3af99c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0129f),
	.w1(32'h3bdc1a0d),
	.w2(32'hbb991e2e),
	.w3(32'hbd00c2af),
	.w4(32'hbba5184a),
	.w5(32'h3a78bc99),
	.w6(32'h3b85a6c5),
	.w7(32'h3bee4c40),
	.w8(32'hbbf4c2d9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb69425),
	.w1(32'hbd023fcc),
	.w2(32'hbd05f1ef),
	.w3(32'hbb10b43e),
	.w4(32'h3b74cc09),
	.w5(32'hbc1d81fc),
	.w6(32'hbca01c36),
	.w7(32'hbc73068a),
	.w8(32'hbc8ca38c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac425b9),
	.w1(32'hbbca7545),
	.w2(32'hbbc97589),
	.w3(32'h3cb750e1),
	.w4(32'hbd281550),
	.w5(32'h3ba14730),
	.w6(32'hbbf913b7),
	.w7(32'hbbec7b79),
	.w8(32'hbb76ddd1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c718ea5),
	.w1(32'h3a372c38),
	.w2(32'h3bfbb92b),
	.w3(32'h3bbbcdec),
	.w4(32'hbba5da87),
	.w5(32'h3a0ec1c8),
	.w6(32'h3bdf6f93),
	.w7(32'hbb990598),
	.w8(32'h3be92565),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73673c),
	.w1(32'h3c146324),
	.w2(32'hbc16722a),
	.w3(32'hbb8057af),
	.w4(32'h3ba766b3),
	.w5(32'hbca64b95),
	.w6(32'h3c651461),
	.w7(32'hbca5dd5d),
	.w8(32'hbb54f76d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23fe6c),
	.w1(32'h3a92eab3),
	.w2(32'h3b298925),
	.w3(32'h3c0ca02d),
	.w4(32'h3b95ebe8),
	.w5(32'hbba017a6),
	.w6(32'hbc330439),
	.w7(32'hbca284f0),
	.w8(32'hbb49646e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bd6ad),
	.w1(32'h3b903155),
	.w2(32'h3cac22ea),
	.w3(32'hbce9f67d),
	.w4(32'hb99b0e0e),
	.w5(32'h3b887d16),
	.w6(32'h3a95ea1f),
	.w7(32'hbc035ec9),
	.w8(32'hbc60a07c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3eedc),
	.w1(32'h3af7062e),
	.w2(32'h3c080fc9),
	.w3(32'hbb042fe7),
	.w4(32'hbb272c99),
	.w5(32'hbbcfaf76),
	.w6(32'h398b527e),
	.w7(32'hbb0fa3b9),
	.w8(32'h3b8d7516),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc85a03),
	.w1(32'hba28d1b2),
	.w2(32'h3d253096),
	.w3(32'h39a96ff0),
	.w4(32'hbc96d99e),
	.w5(32'h3c2af800),
	.w6(32'h3bfe1137),
	.w7(32'h3c48123c),
	.w8(32'h3bfd49ed),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967c6d),
	.w1(32'hbb13e5b0),
	.w2(32'h3a2b4af1),
	.w3(32'h3bee9cff),
	.w4(32'hbc89f3c4),
	.w5(32'h3d044169),
	.w6(32'hbc86a67e),
	.w7(32'h3bd9a82a),
	.w8(32'h3886c5d0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bb795),
	.w1(32'hbac7326e),
	.w2(32'h3ccc0831),
	.w3(32'hbadb801e),
	.w4(32'h3c8081de),
	.w5(32'hbbba7ca6),
	.w6(32'hba33b00d),
	.w7(32'hbc48a0c9),
	.w8(32'h3c875680),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfce379),
	.w1(32'h3b67b69b),
	.w2(32'hbc487fcf),
	.w3(32'hbc42bb8f),
	.w4(32'h3b796e54),
	.w5(32'hbbba70e9),
	.w6(32'hbcfaf804),
	.w7(32'hbba857b6),
	.w8(32'hbc3d8a22),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba334b0),
	.w1(32'hbbe94271),
	.w2(32'hbbfe8c48),
	.w3(32'hbb9cfee8),
	.w4(32'hbc0608bb),
	.w5(32'hbc84081b),
	.w6(32'hbb2a35a0),
	.w7(32'hbaee5d59),
	.w8(32'hbc396d66),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76f441),
	.w1(32'hbbf04782),
	.w2(32'h3ad065fc),
	.w3(32'h3d050280),
	.w4(32'h3c042625),
	.w5(32'hb9b55dc0),
	.w6(32'h3c63cf7b),
	.w7(32'h3c5ee2a9),
	.w8(32'h3cb02137),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce6ca8),
	.w1(32'h3bb1d782),
	.w2(32'h3b68c28b),
	.w3(32'hbbed5309),
	.w4(32'hbbc8d81e),
	.w5(32'h3b0f2766),
	.w6(32'h3b381093),
	.w7(32'h3c19d672),
	.w8(32'hbb0b2a19),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951fa5f),
	.w1(32'hbba93692),
	.w2(32'h3b05d5bc),
	.w3(32'hbb792881),
	.w4(32'hb9def8bb),
	.w5(32'h3aef9875),
	.w6(32'hbc95c740),
	.w7(32'h3bff7774),
	.w8(32'hbb127aba),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdad753),
	.w1(32'hbb009f3f),
	.w2(32'h3b4471e8),
	.w3(32'hbbbd662c),
	.w4(32'hba34be3f),
	.w5(32'h3b6915f5),
	.w6(32'hbab90698),
	.w7(32'hbb58a028),
	.w8(32'h3c726036),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159665),
	.w1(32'hbc7e70b3),
	.w2(32'h3c2a88a7),
	.w3(32'h3c48a565),
	.w4(32'hbb2b77dc),
	.w5(32'hbc0c5051),
	.w6(32'hba786a20),
	.w7(32'hbc02322e),
	.w8(32'hbbce717a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10cae1),
	.w1(32'h39098d97),
	.w2(32'hbbc560ff),
	.w3(32'h3ca8098e),
	.w4(32'hbc1e2287),
	.w5(32'hba309cfe),
	.w6(32'h3b46900e),
	.w7(32'hbd46bee6),
	.w8(32'hbc22d04f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80139),
	.w1(32'h3b8a9573),
	.w2(32'h3829c338),
	.w3(32'h3caf67db),
	.w4(32'h3bb445a0),
	.w5(32'hbb959599),
	.w6(32'h39be58e7),
	.w7(32'hba9b23c5),
	.w8(32'h3a1143a1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4066aa),
	.w1(32'hbc325ce3),
	.w2(32'h3b07ce4a),
	.w3(32'h3ba13b95),
	.w4(32'hbb95e5b6),
	.w5(32'h3a0fa269),
	.w6(32'hbabd3f6a),
	.w7(32'h3be281f5),
	.w8(32'hbb4441fb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ddfb3),
	.w1(32'hb8e22ea4),
	.w2(32'h3c6b9f78),
	.w3(32'h3c3287dc),
	.w4(32'h3ae10fce),
	.w5(32'hbaebf44f),
	.w6(32'hbaf9247f),
	.w7(32'hbb9e74e2),
	.w8(32'hbbfe7e54),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc8f27),
	.w1(32'hbc38cdae),
	.w2(32'hbc6d467c),
	.w3(32'hbb27cdfd),
	.w4(32'h3a86561e),
	.w5(32'hba9e35fc),
	.w6(32'hb9b5a4c3),
	.w7(32'hbb48ea39),
	.w8(32'hb9fe54fe),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77cbe1),
	.w1(32'hbb955c39),
	.w2(32'hbbc8817f),
	.w3(32'hbbf54115),
	.w4(32'h3c1ff209),
	.w5(32'hbc183f94),
	.w6(32'hbb98341b),
	.w7(32'hbbaa5c03),
	.w8(32'h3b96f2e0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce962bd),
	.w1(32'hbc4bbe65),
	.w2(32'hbae2e5c9),
	.w3(32'h3a304033),
	.w4(32'hbc4be344),
	.w5(32'hbc86360a),
	.w6(32'hbba1d43d),
	.w7(32'hbc90f2ff),
	.w8(32'h3a457d9b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae604b),
	.w1(32'hbbd306ad),
	.w2(32'h3b0bc09b),
	.w3(32'hbc5c747c),
	.w4(32'hbb92a23c),
	.w5(32'hbcdd24fc),
	.w6(32'h3aa5a11b),
	.w7(32'h3c6a9668),
	.w8(32'hbc4ec642),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c7e9b),
	.w1(32'hba6c1247),
	.w2(32'h3b52047b),
	.w3(32'hbc1ef5c9),
	.w4(32'h3b5621c5),
	.w5(32'hbb555545),
	.w6(32'h3b9da982),
	.w7(32'hbcaf779a),
	.w8(32'h3c54f169),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule