module layer_10_featuremap_349(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6234a),
	.w1(32'hbbc912ee),
	.w2(32'hbb70edcd),
	.w3(32'hba3b4593),
	.w4(32'hb9929210),
	.w5(32'h3b119ef3),
	.w6(32'h39bfdbce),
	.w7(32'hbb2acd3b),
	.w8(32'hbb134ef5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae45a1f),
	.w1(32'hbbbbf230),
	.w2(32'h3b62513e),
	.w3(32'hbb936c05),
	.w4(32'hbb47500d),
	.w5(32'hbb5196b0),
	.w6(32'hbbcf226a),
	.w7(32'hbb544477),
	.w8(32'hbc26f33b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bdbe7),
	.w1(32'h3ab7701c),
	.w2(32'hbc1df230),
	.w3(32'hbc19a8d6),
	.w4(32'hbb9e4f0c),
	.w5(32'h3b0ba0c4),
	.w6(32'h3ab6793c),
	.w7(32'hb9acddcf),
	.w8(32'h3aef1d96),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8d965),
	.w1(32'h3b8f5eb6),
	.w2(32'h3c31a6b1),
	.w3(32'h3ba40d23),
	.w4(32'h3bebf623),
	.w5(32'hba2853ce),
	.w6(32'h3b260921),
	.w7(32'h3b98ac42),
	.w8(32'h3c565c40),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba444),
	.w1(32'h3bafe23f),
	.w2(32'hbb9aacda),
	.w3(32'h3ac8970d),
	.w4(32'hbb1bec1a),
	.w5(32'hbacc21f8),
	.w6(32'h3c2ee59c),
	.w7(32'h3bfe2cf8),
	.w8(32'hbaedd7c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2499c5),
	.w1(32'hbb8fedd6),
	.w2(32'hba9d5310),
	.w3(32'hb94ee861),
	.w4(32'hbaf9efae),
	.w5(32'hbbe1995a),
	.w6(32'h3b4af1f1),
	.w7(32'hbb90f2d1),
	.w8(32'hbb95196e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb233e2),
	.w1(32'hbbebbfcf),
	.w2(32'hbbd5ddcf),
	.w3(32'hbb446bbf),
	.w4(32'hbb886f13),
	.w5(32'hbc406c24),
	.w6(32'h3a23c9f2),
	.w7(32'hbc1c932e),
	.w8(32'hbbbca11c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2687ac),
	.w1(32'hba9d64c3),
	.w2(32'hbba099a6),
	.w3(32'hbbd6cc62),
	.w4(32'hbacd461f),
	.w5(32'hbc778d2e),
	.w6(32'h3b529db8),
	.w7(32'hb9599724),
	.w8(32'hbc5327c6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc460d9c),
	.w1(32'hbc1b9d6f),
	.w2(32'hbc23b772),
	.w3(32'hbc0d5933),
	.w4(32'hbc2d4244),
	.w5(32'h3b61139f),
	.w6(32'hbb7bac8f),
	.w7(32'hbc174d3d),
	.w8(32'h3ae19140),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00854c),
	.w1(32'hb8e5f8bc),
	.w2(32'hbb38778f),
	.w3(32'h3b5ea9d9),
	.w4(32'h3add3cf4),
	.w5(32'hbbdcdf3c),
	.w6(32'h3b6c0c3c),
	.w7(32'hbb0ceff9),
	.w8(32'hbb80007b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a594daa),
	.w1(32'hbb1f5e8a),
	.w2(32'h3b2e0c27),
	.w3(32'h3afb7283),
	.w4(32'h3ad49485),
	.w5(32'hbb466cee),
	.w6(32'h3be064ad),
	.w7(32'hbadb309c),
	.w8(32'hbc2baaa0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56bb08),
	.w1(32'h3c21785b),
	.w2(32'hbc68cc75),
	.w3(32'hbc2d87ae),
	.w4(32'hbb895131),
	.w5(32'hbac50153),
	.w6(32'hba4e3cfe),
	.w7(32'h3bab681f),
	.w8(32'h3c2b6b3c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63766),
	.w1(32'h3ae316b2),
	.w2(32'hbc27789a),
	.w3(32'hba806283),
	.w4(32'hbbdd0c53),
	.w5(32'hbc08a11c),
	.w6(32'h3c95ff3b),
	.w7(32'h3bf85556),
	.w8(32'hbbe65dd4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c195db),
	.w1(32'hba8e30ca),
	.w2(32'hbbfcc9b7),
	.w3(32'h3850c9ff),
	.w4(32'hbb5377af),
	.w5(32'h3a9c623d),
	.w6(32'h3c0403e5),
	.w7(32'h3a870957),
	.w8(32'hbb587bd3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0158eb),
	.w1(32'hbac22219),
	.w2(32'h3b188500),
	.w3(32'h3bac1dce),
	.w4(32'h3bbf3a17),
	.w5(32'hbaa4a9e7),
	.w6(32'h3be9f84d),
	.w7(32'h3af1edbe),
	.w8(32'hbac8c74b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39204d22),
	.w1(32'hbbc75e49),
	.w2(32'hbaf6b436),
	.w3(32'hbb54d7a2),
	.w4(32'h3ad9fffa),
	.w5(32'hbc226041),
	.w6(32'h3b7b0373),
	.w7(32'h3a9caad3),
	.w8(32'hbb655d66),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd6267),
	.w1(32'hbc3b698b),
	.w2(32'hbc03a9b5),
	.w3(32'hbb7e0400),
	.w4(32'hbaf7e98e),
	.w5(32'h392d8881),
	.w6(32'h3c4c7a26),
	.w7(32'hbb917df8),
	.w8(32'hbb480491),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902eed9),
	.w1(32'hb9984efa),
	.w2(32'hbb26027c),
	.w3(32'h3b56d663),
	.w4(32'hbaeb6366),
	.w5(32'hb8b5eecc),
	.w6(32'hbb6a1ce8),
	.w7(32'h3b0fba5a),
	.w8(32'h3bc678ab),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07ea51),
	.w1(32'h3b86a44d),
	.w2(32'h3beddd75),
	.w3(32'h3c37721e),
	.w4(32'h3bcf6d4c),
	.w5(32'hba858074),
	.w6(32'h3c280c1f),
	.w7(32'h3c12bba6),
	.w8(32'h39939bd8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fcd5d),
	.w1(32'h3a1b0ae1),
	.w2(32'h3b0d36f9),
	.w3(32'h3ab33852),
	.w4(32'hbb9bd37d),
	.w5(32'h3b3b778a),
	.w6(32'h3b81ed0d),
	.w7(32'hbb02632d),
	.w8(32'hbb626e51),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac72ed0),
	.w1(32'hbaaab17c),
	.w2(32'h3a2ec390),
	.w3(32'hba84ec59),
	.w4(32'hbae405d1),
	.w5(32'h3a40ac3b),
	.w6(32'h3b803f72),
	.w7(32'h3abdfccd),
	.w8(32'hbab9e985),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9098271),
	.w1(32'hba868660),
	.w2(32'hba58b909),
	.w3(32'hbb197405),
	.w4(32'hbac46586),
	.w5(32'hbb03948d),
	.w6(32'hbc01cb11),
	.w7(32'hbb208708),
	.w8(32'hbbdfd28f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8cf85),
	.w1(32'h3b88579d),
	.w2(32'hbbddc5ba),
	.w3(32'hbb5fc5c3),
	.w4(32'h3b646b3b),
	.w5(32'hbb247a61),
	.w6(32'hbb9c11b8),
	.w7(32'h3b08914b),
	.w8(32'h3b6d7e58),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e6016),
	.w1(32'hbb82f720),
	.w2(32'h3b796a85),
	.w3(32'h3b6c3a0a),
	.w4(32'h3ad9e271),
	.w5(32'hbac74ef4),
	.w6(32'h3bab1379),
	.w7(32'h3a36b919),
	.w8(32'hbaba6ca6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34bfca),
	.w1(32'hba96643a),
	.w2(32'hbbbae678),
	.w3(32'hb91bc97f),
	.w4(32'h3abf6265),
	.w5(32'hba05fb6d),
	.w6(32'hbc340176),
	.w7(32'h3c3be86d),
	.w8(32'hbb04ff6b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb427466),
	.w1(32'hbbbb7f83),
	.w2(32'h3b4a3a4d),
	.w3(32'hbb4f472a),
	.w4(32'h3b0cbfbf),
	.w5(32'h3ba0db69),
	.w6(32'h3c1c75d0),
	.w7(32'hbb6c25a9),
	.w8(32'h3bceafa0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6b41),
	.w1(32'hbb9190f7),
	.w2(32'hbbe8d38d),
	.w3(32'h3a1d10b6),
	.w4(32'h3b397223),
	.w5(32'h3a0f9d62),
	.w6(32'h3b9a88e9),
	.w7(32'hbb81057f),
	.w8(32'h39ce154a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d90cd8),
	.w1(32'hbbcada2a),
	.w2(32'hbbf60ba7),
	.w3(32'hbb0b4404),
	.w4(32'hbba0ed1c),
	.w5(32'hbaa34665),
	.w6(32'hb8bce603),
	.w7(32'hbbd2677f),
	.w8(32'h3bf3c7ae),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75dd3e),
	.w1(32'h3bf24c93),
	.w2(32'h3c024605),
	.w3(32'hbac2392e),
	.w4(32'hb8487753),
	.w5(32'h3a6e353f),
	.w6(32'hba8697e8),
	.w7(32'h3b594b83),
	.w8(32'hbb470a2b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b419fbb),
	.w1(32'h3ab984aa),
	.w2(32'hb8db1d7c),
	.w3(32'h3bbe4d24),
	.w4(32'h3b242b91),
	.w5(32'h3a764fc5),
	.w6(32'h3bb899ae),
	.w7(32'h3b9f732d),
	.w8(32'hbc2cefdf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae0e9c),
	.w1(32'hbbef1f7f),
	.w2(32'hbc082b1c),
	.w3(32'h3c0fdc2a),
	.w4(32'h3b9e9149),
	.w5(32'hbbb590fc),
	.w6(32'hbc18b74c),
	.w7(32'hbb531fbe),
	.w8(32'h3bef966a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001b79),
	.w1(32'hb8c86ae3),
	.w2(32'h3b146484),
	.w3(32'hbc552d47),
	.w4(32'hbc18a040),
	.w5(32'h37e42ecf),
	.w6(32'h3a9ee8e9),
	.w7(32'hbaa88b71),
	.w8(32'hbbbc5d94),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c99f4),
	.w1(32'hbb9ca1c1),
	.w2(32'hbb9bcc19),
	.w3(32'hbb687eec),
	.w4(32'hb9f80d4d),
	.w5(32'hbbbf9ba4),
	.w6(32'hbc5bc918),
	.w7(32'hbaaf497d),
	.w8(32'hbc3cf924),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1709d0),
	.w1(32'hba9a4a99),
	.w2(32'hbba7401a),
	.w3(32'h39793283),
	.w4(32'hbb17a074),
	.w5(32'hbb319293),
	.w6(32'hbabb3cdf),
	.w7(32'hbaa98f94),
	.w8(32'h3a5cc2cb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08abe9),
	.w1(32'hbb51691f),
	.w2(32'h3b195ff2),
	.w3(32'hbb2182a5),
	.w4(32'hb98f8f35),
	.w5(32'h3c6abe45),
	.w6(32'h3c143f7f),
	.w7(32'hbaddc4e8),
	.w8(32'h3a5dfb90),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa8cd),
	.w1(32'hbb5e637d),
	.w2(32'hbbca641c),
	.w3(32'h3b592028),
	.w4(32'hbb3f32d9),
	.w5(32'hbbca0884),
	.w6(32'hbbbfd24b),
	.w7(32'hbb8ff9ff),
	.w8(32'hbb1fa0a9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9782a3),
	.w1(32'hbb265881),
	.w2(32'hbbe45b9e),
	.w3(32'hbbf97346),
	.w4(32'hbb5e66c3),
	.w5(32'hbb2a10ba),
	.w6(32'hbbda9930),
	.w7(32'hbc16daed),
	.w8(32'hbb33c3b0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9e28),
	.w1(32'hbc020e9f),
	.w2(32'hbbf09ce6),
	.w3(32'hbba0dfb9),
	.w4(32'h3ba43a89),
	.w5(32'hbbbf802e),
	.w6(32'h3bb10624),
	.w7(32'hbb65446b),
	.w8(32'hbb47d13e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373a56),
	.w1(32'hb96c8a53),
	.w2(32'hbb5b9b94),
	.w3(32'hbafca204),
	.w4(32'hbbf756bd),
	.w5(32'h3c09d787),
	.w6(32'hbac45784),
	.w7(32'hbbba5985),
	.w8(32'h3c0fa0c0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fb78e),
	.w1(32'h3c194d2d),
	.w2(32'h3b9c6cea),
	.w3(32'h3c88bd47),
	.w4(32'h3c042373),
	.w5(32'h3b6f4c93),
	.w6(32'h3ba4ab58),
	.w7(32'h3c1d8d90),
	.w8(32'hbb768f42),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6227d9),
	.w1(32'h3bb28a6b),
	.w2(32'hbb313da2),
	.w3(32'h3ab3dab5),
	.w4(32'h3b35df0c),
	.w5(32'h3baa550f),
	.w6(32'hbbda627a),
	.w7(32'h3a78ed01),
	.w8(32'h3b50af81),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391188e5),
	.w1(32'hbbe998f3),
	.w2(32'hbb455942),
	.w3(32'h3aef0156),
	.w4(32'h3a5cab02),
	.w5(32'h3b49aa4a),
	.w6(32'h3c2faba4),
	.w7(32'hbb4547ac),
	.w8(32'hbb66d835),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae447ea),
	.w1(32'hbb161329),
	.w2(32'h3c5c663c),
	.w3(32'h3c2a325d),
	.w4(32'h3ca8e332),
	.w5(32'h3bc91e7d),
	.w6(32'hbbfce44d),
	.w7(32'h3c381cef),
	.w8(32'h3c92a272),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fce85),
	.w1(32'hbbeb174e),
	.w2(32'hbbe815f6),
	.w3(32'hba1b462e),
	.w4(32'h3a81728b),
	.w5(32'hbb81ab5c),
	.w6(32'h3ca0069d),
	.w7(32'hbc2ce662),
	.w8(32'hbc1e639a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb62c6c),
	.w1(32'h38a1a949),
	.w2(32'hbb34ad07),
	.w3(32'h3bbc8b0b),
	.w4(32'h3becc78a),
	.w5(32'hbc32cc4a),
	.w6(32'hbbc5ff46),
	.w7(32'hba9f9922),
	.w8(32'hbc4d3f28),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28e1f5),
	.w1(32'hbc77c55f),
	.w2(32'hbc8e7ba6),
	.w3(32'hbbdb9079),
	.w4(32'hbc05183b),
	.w5(32'hbbf9da7f),
	.w6(32'hbb89d503),
	.w7(32'hbc74f9b0),
	.w8(32'hbc10292f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab5f13),
	.w1(32'hbc2b28ac),
	.w2(32'hbc04b6e2),
	.w3(32'hbc275404),
	.w4(32'hbc0ecccb),
	.w5(32'hbc19c57f),
	.w6(32'hbba0ff27),
	.w7(32'hbc050108),
	.w8(32'hbbd09bc9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea4143),
	.w1(32'hbbbd3865),
	.w2(32'hbb9604af),
	.w3(32'hbc258938),
	.w4(32'hbbd64e13),
	.w5(32'hbc0007e9),
	.w6(32'hbc54a9e0),
	.w7(32'hbc01b6f5),
	.w8(32'hbb9df09b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a0c4c),
	.w1(32'hbb247af7),
	.w2(32'hbc047715),
	.w3(32'h3b6b1b05),
	.w4(32'h3b4f6db4),
	.w5(32'h3b594571),
	.w6(32'h3c047cf2),
	.w7(32'hbb288ca7),
	.w8(32'h3a821c31),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d85d5),
	.w1(32'h3af04235),
	.w2(32'h39b38120),
	.w3(32'h39a80283),
	.w4(32'h39f6ff89),
	.w5(32'h3bb7f63c),
	.w6(32'hba13dfcc),
	.w7(32'hbb0e1eb0),
	.w8(32'h3ba6be70),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaee04),
	.w1(32'h3ac53ec4),
	.w2(32'hbada2b58),
	.w3(32'hbb8b39e3),
	.w4(32'h39bdfb01),
	.w5(32'hbc86a3ec),
	.w6(32'hbc763454),
	.w7(32'h3ab6365e),
	.w8(32'hbc149e89),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc541936),
	.w1(32'hbc8a2a83),
	.w2(32'hbc9c821f),
	.w3(32'hbc852bf4),
	.w4(32'hbc058bc3),
	.w5(32'hba9d93e7),
	.w6(32'hbc859d6f),
	.w7(32'hbca79e20),
	.w8(32'hbbd97f3b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70278c),
	.w1(32'h3ae93600),
	.w2(32'hbc08a5c5),
	.w3(32'hbb0e3433),
	.w4(32'h3b1789dd),
	.w5(32'h3a838f73),
	.w6(32'hbaf2aa34),
	.w7(32'h3a1072f0),
	.w8(32'hbba7b4cb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95fb85),
	.w1(32'hbc022865),
	.w2(32'hbbed25b0),
	.w3(32'hbc0e5e60),
	.w4(32'h3c048850),
	.w5(32'hbbc3f7b6),
	.w6(32'hbc8ace7f),
	.w7(32'h3c0b0cd7),
	.w8(32'hbb6e20f6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad78afe),
	.w1(32'hbaf5933a),
	.w2(32'h3a6ed563),
	.w3(32'hb9ddcfb5),
	.w4(32'hbb02ddab),
	.w5(32'hbb276d62),
	.w6(32'h3a862898),
	.w7(32'hb80c20b7),
	.w8(32'h3bbaedb3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e45e73),
	.w1(32'h3ac264b4),
	.w2(32'hbae4ae49),
	.w3(32'hba8fd223),
	.w4(32'hbb494718),
	.w5(32'h3a8dac7a),
	.w6(32'h3b21863d),
	.w7(32'hbb7a6377),
	.w8(32'h3b90c0ab),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faa0a),
	.w1(32'h3bae0bfe),
	.w2(32'hbad9c8b3),
	.w3(32'h3af83ce4),
	.w4(32'h3a9e3a01),
	.w5(32'hba7d87ec),
	.w6(32'h3b493bbb),
	.w7(32'hbaa789ed),
	.w8(32'hbc093eb3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31f31f),
	.w1(32'h39b5a89d),
	.w2(32'h3b98b0e9),
	.w3(32'h3c1cde2e),
	.w4(32'h3c3d385e),
	.w5(32'h3adaf8e1),
	.w6(32'h3c0219ed),
	.w7(32'h3c449ec8),
	.w8(32'hba60db0c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b483a39),
	.w1(32'h3a024838),
	.w2(32'h391b8d94),
	.w3(32'hba979a73),
	.w4(32'hbaa57f9f),
	.w5(32'h3a2d68ae),
	.w6(32'h3b4dc344),
	.w7(32'hbad3f05d),
	.w8(32'h3c5cc21e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96201f),
	.w1(32'h3b8d5e5b),
	.w2(32'h3b8fe893),
	.w3(32'hbaab7607),
	.w4(32'hb8ce9a84),
	.w5(32'hba9f87a2),
	.w6(32'h3c777165),
	.w7(32'h3c05aab4),
	.w8(32'hb988adfe),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb561ab0),
	.w1(32'hbad97de8),
	.w2(32'hbb8ca4af),
	.w3(32'h3b729043),
	.w4(32'hbaeaddcc),
	.w5(32'hbb13f92f),
	.w6(32'h3b51928c),
	.w7(32'hbb95bb2f),
	.w8(32'h3b00c4a6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392da343),
	.w1(32'hbbb8cc59),
	.w2(32'hbaf497d7),
	.w3(32'hba5ccdc0),
	.w4(32'hba420c74),
	.w5(32'hbbee78df),
	.w6(32'h3c255079),
	.w7(32'hbba9dfc2),
	.w8(32'h3bb856e5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53a66f),
	.w1(32'h39c1cf0b),
	.w2(32'hba402f02),
	.w3(32'hbc3bd6b5),
	.w4(32'hb91e1df9),
	.w5(32'h3b08c9dd),
	.w6(32'hbb1a5b28),
	.w7(32'h3ba3da1b),
	.w8(32'hb9f36660),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389666e3),
	.w1(32'h3b17b856),
	.w2(32'hbb96e1fc),
	.w3(32'hba2cad1d),
	.w4(32'hbb719316),
	.w5(32'h3b8d5ad1),
	.w6(32'h3b26a352),
	.w7(32'hbc2f2c07),
	.w8(32'h3b6ab328),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37711e),
	.w1(32'hb87d3c09),
	.w2(32'h3bdf85f8),
	.w3(32'h3a7c7c1e),
	.w4(32'h3ac36dd7),
	.w5(32'hbaa67a86),
	.w6(32'h3adceee9),
	.w7(32'hb91ebae0),
	.w8(32'hbb319f4f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48604),
	.w1(32'hba9f3ba5),
	.w2(32'h3a42476b),
	.w3(32'hbb55a236),
	.w4(32'h3af288d3),
	.w5(32'hbbdafde5),
	.w6(32'hbc13eeb6),
	.w7(32'h3b97b0be),
	.w8(32'hbb633730),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcef9c3),
	.w1(32'hbb71301e),
	.w2(32'hbc0c0210),
	.w3(32'hb617da3c),
	.w4(32'hbb674751),
	.w5(32'hbc3eb4ff),
	.w6(32'h3c028d40),
	.w7(32'hbbc8b5d4),
	.w8(32'hbc8254e7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb972509),
	.w1(32'hbb2b2447),
	.w2(32'hbbf0f880),
	.w3(32'h3aec9082),
	.w4(32'hba5ce3f6),
	.w5(32'hbb1276a7),
	.w6(32'h3b5c01cb),
	.w7(32'hbc06ff53),
	.w8(32'h3aa9b77d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b97a6),
	.w1(32'hbb1bde3b),
	.w2(32'hba130b39),
	.w3(32'hbb895862),
	.w4(32'h3a5ba408),
	.w5(32'h3c1eb886),
	.w6(32'hbba11e42),
	.w7(32'hbb2a78aa),
	.w8(32'h3c68d27c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4719d0),
	.w1(32'hbc061826),
	.w2(32'hbc4b7ace),
	.w3(32'h3c604018),
	.w4(32'h3c125400),
	.w5(32'h3a9a8789),
	.w6(32'h3ce96610),
	.w7(32'h3a7cdc6a),
	.w8(32'hba93928a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d6054),
	.w1(32'hba6784e1),
	.w2(32'h3a3d1934),
	.w3(32'h3bc5592e),
	.w4(32'h3be42a1c),
	.w5(32'hbb2fbd2e),
	.w6(32'hbbd6a1e3),
	.w7(32'hbb4e17d1),
	.w8(32'hbbd1298f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65d1c5),
	.w1(32'h3b871a94),
	.w2(32'hbbce10ad),
	.w3(32'h3993d348),
	.w4(32'hbbda4917),
	.w5(32'hbc048341),
	.w6(32'h3bf7e985),
	.w7(32'hbb9796de),
	.w8(32'hbbb4465f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462941),
	.w1(32'hbbddc60f),
	.w2(32'hbc21aaf2),
	.w3(32'hbbeb697b),
	.w4(32'hbc2bdd31),
	.w5(32'h3b2e332c),
	.w6(32'h3bafa38e),
	.w7(32'hbbc9a2d8),
	.w8(32'hbbcc56d8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2294ca),
	.w1(32'hbaa79d41),
	.w2(32'h3ba8adf0),
	.w3(32'h3bafffa3),
	.w4(32'h3bae5077),
	.w5(32'hbba32a1c),
	.w6(32'hbbb46956),
	.w7(32'hbaa8392e),
	.w8(32'hbad7b459),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907eed),
	.w1(32'hbbd88b9a),
	.w2(32'hbbbfe914),
	.w3(32'hba3578ef),
	.w4(32'hbb02b42d),
	.w5(32'h3aa08f53),
	.w6(32'h3c10f70e),
	.w7(32'hbb9227eb),
	.w8(32'h391831a6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf99aa),
	.w1(32'h3b6abad2),
	.w2(32'hbbb36fcc),
	.w3(32'h3bcf9a34),
	.w4(32'h39401816),
	.w5(32'h392358a5),
	.w6(32'h3bc00e45),
	.w7(32'h3c13f79b),
	.w8(32'hbb8b6326),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39c849),
	.w1(32'h3aaf20a7),
	.w2(32'hbba21115),
	.w3(32'hbb5b6707),
	.w4(32'hbb916fbb),
	.w5(32'hbc2298fb),
	.w6(32'hbba0a279),
	.w7(32'hb9c3c62a),
	.w8(32'hbbd4a48b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1712a),
	.w1(32'hbc4a18df),
	.w2(32'hbc5b09b5),
	.w3(32'h3ab94cb5),
	.w4(32'hbb07d416),
	.w5(32'hbbe1b3e4),
	.w6(32'hbbbaedab),
	.w7(32'hbbd73f22),
	.w8(32'hbbfce3e9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fc1e7),
	.w1(32'h3c47cd69),
	.w2(32'h3b991255),
	.w3(32'h3bb16eb8),
	.w4(32'h3c22e8f8),
	.w5(32'hbc51ad70),
	.w6(32'h3c022934),
	.w7(32'h3c929509),
	.w8(32'hbc14f1a7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f54b9),
	.w1(32'hbbfa6aaa),
	.w2(32'hbc2ba6f8),
	.w3(32'hbc010834),
	.w4(32'hbbd922c8),
	.w5(32'h3c010cc3),
	.w6(32'h3b0154a7),
	.w7(32'hbc3fa196),
	.w8(32'hbb31af06),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc46bb2),
	.w1(32'h3c6eb09c),
	.w2(32'h3b86688a),
	.w3(32'h3c833add),
	.w4(32'h3c9fcdcf),
	.w5(32'h3baff3cb),
	.w6(32'hba2dbf12),
	.w7(32'h3c8d92d5),
	.w8(32'hbb788497),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa535),
	.w1(32'hbadca12c),
	.w2(32'hbb3ea076),
	.w3(32'h3c6de086),
	.w4(32'h3c244d9a),
	.w5(32'hbac1b4ea),
	.w6(32'hbaaba56d),
	.w7(32'h3bf55bbe),
	.w8(32'hbb83ce9a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fdc51),
	.w1(32'hbb14f664),
	.w2(32'h3b1ec900),
	.w3(32'h3b55859d),
	.w4(32'h3b525a1f),
	.w5(32'h3a892457),
	.w6(32'hbbc92fea),
	.w7(32'hbb67b22b),
	.w8(32'h3bcf3c5b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c728c),
	.w1(32'h3c4df694),
	.w2(32'h3ba3fa73),
	.w3(32'h3c34dce1),
	.w4(32'hb9831a41),
	.w5(32'h3a9bc18e),
	.w6(32'h3cc01296),
	.w7(32'h3bcc432e),
	.w8(32'h395edea6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e483f),
	.w1(32'hbbade768),
	.w2(32'hbc1ae831),
	.w3(32'h3b3ea097),
	.w4(32'h3b1aadd3),
	.w5(32'hbb7407ff),
	.w6(32'hbbf29763),
	.w7(32'hbb36aa46),
	.w8(32'h3a9d5380),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e4ee4),
	.w1(32'hbb0afcb7),
	.w2(32'hbc0d8703),
	.w3(32'hb9a36e92),
	.w4(32'h3a44eeb6),
	.w5(32'hbb0ecd68),
	.w6(32'h3c34d29d),
	.w7(32'hbc07e45d),
	.w8(32'hbbe52823),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f560),
	.w1(32'hbb3ae3ac),
	.w2(32'hbbb79046),
	.w3(32'hbc195aa4),
	.w4(32'h3a259e7f),
	.w5(32'hbbb0988f),
	.w6(32'h3acd0ea7),
	.w7(32'hba26b501),
	.w8(32'h3a94d1ed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67d5e),
	.w1(32'hba1e80bd),
	.w2(32'h3b9bf979),
	.w3(32'hbb638a28),
	.w4(32'hbb3e30b9),
	.w5(32'hbbde1acb),
	.w6(32'hba3e3a1b),
	.w7(32'hbaa63f2c),
	.w8(32'hbb956eae),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc212c3f),
	.w1(32'hbc2e835f),
	.w2(32'hbc392d45),
	.w3(32'hbb2b91a1),
	.w4(32'hbb68e875),
	.w5(32'hba5d57ce),
	.w6(32'h3a009751),
	.w7(32'hbbf008db),
	.w8(32'hbab3be26),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88cb5b),
	.w1(32'hbb4987cd),
	.w2(32'hbadb52b9),
	.w3(32'hbbd7b188),
	.w4(32'hbba6579a),
	.w5(32'h39990c33),
	.w6(32'h3c039751),
	.w7(32'hbbcbd161),
	.w8(32'h3b29896f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b071fa0),
	.w1(32'h39dc155b),
	.w2(32'h3c21a8be),
	.w3(32'hbb82dcad),
	.w4(32'h3bb948f9),
	.w5(32'h39b89a2d),
	.w6(32'h3a4afed9),
	.w7(32'h3bc745e6),
	.w8(32'hba61e22a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84be94),
	.w1(32'hb9892121),
	.w2(32'h3ba478c7),
	.w3(32'h3a0ab56a),
	.w4(32'h3b57f7ee),
	.w5(32'hbb9a4a98),
	.w6(32'h3b89e77f),
	.w7(32'h3b912b00),
	.w8(32'h3bfa0fb6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c029aff),
	.w1(32'h3ba30f44),
	.w2(32'hba6bf833),
	.w3(32'hbc190912),
	.w4(32'hbb8e740a),
	.w5(32'h3ab9c201),
	.w6(32'hbbddc8b1),
	.w7(32'hbbe17879),
	.w8(32'hbbb69cdd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077721),
	.w1(32'h3a371f29),
	.w2(32'hbbb43817),
	.w3(32'hba059c51),
	.w4(32'hbb5cc30b),
	.w5(32'h3b17d5fe),
	.w6(32'h3a0320cb),
	.w7(32'hbba87af2),
	.w8(32'h3ad07d15),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acea635),
	.w1(32'hbb22fb93),
	.w2(32'hb9cd09eb),
	.w3(32'h3bc47793),
	.w4(32'h3b834c4e),
	.w5(32'hbc07452b),
	.w6(32'h3c02d45e),
	.w7(32'h39a11e0b),
	.w8(32'hbb4e4375),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcc4fa),
	.w1(32'hbbe67093),
	.w2(32'h39d75ecf),
	.w3(32'hbc123ff1),
	.w4(32'hbba0275a),
	.w5(32'h3c130f97),
	.w6(32'h3c582d22),
	.w7(32'h3b9ca335),
	.w8(32'h3c097257),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7dbd6),
	.w1(32'h3c752af1),
	.w2(32'h3c453ff7),
	.w3(32'h3c8020ba),
	.w4(32'h3c4b42f2),
	.w5(32'hbaf3a64e),
	.w6(32'h3ba0e6f2),
	.w7(32'h3c94882b),
	.w8(32'h3b0885f5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0893d),
	.w1(32'hbbda4ce8),
	.w2(32'hbba1bd7e),
	.w3(32'hbc219a8e),
	.w4(32'hbbd5620f),
	.w5(32'h3b6306e3),
	.w6(32'hbc51e888),
	.w7(32'hbacc77b9),
	.w8(32'h3bb24016),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1470eb),
	.w1(32'h3c0cf43a),
	.w2(32'h3af3d94c),
	.w3(32'h3c216b87),
	.w4(32'h3b302fbb),
	.w5(32'hbbb7e6eb),
	.w6(32'h3c233e38),
	.w7(32'h3b533e31),
	.w8(32'hbb86777d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf1e45),
	.w1(32'hbc2f259c),
	.w2(32'hbc06d6f6),
	.w3(32'hbb57c827),
	.w4(32'hbb2a29f1),
	.w5(32'hba7811e3),
	.w6(32'hbbb6444a),
	.w7(32'hbb9370de),
	.w8(32'hba3c8346),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99683a),
	.w1(32'h3b6f16ad),
	.w2(32'hbac7a96b),
	.w3(32'hbb24cd90),
	.w4(32'h3bfa77a9),
	.w5(32'h3b8ffc03),
	.w6(32'h3b299b41),
	.w7(32'h3bfdfeca),
	.w8(32'h3a8fc01b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183bde),
	.w1(32'h39dfe9a8),
	.w2(32'hbc3bd7ab),
	.w3(32'h398a59e6),
	.w4(32'h3ae677bf),
	.w5(32'hbbbb0f72),
	.w6(32'h3b75eec9),
	.w7(32'hb9b3c584),
	.w8(32'hbb5a1a7e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9475d),
	.w1(32'hbb352df9),
	.w2(32'hbb0a2dbf),
	.w3(32'hbabceab1),
	.w4(32'h3a61cdee),
	.w5(32'hbbd11cd7),
	.w6(32'hba809f91),
	.w7(32'h3aee2576),
	.w8(32'hbc059b12),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e01e),
	.w1(32'hbb9d67a5),
	.w2(32'hbb89d4ea),
	.w3(32'hbbfc572e),
	.w4(32'hbba930f4),
	.w5(32'hbbd0bdbc),
	.w6(32'hbc165ece),
	.w7(32'hbbce9670),
	.w8(32'h3a1e314d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954ce28),
	.w1(32'h3ace406d),
	.w2(32'hbb23542d),
	.w3(32'h3c1dcc82),
	.w4(32'h3b87ca7e),
	.w5(32'h3b2c3e60),
	.w6(32'h3ab0efd5),
	.w7(32'h3a93ced7),
	.w8(32'hbba321b8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e851e),
	.w1(32'hba920e8a),
	.w2(32'hb866daa6),
	.w3(32'h3aedc200),
	.w4(32'h3b8e3b9c),
	.w5(32'h3ad42604),
	.w6(32'hbb44d00b),
	.w7(32'hba643a20),
	.w8(32'hb9ae4eea),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a431dda),
	.w1(32'hbb775680),
	.w2(32'hbb02ad51),
	.w3(32'hbb748164),
	.w4(32'hbb8f0544),
	.w5(32'hbad6735a),
	.w6(32'hbba0e1ff),
	.w7(32'hbb6e5aa7),
	.w8(32'h3b71ec4d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67b143),
	.w1(32'h3b91261d),
	.w2(32'h3bd4f17c),
	.w3(32'hbbed193c),
	.w4(32'h3aea2b3b),
	.w5(32'h3ac8cf86),
	.w6(32'h3bb89618),
	.w7(32'h3bb45083),
	.w8(32'h3ab616b2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8568ef),
	.w1(32'hba9bb7f0),
	.w2(32'hbb7c3db0),
	.w3(32'hb9961291),
	.w4(32'hbb91ac1e),
	.w5(32'h3bb39ed3),
	.w6(32'hbae8b401),
	.w7(32'hbba80490),
	.w8(32'h3c0982aa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb97206),
	.w1(32'h3ca2a914),
	.w2(32'h3c62d7fd),
	.w3(32'h3c412261),
	.w4(32'h3bfc1ae4),
	.w5(32'hbc792de5),
	.w6(32'h3c977f72),
	.w7(32'h3c54d314),
	.w8(32'hbc1d81a9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1399e1),
	.w1(32'hbbd915e5),
	.w2(32'hbc6afe01),
	.w3(32'hbc059d0c),
	.w4(32'hbc2869b1),
	.w5(32'hba07506f),
	.w6(32'h3b44c381),
	.w7(32'hbc15cfc8),
	.w8(32'h39d16301),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4f1db),
	.w1(32'h3a74c8f4),
	.w2(32'hba4e0161),
	.w3(32'h38f432f2),
	.w4(32'h3af286b6),
	.w5(32'h3c08f5e6),
	.w6(32'h3a41820a),
	.w7(32'h3af88233),
	.w8(32'h3bb579b8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bc8e6),
	.w1(32'h3ae3abae),
	.w2(32'hbb303e78),
	.w3(32'h3c7f5801),
	.w4(32'h3bc0fb44),
	.w5(32'h3ba5fc52),
	.w6(32'h3ba99e36),
	.w7(32'hba790ac9),
	.w8(32'h3b351a05),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9d9b4),
	.w1(32'h3afbf562),
	.w2(32'hba7b7246),
	.w3(32'h3bd4f45a),
	.w4(32'h3be5513b),
	.w5(32'h3b84170d),
	.w6(32'h3b42e5a4),
	.w7(32'h3bcbc38e),
	.w8(32'h392fa7a1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b5285),
	.w1(32'hbb450817),
	.w2(32'hbb942269),
	.w3(32'h3ba09be0),
	.w4(32'h3b935305),
	.w5(32'hbb68e37a),
	.w6(32'hbb5db62a),
	.w7(32'hbb184be3),
	.w8(32'hbb887e87),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ff1f4),
	.w1(32'hba0ed50f),
	.w2(32'hbb581f5c),
	.w3(32'hbaa30789),
	.w4(32'h3ad7aa69),
	.w5(32'h3bcf2eb8),
	.w6(32'h3b8f09c0),
	.w7(32'hb8236ff8),
	.w8(32'h3b9539ca),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ba5f4),
	.w1(32'h3c1849d0),
	.w2(32'h3c6876bc),
	.w3(32'h3c14422d),
	.w4(32'h3c1963eb),
	.w5(32'hbb41cad6),
	.w6(32'h3ba30b8b),
	.w7(32'h3c558f77),
	.w8(32'hbb134cad),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ae28b),
	.w1(32'hbbdc05aa),
	.w2(32'hbb6345fe),
	.w3(32'hba8effbb),
	.w4(32'hbbcd076a),
	.w5(32'hbb4d3722),
	.w6(32'hb9009aaf),
	.w7(32'h3b83c290),
	.w8(32'h3b69cc0c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb605634),
	.w1(32'hbc5a3fb7),
	.w2(32'hbc3a2ed1),
	.w3(32'hbbcdbbe7),
	.w4(32'hbc3ae1e0),
	.w5(32'h3bd037de),
	.w6(32'hbb986771),
	.w7(32'hbbc0bafb),
	.w8(32'h3c2042bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c307775),
	.w1(32'h3c51d14d),
	.w2(32'h3b5f90bf),
	.w3(32'h3c668406),
	.w4(32'h3c1026ca),
	.w5(32'hbacece2b),
	.w6(32'h3c8182b8),
	.w7(32'h3bf30f26),
	.w8(32'hba41a1d8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b608a60),
	.w1(32'h3a861531),
	.w2(32'hbb3a2a88),
	.w3(32'hbb386258),
	.w4(32'h3b63a9be),
	.w5(32'h3a8a7318),
	.w6(32'hbb6158bb),
	.w7(32'hbb036748),
	.w8(32'h3ad0684e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59f8f6),
	.w1(32'hbc265ac2),
	.w2(32'hbbe96e8a),
	.w3(32'h3a1eda06),
	.w4(32'hba291702),
	.w5(32'hbbe4bbe2),
	.w6(32'hb9922c03),
	.w7(32'hba15e49b),
	.w8(32'h3a28cbe3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c83a4),
	.w1(32'h3a2ebedd),
	.w2(32'hbbbf453f),
	.w3(32'hbc8b2c22),
	.w4(32'hbc3429b2),
	.w5(32'hbbabb128),
	.w6(32'h3c714042),
	.w7(32'h3b154100),
	.w8(32'h3a237b78),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc256c2),
	.w1(32'hbb2082cf),
	.w2(32'hbbbd93fd),
	.w3(32'hba1ab312),
	.w4(32'hbb86f25a),
	.w5(32'hbc63f06d),
	.w6(32'h3b57947e),
	.w7(32'hbbbc93b4),
	.w8(32'hbbd92cf3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25fa00),
	.w1(32'h3b21e3d2),
	.w2(32'hbbceb7b3),
	.w3(32'hbca90def),
	.w4(32'hbc9386e4),
	.w5(32'hb9114b9a),
	.w6(32'h3b9bde8f),
	.w7(32'hbc32700d),
	.w8(32'hbaed72d1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880059),
	.w1(32'hbaf7d752),
	.w2(32'hbb91a4ff),
	.w3(32'hba25e854),
	.w4(32'hb9bc03ae),
	.w5(32'hbc769d67),
	.w6(32'hb986ae59),
	.w7(32'h39d09185),
	.w8(32'hbbc3b9b7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfca7c4),
	.w1(32'h3b1bf2f7),
	.w2(32'h3a8e899a),
	.w3(32'hbc8a6220),
	.w4(32'hbbb6e58a),
	.w5(32'h3b9fa6e9),
	.w6(32'h3a6bac81),
	.w7(32'h392c7852),
	.w8(32'h3b3d8d4c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e964),
	.w1(32'hbb44157c),
	.w2(32'hbb9a11e3),
	.w3(32'h3ba311b7),
	.w4(32'h3b869b9a),
	.w5(32'hbbeab9c3),
	.w6(32'h3b3c88db),
	.w7(32'h3aa03e6a),
	.w8(32'hbb11b541),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39212a),
	.w1(32'h3b1e69a2),
	.w2(32'h3a8c4901),
	.w3(32'h3b07a70c),
	.w4(32'hbb087d1a),
	.w5(32'hbca40866),
	.w6(32'h3be15493),
	.w7(32'h3b92dc08),
	.w8(32'hbc2e699a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80cf2e),
	.w1(32'hbc63ee22),
	.w2(32'hbc9ced04),
	.w3(32'hbc611fcc),
	.w4(32'hbc3c0bff),
	.w5(32'h3bf07eca),
	.w6(32'hbbd547d2),
	.w7(32'hbc6df9cd),
	.w8(32'hbbee2ea3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53ab3e),
	.w1(32'h39ac2563),
	.w2(32'hbaff2c56),
	.w3(32'h3a7a9d34),
	.w4(32'h3b858cf7),
	.w5(32'hbc387df0),
	.w6(32'hbabf29b7),
	.w7(32'hba910c7d),
	.w8(32'hbc417d28),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff2d3e),
	.w1(32'hbc0e17f2),
	.w2(32'hbbfd610d),
	.w3(32'hbc2b73b2),
	.w4(32'hbc3039cb),
	.w5(32'h3b86bb80),
	.w6(32'hbc36e634),
	.w7(32'hbc21b046),
	.w8(32'hbbc5a91c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b30719),
	.w1(32'hbaaf61a1),
	.w2(32'hbba91b75),
	.w3(32'h3b2be3e2),
	.w4(32'h3c0e6e55),
	.w5(32'hbaf10dbc),
	.w6(32'h3b20c3b6),
	.w7(32'hbb57be09),
	.w8(32'h3a4033f8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be70be6),
	.w1(32'h3b27e2b0),
	.w2(32'h3b1e0de3),
	.w3(32'h38985138),
	.w4(32'h3b6148ca),
	.w5(32'hbc49080f),
	.w6(32'h3b97c4c1),
	.w7(32'h3b799508),
	.w8(32'hbc05911f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9336a),
	.w1(32'hbb494053),
	.w2(32'hbbe2b51a),
	.w3(32'hbbd92312),
	.w4(32'hbc00ee45),
	.w5(32'h3b6cfaa9),
	.w6(32'h3b2ecbe7),
	.w7(32'hbb9775a2),
	.w8(32'h3a216114),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a045),
	.w1(32'hb9e175a6),
	.w2(32'h3b91389b),
	.w3(32'h3c0b2cf2),
	.w4(32'h3c01d620),
	.w5(32'hbb9f6678),
	.w6(32'h3b0759c3),
	.w7(32'h3c229f3b),
	.w8(32'hbbcd94a0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab6dc6),
	.w1(32'h3a464c26),
	.w2(32'h395fd8fc),
	.w3(32'h3bd78423),
	.w4(32'h3a4d3c20),
	.w5(32'h3b06a1cb),
	.w6(32'h3b7348e4),
	.w7(32'h3b5631cd),
	.w8(32'h3b90cc1b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c451d7c),
	.w1(32'h3bc2a0e7),
	.w2(32'h3bc67184),
	.w3(32'h3b43acc1),
	.w4(32'h3b8a98e5),
	.w5(32'hbbc883a9),
	.w6(32'h3c026142),
	.w7(32'h3b81f60f),
	.w8(32'hbbd7777a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae26234),
	.w1(32'hbb7e28bd),
	.w2(32'hbb349cde),
	.w3(32'hbb9a9d70),
	.w4(32'hbb05afe6),
	.w5(32'h3b9068c0),
	.w6(32'hba83c6c2),
	.w7(32'hb90c66d8),
	.w8(32'h3c07c677),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1010),
	.w1(32'hbb010c1c),
	.w2(32'hbb21ad0a),
	.w3(32'h3acce37a),
	.w4(32'h3b8dba0b),
	.w5(32'h3bf60381),
	.w6(32'h3b9b37bd),
	.w7(32'h399a7bda),
	.w8(32'h3b775bac),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b321),
	.w1(32'h3c27f4ee),
	.w2(32'h3c3ee432),
	.w3(32'h3be4dbef),
	.w4(32'h3c6155cd),
	.w5(32'hbb5e8b58),
	.w6(32'hbbaf7f84),
	.w7(32'h3c05dee1),
	.w8(32'hbb9ea8cc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3130d4),
	.w1(32'hbad6861f),
	.w2(32'hba7b2edc),
	.w3(32'hbae3c88f),
	.w4(32'h3828914f),
	.w5(32'hbc8a683c),
	.w6(32'hbb77d1c1),
	.w7(32'hbb3237fa),
	.w8(32'hbc821fe9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6027ad),
	.w1(32'hbc39f8f5),
	.w2(32'hbc6da2ee),
	.w3(32'hbc68897f),
	.w4(32'hbc7c702f),
	.w5(32'h3a9da677),
	.w6(32'hbbcbf3f6),
	.w7(32'hbc7dc59e),
	.w8(32'hb9fbcbd3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9a43),
	.w1(32'hbaaa107e),
	.w2(32'hbaf04658),
	.w3(32'h3b38387f),
	.w4(32'hb9dec548),
	.w5(32'hbc22bba0),
	.w6(32'h3be4bb6a),
	.w7(32'h39cab5fa),
	.w8(32'hbb13b6a7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f7977),
	.w1(32'hbb3225db),
	.w2(32'hbb80dd07),
	.w3(32'hbc17d2a7),
	.w4(32'hbba0b68d),
	.w5(32'hbaa2c48d),
	.w6(32'hbaec47af),
	.w7(32'hb9863f01),
	.w8(32'hbb1d9368),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530b12),
	.w1(32'hbb129b82),
	.w2(32'hbb4a1245),
	.w3(32'hbaa62f8b),
	.w4(32'hba8a9746),
	.w5(32'hbbccb94a),
	.w6(32'hbaf129c3),
	.w7(32'hbb2b86f3),
	.w8(32'hbb02f16f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5c0cd),
	.w1(32'hbb8b7bfb),
	.w2(32'hbbeb9dfc),
	.w3(32'hbb457930),
	.w4(32'hbbadd2cf),
	.w5(32'h3a231df3),
	.w6(32'hbb254bfb),
	.w7(32'hba05e8f9),
	.w8(32'h3a80d8a4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1735c8),
	.w1(32'hbb256c78),
	.w2(32'hbbeb1649),
	.w3(32'hbac0056a),
	.w4(32'h390ced79),
	.w5(32'hbb010fb2),
	.w6(32'hbba652ec),
	.w7(32'hbb901543),
	.w8(32'hbbd3d524),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb879cc6),
	.w1(32'hbb943a74),
	.w2(32'hbb8e9eb8),
	.w3(32'h3bfd8d6b),
	.w4(32'h38800b23),
	.w5(32'hba8082cb),
	.w6(32'h3bb46e2d),
	.w7(32'hbb171aef),
	.w8(32'h3b573f1b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842862),
	.w1(32'h3bbca13d),
	.w2(32'h3bbdfca8),
	.w3(32'hba4a299b),
	.w4(32'h3b151db6),
	.w5(32'hbb5c8f5b),
	.w6(32'hb9802dfd),
	.w7(32'h3b9c6ecf),
	.w8(32'hbb7dc881),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb482d82),
	.w1(32'hbb744e5d),
	.w2(32'hbb0e291f),
	.w3(32'hb82d3e76),
	.w4(32'h3b393215),
	.w5(32'hbb7a0f93),
	.w6(32'hbb929dac),
	.w7(32'h3a62fd23),
	.w8(32'hbc2573d1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc7fec),
	.w1(32'hba741ae7),
	.w2(32'hbb9316cd),
	.w3(32'h3a9dc014),
	.w4(32'hbb231cac),
	.w5(32'hbb498b2b),
	.w6(32'h3b72e1c2),
	.w7(32'hbafcde5d),
	.w8(32'hbb9224a1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc95ac8),
	.w1(32'h3bb7815c),
	.w2(32'hba8cf608),
	.w3(32'hba4f9706),
	.w4(32'h3afc9387),
	.w5(32'hbc1eea6e),
	.w6(32'h3b8cf5dd),
	.w7(32'h3ba14212),
	.w8(32'hbb74a4f5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bad384),
	.w1(32'h3b3ba037),
	.w2(32'h3b6c981d),
	.w3(32'hbb0efbde),
	.w4(32'hbb85f873),
	.w5(32'hbbba3650),
	.w6(32'h3bbe6da5),
	.w7(32'hbb4258be),
	.w8(32'hbb8da0c2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a5d5c),
	.w1(32'hbb02f171),
	.w2(32'hbba51e54),
	.w3(32'hbb2b8d41),
	.w4(32'hbbd59de4),
	.w5(32'hb9cd622d),
	.w6(32'hba4d5f9d),
	.w7(32'hbb8661cd),
	.w8(32'h3bc70b02),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3afe8d),
	.w1(32'h3c655403),
	.w2(32'h3c1ac3e4),
	.w3(32'h3b9a418d),
	.w4(32'h3b4d8088),
	.w5(32'hbbea394e),
	.w6(32'h3c4672db),
	.w7(32'h3c1d8311),
	.w8(32'hbbf3618e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaee86),
	.w1(32'hbadc56a8),
	.w2(32'hbb31b2bc),
	.w3(32'hb98268ca),
	.w4(32'hbb1a93d3),
	.w5(32'h3ac0ac63),
	.w6(32'h3a164ad8),
	.w7(32'hbae0c21e),
	.w8(32'h3b31c786),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdf3c9),
	.w1(32'hbb3f6909),
	.w2(32'hbb534d0e),
	.w3(32'h3a0160e0),
	.w4(32'h3b6db51e),
	.w5(32'h3c3a9d28),
	.w6(32'h3b823f16),
	.w7(32'h3a5b6eb5),
	.w8(32'h3b902910),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdcdd2),
	.w1(32'h3c3d091c),
	.w2(32'h3c0ac2ba),
	.w3(32'hba6de85a),
	.w4(32'h3baab33d),
	.w5(32'h3c917fea),
	.w6(32'h3c58dd3c),
	.w7(32'h3bb57fa0),
	.w8(32'h3c83e53e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019256),
	.w1(32'h3ba4fc55),
	.w2(32'h3c2503f8),
	.w3(32'h3ca2dcb4),
	.w4(32'h3c8793c0),
	.w5(32'h3b21ae8c),
	.w6(32'h3c4f9121),
	.w7(32'h3c702de2),
	.w8(32'h3af40114),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393620e4),
	.w1(32'hbbf3addc),
	.w2(32'hbbb7f18a),
	.w3(32'h3ba15d08),
	.w4(32'h39c15df7),
	.w5(32'h3bf02b5a),
	.w6(32'hbba7a275),
	.w7(32'hbb06b310),
	.w8(32'h3b2b78a8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba969b97),
	.w1(32'hbb59ea3c),
	.w2(32'hbb677bda),
	.w3(32'h39b841ec),
	.w4(32'h3bbf2af1),
	.w5(32'h3b238719),
	.w6(32'hb7b6d950),
	.w7(32'hbaa6be08),
	.w8(32'hba9a98b4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dfe72),
	.w1(32'h3b01e7ca),
	.w2(32'hbb1b4193),
	.w3(32'h3abe56a2),
	.w4(32'h3b4b5364),
	.w5(32'hbb0dc9cc),
	.w6(32'hba76e1cc),
	.w7(32'hbac5d84f),
	.w8(32'hbbd7f778),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7431),
	.w1(32'hbb90a63b),
	.w2(32'hba67f8dd),
	.w3(32'hbb964ace),
	.w4(32'h37979e61),
	.w5(32'h3bcb9d12),
	.w6(32'hbb3999c1),
	.w7(32'h3b807733),
	.w8(32'hbbc4f084),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfafca),
	.w1(32'h3aaecfb5),
	.w2(32'hbb14ff26),
	.w3(32'h3c12e919),
	.w4(32'h3b6e2aa5),
	.w5(32'hbbd8380c),
	.w6(32'hbb6087c2),
	.w7(32'hbad46ee4),
	.w8(32'hbb5d048a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b8ff),
	.w1(32'h3c3bd7ca),
	.w2(32'h39a69024),
	.w3(32'h3cba22f8),
	.w4(32'h3be28bb4),
	.w5(32'hbc58fda9),
	.w6(32'h3c9d088f),
	.w7(32'h3aa9681a),
	.w8(32'hbb9ae5b7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeeef0),
	.w1(32'h3b5956f6),
	.w2(32'hbb2681fa),
	.w3(32'hbc95190b),
	.w4(32'hbc42518e),
	.w5(32'hbbc9cc1a),
	.w6(32'h3c158cba),
	.w7(32'hbb015e1a),
	.w8(32'hbb58d897),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff94b),
	.w1(32'hbb2a0c97),
	.w2(32'hba4921fd),
	.w3(32'hbb9e6764),
	.w4(32'h3ad2b0f1),
	.w5(32'h39792175),
	.w6(32'hbb0be03d),
	.w7(32'h3b326529),
	.w8(32'h3a05a899),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e6a8a),
	.w1(32'hbaf91b49),
	.w2(32'hbb25b442),
	.w3(32'h3b170554),
	.w4(32'h3b876214),
	.w5(32'hbc749b92),
	.w6(32'hbb335584),
	.w7(32'h3a27bf39),
	.w8(32'hbbd1cbe6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39fdaa),
	.w1(32'hba21153b),
	.w2(32'h3b47d121),
	.w3(32'hbbdf5c2c),
	.w4(32'hbb06b359),
	.w5(32'h3b824906),
	.w6(32'h3bb13f51),
	.w7(32'h3b180a1c),
	.w8(32'h3b9d31b7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20079a),
	.w1(32'h3c0d2e63),
	.w2(32'h3bce3b38),
	.w3(32'h3ca1f94a),
	.w4(32'h3c28027a),
	.w5(32'hbbf321e4),
	.w6(32'h3c362a01),
	.w7(32'h3c27c25f),
	.w8(32'hbc2324ec),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaab05),
	.w1(32'hbc1a2d39),
	.w2(32'hbc12f62b),
	.w3(32'hbbd4767a),
	.w4(32'hbbdbd69f),
	.w5(32'hbba0a4b9),
	.w6(32'hbabe835f),
	.w7(32'hbb90d296),
	.w8(32'hbb932efd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b4b9d),
	.w1(32'hba964d8e),
	.w2(32'h384714c5),
	.w3(32'hbb9a4d6e),
	.w4(32'hbbb985c8),
	.w5(32'hbbc59879),
	.w6(32'hbbba1c88),
	.w7(32'hbb98a409),
	.w8(32'h3bf880fd),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6da95c),
	.w1(32'h3c5d15f4),
	.w2(32'h3c1c3c87),
	.w3(32'hbcb412e6),
	.w4(32'hbaa8fc25),
	.w5(32'hbacbc12e),
	.w6(32'h3c1b0e41),
	.w7(32'h3bf00091),
	.w8(32'h3a81a39e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a8fe),
	.w1(32'hba1dbb6a),
	.w2(32'hbbc91d82),
	.w3(32'h3b18922d),
	.w4(32'hb9176721),
	.w5(32'hbb679a65),
	.w6(32'h39c7dd4e),
	.w7(32'hbb4082aa),
	.w8(32'hbaa7cdb7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991bcf),
	.w1(32'h3bb4e8f6),
	.w2(32'h3bd48786),
	.w3(32'h3bb0b00d),
	.w4(32'h3a572324),
	.w5(32'hbc66a30b),
	.w6(32'h3b1a63bb),
	.w7(32'h3b503bf0),
	.w8(32'hbc485705),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf26d6),
	.w1(32'hbbaf585d),
	.w2(32'hbb822eb8),
	.w3(32'hbc7ee5b4),
	.w4(32'hbbd8f426),
	.w5(32'hbc437c41),
	.w6(32'hbc08405c),
	.w7(32'hbb5472dc),
	.w8(32'hbb38f3e8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5614b),
	.w1(32'h3b3f5b8f),
	.w2(32'hba6e4670),
	.w3(32'hb8f7647f),
	.w4(32'hbba1af5e),
	.w5(32'h3b87ceb2),
	.w6(32'h3be5b17f),
	.w7(32'hba78ebb9),
	.w8(32'h3b4127d2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211141),
	.w1(32'h3aba2085),
	.w2(32'h3af2fa54),
	.w3(32'hba99b91a),
	.w4(32'hbb001f51),
	.w5(32'hbb62f5ac),
	.w6(32'h3b18ee46),
	.w7(32'hba84a621),
	.w8(32'hbbc20350),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9dbb3),
	.w1(32'hbbdc3dd6),
	.w2(32'hbb924f97),
	.w3(32'h3a586d55),
	.w4(32'hbb1c3d97),
	.w5(32'h3a1ff639),
	.w6(32'hbb5e4c2b),
	.w7(32'hbb4284ea),
	.w8(32'hbb90e1a2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122ded),
	.w1(32'hba13fb33),
	.w2(32'hbb255e2f),
	.w3(32'hbb7e0e23),
	.w4(32'hbb34f267),
	.w5(32'h3be1b4f7),
	.w6(32'hbbdbf4fc),
	.w7(32'hbbc228e7),
	.w8(32'h3ba5a014),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c3e1),
	.w1(32'hbb5e4c45),
	.w2(32'hba55eb58),
	.w3(32'h3ba6ee91),
	.w4(32'h3bee4d88),
	.w5(32'hbb01aa97),
	.w6(32'h3a091fdb),
	.w7(32'h3b232115),
	.w8(32'h3a32cbd6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf63d),
	.w1(32'h3ad3d66d),
	.w2(32'h3aec59ce),
	.w3(32'h3b86f3bc),
	.w4(32'h3be9d9c2),
	.w5(32'hbbe190bf),
	.w6(32'h3adda827),
	.w7(32'h3afa6581),
	.w8(32'hbb8333b2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baae50),
	.w1(32'h3b068f20),
	.w2(32'h3b17088f),
	.w3(32'hbb20f787),
	.w4(32'h3af8da00),
	.w5(32'h3bc86173),
	.w6(32'hba4ebd17),
	.w7(32'hbb8dafe1),
	.w8(32'h3be00340),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900a8b),
	.w1(32'h3bd16233),
	.w2(32'h3bea0328),
	.w3(32'h39b16be6),
	.w4(32'h3b3bb013),
	.w5(32'h3b0e074d),
	.w6(32'hbac3fdcf),
	.w7(32'h3b99085e),
	.w8(32'h3b179783),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee09d4),
	.w1(32'h3b5f7348),
	.w2(32'hb902da34),
	.w3(32'h3ad74f96),
	.w4(32'h3b0ef01b),
	.w5(32'hbc455ab7),
	.w6(32'h3b6f6455),
	.w7(32'h3b15a32c),
	.w8(32'hbbe7a7b6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc4979),
	.w1(32'h3a2aa4d2),
	.w2(32'hbb1835db),
	.w3(32'h3ba5001a),
	.w4(32'hbba97ff5),
	.w5(32'hbc33724f),
	.w6(32'h3c3c8ff9),
	.w7(32'h3a238d74),
	.w8(32'hbc01e3a3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cef97e),
	.w1(32'h3b35accc),
	.w2(32'hbb08c516),
	.w3(32'hbcc61d62),
	.w4(32'hbbfe3627),
	.w5(32'hbc585694),
	.w6(32'hbc97bb03),
	.w7(32'hbbec4964),
	.w8(32'hbc060404),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac754e),
	.w1(32'h3a40991a),
	.w2(32'hbaf45ae2),
	.w3(32'hbc2fb026),
	.w4(32'hbbb58df4),
	.w5(32'hbc4d117f),
	.w6(32'h3bd768c2),
	.w7(32'hba5eab02),
	.w8(32'hbb2eadc4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abba7a8),
	.w1(32'hbafafad8),
	.w2(32'hbafc9264),
	.w3(32'hbc58ddc5),
	.w4(32'hbb4dc236),
	.w5(32'hba1da411),
	.w6(32'hbaea83bf),
	.w7(32'hbb1f7a0f),
	.w8(32'hbb17fee7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e397e),
	.w1(32'h38c908bf),
	.w2(32'hba3c7d1a),
	.w3(32'hbb00c754),
	.w4(32'h3b64ca3b),
	.w5(32'h3afee4bc),
	.w6(32'h3ba72aed),
	.w7(32'h3abb6e0b),
	.w8(32'h3abf810e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa858a8),
	.w1(32'hb903d70e),
	.w2(32'hb8aa7554),
	.w3(32'hba540a49),
	.w4(32'hbadb84e0),
	.w5(32'hbb8e3b8e),
	.w6(32'h3a150398),
	.w7(32'hbb26731d),
	.w8(32'hbad45e88),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ff39e),
	.w1(32'hba754c44),
	.w2(32'hbb067c7a),
	.w3(32'hbb804b08),
	.w4(32'hbaf9a196),
	.w5(32'hbba11b16),
	.w6(32'hbba88c52),
	.w7(32'hbc1fa94f),
	.w8(32'hbba95b80),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab45cc5),
	.w1(32'hbb7d7c18),
	.w2(32'hbbe9225a),
	.w3(32'hbb48e617),
	.w4(32'h3ad2a49f),
	.w5(32'h3b480202),
	.w6(32'h39364c6f),
	.w7(32'hbba39e2c),
	.w8(32'h391edaed),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c8cd3),
	.w1(32'hbaea79b4),
	.w2(32'hbbbfacac),
	.w3(32'hbaa42f63),
	.w4(32'h3b1eca56),
	.w5(32'hbb386ac8),
	.w6(32'h3bc253e3),
	.w7(32'h3ae65957),
	.w8(32'hbb99e5ac),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030b82),
	.w1(32'hbbfc1b7c),
	.w2(32'hbc14d182),
	.w3(32'hbb658f91),
	.w4(32'hbc475e98),
	.w5(32'hbbfc3bf5),
	.w6(32'hb9800559),
	.w7(32'hbbe1b1d2),
	.w8(32'hbb61270f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09daa8),
	.w1(32'hbbda0eb0),
	.w2(32'hbbd51191),
	.w3(32'hbb0682d8),
	.w4(32'hbbd5b193),
	.w5(32'hbb3dcaa8),
	.w6(32'hbad91cef),
	.w7(32'hbbfa6e49),
	.w8(32'hbc2172a1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a77df),
	.w1(32'hbc3eb05b),
	.w2(32'hbc0d099f),
	.w3(32'hbb51afa1),
	.w4(32'hbb1222b9),
	.w5(32'hbbc91c11),
	.w6(32'hbc63d958),
	.w7(32'hbbdc90a7),
	.w8(32'hbbdd0bc7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891201),
	.w1(32'hb8481bb9),
	.w2(32'hbb2261eb),
	.w3(32'h3b9941b3),
	.w4(32'hbaf99bad),
	.w5(32'hba945748),
	.w6(32'h3aa81dde),
	.w7(32'hba6b9ee0),
	.w8(32'hbb4e3703),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb433ce8),
	.w1(32'hbbe0b7a9),
	.w2(32'hbbb65282),
	.w3(32'h3b5b2cd6),
	.w4(32'hbb3cb1e5),
	.w5(32'hbc023576),
	.w6(32'h3ba7ed46),
	.w7(32'hba3a6373),
	.w8(32'hbc153954),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8734),
	.w1(32'hbbbaf7d6),
	.w2(32'hbba79773),
	.w3(32'hbbbad3e0),
	.w4(32'hbc2b30c1),
	.w5(32'h3b33b9fa),
	.w6(32'hbb18c6eb),
	.w7(32'hbb9dbffb),
	.w8(32'h3bb52775),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59cd3d),
	.w1(32'h3b2efe35),
	.w2(32'h3b4da5d3),
	.w3(32'hb9886ad9),
	.w4(32'h3b020a21),
	.w5(32'h3bb9724d),
	.w6(32'h3b2d5876),
	.w7(32'hbb036fa7),
	.w8(32'h3bf8a3bc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b524f7a),
	.w1(32'h3b2259ba),
	.w2(32'hbb30e952),
	.w3(32'h3bba1831),
	.w4(32'h3ae1e104),
	.w5(32'h3bb0653a),
	.w6(32'h3c025a61),
	.w7(32'h3b19a165),
	.w8(32'h3b17d35c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7d145),
	.w1(32'h3be89111),
	.w2(32'h3c2b59c2),
	.w3(32'h3adc0aef),
	.w4(32'h3c21dd28),
	.w5(32'hba7ddeca),
	.w6(32'hbb0dec69),
	.w7(32'h3bf12269),
	.w8(32'hbb2740a1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede2b8),
	.w1(32'hbac6b41f),
	.w2(32'hbb3b52d4),
	.w3(32'hb9c52321),
	.w4(32'h3b290e5d),
	.w5(32'hbbb66eba),
	.w6(32'hbb8c9810),
	.w7(32'hba0d830f),
	.w8(32'hbbc7dcd4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92311f),
	.w1(32'hbbb26500),
	.w2(32'hbbbfb5dd),
	.w3(32'hbbfd0d73),
	.w4(32'hbc3d71d2),
	.w5(32'h3a2a9767),
	.w6(32'hbc02f878),
	.w7(32'hbbef0930),
	.w8(32'hbb9207ed),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6aa71),
	.w1(32'hbc1a79f3),
	.w2(32'hbc3142f7),
	.w3(32'hbbc75fb3),
	.w4(32'hba890aed),
	.w5(32'hbb474fb4),
	.w6(32'hbc02da18),
	.w7(32'hbb6b9a48),
	.w8(32'hbb2c81bd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec5d49),
	.w1(32'h3b3d0af4),
	.w2(32'hb9fa0953),
	.w3(32'hbc0b1ff1),
	.w4(32'hb9cc15f0),
	.w5(32'h3c604ff1),
	.w6(32'h3b5ee8f5),
	.w7(32'h3b1b22ce),
	.w8(32'hbb2e8a1f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149a58),
	.w1(32'hbc642e67),
	.w2(32'hbc5458a7),
	.w3(32'h3c47d6c0),
	.w4(32'h3ba14d0c),
	.w5(32'hbc1fee09),
	.w6(32'hbbf0ec7d),
	.w7(32'hbb8e1fd4),
	.w8(32'hbbdabecc),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8317f),
	.w1(32'h3988d8c1),
	.w2(32'h3ad6dee0),
	.w3(32'hbbe7cba7),
	.w4(32'hbb60d91f),
	.w5(32'hba51b0b1),
	.w6(32'hbb2c8743),
	.w7(32'h3a119d2f),
	.w8(32'h3b89fcf5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde35aa),
	.w1(32'h3addb4ac),
	.w2(32'hbb92ad50),
	.w3(32'hbb8f5099),
	.w4(32'hbbc48ef5),
	.w5(32'hbbf7d5c9),
	.w6(32'h3b11f90d),
	.w7(32'hb9ca4346),
	.w8(32'hbbe4cc35),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c522c),
	.w1(32'hbbedbed6),
	.w2(32'hbc3a7622),
	.w3(32'hbb2f24b1),
	.w4(32'hbc1befc1),
	.w5(32'hbb2237cb),
	.w6(32'h3a2d9668),
	.w7(32'hbb7d7c07),
	.w8(32'hb9326c2b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba068a22),
	.w1(32'h399a5ac3),
	.w2(32'hbb9d1ac1),
	.w3(32'h3977a7d5),
	.w4(32'h3a80e996),
	.w5(32'hbc08a79f),
	.w6(32'h3a0ac261),
	.w7(32'h3bb61972),
	.w8(32'h399497d9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ccdd),
	.w1(32'h3ab1a322),
	.w2(32'hba28bf61),
	.w3(32'hbcafeabf),
	.w4(32'hbbb2df5a),
	.w5(32'hbb231f91),
	.w6(32'h3c11628c),
	.w7(32'h3bdd0601),
	.w8(32'hb91e3c80),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e3e59),
	.w1(32'hbb84138f),
	.w2(32'hbba647e5),
	.w3(32'hbbdc8fad),
	.w4(32'hbb3882b2),
	.w5(32'hbb82bff6),
	.w6(32'h3bcc261c),
	.w7(32'hba85b911),
	.w8(32'h3838a095),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd2e69),
	.w1(32'h3b2d0f6d),
	.w2(32'h392ccadd),
	.w3(32'hba6bd7ef),
	.w4(32'h3a27ed36),
	.w5(32'hbc1aace5),
	.w6(32'h3b914334),
	.w7(32'h3b592939),
	.w8(32'hbba11ac0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cd85f),
	.w1(32'h3a1d039a),
	.w2(32'h3a4bb1b9),
	.w3(32'h3b115160),
	.w4(32'h3a1cfec5),
	.w5(32'h3b958b23),
	.w6(32'hba13d3d9),
	.w7(32'h3a86f898),
	.w8(32'h3b86f946),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba722774),
	.w1(32'hbadd45e1),
	.w2(32'h38ae8625),
	.w3(32'h3c04ce9d),
	.w4(32'hbb3f7f65),
	.w5(32'h3b4016b2),
	.w6(32'h3c126fea),
	.w7(32'hbabd2786),
	.w8(32'hbbe4ea27),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3453e7),
	.w1(32'hbbc2e2f4),
	.w2(32'hbbaa4f07),
	.w3(32'h3ba96890),
	.w4(32'h3ae9e985),
	.w5(32'hbb1611dd),
	.w6(32'hbb7f00be),
	.w7(32'h3b38bf15),
	.w8(32'hbb437d70),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39837),
	.w1(32'hbc212811),
	.w2(32'hbc4017ed),
	.w3(32'hba8cf088),
	.w4(32'hbc0877ca),
	.w5(32'h397b4aab),
	.w6(32'hbc05e3cf),
	.w7(32'hbc35a71f),
	.w8(32'hba0b258a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91553f),
	.w1(32'hbb4094d4),
	.w2(32'hbb099117),
	.w3(32'h3bc2ec59),
	.w4(32'h3ad35bc2),
	.w5(32'h3b1060db),
	.w6(32'h3c300d65),
	.w7(32'h3b8dc418),
	.w8(32'h3b5a8319),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5c51),
	.w1(32'h3b2ea7b2),
	.w2(32'hbc3253c9),
	.w3(32'h3c10ae75),
	.w4(32'h39c79bc7),
	.w5(32'h3afe13fc),
	.w6(32'h3c388ff5),
	.w7(32'h3b25fcaf),
	.w8(32'h3baa37d9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139f49),
	.w1(32'h3c1980a3),
	.w2(32'h3b93b7af),
	.w3(32'h3cabb2f9),
	.w4(32'h3c06eba7),
	.w5(32'h3c04981e),
	.w6(32'h3c9ff781),
	.w7(32'h3be58072),
	.w8(32'hbb5783cd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa2b8b),
	.w1(32'h3b558289),
	.w2(32'h3b6f8fe2),
	.w3(32'h3cbcad49),
	.w4(32'h3bde6f50),
	.w5(32'hbbcd75c7),
	.w6(32'h3bbab1b8),
	.w7(32'hbb8f13a7),
	.w8(32'hbbb6ceda),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfabd75),
	.w1(32'hbc0e9682),
	.w2(32'hbbd4674a),
	.w3(32'hbc7e05ca),
	.w4(32'hbc003db7),
	.w5(32'h3b05e3b8),
	.w6(32'hbc43fee6),
	.w7(32'hbbff0918),
	.w8(32'hba777747),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf676),
	.w1(32'hbb635791),
	.w2(32'h3aa526ab),
	.w3(32'h3bbcdf2a),
	.w4(32'h3bb0aa21),
	.w5(32'h3b40ba81),
	.w6(32'h3b19208e),
	.w7(32'h3afc680e),
	.w8(32'h3ab89bc6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9933a),
	.w1(32'h3ae9f942),
	.w2(32'hba1cfe3c),
	.w3(32'hb8e95249),
	.w4(32'hbbb49329),
	.w5(32'hbaf4ff39),
	.w6(32'hbba991db),
	.w7(32'hb9b51207),
	.w8(32'hbb59bcad),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e2b6),
	.w1(32'h3af93352),
	.w2(32'hbaf20e6b),
	.w3(32'h3b9e803d),
	.w4(32'hbba53413),
	.w5(32'hbc495e28),
	.w6(32'h3be1ef36),
	.w7(32'hbc2fac07),
	.w8(32'h3a8ea9d3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24720d),
	.w1(32'h3cae308a),
	.w2(32'h3b2102be),
	.w3(32'hbca217eb),
	.w4(32'hbc368b00),
	.w5(32'hbb7d812e),
	.w6(32'hbbc66ebb),
	.w7(32'hbc4af3f9),
	.w8(32'hbb1746da),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0788),
	.w1(32'h3bf4dcb6),
	.w2(32'h3a99f15d),
	.w3(32'hba4a1ea8),
	.w4(32'hba95c131),
	.w5(32'hb9ca9471),
	.w6(32'h3bb47233),
	.w7(32'hbbb1c66f),
	.w8(32'h3a762f76),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90dfdf),
	.w1(32'h3a2b687c),
	.w2(32'hbba5f56b),
	.w3(32'hb8aa6890),
	.w4(32'hbafe2b09),
	.w5(32'hbb93e644),
	.w6(32'hbb54d958),
	.w7(32'hbb01c13e),
	.w8(32'hbc898ad1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c9fd0),
	.w1(32'hbd0cb556),
	.w2(32'hbbcd6788),
	.w3(32'h3d06b592),
	.w4(32'h3ca267f1),
	.w5(32'hbad78c36),
	.w6(32'h3bcecbf7),
	.w7(32'h3c642565),
	.w8(32'h3c0151ea),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77ad53),
	.w1(32'h3c561bfd),
	.w2(32'h3b1f227f),
	.w3(32'hbc96844b),
	.w4(32'hbc88d3f2),
	.w5(32'h3aa1538d),
	.w6(32'hbb45d348),
	.w7(32'hbc0df386),
	.w8(32'h3b42cdeb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8085fa),
	.w1(32'hbb985784),
	.w2(32'hbbd41ae7),
	.w3(32'h3c2a91bf),
	.w4(32'h3c1f36ff),
	.w5(32'hbc0925de),
	.w6(32'h3ae56fe4),
	.w7(32'h3b730aff),
	.w8(32'h3b919e79),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2da900),
	.w1(32'h3c17a18f),
	.w2(32'hbb7bdc1f),
	.w3(32'hbc963636),
	.w4(32'h3b2f26da),
	.w5(32'h3b115b14),
	.w6(32'h3b395c20),
	.w7(32'h3c29c5c9),
	.w8(32'h3a993f54),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4df681),
	.w1(32'h3bd5daf4),
	.w2(32'hbbc01126),
	.w3(32'hba50c34e),
	.w4(32'hbb334e73),
	.w5(32'h3b86773e),
	.w6(32'h3b99bc2d),
	.w7(32'hbbc46233),
	.w8(32'h3bc23999),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b932d),
	.w1(32'h3bc17e94),
	.w2(32'h3b880416),
	.w3(32'hbbd0eb79),
	.w4(32'hbc51b744),
	.w5(32'hba4fa56d),
	.w6(32'hbb470177),
	.w7(32'hba975057),
	.w8(32'h3b41466a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba185f85),
	.w1(32'h3a124025),
	.w2(32'hbb119c6e),
	.w3(32'hbbd9827e),
	.w4(32'hbbbffdc1),
	.w5(32'h3ae3babb),
	.w6(32'hba487bca),
	.w7(32'hbb17c532),
	.w8(32'hb9c78729),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192696),
	.w1(32'h3bad35a8),
	.w2(32'h3c13979b),
	.w3(32'hbc015b49),
	.w4(32'hbc1e8833),
	.w5(32'h3a56f0e9),
	.w6(32'hbb837c0e),
	.w7(32'h3b5db15f),
	.w8(32'hbb6f3111),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb628602),
	.w1(32'hbb769ebe),
	.w2(32'hbc66c71c),
	.w3(32'hbbdd582e),
	.w4(32'hbbc8d9aa),
	.w5(32'hbb108195),
	.w6(32'hbaecc9f8),
	.w7(32'hbbee5d63),
	.w8(32'hbb35a319),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023532),
	.w1(32'hbaa9e5d8),
	.w2(32'hbc10532d),
	.w3(32'hb9ce0249),
	.w4(32'hbb8125d3),
	.w5(32'h3bee8981),
	.w6(32'hbaf9c974),
	.w7(32'hbb470bad),
	.w8(32'h3b7e283a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b847f4f),
	.w1(32'h3a533815),
	.w2(32'hbb818d8b),
	.w3(32'hbb47b2da),
	.w4(32'hbb2e65ba),
	.w5(32'h3ae09d80),
	.w6(32'h3bf80480),
	.w7(32'hbb82d4a5),
	.w8(32'h3be923b7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6563),
	.w1(32'h3cd2ef0f),
	.w2(32'h3c02e8c6),
	.w3(32'hb9e1d722),
	.w4(32'hbc45f720),
	.w5(32'h39e7755f),
	.w6(32'h3c8f2a29),
	.w7(32'hbb17dad6),
	.w8(32'hb8283eb2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cc2e5),
	.w1(32'hbaae4791),
	.w2(32'h3a4e4d05),
	.w3(32'hbaf073f7),
	.w4(32'h3b2304bc),
	.w5(32'hbb1c6460),
	.w6(32'hb963d815),
	.w7(32'hbaa3be0a),
	.w8(32'hbb379588),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20f0e),
	.w1(32'h3abcc826),
	.w2(32'h3aaf192f),
	.w3(32'h36d36ec5),
	.w4(32'hbb1aacf9),
	.w5(32'hbbc271ae),
	.w6(32'hbb8728c6),
	.w7(32'hba74b7ba),
	.w8(32'h3ad123f1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39609966),
	.w1(32'h3c22a71d),
	.w2(32'hbbf31a04),
	.w3(32'hbc5cd682),
	.w4(32'hbb288ca2),
	.w5(32'h3bb5f686),
	.w6(32'hbc84b9ee),
	.w7(32'hbc05cb00),
	.w8(32'hba5a5a23),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17073),
	.w1(32'hbc09c3e9),
	.w2(32'hbb7cba00),
	.w3(32'hbb894e67),
	.w4(32'h3ac85c3c),
	.w5(32'h3b71cdd6),
	.w6(32'hbc1a69b8),
	.w7(32'hbb663eea),
	.w8(32'h3c2ce289),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c53cd),
	.w1(32'hbbec6cb7),
	.w2(32'h3bac601c),
	.w3(32'h3c06bece),
	.w4(32'h3b5651fb),
	.w5(32'h3aa7dd8a),
	.w6(32'h3bc296ac),
	.w7(32'h3aee0e4d),
	.w8(32'h3bc8e75e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59f027),
	.w1(32'h3be07ac8),
	.w2(32'h3b3746f8),
	.w3(32'h3b848025),
	.w4(32'hbb2b74ac),
	.w5(32'h3b2645b7),
	.w6(32'hbb8fd119),
	.w7(32'h3b0a1941),
	.w8(32'hbad50c67),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104278),
	.w1(32'hbb9e6e06),
	.w2(32'h39efb276),
	.w3(32'hb697035a),
	.w4(32'hbb348b2b),
	.w5(32'hbb26eb5b),
	.w6(32'h3aaacf25),
	.w7(32'h3b95b4fe),
	.w8(32'hbbd03aa1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2ceb0),
	.w1(32'hba91dfc0),
	.w2(32'h3b96a6b4),
	.w3(32'h3b94aaa5),
	.w4(32'h3b74dc50),
	.w5(32'h3a98a8aa),
	.w6(32'hbaee82e9),
	.w7(32'hbbd9a93a),
	.w8(32'hbbb56d8c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18298e),
	.w1(32'hbafd851d),
	.w2(32'hbb940af8),
	.w3(32'h3c319b1a),
	.w4(32'h3bdeda8e),
	.w5(32'hbbc47a72),
	.w6(32'hba15904b),
	.w7(32'h3b8265bf),
	.w8(32'hbbc97bb5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff9b6e),
	.w1(32'hbc265af7),
	.w2(32'hbbb232b0),
	.w3(32'hbc0ae043),
	.w4(32'hbc1f13e2),
	.w5(32'h3aae6615),
	.w6(32'hbb77abd1),
	.w7(32'hbbb4e81a),
	.w8(32'h3c102b76),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4d02),
	.w1(32'h3a7db695),
	.w2(32'h3b052150),
	.w3(32'hb7b0134f),
	.w4(32'hbc16de89),
	.w5(32'hbba8c930),
	.w6(32'h3d2b6e17),
	.w7(32'hbb5b310e),
	.w8(32'h3ba8b4a5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5c1a9),
	.w1(32'h3c06ab48),
	.w2(32'h39b4b566),
	.w3(32'hbbb0441c),
	.w4(32'hbbd502a2),
	.w5(32'h3c5c8ac8),
	.w6(32'hbab28d5d),
	.w7(32'hbb9473fd),
	.w8(32'h3be5370b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272296),
	.w1(32'hbc0132f1),
	.w2(32'hbb354b3e),
	.w3(32'hbb218d90),
	.w4(32'hb94d5540),
	.w5(32'hbb14c019),
	.w6(32'h3b69a8d1),
	.w7(32'hbb05d74a),
	.w8(32'hba0a57f6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule