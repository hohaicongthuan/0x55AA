module layer_8_featuremap_74(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9538b49),
	.w1(32'h3623a22c),
	.w2(32'h39931101),
	.w3(32'hb846ebf7),
	.w4(32'hb7a52f02),
	.w5(32'h39591eb6),
	.w6(32'hb9ba66a7),
	.w7(32'h39b2e0bb),
	.w8(32'hba56a1bd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf243f),
	.w1(32'hb9e245b4),
	.w2(32'hb8fb9385),
	.w3(32'hb9337f95),
	.w4(32'hb93eb5d7),
	.w5(32'hb94a7cc2),
	.w6(32'hba18eebb),
	.w7(32'hb980a980),
	.w8(32'hb9bfccf4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb687eadb),
	.w1(32'hb9703d1c),
	.w2(32'hb863a3da),
	.w3(32'h397838f2),
	.w4(32'hb9181ab1),
	.w5(32'hb99c15d3),
	.w6(32'hb9c3bb03),
	.w7(32'h373f3732),
	.w8(32'h39cc44c9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa2f20),
	.w1(32'hbaca7136),
	.w2(32'hbb13c449),
	.w3(32'hba72b59a),
	.w4(32'hb99a12b1),
	.w5(32'h392c56b5),
	.w6(32'hb943a86a),
	.w7(32'hbab2628c),
	.w8(32'hb983c870),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39411d38),
	.w1(32'h3692b318),
	.w2(32'h3a2ba201),
	.w3(32'h3995b2e5),
	.w4(32'h3a432e7e),
	.w5(32'h3aa49099),
	.w6(32'hba14f702),
	.w7(32'h39b5d944),
	.w8(32'hbb1192cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35def6),
	.w1(32'hbace5fda),
	.w2(32'hba4b4edd),
	.w3(32'hba1f2cb8),
	.w4(32'h395769e9),
	.w5(32'h3acd4d4e),
	.w6(32'hba3c76a8),
	.w7(32'hb8ddf574),
	.w8(32'hbaadf1f7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df1a6f),
	.w1(32'hb9e978b8),
	.w2(32'h393076b8),
	.w3(32'hb9395b8d),
	.w4(32'hb857d979),
	.w5(32'h37ff420a),
	.w6(32'hba93ce8b),
	.w7(32'hb8e7ac98),
	.w8(32'hb945f4b4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956039e),
	.w1(32'hb95f7ba8),
	.w2(32'h39c1e22e),
	.w3(32'h39c64b3c),
	.w4(32'h3a7fb776),
	.w5(32'h3ac16090),
	.w6(32'hba15bc63),
	.w7(32'h39d0a005),
	.w8(32'hbab3032f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29cfa8),
	.w1(32'hba319d8c),
	.w2(32'h3920c1d0),
	.w3(32'hb8b8f971),
	.w4(32'hb6a6edd3),
	.w5(32'hb803458a),
	.w6(32'hbacd4534),
	.w7(32'hb95a9369),
	.w8(32'hbb1be800),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9612f9c),
	.w1(32'hba14b4a8),
	.w2(32'hb9bfafdd),
	.w3(32'hbb43ddb1),
	.w4(32'hbb381f32),
	.w5(32'hbaa000bf),
	.w6(32'hbafe1bfc),
	.w7(32'hbb301686),
	.w8(32'h3a3065f2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82396b),
	.w1(32'h39a5d1a6),
	.w2(32'h3a316da5),
	.w3(32'h3a852487),
	.w4(32'h3a257c1a),
	.w5(32'h39e3f098),
	.w6(32'hb890489a),
	.w7(32'h39e67b4a),
	.w8(32'hba4ce526),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3779cca8),
	.w1(32'hb922d764),
	.w2(32'h37cde65f),
	.w3(32'hb9045e41),
	.w4(32'hb769978e),
	.w5(32'hb8a62c77),
	.w6(32'hba344205),
	.w7(32'hb7b5517f),
	.w8(32'h38bfdd96),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39012ff2),
	.w1(32'h37c2e573),
	.w2(32'h39d786be),
	.w3(32'h37c34c34),
	.w4(32'h39bcd46f),
	.w5(32'h39b1cf04),
	.w6(32'hba0638b1),
	.w7(32'h39167aad),
	.w8(32'hbb31dbd4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb459fac),
	.w1(32'hbabddd67),
	.w2(32'hba420e4a),
	.w3(32'hba2ea382),
	.w4(32'h39af199a),
	.w5(32'h3b0382e0),
	.w6(32'hb9d63b30),
	.w7(32'h39656477),
	.w8(32'hbaa8bcee),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bdd00),
	.w1(32'hba1f3253),
	.w2(32'hb9e3d0d4),
	.w3(32'h38f31b60),
	.w4(32'h3993f237),
	.w5(32'h3a77a211),
	.w6(32'hba2303d6),
	.w7(32'hb8680610),
	.w8(32'hba2f1da0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b70346),
	.w1(32'h39158477),
	.w2(32'h3a1885b6),
	.w3(32'hb9bb84d4),
	.w4(32'hb90ed537),
	.w5(32'h3888c6e8),
	.w6(32'h39325733),
	.w7(32'hb92ae59f),
	.w8(32'h3a89f275),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894f4d),
	.w1(32'h3c058ed5),
	.w2(32'h3be60847),
	.w3(32'hb9ac8107),
	.w4(32'hb986742e),
	.w5(32'h3affaaf0),
	.w6(32'h39c57dab),
	.w7(32'hbaf325f4),
	.w8(32'h38e70674),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39504a2c),
	.w1(32'h38d0cd7f),
	.w2(32'h3a5b84a9),
	.w3(32'h390c643c),
	.w4(32'h39c782f5),
	.w5(32'h3a7193a2),
	.w6(32'h37a1df23),
	.w7(32'h3912ecc6),
	.w8(32'hb903d670),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14277c),
	.w1(32'hba370f8d),
	.w2(32'h39bdeea3),
	.w3(32'h3908f429),
	.w4(32'h3a824fae),
	.w5(32'h3ad961c9),
	.w6(32'hb9cfb87d),
	.w7(32'h39aaf835),
	.w8(32'hbb2687df),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d717e),
	.w1(32'h3a003d03),
	.w2(32'hba0a8718),
	.w3(32'hbb736b0c),
	.w4(32'hbb8195da),
	.w5(32'hbb810c02),
	.w6(32'h3a622307),
	.w7(32'hba3872da),
	.w8(32'h3a817345),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab779e0),
	.w1(32'h3ab9a335),
	.w2(32'h3a0422d8),
	.w3(32'h3a477aff),
	.w4(32'h39342d4f),
	.w5(32'hbaa4bef9),
	.w6(32'h3a6707de),
	.w7(32'h388641b8),
	.w8(32'hb8f8ff5a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995f406),
	.w1(32'h38290449),
	.w2(32'h3a104743),
	.w3(32'hb8fa8b3e),
	.w4(32'hb8bf5881),
	.w5(32'h3a778576),
	.w6(32'hb9eb570f),
	.w7(32'hb82ea323),
	.w8(32'h3b12fabf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa8f08),
	.w1(32'h3a5b14d5),
	.w2(32'h3819bd36),
	.w3(32'hb9b22999),
	.w4(32'h39e18285),
	.w5(32'hba2cf810),
	.w6(32'h3aa0b39c),
	.w7(32'h38617725),
	.w8(32'hbaa7badb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1f789),
	.w1(32'hb9f9bac8),
	.w2(32'h37b93abf),
	.w3(32'hb9ea0313),
	.w4(32'h38dc8dd7),
	.w5(32'h3a82090d),
	.w6(32'hba2f102b),
	.w7(32'h396e754f),
	.w8(32'hbb0d9335),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaededd),
	.w1(32'h3a0f6389),
	.w2(32'hbaf857c9),
	.w3(32'hbaf43457),
	.w4(32'h39adef82),
	.w5(32'hbb72e189),
	.w6(32'hbb275681),
	.w7(32'hbb69d22d),
	.w8(32'h3aaf95c0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c93bd),
	.w1(32'h3a8511b7),
	.w2(32'h39858161),
	.w3(32'hb90d5750),
	.w4(32'h3a016e70),
	.w5(32'hba1e6812),
	.w6(32'h3adf092c),
	.w7(32'h39f2ed7a),
	.w8(32'h3af1e6ff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a939fb8),
	.w1(32'h3a7fffb7),
	.w2(32'h39a41714),
	.w3(32'h391c0ceb),
	.w4(32'h3a0b53e8),
	.w5(32'hba237332),
	.w6(32'h3ae30d3e),
	.w7(32'h3a15feec),
	.w8(32'h3a25e361),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1c3f),
	.w1(32'h3a584077),
	.w2(32'hbb06f866),
	.w3(32'hb9d10565),
	.w4(32'hba9a197e),
	.w5(32'hbb477988),
	.w6(32'hba5fd8d2),
	.w7(32'hbab0a614),
	.w8(32'hbb093681),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e82e2),
	.w1(32'hbae27919),
	.w2(32'hba51a099),
	.w3(32'hbb9d2ee4),
	.w4(32'hbb78f3db),
	.w5(32'hba956253),
	.w6(32'h3b3ac35f),
	.w7(32'hb9dfb242),
	.w8(32'hb9b68edf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7f8f4),
	.w1(32'hb87f97e1),
	.w2(32'h3988f88e),
	.w3(32'h39ebb8d1),
	.w4(32'h38fcc6b8),
	.w5(32'h3912963d),
	.w6(32'h3913f660),
	.w7(32'h39a312d3),
	.w8(32'hbad4c198),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb521128),
	.w1(32'hbab44b75),
	.w2(32'hbb4b1fda),
	.w3(32'hbbd39b93),
	.w4(32'hbba4754c),
	.w5(32'hbb60d27b),
	.w6(32'hba13997c),
	.w7(32'hbbb91526),
	.w8(32'hb9b15621),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd8542),
	.w1(32'h3b312c47),
	.w2(32'h3a1df6a3),
	.w3(32'h3a793c8c),
	.w4(32'h39f99e3c),
	.w5(32'hbb8c5528),
	.w6(32'h39943419),
	.w7(32'hbaf86ac2),
	.w8(32'hbb2c0af6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270409),
	.w1(32'hbb490bf9),
	.w2(32'hbb7ad658),
	.w3(32'hbb8c195e),
	.w4(32'hbae18565),
	.w5(32'h391e70f2),
	.w6(32'hbb359ae4),
	.w7(32'hbb3c682d),
	.w8(32'h397c25f0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41810e),
	.w1(32'hbb7eade0),
	.w2(32'hbb448810),
	.w3(32'hbb2bddc3),
	.w4(32'hbb1f8565),
	.w5(32'h3a5dee43),
	.w6(32'h3a150311),
	.w7(32'hbb6b3eea),
	.w8(32'hbb13cd92),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3591),
	.w1(32'hbaa17dfb),
	.w2(32'hba115bef),
	.w3(32'hb9e880e1),
	.w4(32'h39d00182),
	.w5(32'h3af69a9e),
	.w6(32'hb96dc046),
	.w7(32'h39a348f5),
	.w8(32'hba1b9b6e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818efc4),
	.w1(32'hb98785aa),
	.w2(32'h39b8eed2),
	.w3(32'hb9ca0c94),
	.w4(32'h3a19ee22),
	.w5(32'h3a913580),
	.w6(32'hba6b75f6),
	.w7(32'h3918ab79),
	.w8(32'hba5e6390),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5feda),
	.w1(32'h3b665971),
	.w2(32'hba0373bb),
	.w3(32'hb986d2f6),
	.w4(32'hba2c12a1),
	.w5(32'hbaff691e),
	.w6(32'hb98ace2b),
	.w7(32'hbaf5b39c),
	.w8(32'hb9b41c82),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396aa992),
	.w1(32'h38da48f9),
	.w2(32'h3991c689),
	.w3(32'h3a11164e),
	.w4(32'h38a6e990),
	.w5(32'hb92cfa78),
	.w6(32'hb97130fe),
	.w7(32'h39b8fbe0),
	.w8(32'hbaee95fb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20ac2),
	.w1(32'hba654d27),
	.w2(32'hba9071bd),
	.w3(32'h3a025b3d),
	.w4(32'h3a4b92b2),
	.w5(32'h3ae0016c),
	.w6(32'hba952be1),
	.w7(32'hb8fc447b),
	.w8(32'hba42cee8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1965ec),
	.w1(32'h3ab88e91),
	.w2(32'hba5abbd6),
	.w3(32'hb919591e),
	.w4(32'hba509ea9),
	.w5(32'hbb58ff26),
	.w6(32'hba1f0341),
	.w7(32'hbacbd345),
	.w8(32'h3a5a485e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dfe1e),
	.w1(32'h393ee396),
	.w2(32'hb9a99570),
	.w3(32'hb5ac21ae),
	.w4(32'h38a35617),
	.w5(32'hba1af56c),
	.w6(32'h3a10334b),
	.w7(32'hb8345247),
	.w8(32'hb98e8b8f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a723a),
	.w1(32'hbafaa951),
	.w2(32'hbab8dc46),
	.w3(32'hb9af1907),
	.w4(32'hba3e59d0),
	.w5(32'hbab1c20d),
	.w6(32'hba0905a7),
	.w7(32'hba1abaca),
	.w8(32'h3af8ec48),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af083),
	.w1(32'h3c383951),
	.w2(32'h3b6f64bd),
	.w3(32'h3afe1865),
	.w4(32'h3c0c174b),
	.w5(32'h3b641d51),
	.w6(32'h3bcba8ba),
	.w7(32'hba209a00),
	.w8(32'hb9dcc552),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fac7),
	.w1(32'hbacc03cf),
	.w2(32'hba9ec6f3),
	.w3(32'hb99c46f8),
	.w4(32'hba70f178),
	.w5(32'hbaa1fc33),
	.w6(32'hbaad1e27),
	.w7(32'hba94eec5),
	.w8(32'h3a2d25ee),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf412d),
	.w1(32'hb7c2c02c),
	.w2(32'hb996abfc),
	.w3(32'h3a8a8234),
	.w4(32'h3a25900e),
	.w5(32'h37726ec3),
	.w6(32'h3a9291b2),
	.w7(32'h396506f4),
	.w8(32'hb8a0e7b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991eac2),
	.w1(32'h3a98a034),
	.w2(32'h39125666),
	.w3(32'h3a02ee72),
	.w4(32'h3abe6b21),
	.w5(32'h39a06042),
	.w6(32'h39fb4da4),
	.w7(32'hba040255),
	.w8(32'hbb7067df),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9724c93),
	.w1(32'hbb98ac97),
	.w2(32'hbb8cda9a),
	.w3(32'hb9c39e7f),
	.w4(32'hbc04d8d8),
	.w5(32'hbb757ecc),
	.w6(32'hbbb1a9c8),
	.w7(32'hbbb7ad57),
	.w8(32'hb928ca98),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d19ad),
	.w1(32'hb9b53266),
	.w2(32'hba99332a),
	.w3(32'hb9a388a1),
	.w4(32'h39d0fd60),
	.w5(32'hb99bfa6d),
	.w6(32'h39df5cad),
	.w7(32'hb9dc9b30),
	.w8(32'h3a027325),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a040ce1),
	.w1(32'hba83c7e4),
	.w2(32'h3910b174),
	.w3(32'h3a1e5621),
	.w4(32'hb9294714),
	.w5(32'h3b03cfcb),
	.w6(32'hbaac3282),
	.w7(32'h39f5be79),
	.w8(32'h39e2be8f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc49d1),
	.w1(32'hba014281),
	.w2(32'hba3b0702),
	.w3(32'h3a5082ca),
	.w4(32'h39fea2b2),
	.w5(32'hb997babe),
	.w6(32'h3a4ac526),
	.w7(32'h37248d70),
	.w8(32'h3a16fe45),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f70f74),
	.w1(32'h3999f942),
	.w2(32'h3802e6a2),
	.w3(32'h39d978ce),
	.w4(32'h3a6b4dec),
	.w5(32'h3904980d),
	.w6(32'h39f698d5),
	.w7(32'h362e4662),
	.w8(32'h39894e26),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a88a79),
	.w1(32'hb9bb548a),
	.w2(32'hbac69a20),
	.w3(32'h3a8774a2),
	.w4(32'h3a852bbd),
	.w5(32'hba61dc8d),
	.w6(32'h3a343d92),
	.w7(32'hba5bbd1b),
	.w8(32'h3b4aa52d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b1a9),
	.w1(32'h39317b4e),
	.w2(32'h3b4de705),
	.w3(32'h3b936758),
	.w4(32'hba886d90),
	.w5(32'h3b5e7335),
	.w6(32'hbad9bdf5),
	.w7(32'h3b34e493),
	.w8(32'h3b28f8c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334d13),
	.w1(32'h3b5db0b3),
	.w2(32'h3b8140ea),
	.w3(32'h3b5c4d95),
	.w4(32'h3b7d11b3),
	.w5(32'h3b9fcd85),
	.w6(32'h3b8b39cb),
	.w7(32'h3b973eff),
	.w8(32'hbab5ad42),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1395af),
	.w1(32'h3b8a5a72),
	.w2(32'h3ba4d56a),
	.w3(32'h399f309a),
	.w4(32'h3b3eae0c),
	.w5(32'h3b855df2),
	.w6(32'h3a3ea113),
	.w7(32'h3a4f997b),
	.w8(32'hbb423e38),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82bcc8),
	.w1(32'h391123d3),
	.w2(32'hba8c732f),
	.w3(32'hb9919b12),
	.w4(32'h3a654cd0),
	.w5(32'h3b1ccbae),
	.w6(32'hba72666a),
	.w7(32'hbaade95f),
	.w8(32'h399881fc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e4186),
	.w1(32'h3b3f03de),
	.w2(32'h3a4df4ef),
	.w3(32'h3a3b6700),
	.w4(32'h39dd2639),
	.w5(32'hbafd163b),
	.w6(32'hbaf02b5d),
	.w7(32'h3a9e06e7),
	.w8(32'h3ae39341),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b386e0a),
	.w1(32'h3ad2bf7d),
	.w2(32'hba2bf31d),
	.w3(32'hbb257677),
	.w4(32'h3a0c0192),
	.w5(32'h3b06250b),
	.w6(32'h3a3c70c7),
	.w7(32'hbab818e1),
	.w8(32'h3abe9d4f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad864a3),
	.w1(32'hb941006c),
	.w2(32'h396d8d38),
	.w3(32'h3b024590),
	.w4(32'h39af121d),
	.w5(32'h39d3c06b),
	.w6(32'hb9ea1b68),
	.w7(32'hb71fd44e),
	.w8(32'hbba1ae94),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaeb74),
	.w1(32'hbbcde526),
	.w2(32'hbb9363a7),
	.w3(32'hbbb430fd),
	.w4(32'hbbfefbbe),
	.w5(32'hbb9c9462),
	.w6(32'hbbfb2aeb),
	.w7(32'hbbadda6b),
	.w8(32'h3a2a2f57),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d9e10),
	.w1(32'h3b9e1def),
	.w2(32'h3af46129),
	.w3(32'h3b49ceca),
	.w4(32'h3ba7ad60),
	.w5(32'hb982c111),
	.w6(32'hbb7a90b8),
	.w7(32'hba27fe43),
	.w8(32'hb93ec789),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842b8b3),
	.w1(32'h3a374d03),
	.w2(32'hb9d912f7),
	.w3(32'hb92b9d1b),
	.w4(32'h3994ffbe),
	.w5(32'hba3bbff3),
	.w6(32'h3aa9cca9),
	.w7(32'h39437163),
	.w8(32'h3ae1894f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b21b9),
	.w1(32'hba5766c2),
	.w2(32'hbad6f510),
	.w3(32'h3a9e7ea0),
	.w4(32'h389e40bf),
	.w5(32'hbabd5787),
	.w6(32'h3a3e9cca),
	.w7(32'hb97f77ab),
	.w8(32'h3a3649fa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8ca3),
	.w1(32'hbb0c6af4),
	.w2(32'hbb459911),
	.w3(32'hba93458b),
	.w4(32'hbb9ea7d8),
	.w5(32'hbb54b108),
	.w6(32'h38a4ea8f),
	.w7(32'hbb734acc),
	.w8(32'h3a053e1d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da8b91),
	.w1(32'hba96143a),
	.w2(32'hba640b35),
	.w3(32'h3884e45a),
	.w4(32'hba5ce55f),
	.w5(32'hba95541f),
	.w6(32'hba41fa38),
	.w7(32'hba2a506e),
	.w8(32'hba4e6471),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b99e7),
	.w1(32'hba854d38),
	.w2(32'hba92316c),
	.w3(32'hba359703),
	.w4(32'hba3fd778),
	.w5(32'hba93c829),
	.w6(32'hba8522cb),
	.w7(32'hba845306),
	.w8(32'h39af4210),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d48ba),
	.w1(32'hb9fbdc2a),
	.w2(32'hba573cf0),
	.w3(32'hb6c5e4f1),
	.w4(32'h38882e2e),
	.w5(32'hba20ab5e),
	.w6(32'hb96c4512),
	.w7(32'hba22a6e7),
	.w8(32'h3ad28d51),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8950a5),
	.w1(32'h3b63dd64),
	.w2(32'h3b7846ed),
	.w3(32'h3ac48442),
	.w4(32'h3a91b86a),
	.w5(32'h3a52103e),
	.w6(32'h3b4b1426),
	.w7(32'h3af709a2),
	.w8(32'h3a8660c8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dadbd6),
	.w1(32'hb80b6106),
	.w2(32'hb966bffa),
	.w3(32'h394101c7),
	.w4(32'h39ae4b99),
	.w5(32'hb98b7a0b),
	.w6(32'h39aff935),
	.w7(32'hb8843e45),
	.w8(32'h3ae7dc17),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b249af3),
	.w1(32'h3aabeb1c),
	.w2(32'h3a0544c0),
	.w3(32'h3b3492a7),
	.w4(32'h3aa03897),
	.w5(32'hba6ce93e),
	.w6(32'h3a92de00),
	.w7(32'hb9ec783a),
	.w8(32'hb790553f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba563fc5),
	.w1(32'hbacec631),
	.w2(32'hbabf9a31),
	.w3(32'hb9aee6bd),
	.w4(32'hba66f074),
	.w5(32'hbac1d37e),
	.w6(32'hba2a9eb0),
	.w7(32'hba78525a),
	.w8(32'h39e34cab),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d503c),
	.w1(32'hb91747a5),
	.w2(32'hb9a5baed),
	.w3(32'h39b16c39),
	.w4(32'h3a3b0e87),
	.w5(32'hb822d921),
	.w6(32'h3a393ca3),
	.w7(32'h37a8ca24),
	.w8(32'h37ee373b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abbe7),
	.w1(32'hbad33b0c),
	.w2(32'hbac48435),
	.w3(32'h3917bcb1),
	.w4(32'hba23eede),
	.w5(32'hbac1ca38),
	.w6(32'hb9ede1d5),
	.w7(32'hba4a7321),
	.w8(32'hba98caf6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a813156),
	.w1(32'h3964add8),
	.w2(32'hbb305fba),
	.w3(32'hbb9f2701),
	.w4(32'hbb8d5648),
	.w5(32'hbb45fdcb),
	.w6(32'h3b079fab),
	.w7(32'hbb25479c),
	.w8(32'h3aadb706),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a2b5),
	.w1(32'h3aad164c),
	.w2(32'h39dadd7a),
	.w3(32'h3aa440d7),
	.w4(32'h3b0d9915),
	.w5(32'h3a2706e9),
	.w6(32'h3b0520f7),
	.w7(32'h3a7ae444),
	.w8(32'hb93c4f21),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e8582),
	.w1(32'hba591569),
	.w2(32'hba5e5305),
	.w3(32'hb998339f),
	.w4(32'hb9d8ffc7),
	.w5(32'hba856740),
	.w6(32'hba24b38e),
	.w7(32'hba4d7acb),
	.w8(32'h3a33a21f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d83ae),
	.w1(32'hb9b4394d),
	.w2(32'hba80e376),
	.w3(32'h3a099fd4),
	.w4(32'h39abdcad),
	.w5(32'hba4f9e8b),
	.w6(32'h3a148cc2),
	.w7(32'hb95ce2ae),
	.w8(32'h3b18d31e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2faf64),
	.w1(32'h3a9676b8),
	.w2(32'h3a0dcdf7),
	.w3(32'h3b47e9fd),
	.w4(32'h3a86bf08),
	.w5(32'hbaa8c433),
	.w6(32'h3a6668bc),
	.w7(32'hba17e39b),
	.w8(32'h3a3bf0c0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60ab57),
	.w1(32'h3a0f28ae),
	.w2(32'hb89f60d7),
	.w3(32'h3a91b9cb),
	.w4(32'h3a4b8a59),
	.w5(32'hba8c4e67),
	.w6(32'h3a6ea031),
	.w7(32'hb99dd849),
	.w8(32'hb8c794d9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fcd20),
	.w1(32'hba4a6cf0),
	.w2(32'hb9e587a8),
	.w3(32'hba05216c),
	.w4(32'hba8cb952),
	.w5(32'hb9b877ef),
	.w6(32'hba038805),
	.w7(32'hba23514a),
	.w8(32'h3b8cfd34),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0931be),
	.w1(32'h3b828b0f),
	.w2(32'h3b684d6f),
	.w3(32'h3b6ad8ea),
	.w4(32'h3b31f539),
	.w5(32'h3b1da610),
	.w6(32'h3b06f968),
	.w7(32'h3b01626f),
	.w8(32'h3a23dc01),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aee7d8),
	.w1(32'h395cb029),
	.w2(32'hb9d8062b),
	.w3(32'h3a73c40c),
	.w4(32'h3a6cc1a0),
	.w5(32'hb96696eb),
	.w6(32'h3a82cf96),
	.w7(32'h39248053),
	.w8(32'h39e51f17),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e34dd0),
	.w1(32'h3a37c60a),
	.w2(32'h392f6c38),
	.w3(32'h39f27e5e),
	.w4(32'h39ae84c4),
	.w5(32'h3a0d003e),
	.w6(32'h39820a03),
	.w7(32'hba383cd5),
	.w8(32'hbb2166ee),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2eca78),
	.w1(32'hb9c32c48),
	.w2(32'hbb4b0789),
	.w3(32'hb8deef8d),
	.w4(32'hbb07ac85),
	.w5(32'hbab064a9),
	.w6(32'hbbb3f02c),
	.w7(32'hbb2aa9d2),
	.w8(32'h3a25e8e5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a743d32),
	.w1(32'h3b090efe),
	.w2(32'h3b413ae6),
	.w3(32'h3a42c335),
	.w4(32'h3b3e09f9),
	.w5(32'h3b567740),
	.w6(32'h3ae8e82a),
	.w7(32'h3b41237f),
	.w8(32'h3a7d67b4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c74f3),
	.w1(32'hba0beef4),
	.w2(32'hba4f8f4f),
	.w3(32'h3a5d615d),
	.w4(32'h3a0a923c),
	.w5(32'hba07482d),
	.w6(32'h3a2d7914),
	.w7(32'h388eac3b),
	.w8(32'h38742ddc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a246faf),
	.w1(32'hbab28a42),
	.w2(32'h39016e6c),
	.w3(32'h3a483179),
	.w4(32'hb985513b),
	.w5(32'h3b2bbb16),
	.w6(32'hbaecc2f6),
	.w7(32'h3a14dbe2),
	.w8(32'h3a4be04d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd06e8),
	.w1(32'h39b49df7),
	.w2(32'hba0c779a),
	.w3(32'h3a139eff),
	.w4(32'h39fd263a),
	.w5(32'hbadfea38),
	.w6(32'h39ae3640),
	.w7(32'hba3469b8),
	.w8(32'hbbda8e5d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe008b9),
	.w1(32'hbbcf3324),
	.w2(32'hbbc3cb8b),
	.w3(32'hbbd92578),
	.w4(32'hbbe3878a),
	.w5(32'hbbb46b99),
	.w6(32'hbbdedbb1),
	.w7(32'hbbcd4765),
	.w8(32'h3998d03b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000e1b),
	.w1(32'hbaa4170b),
	.w2(32'h39548b28),
	.w3(32'h3a214127),
	.w4(32'hb94ea870),
	.w5(32'h3b2637f0),
	.w6(32'hbaf0ca5f),
	.w7(32'h3a02609c),
	.w8(32'h38b7f3b6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13a9a6),
	.w1(32'hba888629),
	.w2(32'h3898d096),
	.w3(32'h3a39324c),
	.w4(32'hb88510cd),
	.w5(32'h3b0a05f6),
	.w6(32'hbaad8936),
	.w7(32'h3a1af4d0),
	.w8(32'h3963584b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e365d7),
	.w1(32'h3a7b2cbc),
	.w2(32'h3ad3b4d4),
	.w3(32'hb9989b9f),
	.w4(32'h3a58443f),
	.w5(32'h3aeaeb30),
	.w6(32'h3a453cf5),
	.w7(32'h3ae05c64),
	.w8(32'h3b654736),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474c81),
	.w1(32'h3c04c68e),
	.w2(32'h3b2eb0d9),
	.w3(32'h3b21029c),
	.w4(32'h3b604379),
	.w5(32'h3b3aebb3),
	.w6(32'h3b8c8dd5),
	.w7(32'hba257065),
	.w8(32'h37ce093a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39984f25),
	.w1(32'h39bb08b4),
	.w2(32'h3a15c91c),
	.w3(32'h3a7f903e),
	.w4(32'h3a88e8ad),
	.w5(32'h3a369d74),
	.w6(32'h3ac2fb6d),
	.w7(32'h3a6e9afc),
	.w8(32'hba47a77d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70a9e5),
	.w1(32'h3a9942d2),
	.w2(32'h3a15ed07),
	.w3(32'hb9cde250),
	.w4(32'h395f788e),
	.w5(32'hb9ba6072),
	.w6(32'hb98fd2ee),
	.w7(32'h3ab871e2),
	.w8(32'hbaa613ea),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb525cd3),
	.w1(32'hbb2c2437),
	.w2(32'hba1e0cf0),
	.w3(32'hbb4605f0),
	.w4(32'hbae205b7),
	.w5(32'hb85ff8ce),
	.w6(32'hb9cf9a86),
	.w7(32'h3a97011f),
	.w8(32'h3b236fd2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac09107),
	.w1(32'hbaa49512),
	.w2(32'hb885e4d4),
	.w3(32'h3aa308a4),
	.w4(32'h3a90a489),
	.w5(32'hba39a444),
	.w6(32'h3a4d4403),
	.w7(32'hb7b4efc6),
	.w8(32'hba30a5d9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e8fd0),
	.w1(32'h3b9ada55),
	.w2(32'h3b628502),
	.w3(32'h3ad08908),
	.w4(32'h3a0a28e4),
	.w5(32'h3b39e7c6),
	.w6(32'h3b96542f),
	.w7(32'h3b8eb3a9),
	.w8(32'h3b068cb8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1030cb),
	.w1(32'h3a727878),
	.w2(32'h39efba4c),
	.w3(32'h3b35bdb1),
	.w4(32'h3a6cfad2),
	.w5(32'hba99e109),
	.w6(32'h3a6cae19),
	.w7(32'hb9c9dbc9),
	.w8(32'h39c8e575),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e65f3),
	.w1(32'hb9905f5e),
	.w2(32'hb99f5cd5),
	.w3(32'h39588f52),
	.w4(32'hb9aba3aa),
	.w5(32'hba90daa3),
	.w6(32'hb9972f41),
	.w7(32'hb9d30823),
	.w8(32'hb9fc2970),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba7aa),
	.w1(32'hba88cb61),
	.w2(32'hbac8508d),
	.w3(32'hbade7352),
	.w4(32'hbb185817),
	.w5(32'hbaafb756),
	.w6(32'hbad546c1),
	.w7(32'hba77080d),
	.w8(32'h3a111be6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891c43a),
	.w1(32'hb9361096),
	.w2(32'hba07c999),
	.w3(32'h39a2deec),
	.w4(32'h39fd9434),
	.w5(32'hb9f5df79),
	.w6(32'h39c98771),
	.w7(32'hb9eaa74c),
	.w8(32'h3a473e41),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b675ca),
	.w1(32'h39ff8d5b),
	.w2(32'h39e7a379),
	.w3(32'h3ac3c547),
	.w4(32'h3a4b1bb6),
	.w5(32'hbae463c8),
	.w6(32'h3acd7ff7),
	.w7(32'hb9b33063),
	.w8(32'hbaa0c01a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadce716),
	.w1(32'h389dc3b3),
	.w2(32'h3996ecc4),
	.w3(32'hba9a8c38),
	.w4(32'hb606d4a6),
	.w5(32'h3a15b9f9),
	.w6(32'h3924c2eb),
	.w7(32'h39aecf1f),
	.w8(32'hb879263d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c4146),
	.w1(32'hba164cf4),
	.w2(32'hb446a8e9),
	.w3(32'h391ef1bc),
	.w4(32'hb935e955),
	.w5(32'h3a765b2b),
	.w6(32'hba323d6b),
	.w7(32'h396026d1),
	.w8(32'hb9f4e4f7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c835b),
	.w1(32'hba0623f2),
	.w2(32'hb9164ae8),
	.w3(32'hb9c168fd),
	.w4(32'hb99155f4),
	.w5(32'h390816ea),
	.w6(32'hba082010),
	.w7(32'hb9582fcc),
	.w8(32'h388dd720),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba147370),
	.w1(32'hb96d00b3),
	.w2(32'h3a856c5b),
	.w3(32'hb971e9c5),
	.w4(32'hb947e1c3),
	.w5(32'h3a2fe3b1),
	.w6(32'hb9f57f89),
	.w7(32'h3a947f61),
	.w8(32'hb9f6f982),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f43fa9),
	.w1(32'hba28156f),
	.w2(32'hb996abb8),
	.w3(32'hb9e7f955),
	.w4(32'hba2d6b55),
	.w5(32'hb98387dc),
	.w6(32'hba693a26),
	.w7(32'hba29ac83),
	.w8(32'hb964de4d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c040e8),
	.w1(32'hb9b1cfc9),
	.w2(32'h37f5c838),
	.w3(32'h39209177),
	.w4(32'h38e70628),
	.w5(32'h3944e301),
	.w6(32'h39b50638),
	.w7(32'h39d9ba13),
	.w8(32'h39ba1bb6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f52e2),
	.w1(32'hb7bf2ecd),
	.w2(32'h37d26c68),
	.w3(32'hb90c9801),
	.w4(32'h39924281),
	.w5(32'h3929c4b4),
	.w6(32'hb98f0047),
	.w7(32'hb953a2b9),
	.w8(32'hb9527bc7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef21d2),
	.w1(32'hba162d44),
	.w2(32'hb90889e3),
	.w3(32'hb90795c2),
	.w4(32'hba31fc84),
	.w5(32'hba205875),
	.w6(32'hb9aec7e6),
	.w7(32'hb7a83bcd),
	.w8(32'hb9e3ca82),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92de1d3),
	.w1(32'h39762603),
	.w2(32'hb83a6681),
	.w3(32'h398e9aa8),
	.w4(32'h394c0346),
	.w5(32'hb96a916b),
	.w6(32'h399cbb01),
	.w7(32'h39765b27),
	.w8(32'h3b236b14),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6009b),
	.w1(32'h3a4028a1),
	.w2(32'h3a371487),
	.w3(32'h3acf7b77),
	.w4(32'h3a373d7d),
	.w5(32'h3a295757),
	.w6(32'h3a8cdb7b),
	.w7(32'h3aba8da5),
	.w8(32'hb9ae6e02),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a53c9),
	.w1(32'hb98127ea),
	.w2(32'hb965a915),
	.w3(32'hb9733826),
	.w4(32'hb95171fd),
	.w5(32'hb966f7e3),
	.w6(32'hb9cbffd8),
	.w7(32'hb9e0f2d7),
	.w8(32'hb9af9878),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dc85d),
	.w1(32'hb983cc5c),
	.w2(32'hb9667684),
	.w3(32'hb9a0f5b2),
	.w4(32'hb8ee1ebb),
	.w5(32'hb8f608c7),
	.w6(32'hb9581dbb),
	.w7(32'hb9657dce),
	.w8(32'hba838a87),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8661e8),
	.w1(32'hba4aad59),
	.w2(32'hba196fdd),
	.w3(32'hba8162d2),
	.w4(32'hba2707aa),
	.w5(32'hba06a937),
	.w6(32'hba4318c7),
	.w7(32'hba435e14),
	.w8(32'hb92379d0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a35154),
	.w1(32'h39debfa6),
	.w2(32'h3a2d4d92),
	.w3(32'h39647f21),
	.w4(32'h396aa121),
	.w5(32'h3a3ff481),
	.w6(32'h39a951f5),
	.w7(32'h3a5e80ed),
	.w8(32'h3a8d2c19),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c865d),
	.w1(32'h3a883efd),
	.w2(32'h3a3651d5),
	.w3(32'h3a6aadd3),
	.w4(32'h3a7be5fa),
	.w5(32'h3a1e3b38),
	.w6(32'h3a97f7e1),
	.w7(32'h3a5b55a9),
	.w8(32'h38a0ece9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc129a),
	.w1(32'hb87e293d),
	.w2(32'h39af3ce5),
	.w3(32'hb6d10b68),
	.w4(32'hb9bdfd63),
	.w5(32'h37d0df41),
	.w6(32'hb99f4e4e),
	.w7(32'h39f9ee1a),
	.w8(32'hb91c97d0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37356ce3),
	.w1(32'hba037934),
	.w2(32'hba42bf60),
	.w3(32'hb901eb65),
	.w4(32'hb942efe2),
	.w5(32'hba05c12a),
	.w6(32'hba38ef41),
	.w7(32'hba482bdc),
	.w8(32'h399cbf26),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861ef90),
	.w1(32'hb9d5aac0),
	.w2(32'h3892c3d7),
	.w3(32'h39195c70),
	.w4(32'hb9df06a9),
	.w5(32'h398f2520),
	.w6(32'hb8c32d09),
	.w7(32'hb94a6bef),
	.w8(32'h39b5333a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b717a),
	.w1(32'h38f3bcc8),
	.w2(32'h390299b0),
	.w3(32'h3990f240),
	.w4(32'hba0a3ad1),
	.w5(32'hb954c45b),
	.w6(32'h395f5c64),
	.w7(32'h3a15ec81),
	.w8(32'h3ad5acf3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38b113),
	.w1(32'hba0a778b),
	.w2(32'hb99955ba),
	.w3(32'h3a5a98c6),
	.w4(32'hb9f4a795),
	.w5(32'hb99aa88c),
	.w6(32'hb82aebd4),
	.w7(32'h39afb990),
	.w8(32'h3941d1ca),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1decaa),
	.w1(32'hbae1cfb4),
	.w2(32'hb982af0f),
	.w3(32'h38179399),
	.w4(32'hba815418),
	.w5(32'hb94c1199),
	.w6(32'hba36cee1),
	.w7(32'h39b56458),
	.w8(32'hba041d1c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47412b),
	.w1(32'hba2c6704),
	.w2(32'h383513c8),
	.w3(32'hba8d4743),
	.w4(32'hba6ec299),
	.w5(32'hb9c53f0c),
	.w6(32'hba8b4165),
	.w7(32'hbaa8e448),
	.w8(32'hb93b6c74),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390255f8),
	.w1(32'h39df03b0),
	.w2(32'hb9839fd4),
	.w3(32'hb9d46524),
	.w4(32'hb91dcd68),
	.w5(32'hb9825a1e),
	.w6(32'h39bace2c),
	.w7(32'hb948f10a),
	.w8(32'hba6136ae),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aef56),
	.w1(32'hba4d30a8),
	.w2(32'hba94b62e),
	.w3(32'hbab393b2),
	.w4(32'hba77f36b),
	.w5(32'hba932b70),
	.w6(32'hba90b541),
	.w7(32'hbae72148),
	.w8(32'h3945f0e1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59dc43),
	.w1(32'h39d0df15),
	.w2(32'h38eddd13),
	.w3(32'h39ed3ca9),
	.w4(32'h37487c96),
	.w5(32'hb965fc8e),
	.w6(32'h39d9eaff),
	.w7(32'h3988f3d6),
	.w8(32'hb8381a16),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule