module layer_10_featuremap_294(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62355c),
	.w1(32'h3ad1f22c),
	.w2(32'hbb7e1704),
	.w3(32'hbb311070),
	.w4(32'hba311abe),
	.w5(32'h3aaa5bf7),
	.w6(32'h3b42b72f),
	.w7(32'h39f31832),
	.w8(32'h3b10aa63),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57b593),
	.w1(32'h3a59d6ef),
	.w2(32'h3b86576e),
	.w3(32'h3becf778),
	.w4(32'h3bee7239),
	.w5(32'h3a1b46ce),
	.w6(32'hbb6b2d60),
	.w7(32'h3ba9d01f),
	.w8(32'h3a2e9d30),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b946f36),
	.w1(32'h3b8a6d2c),
	.w2(32'hbb220912),
	.w3(32'h3a150b74),
	.w4(32'hbb8d9522),
	.w5(32'h3972c734),
	.w6(32'hbab330b7),
	.w7(32'hbb94e009),
	.w8(32'hba3917ab),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bd58b),
	.w1(32'hbb9bc44b),
	.w2(32'hbb110383),
	.w3(32'h3b8c4578),
	.w4(32'h3b1f41d3),
	.w5(32'h3ad519a3),
	.w6(32'hb9c0e3f7),
	.w7(32'h3a9364b0),
	.w8(32'hbc02e96e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446b62),
	.w1(32'hbc1faf0e),
	.w2(32'hbbbdd890),
	.w3(32'h3c4fc6de),
	.w4(32'h3bcef6c9),
	.w5(32'hba3c85d0),
	.w6(32'hbb96fd23),
	.w7(32'hb88a51dc),
	.w8(32'hb9386e61),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7575),
	.w1(32'hbb746b54),
	.w2(32'hbba37d39),
	.w3(32'h3a54c243),
	.w4(32'hbb11d9d7),
	.w5(32'hb9d02ea3),
	.w6(32'h3b0ed5a7),
	.w7(32'hbb1cf871),
	.w8(32'hbac22c2e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab98c66),
	.w1(32'hbb15d2b1),
	.w2(32'h38c1e811),
	.w3(32'hba2e955e),
	.w4(32'h39b3bb5a),
	.w5(32'hbbae55b9),
	.w6(32'hb9fa1317),
	.w7(32'hba835fc1),
	.w8(32'hba3dbbcc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0999e3),
	.w1(32'hbb19ec0d),
	.w2(32'hbc7bff08),
	.w3(32'hbc71f33c),
	.w4(32'hbc1f2adf),
	.w5(32'hba2ffc1a),
	.w6(32'h3ae0b43b),
	.w7(32'hbb92d879),
	.w8(32'hbb4ad6a0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04d588),
	.w1(32'hbaf42d0b),
	.w2(32'hbb63071d),
	.w3(32'h3607e713),
	.w4(32'hba9de78f),
	.w5(32'h39a1b46b),
	.w6(32'h3b4e834c),
	.w7(32'h3b3d868a),
	.w8(32'hb9704d72),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd29a2),
	.w1(32'hbb479d38),
	.w2(32'h3aae77fe),
	.w3(32'h3b1e82bb),
	.w4(32'hb9857c4f),
	.w5(32'hb9e47ce4),
	.w6(32'h39d3e030),
	.w7(32'hbb91550f),
	.w8(32'hbb15fc60),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a517),
	.w1(32'hbb411ff6),
	.w2(32'hbba5fec8),
	.w3(32'hba2791d4),
	.w4(32'hbaed1426),
	.w5(32'hbbaf5de0),
	.w6(32'h3af101ae),
	.w7(32'hbb49b74d),
	.w8(32'hbb4f85d1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2614a),
	.w1(32'h3c089d6a),
	.w2(32'h3b6d21ad),
	.w3(32'hbba62a3f),
	.w4(32'hb9230f7f),
	.w5(32'hbc088535),
	.w6(32'hbab16ad2),
	.w7(32'hbb8d4177),
	.w8(32'h3b3b5dd2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27f641),
	.w1(32'h3c6e957a),
	.w2(32'h3c697512),
	.w3(32'hbc00cfe4),
	.w4(32'hbc3107e3),
	.w5(32'h3a8cfb45),
	.w6(32'h3b85345e),
	.w7(32'hbaa1389a),
	.w8(32'h3b1f3be5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71bc68),
	.w1(32'hbad177d7),
	.w2(32'hbb97e4de),
	.w3(32'hbb18cb14),
	.w4(32'h3b6ea4a0),
	.w5(32'hbadead2d),
	.w6(32'hbad03376),
	.w7(32'hbb65348b),
	.w8(32'hbba7ac8c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d8147),
	.w1(32'hbb2895e4),
	.w2(32'h3a8d385a),
	.w3(32'hbab40f4f),
	.w4(32'hbb82c613),
	.w5(32'h3aab5b85),
	.w6(32'hba3d56f8),
	.w7(32'hbb234e1d),
	.w8(32'h382fbff2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2c17),
	.w1(32'hbacfe3d9),
	.w2(32'h3b71f078),
	.w3(32'hbac178dc),
	.w4(32'hb9523f6a),
	.w5(32'h3a7dcbd4),
	.w6(32'hbba2e8d0),
	.w7(32'hbb7aacb2),
	.w8(32'hb9c4762b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bccea),
	.w1(32'hbb960cce),
	.w2(32'hb9d1ceca),
	.w3(32'hba6d2dd1),
	.w4(32'hb87f777b),
	.w5(32'hbba75bc8),
	.w6(32'hbb36a15a),
	.w7(32'hbb4732b5),
	.w8(32'hbb37c3f9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9fe8),
	.w1(32'hbc050eb2),
	.w2(32'hbc3cb0a1),
	.w3(32'hbc8ad05f),
	.w4(32'hbc387b64),
	.w5(32'hba9bf92c),
	.w6(32'hbc526ea7),
	.w7(32'hbc51629e),
	.w8(32'hbb0504ea),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78ffc4),
	.w1(32'hb9dfa012),
	.w2(32'h3a8f478f),
	.w3(32'hbbace2e2),
	.w4(32'hbb49680f),
	.w5(32'h384f6865),
	.w6(32'h3b60290e),
	.w7(32'hbb8fb182),
	.w8(32'hbb405e09),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e2d3),
	.w1(32'hbb9fa704),
	.w2(32'hbb5a57de),
	.w3(32'h39dc33f7),
	.w4(32'h39a327db),
	.w5(32'hba64984e),
	.w6(32'hbb7d8d27),
	.w7(32'hbb27df4a),
	.w8(32'hba53a8cd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88dfc),
	.w1(32'h3a731a5b),
	.w2(32'h38c166d5),
	.w3(32'hbb7e698e),
	.w4(32'hbb1a89f9),
	.w5(32'hba3b704f),
	.w6(32'h3a3b7abd),
	.w7(32'hbb06fba5),
	.w8(32'hbad02835),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb0555),
	.w1(32'hbb9bee56),
	.w2(32'hbb9c2c3e),
	.w3(32'h3b7abecd),
	.w4(32'hb78703bc),
	.w5(32'h3b866826),
	.w6(32'hba412946),
	.w7(32'hbb17b4f8),
	.w8(32'h3acba31a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80d44),
	.w1(32'hbba08a58),
	.w2(32'h38b39896),
	.w3(32'hbc3492be),
	.w4(32'hbb2ef6c5),
	.w5(32'hbc4a200c),
	.w6(32'hbc4d8cfa),
	.w7(32'hbc3391b5),
	.w8(32'hbbdbd687),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e4da),
	.w1(32'h3aa09119),
	.w2(32'h3bf73320),
	.w3(32'hbb8acaed),
	.w4(32'hbb78a949),
	.w5(32'h3c19ab00),
	.w6(32'h3bdc5d6a),
	.w7(32'hbb689e0b),
	.w8(32'hbb7c9dd2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dab0a),
	.w1(32'hb8d9b13d),
	.w2(32'hb9f1a411),
	.w3(32'h3c843409),
	.w4(32'h3b03f2e0),
	.w5(32'h3b3e8d69),
	.w6(32'h3b0636f7),
	.w7(32'h3bd91cee),
	.w8(32'hbab279e7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe23bdc),
	.w1(32'hbb687d15),
	.w2(32'h39461be3),
	.w3(32'hbaf64a74),
	.w4(32'hb93a33e7),
	.w5(32'h3ac7f886),
	.w6(32'h3b188c4f),
	.w7(32'hbaeb6835),
	.w8(32'h3a616700),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac20478),
	.w1(32'hba80be94),
	.w2(32'h39a4d940),
	.w3(32'h3a89a770),
	.w4(32'h3b812d7a),
	.w5(32'h3b8abe9a),
	.w6(32'hb9b5e4e7),
	.w7(32'hbb286914),
	.w8(32'h3b7605b5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47abf8),
	.w1(32'h3b083a97),
	.w2(32'hb9aba6ae),
	.w3(32'h3ba4ea7a),
	.w4(32'h3bdc473a),
	.w5(32'h3ae3bd2b),
	.w6(32'h3bc7012b),
	.w7(32'h3ace4868),
	.w8(32'hba804c06),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f155),
	.w1(32'hbb73e35c),
	.w2(32'hbb9548be),
	.w3(32'h3b8564c5),
	.w4(32'h3b19cca8),
	.w5(32'h3aba0ada),
	.w6(32'hb860545d),
	.w7(32'h3ad5ce29),
	.w8(32'h3acd4b6d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934de63),
	.w1(32'hbb4ca1cc),
	.w2(32'hbb42c5c1),
	.w3(32'h3c289b5b),
	.w4(32'h3bf1cb44),
	.w5(32'h3c04ebcb),
	.w6(32'h3ba45c34),
	.w7(32'h3ba5d47d),
	.w8(32'hbaafbcea),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56ecb3),
	.w1(32'hbba4f863),
	.w2(32'h39c065ed),
	.w3(32'h3baacffb),
	.w4(32'hbb2af239),
	.w5(32'hbbeb6d8b),
	.w6(32'h3afd01cd),
	.w7(32'hba9b2966),
	.w8(32'hbbb6d259),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26a70d),
	.w1(32'h3c0c5378),
	.w2(32'hb9ffa26e),
	.w3(32'hbbe44283),
	.w4(32'hbb847ab3),
	.w5(32'h399c9e1a),
	.w6(32'hbc37b052),
	.w7(32'hbbcbfb70),
	.w8(32'hbaed430e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6b5c),
	.w1(32'hbb6a0396),
	.w2(32'h3b1ef7b3),
	.w3(32'hbbdff98c),
	.w4(32'hbb055c75),
	.w5(32'hbb97816c),
	.w6(32'hbb3bcd6a),
	.w7(32'hbb797e46),
	.w8(32'hbba2976f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb476ca0),
	.w1(32'h3b933eaa),
	.w2(32'h3a1e4092),
	.w3(32'hbbe140a0),
	.w4(32'hbb30dd6d),
	.w5(32'h3a5a59a2),
	.w6(32'hbb03308e),
	.w7(32'h3a9f900d),
	.w8(32'hbb357155),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3808fe),
	.w1(32'hbafe23ab),
	.w2(32'hba2de44d),
	.w3(32'h3bb0299f),
	.w4(32'h3af9d7bf),
	.w5(32'hb9e64b4a),
	.w6(32'hbb21c7a9),
	.w7(32'h3b598f36),
	.w8(32'hb8f9fe67),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42c770),
	.w1(32'h3a833b3c),
	.w2(32'h3a76652a),
	.w3(32'hbbca9b24),
	.w4(32'hbb63b617),
	.w5(32'h3ae8cd01),
	.w6(32'h3ba5947f),
	.w7(32'hbba3a574),
	.w8(32'hbc061bd8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb29dc),
	.w1(32'hbc3d7dcd),
	.w2(32'hbb5d1a39),
	.w3(32'hbb02fe9c),
	.w4(32'hbbc3efec),
	.w5(32'h3c0821e9),
	.w6(32'hbc138be2),
	.w7(32'hbac5fdd3),
	.w8(32'h3b22b19b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d4c18),
	.w1(32'h3bba5fe6),
	.w2(32'h3bf354f7),
	.w3(32'h3c979d10),
	.w4(32'h3c26c995),
	.w5(32'h3bb66019),
	.w6(32'h3c5d10db),
	.w7(32'h3c046271),
	.w8(32'h3b7db436),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c631751),
	.w1(32'h3c205832),
	.w2(32'h3c14f56b),
	.w3(32'h3ca84df5),
	.w4(32'h3bda62de),
	.w5(32'h3b176ffd),
	.w6(32'h3c217805),
	.w7(32'h3c091453),
	.w8(32'h3bb668ba),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92870b),
	.w1(32'hbc159e59),
	.w2(32'hbc0a88b8),
	.w3(32'h3b77b911),
	.w4(32'hbb11284d),
	.w5(32'hbb9859ab),
	.w6(32'h3b3bd442),
	.w7(32'h3aad6e75),
	.w8(32'hbbd54950),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd15589),
	.w1(32'h3a631720),
	.w2(32'hbb83c7c0),
	.w3(32'hbb9d6be7),
	.w4(32'h38a1c966),
	.w5(32'h3aebce07),
	.w6(32'hbb988c3d),
	.w7(32'hbba54d00),
	.w8(32'hbacdc702),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a767),
	.w1(32'hbb9f90de),
	.w2(32'hbb4dc053),
	.w3(32'h3adcf00e),
	.w4(32'h3aa86243),
	.w5(32'h3c1273fa),
	.w6(32'h39c40870),
	.w7(32'hbb2f2fdb),
	.w8(32'h3b78a52f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d73ac),
	.w1(32'h3b3ed61e),
	.w2(32'h3ba4b999),
	.w3(32'h3bc354a6),
	.w4(32'h3b86bba6),
	.w5(32'hba71a50b),
	.w6(32'h3b9650cc),
	.w7(32'h3be43c94),
	.w8(32'hbbde11ee),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db98e),
	.w1(32'h3aac4e90),
	.w2(32'h3c2ad78f),
	.w3(32'hbb897b3f),
	.w4(32'h3b89a685),
	.w5(32'hbb11524f),
	.w6(32'h3b90f7a8),
	.w7(32'hbaf9ea18),
	.w8(32'hbb42685b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf89334),
	.w1(32'hbb79886d),
	.w2(32'hba2bf6bf),
	.w3(32'h3b500616),
	.w4(32'h3b582e65),
	.w5(32'hbb7855b1),
	.w6(32'hb888aca6),
	.w7(32'hba05aa58),
	.w8(32'h3a211c81),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b4d34),
	.w1(32'h3b241647),
	.w2(32'h3b844203),
	.w3(32'hbb092f28),
	.w4(32'hb8c67b75),
	.w5(32'h3ab2f112),
	.w6(32'h39384e3b),
	.w7(32'hbbb471c5),
	.w8(32'hba82ea84),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782d7d),
	.w1(32'hbbac6fd2),
	.w2(32'hbb0256b1),
	.w3(32'hbbb16d1e),
	.w4(32'hba6a55f9),
	.w5(32'h3bb6573a),
	.w6(32'hbb7aa9da),
	.w7(32'hbb9be879),
	.w8(32'h3bc6a629),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510843),
	.w1(32'hbba706ca),
	.w2(32'hbbbd5a24),
	.w3(32'hbbed4d60),
	.w4(32'hbc0d788f),
	.w5(32'hbbcfac81),
	.w6(32'hbbddc9f6),
	.w7(32'hbbf54f48),
	.w8(32'hbaf8d93a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cc32e),
	.w1(32'h3c6a4394),
	.w2(32'h3c1efecc),
	.w3(32'hbad10934),
	.w4(32'hbb9a4364),
	.w5(32'h3b8f3810),
	.w6(32'h3c456fcc),
	.w7(32'h3b90a62c),
	.w8(32'h38bfcde0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a8f69),
	.w1(32'hbbd6e393),
	.w2(32'hbbc1d1a8),
	.w3(32'h3acd8749),
	.w4(32'h3a45151c),
	.w5(32'h3bae45a3),
	.w6(32'hbbc6f843),
	.w7(32'hbba6ab20),
	.w8(32'h3bcf3379),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad153),
	.w1(32'hbbd2bb57),
	.w2(32'hbb92357f),
	.w3(32'hbb2b2555),
	.w4(32'hbb5903dd),
	.w5(32'hbba44ed5),
	.w6(32'hbbb526b1),
	.w7(32'hbbb5ad29),
	.w8(32'hbc0bbdaa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf36757),
	.w1(32'hbbbf4862),
	.w2(32'hbb41045e),
	.w3(32'h3ac1b387),
	.w4(32'h3b2f9565),
	.w5(32'h3a7d8e2d),
	.w6(32'hbb9f4468),
	.w7(32'h39afabfe),
	.w8(32'hbb20afca),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890f0d),
	.w1(32'hbaabe465),
	.w2(32'hbba44dd0),
	.w3(32'h3b3866a2),
	.w4(32'h3ba42345),
	.w5(32'h3a68df28),
	.w6(32'h3b5cbd80),
	.w7(32'hbbd05d55),
	.w8(32'hba139421),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa4bb),
	.w1(32'hb9ed89e8),
	.w2(32'h3b035c3f),
	.w3(32'hbc796d83),
	.w4(32'hbbef6a6f),
	.w5(32'hbac26b5b),
	.w6(32'hbc54452d),
	.w7(32'hbb5035fe),
	.w8(32'hbb4ddc50),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92852a),
	.w1(32'hba32f981),
	.w2(32'hbb404ea3),
	.w3(32'h3a380d43),
	.w4(32'h3912f3d9),
	.w5(32'h3aa9e899),
	.w6(32'hbac3c22b),
	.w7(32'hbafc3d4e),
	.w8(32'hbb1689cd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982183),
	.w1(32'h376c6c3a),
	.w2(32'hbb8325ed),
	.w3(32'h3b81b167),
	.w4(32'h3b907a96),
	.w5(32'h3ac997b0),
	.w6(32'hbbcfe2c2),
	.w7(32'hba3d1020),
	.w8(32'hbb7c66f9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabffc43),
	.w1(32'hb9f8caa0),
	.w2(32'hbb0509cf),
	.w3(32'hbad6126f),
	.w4(32'hba3ba4b0),
	.w5(32'hbb2689c4),
	.w6(32'hbb110af5),
	.w7(32'hbb494f67),
	.w8(32'hba864321),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031382),
	.w1(32'hbb1eefeb),
	.w2(32'h3abd726a),
	.w3(32'h3a87afab),
	.w4(32'h3b81fecc),
	.w5(32'h3baf1ff6),
	.w6(32'h39435635),
	.w7(32'h3b4b47dc),
	.w8(32'h3a6965a3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0ae2c),
	.w1(32'hbb90e33e),
	.w2(32'hbb6edd02),
	.w3(32'h3b13bf99),
	.w4(32'h3b804367),
	.w5(32'hbc055b38),
	.w6(32'hbb62ab93),
	.w7(32'hbacc509e),
	.w8(32'hbb7ad9d6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c1cef),
	.w1(32'hbb1f5b79),
	.w2(32'h3a967f35),
	.w3(32'hbb9ad7bb),
	.w4(32'hbc37637c),
	.w5(32'hbaf03d2f),
	.w6(32'hbbb650c1),
	.w7(32'hbc6858a2),
	.w8(32'hb99c2cc1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb463778),
	.w1(32'hbb7d4884),
	.w2(32'hbb7725d4),
	.w3(32'hbb1cbf79),
	.w4(32'hbb02f619),
	.w5(32'hbb483063),
	.w6(32'hbb9ffb8f),
	.w7(32'hbb9d6701),
	.w8(32'hbba7e770),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4616),
	.w1(32'hbc10bf84),
	.w2(32'hbb8654aa),
	.w3(32'hbbb38202),
	.w4(32'h3ab2d80e),
	.w5(32'h3b54306a),
	.w6(32'hbbd61ab5),
	.w7(32'hbbda4d82),
	.w8(32'hbc0640dc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136265),
	.w1(32'hbbd17016),
	.w2(32'hbbc4ad0b),
	.w3(32'h3c2a92c7),
	.w4(32'h3b205ca5),
	.w5(32'h3b07aa92),
	.w6(32'hbae61080),
	.w7(32'hbae45644),
	.w8(32'hba209679),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba060f53),
	.w1(32'h38830e8f),
	.w2(32'h3a015440),
	.w3(32'h3ab36029),
	.w4(32'h3bb7e106),
	.w5(32'h3a96298d),
	.w6(32'hba396002),
	.w7(32'h3b88e7ed),
	.w8(32'hba999631),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4533b1),
	.w1(32'h396ed2ec),
	.w2(32'h3b67e0eb),
	.w3(32'h3bc90552),
	.w4(32'h3af4cd60),
	.w5(32'h3b522f41),
	.w6(32'h3a9660b9),
	.w7(32'h3b1fce52),
	.w8(32'hbb1ca5b9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf40179),
	.w1(32'hbaab0a35),
	.w2(32'hba97f411),
	.w3(32'h3bbea329),
	.w4(32'h3b2a68f0),
	.w5(32'hbb47e2eb),
	.w6(32'h39cfd98e),
	.w7(32'hb9735d77),
	.w8(32'hbb04bb18),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988770),
	.w1(32'hba100d8b),
	.w2(32'hbb6621b8),
	.w3(32'hbb377e99),
	.w4(32'hbb44070d),
	.w5(32'h3ba6c7b1),
	.w6(32'hbafacacd),
	.w7(32'hbab3d508),
	.w8(32'h3b0a2d27),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995e2c),
	.w1(32'hbb886dd0),
	.w2(32'h3babf41d),
	.w3(32'h3c0e62c2),
	.w4(32'hbb54eb86),
	.w5(32'h3afda193),
	.w6(32'h3c5a2388),
	.w7(32'h3bae37d7),
	.w8(32'h3b819438),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39845a33),
	.w1(32'hbb9adfec),
	.w2(32'hbb84eace),
	.w3(32'hbbcb8867),
	.w4(32'h39d6454e),
	.w5(32'hbc04e9ec),
	.w6(32'hbb8b786d),
	.w7(32'hbbdc35d2),
	.w8(32'hbc0d9871),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83fbbe),
	.w1(32'h3b260b15),
	.w2(32'h3bde7f9a),
	.w3(32'h3ba4c395),
	.w4(32'hb8de2df4),
	.w5(32'h3bf328a4),
	.w6(32'h3c0755ab),
	.w7(32'h3b2f8b40),
	.w8(32'h3b76f539),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6e747),
	.w1(32'h3aa6b250),
	.w2(32'h3b78134a),
	.w3(32'h3acb0418),
	.w4(32'h3b9e0c30),
	.w5(32'h3b0e8875),
	.w6(32'h3aec1f04),
	.w7(32'h39346bfd),
	.w8(32'hbbe1ad50),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd4378),
	.w1(32'h3bb1e8e5),
	.w2(32'hba4a4880),
	.w3(32'h3a5f3a28),
	.w4(32'h3b0c174a),
	.w5(32'h3b934864),
	.w6(32'h3c5ad008),
	.w7(32'hbb6e8f97),
	.w8(32'hbb0e4419),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4da0),
	.w1(32'h3b87ca23),
	.w2(32'h3be31ba4),
	.w3(32'h3bb4ba0c),
	.w4(32'h3bcd245f),
	.w5(32'hbbb0f3b7),
	.w6(32'h3a5144c5),
	.w7(32'hbacb4f40),
	.w8(32'h3abd93fc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407c78),
	.w1(32'h3b41c5df),
	.w2(32'h3beea978),
	.w3(32'hbb213fe8),
	.w4(32'hba82154a),
	.w5(32'hbae587d0),
	.w6(32'hba86f4b0),
	.w7(32'h3c286328),
	.w8(32'hba8e67ec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1015e7),
	.w1(32'h3b05bf41),
	.w2(32'hbb7c169e),
	.w3(32'h39d4f8c6),
	.w4(32'hba3efe0b),
	.w5(32'hbb7e6506),
	.w6(32'h3a92174b),
	.w7(32'h3a22b068),
	.w8(32'h3afb221b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc33a17),
	.w1(32'h3c2e3a5e),
	.w2(32'h3b9205d7),
	.w3(32'hbc4ac675),
	.w4(32'hbc4d9d2b),
	.w5(32'hbaff557f),
	.w6(32'h3aad99bd),
	.w7(32'hbb4c7074),
	.w8(32'hbbe7e8d2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64c05),
	.w1(32'hbb300821),
	.w2(32'hbbfb52c6),
	.w3(32'hbc18b4d3),
	.w4(32'hbc007c4c),
	.w5(32'hbb87721c),
	.w6(32'hbc2467ed),
	.w7(32'hbc5ef62b),
	.w8(32'hbc87b294),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8cbdd),
	.w1(32'hbb88fe17),
	.w2(32'hbb558855),
	.w3(32'h3b2e5785),
	.w4(32'h3b3af2fe),
	.w5(32'hbb1790a9),
	.w6(32'hbb81035c),
	.w7(32'hbb2b94f8),
	.w8(32'h3b52971d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaed33),
	.w1(32'hbae29468),
	.w2(32'hbbdcd888),
	.w3(32'hbb850182),
	.w4(32'hbb8a9c51),
	.w5(32'hbb0c7bb0),
	.w6(32'h3bac82e5),
	.w7(32'hba8ec4c6),
	.w8(32'hba7afaf9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29e96d),
	.w1(32'hbb28a1d0),
	.w2(32'hba81b836),
	.w3(32'h386011af),
	.w4(32'hb914ddb8),
	.w5(32'h3b89d5ac),
	.w6(32'h3a8b61e0),
	.w7(32'h39b5485e),
	.w8(32'h3c3feb0f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c684e),
	.w1(32'h3c37be50),
	.w2(32'h3c228c9b),
	.w3(32'h3b942988),
	.w4(32'hb9b419f4),
	.w5(32'h3a8b79a4),
	.w6(32'h3bfa3d85),
	.w7(32'h3b8d1940),
	.w8(32'h3b1254ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71ef42),
	.w1(32'h3ab08260),
	.w2(32'h3a55c366),
	.w3(32'hbbad3527),
	.w4(32'hbbff1af7),
	.w5(32'hbacf101f),
	.w6(32'h3baba6c9),
	.w7(32'h3a0ff7e2),
	.w8(32'hbb08f7f6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41e932),
	.w1(32'hbba3a3c4),
	.w2(32'hbb6b3e5c),
	.w3(32'h3b1813e1),
	.w4(32'hb9d86afb),
	.w5(32'h3b8d2572),
	.w6(32'hb978c42b),
	.w7(32'hbb600b82),
	.w8(32'h3af3a6a3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a1cb8),
	.w1(32'hbad150d5),
	.w2(32'h3be460a0),
	.w3(32'h3c4ef586),
	.w4(32'h3c456029),
	.w5(32'h3a5f28cf),
	.w6(32'h3c1715bd),
	.w7(32'h3ade560d),
	.w8(32'h3812dc37),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38677c),
	.w1(32'hbb5db676),
	.w2(32'hbadb1433),
	.w3(32'h3b820d84),
	.w4(32'h3b149dc3),
	.w5(32'hbb96aab4),
	.w6(32'hb8f22aad),
	.w7(32'hbb3caeaa),
	.w8(32'hbb5d68bb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a4d3e),
	.w1(32'h3b920e12),
	.w2(32'hbae6c820),
	.w3(32'hbb0c58dc),
	.w4(32'hbb39b748),
	.w5(32'h3b46e9a7),
	.w6(32'h3bbdda92),
	.w7(32'hba5c3a61),
	.w8(32'h39977158),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a7c6),
	.w1(32'hbb47a587),
	.w2(32'h3a2c4cf1),
	.w3(32'h3bdee688),
	.w4(32'h3a4fe026),
	.w5(32'h3c0e1047),
	.w6(32'h3b10ee30),
	.w7(32'hbb4903c8),
	.w8(32'hbb1af1c6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c1d36),
	.w1(32'hbb2ab9df),
	.w2(32'h3afc8f7a),
	.w3(32'h3c09e769),
	.w4(32'h3b852b74),
	.w5(32'h3af46708),
	.w6(32'hbb49c128),
	.w7(32'h3b27e98a),
	.w8(32'h3a86a9bb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad1a96),
	.w1(32'hbbc4e96d),
	.w2(32'hbade0c9f),
	.w3(32'hb9a6995f),
	.w4(32'hbb0b406b),
	.w5(32'hba960769),
	.w6(32'hba8c29a7),
	.w7(32'hbb6ba198),
	.w8(32'h3ba617af),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889941),
	.w1(32'hbc06e546),
	.w2(32'hbc982b95),
	.w3(32'hbbe9f7d5),
	.w4(32'h39f9c722),
	.w5(32'hbc30cfd5),
	.w6(32'hbc1e293e),
	.w7(32'hbc23c3e0),
	.w8(32'hbb39ae75),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b2e2d),
	.w1(32'h3bb11e6a),
	.w2(32'hbb42ec2f),
	.w3(32'h39e58d6c),
	.w4(32'h3b3c2c34),
	.w5(32'hba767bdc),
	.w6(32'h3b3009e4),
	.w7(32'h3b474fec),
	.w8(32'hbadc70e1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e79e),
	.w1(32'hbbc73361),
	.w2(32'h3b355025),
	.w3(32'h3ba05175),
	.w4(32'h3c136005),
	.w5(32'h3bbb3cec),
	.w6(32'hbb0f5dcb),
	.w7(32'h3bde6ab7),
	.w8(32'h39c37f03),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07dd33),
	.w1(32'h3b159931),
	.w2(32'h39a06556),
	.w3(32'h3b87b1a6),
	.w4(32'h3c997636),
	.w5(32'hb994dd34),
	.w6(32'hbae40955),
	.w7(32'h3a945256),
	.w8(32'h3b95affd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e6690),
	.w1(32'h3980e68d),
	.w2(32'h3b7cc022),
	.w3(32'hbbc01e9e),
	.w4(32'hbafe98f5),
	.w5(32'h3bbb628f),
	.w6(32'hbb33352f),
	.w7(32'hbacc3594),
	.w8(32'h3b169646),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067628),
	.w1(32'hbabf4a7c),
	.w2(32'h3b495713),
	.w3(32'h3bf660ca),
	.w4(32'h3be70da3),
	.w5(32'h3b1b80c5),
	.w6(32'h3bb5de03),
	.w7(32'h3b0c3792),
	.w8(32'hbb17e432),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954946),
	.w1(32'h3b6b6fd2),
	.w2(32'h3ad742a4),
	.w3(32'h3b484fe1),
	.w4(32'h3b1273e4),
	.w5(32'hbaf01698),
	.w6(32'h3a9488fc),
	.w7(32'h3afdc897),
	.w8(32'h3b998427),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bec89),
	.w1(32'hb9d536ab),
	.w2(32'hbb4768c0),
	.w3(32'h3a53ae7b),
	.w4(32'h3a7c6c61),
	.w5(32'hbb74a044),
	.w6(32'h3b882881),
	.w7(32'h3b8abd13),
	.w8(32'hbb8e3aaf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0f139),
	.w1(32'hbbb1db8a),
	.w2(32'h3b334f22),
	.w3(32'hbbf25ff0),
	.w4(32'hba50ee3f),
	.w5(32'hbafebb12),
	.w6(32'hbbdfd960),
	.w7(32'hbbf76e0f),
	.w8(32'hbb8f4bbb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46c930),
	.w1(32'hbb45c616),
	.w2(32'h3b25a672),
	.w3(32'hba7cef6b),
	.w4(32'h3af8385d),
	.w5(32'hba82c847),
	.w6(32'hbaa5509f),
	.w7(32'hba64ad4c),
	.w8(32'hbb8d39b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9afb0a),
	.w1(32'hbc6d7ff0),
	.w2(32'hbc46856f),
	.w3(32'hbc234960),
	.w4(32'hbc1afc30),
	.w5(32'hbc052914),
	.w6(32'hbc466a75),
	.w7(32'hbc1146f2),
	.w8(32'hbbee99a9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40ff06),
	.w1(32'h3b64debe),
	.w2(32'h3ab89d76),
	.w3(32'h3bfc96ae),
	.w4(32'h3ba0e6ee),
	.w5(32'h3b6e43c0),
	.w6(32'h3bf0e55f),
	.w7(32'h3bae158a),
	.w8(32'h3b23bb78),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f94f7a),
	.w1(32'h3b15035a),
	.w2(32'h3b49e47f),
	.w3(32'h3b00626a),
	.w4(32'hba14b3f5),
	.w5(32'h3b1722c6),
	.w6(32'h3b32ce50),
	.w7(32'h3a0fc24e),
	.w8(32'hb8a9a151),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3c74),
	.w1(32'hbb6f938c),
	.w2(32'h39c4d531),
	.w3(32'hba88841c),
	.w4(32'hba695c3d),
	.w5(32'hbabe4ee2),
	.w6(32'hbb3ed5b5),
	.w7(32'hba8ae85f),
	.w8(32'hbb918e40),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd743b),
	.w1(32'hba2f9cbf),
	.w2(32'hb98f85f0),
	.w3(32'h397c113c),
	.w4(32'h3a9ed930),
	.w5(32'h3ab7f39c),
	.w6(32'h3a52d1e0),
	.w7(32'h3ab48ba6),
	.w8(32'h3b01b359),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad7492),
	.w1(32'hbc77ebba),
	.w2(32'hbc987947),
	.w3(32'hbbf68d1a),
	.w4(32'hbc471273),
	.w5(32'hbc1f575e),
	.w6(32'hbb937f70),
	.w7(32'hbbb2f099),
	.w8(32'hbc2b4723),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73bc682),
	.w1(32'hbb8930b4),
	.w2(32'hb989ae86),
	.w3(32'h3a7dde39),
	.w4(32'hbb00cdb5),
	.w5(32'hbaf3834f),
	.w6(32'h3a9e8839),
	.w7(32'h392ac294),
	.w8(32'h3a38aec0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00cd86),
	.w1(32'hbae82a04),
	.w2(32'hbae804fd),
	.w3(32'hbae7b1bd),
	.w4(32'hb93c7acc),
	.w5(32'hba12875e),
	.w6(32'hb97444ab),
	.w7(32'h3aac3d8f),
	.w8(32'hb9b752ae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba706cc7),
	.w1(32'h3a69d729),
	.w2(32'h3ae4fa8d),
	.w3(32'h3aeed864),
	.w4(32'h3a731a31),
	.w5(32'hbbb79215),
	.w6(32'h3a24e34d),
	.w7(32'h39be59f6),
	.w8(32'hbb8e0b70),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5ba5),
	.w1(32'hbb6a6a1a),
	.w2(32'h3a7977f9),
	.w3(32'hbbcc55c7),
	.w4(32'hbb9e6796),
	.w5(32'h3aa489f0),
	.w6(32'hbbce00b0),
	.w7(32'hbbb1be7d),
	.w8(32'hbab8bf0c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d84c0),
	.w1(32'h3abaf38e),
	.w2(32'h3b68b7a0),
	.w3(32'h3b55485a),
	.w4(32'h3ae8e613),
	.w5(32'h3b2e9123),
	.w6(32'h3ab7857a),
	.w7(32'h3ab12853),
	.w8(32'h3ae25123),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d5811),
	.w1(32'h3a0587de),
	.w2(32'hbb937afd),
	.w3(32'h3b2d558e),
	.w4(32'h3b1e4b33),
	.w5(32'hbb1a2c6b),
	.w6(32'hb984dd23),
	.w7(32'hbb01a7d5),
	.w8(32'h3a11c4f5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c2cf9),
	.w1(32'h399fbb73),
	.w2(32'h3a12bcbb),
	.w3(32'hba450481),
	.w4(32'hba503aa5),
	.w5(32'h3a6b48a3),
	.w6(32'h394f36b9),
	.w7(32'hba58fa2c),
	.w8(32'hba0f85b7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc4eca),
	.w1(32'h3af2d07c),
	.w2(32'h3b3e2cf4),
	.w3(32'hba87ac36),
	.w4(32'h3939c836),
	.w5(32'h3af35a41),
	.w6(32'h3ac9ce4f),
	.w7(32'h3b47ddaf),
	.w8(32'h3abced4b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5bc2d),
	.w1(32'hbacfaaa9),
	.w2(32'h399c0540),
	.w3(32'hbb35aa26),
	.w4(32'hbadb3acb),
	.w5(32'hbab84142),
	.w6(32'hbb6c67c7),
	.w7(32'hbb386c8f),
	.w8(32'hba07b78b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8429fc),
	.w1(32'hbb182da7),
	.w2(32'h38ffe343),
	.w3(32'h3a8caa78),
	.w4(32'hba3a92c5),
	.w5(32'h3a9ad661),
	.w6(32'h3a3d1e7b),
	.w7(32'h39480799),
	.w8(32'h3a8856bf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e38dd),
	.w1(32'hba1fa0c6),
	.w2(32'hba341ac1),
	.w3(32'hbaa0abb7),
	.w4(32'hba545743),
	.w5(32'h3b2f7905),
	.w6(32'hba0752fd),
	.w7(32'hb972a02f),
	.w8(32'h3af75d29),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd0c5),
	.w1(32'h3a990701),
	.w2(32'h3ab69f1f),
	.w3(32'h3b1009ad),
	.w4(32'h3b11065a),
	.w5(32'h3b2b02bf),
	.w6(32'h3aeb31cb),
	.w7(32'h3b003198),
	.w8(32'h399c0d19),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a0754),
	.w1(32'hb9e3f94d),
	.w2(32'h3b268e19),
	.w3(32'h39a884f9),
	.w4(32'h3a067001),
	.w5(32'hbb165faa),
	.w6(32'h37c4af65),
	.w7(32'hba45bff8),
	.w8(32'hbb8f9698),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec511e),
	.w1(32'hbad1114c),
	.w2(32'h3a51861a),
	.w3(32'h3a1fd4b2),
	.w4(32'h3afe8c9e),
	.w5(32'hb9af5af1),
	.w6(32'hbb3519fb),
	.w7(32'hba9a5b16),
	.w8(32'hb9c840cf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bfb38),
	.w1(32'h3a8fa2ac),
	.w2(32'h3b8fe617),
	.w3(32'hbb0f56ef),
	.w4(32'hba56b87e),
	.w5(32'h3ad6451b),
	.w6(32'hbb54cf95),
	.w7(32'hb911dc0c),
	.w8(32'h3b2409e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc6e0),
	.w1(32'h3b1b3036),
	.w2(32'h3a6abcde),
	.w3(32'h39cb2b1f),
	.w4(32'h39149f8d),
	.w5(32'h3937e512),
	.w6(32'h3a0e8dbd),
	.w7(32'h3a00301b),
	.w8(32'h3b1efaf9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02e0b3),
	.w1(32'h3a9f6caa),
	.w2(32'h3a153ea0),
	.w3(32'hbaba7b5b),
	.w4(32'hbab9d006),
	.w5(32'h3b3153c1),
	.w6(32'hba7b4103),
	.w7(32'hbb16891a),
	.w8(32'hb715bec0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a217d),
	.w1(32'h3acfb759),
	.w2(32'hba47d62b),
	.w3(32'h3bf9870c),
	.w4(32'h3b85a530),
	.w5(32'h3a5f9424),
	.w6(32'h3b940001),
	.w7(32'h3a1efba2),
	.w8(32'h3a34bf40),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bb52e),
	.w1(32'h3a93ab90),
	.w2(32'hba175b39),
	.w3(32'h3a2d6318),
	.w4(32'h39aa401c),
	.w5(32'h3a0583cc),
	.w6(32'h3a8ef7e3),
	.w7(32'h3a12f697),
	.w8(32'h3a9f5731),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb799abf8),
	.w1(32'hbb18d96b),
	.w2(32'hbae2e8e5),
	.w3(32'hb9d93bbd),
	.w4(32'hbaad15e7),
	.w5(32'hbad007b7),
	.w6(32'h3969ec51),
	.w7(32'hba2a13b7),
	.w8(32'hbab936c0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9160419),
	.w1(32'hb93278a7),
	.w2(32'hb9eb1ec8),
	.w3(32'hba5b1330),
	.w4(32'h38f0ad2a),
	.w5(32'h3a67fea9),
	.w6(32'hba81680c),
	.w7(32'hba159b74),
	.w8(32'hba4ec66f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e5779),
	.w1(32'hba514e78),
	.w2(32'hb9cb8177),
	.w3(32'h3b10fa94),
	.w4(32'h3a1e0e98),
	.w5(32'hba4580f2),
	.w6(32'h3a91adce),
	.w7(32'h389e4357),
	.w8(32'hb855e1ab),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55bc6a),
	.w1(32'h39365a42),
	.w2(32'h3ae4a37e),
	.w3(32'hbb922bc3),
	.w4(32'hbb8d4e50),
	.w5(32'h3830c712),
	.w6(32'hbb1c7b84),
	.w7(32'hbaf8f467),
	.w8(32'hba5bc0f0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9882b97),
	.w1(32'h3a5ed177),
	.w2(32'h3ba989a1),
	.w3(32'hbb6574d8),
	.w4(32'h3945b2da),
	.w5(32'h3b37fad8),
	.w6(32'hbb806648),
	.w7(32'hb9d9be39),
	.w8(32'h3a98a412),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94edf5d),
	.w1(32'h3a3310ce),
	.w2(32'hb96dc0ab),
	.w3(32'h3a7f7000),
	.w4(32'hb9d85a09),
	.w5(32'hbb0b98eb),
	.w6(32'h3a4551cd),
	.w7(32'hba206e4c),
	.w8(32'hba189f97),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f6ef),
	.w1(32'hba1cd0e0),
	.w2(32'h3a2dcd4c),
	.w3(32'hbb6e7f0d),
	.w4(32'hbb8209ce),
	.w5(32'h3b2ba89d),
	.w6(32'hb9861c7e),
	.w7(32'h3912eb89),
	.w8(32'h3a7853f7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae07173),
	.w1(32'h3ac20789),
	.w2(32'h39612970),
	.w3(32'h3b2eda51),
	.w4(32'h38c4ebbd),
	.w5(32'h3aa86db9),
	.w6(32'h3b045754),
	.w7(32'hb9f8b10f),
	.w8(32'hbbb37704),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780b37),
	.w1(32'hbb981507),
	.w2(32'hbac62642),
	.w3(32'hbaad64dc),
	.w4(32'h39d55584),
	.w5(32'h3ab444e0),
	.w6(32'hbbd6c482),
	.w7(32'hbb80885e),
	.w8(32'h398eb0e7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96966a8),
	.w1(32'h3b0730b3),
	.w2(32'h3b18e91e),
	.w3(32'h3a974ff6),
	.w4(32'h3b0ced5f),
	.w5(32'h3b13a38f),
	.w6(32'h39b893d9),
	.w7(32'h38bdd1d6),
	.w8(32'h3a3b7c3f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f06f),
	.w1(32'hbbc5509e),
	.w2(32'hbb45c280),
	.w3(32'hbbe293ce),
	.w4(32'hbb82e0d4),
	.w5(32'hb7030b17),
	.w6(32'hbbe18718),
	.w7(32'hbc02b40e),
	.w8(32'hbaf5cbe9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f51cd),
	.w1(32'h3b215daa),
	.w2(32'h3b31b650),
	.w3(32'h3b92672f),
	.w4(32'h3b0cc99d),
	.w5(32'h3ab7122c),
	.w6(32'h3b857d01),
	.w7(32'h3adadaa0),
	.w8(32'h3aaedfdc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab4d91),
	.w1(32'h3aa80890),
	.w2(32'h3abc1b43),
	.w3(32'hba32253e),
	.w4(32'h3a2761f1),
	.w5(32'h3a2f2b6f),
	.w6(32'hb9b9b933),
	.w7(32'hba6a1705),
	.w8(32'hbb4bdf6a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eeab6),
	.w1(32'hbb672cbd),
	.w2(32'hbb503064),
	.w3(32'hbbda68a0),
	.w4(32'hbb214deb),
	.w5(32'hbb071b4b),
	.w6(32'hbbbcbce2),
	.w7(32'hbb9cc89e),
	.w8(32'hbb216bcb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1f637),
	.w1(32'h39b8254d),
	.w2(32'h3ae935ac),
	.w3(32'h3b1239dc),
	.w4(32'hba846e92),
	.w5(32'hbb12aecb),
	.w6(32'h3b0b9008),
	.w7(32'h3a310850),
	.w8(32'hba1340fe),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c85b),
	.w1(32'hb93eb59b),
	.w2(32'h3aef2603),
	.w3(32'hbb72c678),
	.w4(32'hbb31f71c),
	.w5(32'h39d5d500),
	.w6(32'hba7b0c13),
	.w7(32'hbb0508d5),
	.w8(32'hba3759cb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae1567),
	.w1(32'hbaf3cfbb),
	.w2(32'hbaa70be4),
	.w3(32'h39a891af),
	.w4(32'h3ab284b3),
	.w5(32'hba036eb5),
	.w6(32'hba0c0436),
	.w7(32'hb7a6877f),
	.w8(32'hba2ae189),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe93c),
	.w1(32'h3b035fd1),
	.w2(32'h3b957b14),
	.w3(32'h3bee144f),
	.w4(32'h3bc32af5),
	.w5(32'h3aca4950),
	.w6(32'h3be4ae26),
	.w7(32'h3bc833cb),
	.w8(32'hba120e4f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238b59),
	.w1(32'hbb61c37c),
	.w2(32'hbbab466d),
	.w3(32'h3a1ee9d1),
	.w4(32'hb898a900),
	.w5(32'hbac418a5),
	.w6(32'hbb085d68),
	.w7(32'hbb725e28),
	.w8(32'hbb5b5ccb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83dee2),
	.w1(32'h39b4b21c),
	.w2(32'h3aaeebdc),
	.w3(32'hb5c195fe),
	.w4(32'h3a01a1fb),
	.w5(32'h3a398fdd),
	.w6(32'hba19518e),
	.w7(32'h3a8eccae),
	.w8(32'h3a1494ec),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4821b),
	.w1(32'h3a722a92),
	.w2(32'h3a47e8d8),
	.w3(32'h3a628487),
	.w4(32'h39b75d1c),
	.w5(32'hba37a876),
	.w6(32'h3a870013),
	.w7(32'hb9fefa1f),
	.w8(32'hbaa337c2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10197a),
	.w1(32'hbb063c76),
	.w2(32'hb9c9b534),
	.w3(32'h39a34ebf),
	.w4(32'hbae3574e),
	.w5(32'hbaa6d3bf),
	.w6(32'hba7962ce),
	.w7(32'hba8fa4c4),
	.w8(32'hbb0d15a1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8feef4),
	.w1(32'hbb4e553a),
	.w2(32'hbbc04361),
	.w3(32'h39106af2),
	.w4(32'hbb260804),
	.w5(32'hb9aaa2d1),
	.w6(32'hba942984),
	.w7(32'hbb74b89e),
	.w8(32'hbb043638),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d96035),
	.w1(32'hb940d482),
	.w2(32'h3b83f46d),
	.w3(32'h3a53da6e),
	.w4(32'h3982b788),
	.w5(32'h3b4d8539),
	.w6(32'h3a43cd7d),
	.w7(32'hb8a3ff23),
	.w8(32'h3a9d632a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945ac0),
	.w1(32'h3ad29f16),
	.w2(32'h3aef0488),
	.w3(32'h3ab1eda3),
	.w4(32'h3b1343a4),
	.w5(32'h3b0f5642),
	.w6(32'h399ea848),
	.w7(32'h3b0b20c4),
	.w8(32'h3aad8856),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e6af0),
	.w1(32'h3a42cc7e),
	.w2(32'h3baf06fe),
	.w3(32'h3a10b3a1),
	.w4(32'h390acc2e),
	.w5(32'h3812b4b9),
	.w6(32'hb9b2f2b1),
	.w7(32'hba922d56),
	.w8(32'hbaef9479),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a884ffc),
	.w1(32'h3a990b44),
	.w2(32'h3b803362),
	.w3(32'h39ad4267),
	.w4(32'hbacbe78b),
	.w5(32'h3b6d44e6),
	.w6(32'hb9ad2f41),
	.w7(32'hba04c77a),
	.w8(32'h3a1cdb5d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b74b89),
	.w1(32'h3ae35334),
	.w2(32'hb9f8ef4c),
	.w3(32'h3a116457),
	.w4(32'h3aa288ca),
	.w5(32'hbb90dd94),
	.w6(32'hbb0ce3af),
	.w7(32'hbb16357d),
	.w8(32'hbba5d4c7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dfc20),
	.w1(32'hbb6db9f2),
	.w2(32'hbb760068),
	.w3(32'h39b7474c),
	.w4(32'h3a3eee23),
	.w5(32'h3aebdee6),
	.w6(32'h3b2a4a15),
	.w7(32'hb9ca1bce),
	.w8(32'hba169709),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7bf65),
	.w1(32'h39bbae92),
	.w2(32'hba7d75c5),
	.w3(32'h3b441779),
	.w4(32'h3ad5fa40),
	.w5(32'hbb4adb13),
	.w6(32'h3ae61e02),
	.w7(32'hb99ed03c),
	.w8(32'hbb285250),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bae76a),
	.w1(32'hba5637ef),
	.w2(32'hba3ae022),
	.w3(32'hbac17678),
	.w4(32'hba0d407d),
	.w5(32'h3ab053b5),
	.w6(32'hbacec8d4),
	.w7(32'hba5f3b1a),
	.w8(32'hb9912ea0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba613ac8),
	.w1(32'hb9469eb8),
	.w2(32'h38c09caa),
	.w3(32'h3a2b158e),
	.w4(32'h3a666b89),
	.w5(32'hbaa82ac2),
	.w6(32'hba372b36),
	.w7(32'h3a3f2b70),
	.w8(32'hbae37aed),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53b247),
	.w1(32'h3acf89da),
	.w2(32'h3b1260cf),
	.w3(32'h3b2d72b3),
	.w4(32'h3afcb4c0),
	.w5(32'h3a5a2d63),
	.w6(32'h3ac1eb26),
	.w7(32'h39ecb86b),
	.w8(32'hb7f84ad9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd514),
	.w1(32'h3ab47e96),
	.w2(32'h3abbcc69),
	.w3(32'h3b2e7f60),
	.w4(32'h3ae56151),
	.w5(32'h3b11e5fd),
	.w6(32'h3b0077a0),
	.w7(32'h3a7ecab2),
	.w8(32'h399fb869),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39dc0f),
	.w1(32'hbb4575eb),
	.w2(32'hbb6a0061),
	.w3(32'hb9d7cb10),
	.w4(32'h39f6abb0),
	.w5(32'hbb8375bb),
	.w6(32'hbb1e506e),
	.w7(32'hbb903387),
	.w8(32'hba777df0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa297ad),
	.w1(32'hbb4e0547),
	.w2(32'hbb11810b),
	.w3(32'hbb636ad4),
	.w4(32'hbb89163a),
	.w5(32'hbaaaae7d),
	.w6(32'hb9bc982d),
	.w7(32'hba0704be),
	.w8(32'hba932401),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c959),
	.w1(32'hbb2f5aa1),
	.w2(32'hbb3ed9b1),
	.w3(32'hbba7589e),
	.w4(32'hbb91d368),
	.w5(32'hb988a6d4),
	.w6(32'hbb84d6f4),
	.w7(32'hbba17556),
	.w8(32'hbb17ce3f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca850),
	.w1(32'hbb4b535e),
	.w2(32'hbaa09122),
	.w3(32'hba4616df),
	.w4(32'h3a9fe077),
	.w5(32'hba599e6b),
	.w6(32'hbb026bea),
	.w7(32'hba94fafa),
	.w8(32'h3ac3d25d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b0823),
	.w1(32'h394aeda0),
	.w2(32'h3b17f07c),
	.w3(32'hba738bc4),
	.w4(32'hbabdaf7f),
	.w5(32'hba8dbe02),
	.w6(32'h3af3c273),
	.w7(32'h3b2715ff),
	.w8(32'hbadda590),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb72d7),
	.w1(32'hbb198f2b),
	.w2(32'hbacc276e),
	.w3(32'hbaff13c2),
	.w4(32'hb9178014),
	.w5(32'hba2bebab),
	.w6(32'hbb2a2ca0),
	.w7(32'hbaed2520),
	.w8(32'hb9585c9e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb75b),
	.w1(32'hba975150),
	.w2(32'hba8fb4d0),
	.w3(32'h3b54ef03),
	.w4(32'hb91f3a42),
	.w5(32'h3a80d895),
	.w6(32'h3b8df889),
	.w7(32'hba42db0f),
	.w8(32'hba1d4132),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e5e8),
	.w1(32'hba307beb),
	.w2(32'h3ac37a57),
	.w3(32'hbb4c24db),
	.w4(32'hbab831bc),
	.w5(32'h3a24c8c3),
	.w6(32'hbac8a6b3),
	.w7(32'hbaa9702f),
	.w8(32'hba9315f3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01cadd),
	.w1(32'hba226dd4),
	.w2(32'hbaee5fc5),
	.w3(32'h39f317f0),
	.w4(32'h3a929ab4),
	.w5(32'h3ad2ca92),
	.w6(32'hb9a55f0b),
	.w7(32'hb9a5e069),
	.w8(32'hb9fc5186),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83c37c),
	.w1(32'h3ad57e38),
	.w2(32'h3a871f76),
	.w3(32'h3b9b8106),
	.w4(32'h3b69320c),
	.w5(32'hbafd48d8),
	.w6(32'h3b13b00b),
	.w7(32'h3b0478cf),
	.w8(32'hbad8fcbb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e3c9),
	.w1(32'hbad1e3ee),
	.w2(32'hb9f1dd77),
	.w3(32'hbc112a98),
	.w4(32'hbbfaa6d3),
	.w5(32'hbad7e0c5),
	.w6(32'hbc2a1c88),
	.w7(32'hbbe21477),
	.w8(32'hbba19f70),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7929e),
	.w1(32'hbab710f8),
	.w2(32'hba734653),
	.w3(32'h3a6cec07),
	.w4(32'h39351d14),
	.w5(32'h39738056),
	.w6(32'h3a941fdd),
	.w7(32'hb9ba3f9e),
	.w8(32'hb9c82aeb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb508375),
	.w1(32'hbbaae41f),
	.w2(32'hbb7c100c),
	.w3(32'h393add23),
	.w4(32'hbb0baad9),
	.w5(32'hbb17dfd3),
	.w6(32'hb98183e8),
	.w7(32'hbb17edcf),
	.w8(32'hbb169432),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca95cf),
	.w1(32'h3ad8ff32),
	.w2(32'h3b0a2e31),
	.w3(32'hba8d6d40),
	.w4(32'hba404f55),
	.w5(32'h3a85174e),
	.w6(32'h39c77118),
	.w7(32'hbac53f45),
	.w8(32'h39ca7c59),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39592af9),
	.w1(32'hb8aaab33),
	.w2(32'h3b65909c),
	.w3(32'h3adf5575),
	.w4(32'hb9fdd794),
	.w5(32'h3b8d1676),
	.w6(32'h3aee1934),
	.w7(32'hba4ebb09),
	.w8(32'h3b5288cf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947ac94),
	.w1(32'hb98d6b73),
	.w2(32'h3a086197),
	.w3(32'h3aff7206),
	.w4(32'h3aa40719),
	.w5(32'hbacf6b23),
	.w6(32'h3a21019f),
	.w7(32'hbaa293fd),
	.w8(32'hbac3b436),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa642),
	.w1(32'hbb0e648a),
	.w2(32'h39f8dd47),
	.w3(32'hbc1e2957),
	.w4(32'hbbbc5d8b),
	.w5(32'h3af5dc21),
	.w6(32'hbbeb9232),
	.w7(32'hbbe083a1),
	.w8(32'hba60a7a3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6304f4),
	.w1(32'h3b474368),
	.w2(32'h3b21f1c9),
	.w3(32'h3b3327a8),
	.w4(32'h3b3e0722),
	.w5(32'h3986ba79),
	.w6(32'h3b0f98e5),
	.w7(32'h3b1bc987),
	.w8(32'h3a465364),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee33c1),
	.w1(32'h38aa4866),
	.w2(32'hb99d1783),
	.w3(32'hba3bdfe9),
	.w4(32'h3a3508a3),
	.w5(32'h3ac1dbfa),
	.w6(32'hbae00fee),
	.w7(32'hbae983b8),
	.w8(32'h3a0d365e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74d42f),
	.w1(32'hb6d936b4),
	.w2(32'h3a82c675),
	.w3(32'h3a25cd51),
	.w4(32'h3a9aaa46),
	.w5(32'hbb04d7a9),
	.w6(32'h3a159f43),
	.w7(32'h3a470cdd),
	.w8(32'hbaf3bd13),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944fb6),
	.w1(32'hbaf4affc),
	.w2(32'h39ca00df),
	.w3(32'hbad20747),
	.w4(32'h398d0ef7),
	.w5(32'h3a094591),
	.w6(32'hbb4d6649),
	.w7(32'hbaeccb66),
	.w8(32'hb933fafc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d8b6b),
	.w1(32'hba20a3fd),
	.w2(32'hb8ba1e0e),
	.w3(32'hba8b808a),
	.w4(32'hba9338ec),
	.w5(32'hb9c3a64d),
	.w6(32'hba8b158b),
	.w7(32'hba8b66b3),
	.w8(32'h38879398),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919a86e),
	.w1(32'h3a48d544),
	.w2(32'h3ad7c95b),
	.w3(32'hb9967d05),
	.w4(32'h3a913ee8),
	.w5(32'hb9aa95c2),
	.w6(32'hb9e2669c),
	.w7(32'hba4e2045),
	.w8(32'hbb3bb2cf),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb15f),
	.w1(32'hba22fe6e),
	.w2(32'h3980f84f),
	.w3(32'h389c460a),
	.w4(32'h3aa45214),
	.w5(32'hb9534908),
	.w6(32'hba95b832),
	.w7(32'h3a9c53f3),
	.w8(32'hba9b48e4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba435323),
	.w1(32'hba9606dd),
	.w2(32'hba31ba49),
	.w3(32'h39b55ebb),
	.w4(32'hb8e70e32),
	.w5(32'hbb1aa44b),
	.w6(32'h3a3de7a5),
	.w7(32'hb8ea09c5),
	.w8(32'hba1d159c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a8f86),
	.w1(32'h39a086b2),
	.w2(32'h3a2fd5f3),
	.w3(32'hbab4a717),
	.w4(32'hbacfb168),
	.w5(32'h39b41659),
	.w6(32'h37452140),
	.w7(32'h3aa106b5),
	.w8(32'h38b6d7ec),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac15345),
	.w1(32'h3a366a19),
	.w2(32'h3b36a7d2),
	.w3(32'h3b692022),
	.w4(32'hb894b2ad),
	.w5(32'hb93994d1),
	.w6(32'h3b3832f8),
	.w7(32'h3a3453e6),
	.w8(32'hbb139293),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d71f6),
	.w1(32'hbae2e51f),
	.w2(32'hba408f7a),
	.w3(32'hbb1bb3a4),
	.w4(32'hba8361d6),
	.w5(32'h3ae5b5e8),
	.w6(32'hbaf5e2d5),
	.w7(32'h391dddcc),
	.w8(32'hbb079845),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f74aae),
	.w1(32'hbb1b8c16),
	.w2(32'hbadf8396),
	.w3(32'hba130151),
	.w4(32'h3a1a8115),
	.w5(32'hbb720bb7),
	.w6(32'hba20e8cf),
	.w7(32'hba4c3eda),
	.w8(32'hbac174ff),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda43e6),
	.w1(32'hbbab1742),
	.w2(32'h3b9e4094),
	.w3(32'hbc209dde),
	.w4(32'hbbd5f8f0),
	.w5(32'hbb0f2005),
	.w6(32'hbb9446fe),
	.w7(32'hbb89acf0),
	.w8(32'hbb735391),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b203c),
	.w1(32'h3b1397ae),
	.w2(32'h3b2fe035),
	.w3(32'h3bd85709),
	.w4(32'h3bb8639c),
	.w5(32'h3b7473ce),
	.w6(32'h3b845cec),
	.w7(32'h3af823ab),
	.w8(32'h3b1a51ab),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398413e7),
	.w1(32'h3925bf58),
	.w2(32'hb91e39ea),
	.w3(32'h3b018a13),
	.w4(32'h3a9c1961),
	.w5(32'hb9c36df3),
	.w6(32'h3b1a2f39),
	.w7(32'h3a58cf54),
	.w8(32'hba656892),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad1545),
	.w1(32'hb9f36325),
	.w2(32'hba080573),
	.w3(32'hb9a3ae0a),
	.w4(32'hba0d8847),
	.w5(32'hbb05eb9c),
	.w6(32'h39b4a425),
	.w7(32'h3a611bd2),
	.w8(32'hbb097e39),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8f43),
	.w1(32'hba9522e9),
	.w2(32'hb9ef0326),
	.w3(32'hbb0973aa),
	.w4(32'hba6c11ec),
	.w5(32'hb9ba17fb),
	.w6(32'hbb27cec0),
	.w7(32'h39cfa075),
	.w8(32'h38524a5a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a806656),
	.w1(32'h3a261527),
	.w2(32'h39b26f2f),
	.w3(32'hbaddc269),
	.w4(32'hbb14c5f9),
	.w5(32'hba5f85f5),
	.w6(32'hbad58f67),
	.w7(32'hba2548f4),
	.w8(32'hbb20eeee),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba928e0f),
	.w1(32'hbac96048),
	.w2(32'hba199aa7),
	.w3(32'hba83978c),
	.w4(32'hb8be85de),
	.w5(32'h3af622f6),
	.w6(32'hba30462c),
	.w7(32'hbac2d365),
	.w8(32'h3a9f11a7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9ab1b),
	.w1(32'h3a241948),
	.w2(32'hb83171c6),
	.w3(32'h3b7219cc),
	.w4(32'h3acded81),
	.w5(32'hba871c09),
	.w6(32'h3b2c5b25),
	.w7(32'hba705634),
	.w8(32'hbab4f641),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48b1d1),
	.w1(32'h3a94017d),
	.w2(32'h3b273ee5),
	.w3(32'h3b26e995),
	.w4(32'h3a5bcdcc),
	.w5(32'h3b2fdeb7),
	.w6(32'h3b12ddda),
	.w7(32'h3a1ad4a8),
	.w8(32'h3b08b814),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f8a1d),
	.w1(32'hbad1e7d8),
	.w2(32'hba87dc13),
	.w3(32'hbb11cd90),
	.w4(32'hbaff9b28),
	.w5(32'hbb079ff0),
	.w6(32'hbb46388a),
	.w7(32'hbb071958),
	.w8(32'hbae7fe93),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de4cf),
	.w1(32'hbb662885),
	.w2(32'hba102258),
	.w3(32'hbb7c7412),
	.w4(32'hbb87051d),
	.w5(32'hbac51f49),
	.w6(32'hbb5b4d6b),
	.w7(32'hbbc4b80c),
	.w8(32'hbb14ad37),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea055a),
	.w1(32'hbb8a282d),
	.w2(32'hbaf9eb91),
	.w3(32'hbb25adfe),
	.w4(32'hbb6544fd),
	.w5(32'h3b48a424),
	.w6(32'hbb15c8ce),
	.w7(32'hbacd3f4c),
	.w8(32'h3b22ff6c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7cc97),
	.w1(32'h3b388181),
	.w2(32'h3b1b683f),
	.w3(32'h3a911a68),
	.w4(32'h3b28bf66),
	.w5(32'hb9f066bc),
	.w6(32'h3adcc888),
	.w7(32'h3afd5f76),
	.w8(32'h3913c258),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a74c1),
	.w1(32'hbb21d4fa),
	.w2(32'hbae8b4ec),
	.w3(32'hbb5e5f80),
	.w4(32'hbb14733c),
	.w5(32'hb8a26b24),
	.w6(32'h3a5fb050),
	.w7(32'h3ad4cade),
	.w8(32'hba7b74a8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b47df5),
	.w1(32'hba5159e1),
	.w2(32'h3ad4db9b),
	.w3(32'h3a11b68a),
	.w4(32'h3af64a78),
	.w5(32'hba24da58),
	.w6(32'h39aec005),
	.w7(32'h3aab828c),
	.w8(32'h3a0cf1c8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ade66),
	.w1(32'h3b040285),
	.w2(32'h3b424670),
	.w3(32'h392c959d),
	.w4(32'hb937c1fa),
	.w5(32'hba4175e9),
	.w6(32'h3a922b18),
	.w7(32'h3a337479),
	.w8(32'hbb0e445f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefdae5),
	.w1(32'h39c40029),
	.w2(32'hb94e49d6),
	.w3(32'h3b9a410a),
	.w4(32'h3b4cc9cf),
	.w5(32'h3a9b7eba),
	.w6(32'h3ab6c298),
	.w7(32'h3a662874),
	.w8(32'hb9984881),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930672b),
	.w1(32'h38ad4cdd),
	.w2(32'h3a9815e9),
	.w3(32'h3b5fc3f3),
	.w4(32'h3acca4d0),
	.w5(32'h3a145a83),
	.w6(32'h3b38317a),
	.w7(32'h3acc660d),
	.w8(32'hba7926b2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac6090),
	.w1(32'hbb025f8c),
	.w2(32'hba616f2e),
	.w3(32'h3a5fa879),
	.w4(32'h3aa0ddf1),
	.w5(32'h3a8ca373),
	.w6(32'h39adf87c),
	.w7(32'h393772d8),
	.w8(32'hb9b305ed),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34c31e),
	.w1(32'h3b1e9662),
	.w2(32'h3b2b2352),
	.w3(32'h3bb306c1),
	.w4(32'h3aa8c63f),
	.w5(32'h3b159978),
	.w6(32'h3b720544),
	.w7(32'h3aad0e34),
	.w8(32'h3ad1e04a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddff83),
	.w1(32'h39378975),
	.w2(32'h3b1d24e0),
	.w3(32'h39201736),
	.w4(32'h3a474d11),
	.w5(32'h3b88ae03),
	.w6(32'hb9812846),
	.w7(32'hbabf2a8b),
	.w8(32'h3b3363cf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370f50),
	.w1(32'h3bac6deb),
	.w2(32'h3c082b66),
	.w3(32'h3b9fbf84),
	.w4(32'h3b9060b0),
	.w5(32'h39cc6ac4),
	.w6(32'h3b83164b),
	.w7(32'h3b847425),
	.w8(32'hba9fb02a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89aa33),
	.w1(32'hbb07865c),
	.w2(32'hbadaf659),
	.w3(32'hb9b151e1),
	.w4(32'h3a535813),
	.w5(32'h3a92fae9),
	.w6(32'hbafd07f3),
	.w7(32'hbaf273a0),
	.w8(32'h3aa0f3ec),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d255),
	.w1(32'h3a542beb),
	.w2(32'hb96cfb55),
	.w3(32'h39da571e),
	.w4(32'hb9ffd1cb),
	.w5(32'hbb8c9ffc),
	.w6(32'hb99da3b2),
	.w7(32'hbaaf3a2b),
	.w8(32'hbb28bc69),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933a787),
	.w1(32'h3afb23f1),
	.w2(32'h3b8a3b18),
	.w3(32'h3993c2f5),
	.w4(32'hbb8f39ff),
	.w5(32'h3b6840d1),
	.w6(32'h3a898b36),
	.w7(32'hba4ad777),
	.w8(32'h3b4e56a9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf4818),
	.w1(32'hbb96c372),
	.w2(32'hb8c3a9e8),
	.w3(32'hbbb9b80b),
	.w4(32'hbbf43977),
	.w5(32'hb9eaab50),
	.w6(32'hbbe77cf8),
	.w7(32'hbbd66fad),
	.w8(32'hbbb26540),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb839bd82),
	.w1(32'h3a56a291),
	.w2(32'h3b41cc69),
	.w3(32'h3b7cf51b),
	.w4(32'h3a91df0d),
	.w5(32'hb9fa07f4),
	.w6(32'h3b3b636d),
	.w7(32'h39e3bcb5),
	.w8(32'hba88fc7d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349514),
	.w1(32'hb9be8c49),
	.w2(32'h3b3c3ed2),
	.w3(32'hbb50f7dd),
	.w4(32'hb9da6a5c),
	.w5(32'h3ac2ff43),
	.w6(32'hbafdbe52),
	.w7(32'hbaae6bce),
	.w8(32'hbabc3185),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bb20a),
	.w1(32'hbac939c3),
	.w2(32'hba8f2664),
	.w3(32'hb9e633c4),
	.w4(32'h3a0d8d32),
	.w5(32'h3a6119b6),
	.w6(32'hb8c42cf2),
	.w7(32'hba1ca281),
	.w8(32'h3a06c41f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba100b9f),
	.w1(32'hba93d93e),
	.w2(32'hba0987f2),
	.w3(32'hb8ef749c),
	.w4(32'h38c10607),
	.w5(32'h3ace231e),
	.w6(32'h391f05de),
	.w7(32'hb9ba4915),
	.w8(32'h3ae36b05),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b1dc6),
	.w1(32'h3abbb7d4),
	.w2(32'hbb00302e),
	.w3(32'hb9bd4aec),
	.w4(32'hbb4cb48f),
	.w5(32'h3a8f834c),
	.w6(32'hbb02f36b),
	.w7(32'hbb210d6e),
	.w8(32'h39b1c8b8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0db47),
	.w1(32'hbb10b1da),
	.w2(32'h38e5f4a3),
	.w3(32'hbb7384b8),
	.w4(32'hbb75807e),
	.w5(32'hbb66bec2),
	.w6(32'hbb1afc18),
	.w7(32'hbbab279c),
	.w8(32'hbb54f71b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecc94),
	.w1(32'hbab2143a),
	.w2(32'hba99f05e),
	.w3(32'hbb98f84a),
	.w4(32'hbbabb1be),
	.w5(32'hbb4c7cea),
	.w6(32'hbbd76016),
	.w7(32'hbbb34b2f),
	.w8(32'hbba2a3b4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a632e78),
	.w1(32'h3a86efd7),
	.w2(32'hb9a87b41),
	.w3(32'h3adbae22),
	.w4(32'h3a53dd4e),
	.w5(32'hb99f9c73),
	.w6(32'h3a3ad197),
	.w7(32'h3ab17da8),
	.w8(32'hbabb2dab),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39382fad),
	.w1(32'h39200681),
	.w2(32'hb91416d3),
	.w3(32'h3ab3b30c),
	.w4(32'h3ac96a44),
	.w5(32'h3a9085f2),
	.w6(32'hba14eb65),
	.w7(32'hbacf7114),
	.w8(32'hb992992c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e83a90),
	.w1(32'hba8a087f),
	.w2(32'hb91086a5),
	.w3(32'hba8f9d5f),
	.w4(32'hb98c8f41),
	.w5(32'hbb0ac474),
	.w6(32'hbaa13687),
	.w7(32'hb9b05f43),
	.w8(32'hbac56976),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf5e3),
	.w1(32'hbb7e90bb),
	.w2(32'hbb163bfa),
	.w3(32'hbb4834cf),
	.w4(32'hbb6a0333),
	.w5(32'h3adca553),
	.w6(32'hbb45cb47),
	.w7(32'hbae7bff5),
	.w8(32'h3ad6614c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fbeb8),
	.w1(32'h3b908370),
	.w2(32'h3b4945c8),
	.w3(32'h3ae2997c),
	.w4(32'h3acee3fe),
	.w5(32'h3a994807),
	.w6(32'h3af9f337),
	.w7(32'h3ad60fe1),
	.w8(32'hb9cae886),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba825953),
	.w1(32'h398745e9),
	.w2(32'hbaafb037),
	.w3(32'h3b042564),
	.w4(32'h3b1be1cd),
	.w5(32'h3827a7ca),
	.w6(32'h39b2371e),
	.w7(32'h3ad32bac),
	.w8(32'h391cb3ac),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a897fc9),
	.w1(32'h399ffd75),
	.w2(32'hba51ed15),
	.w3(32'h39fba467),
	.w4(32'h3924c288),
	.w5(32'hb9a4ab4b),
	.w6(32'h3a2fc6ff),
	.w7(32'hb92e99ac),
	.w8(32'hb9c4485e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50ffa9),
	.w1(32'hbb544312),
	.w2(32'hb9214c92),
	.w3(32'hbb153225),
	.w4(32'hbb77890f),
	.w5(32'hba97ee6a),
	.w6(32'hbb3b3a58),
	.w7(32'hbb522166),
	.w8(32'hbaed7444),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d468a6),
	.w1(32'h3a989788),
	.w2(32'h3a06b78a),
	.w3(32'h3a67f8cc),
	.w4(32'hba20ec57),
	.w5(32'h3a9f1ad6),
	.w6(32'h3a8ba566),
	.w7(32'h39a28c19),
	.w8(32'hbafea0ce),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a27f7),
	.w1(32'h39b39d37),
	.w2(32'h39d40ec4),
	.w3(32'hb9a8509b),
	.w4(32'hb783f73f),
	.w5(32'h3981f122),
	.w6(32'hba713cbc),
	.w7(32'hb9b12d21),
	.w8(32'h371b91e2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c72a9),
	.w1(32'hbb52fec7),
	.w2(32'hbb8c734b),
	.w3(32'hbc0003d0),
	.w4(32'hbbadea54),
	.w5(32'hbaece887),
	.w6(32'hbbe6bcbb),
	.w7(32'hbbe924a6),
	.w8(32'hbb98a6b5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188d9a),
	.w1(32'hbb084c57),
	.w2(32'hb9b339e5),
	.w3(32'hbb76fc00),
	.w4(32'hbb107a8f),
	.w5(32'h38feb754),
	.w6(32'hbb81ef68),
	.w7(32'hbb3ffd0a),
	.w8(32'hba8448a5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a468a2),
	.w1(32'hb9ae4d8c),
	.w2(32'hb9469b07),
	.w3(32'hba141827),
	.w4(32'hba81c64b),
	.w5(32'hb993eb17),
	.w6(32'hba490ea1),
	.w7(32'hb9d5a2c9),
	.w8(32'hba555e64),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb385ca8),
	.w1(32'hbb2cceb4),
	.w2(32'hba9f1cb6),
	.w3(32'hbb81dc75),
	.w4(32'hbb0c123f),
	.w5(32'hba715bae),
	.w6(32'hbb681fca),
	.w7(32'hbb359bb1),
	.w8(32'hbab28697),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0b865),
	.w1(32'hba6248db),
	.w2(32'hbab0e5d8),
	.w3(32'h3a83df28),
	.w4(32'hb8811c75),
	.w5(32'h3a113e61),
	.w6(32'h3aa8bbe8),
	.w7(32'hba4d999b),
	.w8(32'h3a109c3f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b64fb),
	.w1(32'h3a3e88aa),
	.w2(32'h3a5d0261),
	.w3(32'h39c811ca),
	.w4(32'h3a09d6c2),
	.w5(32'h39a06584),
	.w6(32'h39b10da0),
	.w7(32'h39020c5e),
	.w8(32'h39189091),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a18153),
	.w1(32'hb9242aaf),
	.w2(32'hb9ba4901),
	.w3(32'h38f4dce1),
	.w4(32'hb70f97c5),
	.w5(32'h39c1213d),
	.w6(32'h39e976ea),
	.w7(32'h39162bd6),
	.w8(32'h39ea7186),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f225),
	.w1(32'h39f6ca6b),
	.w2(32'hb8779563),
	.w3(32'h39f50a1a),
	.w4(32'h37f61600),
	.w5(32'hba732575),
	.w6(32'h3995bb0b),
	.w7(32'hb8d7be71),
	.w8(32'hba58f2fa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cfd6a),
	.w1(32'hb9d98c0b),
	.w2(32'hb86993b0),
	.w3(32'h3a28b9fd),
	.w4(32'h39e5336c),
	.w5(32'h3a07e0f0),
	.w6(32'h38cd4bf8),
	.w7(32'hb8ccd5bc),
	.w8(32'h3a5c0ca1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd899b),
	.w1(32'h3a9f00c3),
	.w2(32'h3b9f40aa),
	.w3(32'hbb091507),
	.w4(32'h389c9f84),
	.w5(32'h3b00b739),
	.w6(32'hbb442b61),
	.w7(32'hbb274625),
	.w8(32'h39badba8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b78c),
	.w1(32'hbae2175c),
	.w2(32'h390a506b),
	.w3(32'hbb7c13b1),
	.w4(32'hbb174ff0),
	.w5(32'hb9a5360b),
	.w6(32'hbb2c3fd1),
	.w7(32'hbb1af331),
	.w8(32'hb9efaedb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ad47),
	.w1(32'hbab95539),
	.w2(32'h3b08aed5),
	.w3(32'hbb866dfe),
	.w4(32'hbaec55bf),
	.w5(32'h3906a3ed),
	.w6(32'hbb607bd1),
	.w7(32'hbb5a7492),
	.w8(32'hba8959dc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f5ea0),
	.w1(32'hb99a1265),
	.w2(32'h39ada492),
	.w3(32'hb995408a),
	.w4(32'h39df2cca),
	.w5(32'hb9adc90b),
	.w6(32'h37c7f7d0),
	.w7(32'h3989b415),
	.w8(32'hb99d24d9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbd1a4),
	.w1(32'h39500799),
	.w2(32'h39ab677a),
	.w3(32'hba0d9ad1),
	.w4(32'hb9cf3713),
	.w5(32'h3a036476),
	.w6(32'hb827d75d),
	.w7(32'h3998cf1b),
	.w8(32'h3a17b6de),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35d725),
	.w1(32'h39cb0e1a),
	.w2(32'h3a16fc8d),
	.w3(32'h39c6647c),
	.w4(32'h3a5b86db),
	.w5(32'h3998c99d),
	.w6(32'h38b16094),
	.w7(32'h3a18adfb),
	.w8(32'h383984b5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981eaf5),
	.w1(32'h3a0ae3f2),
	.w2(32'h39f6475c),
	.w3(32'hb98c7a26),
	.w4(32'hb920eb9b),
	.w5(32'hb94b3e99),
	.w6(32'h397644bd),
	.w7(32'hb78c27a3),
	.w8(32'hb984e266),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043621),
	.w1(32'hbae13b32),
	.w2(32'hbb0ff81e),
	.w3(32'hbb546179),
	.w4(32'hbb16df02),
	.w5(32'hbb0710d3),
	.w6(32'hbb5091a9),
	.w7(32'hbb53e049),
	.w8(32'hbad7eea7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88597df),
	.w1(32'h39875ac6),
	.w2(32'hb7ba6186),
	.w3(32'hba04d6ca),
	.w4(32'hb913991d),
	.w5(32'hba9c7fd3),
	.w6(32'h3a8429ac),
	.w7(32'h3a2f4709),
	.w8(32'hba8449af),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061a83),
	.w1(32'h3a84ca2d),
	.w2(32'h3980217d),
	.w3(32'h3ad41b4a),
	.w4(32'h3a34336f),
	.w5(32'h3a73025f),
	.w6(32'h3a8c0801),
	.w7(32'h3a86579e),
	.w8(32'h3a14680d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec66ea),
	.w1(32'hba6ec638),
	.w2(32'hb959c174),
	.w3(32'hb90cfdee),
	.w4(32'hb9bef2d3),
	.w5(32'hb9d2d2b8),
	.w6(32'hb7cb8b15),
	.w7(32'hb95c503a),
	.w8(32'hb9abba7c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6456e6),
	.w1(32'hba022f37),
	.w2(32'hb9e79992),
	.w3(32'hbaa7b13d),
	.w4(32'hbab3b56b),
	.w5(32'hb914d68f),
	.w6(32'hba19391f),
	.w7(32'hba21808b),
	.w8(32'hb9c1110e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec1c98),
	.w1(32'h3a0038c6),
	.w2(32'h397e7742),
	.w3(32'h38fdd59e),
	.w4(32'h38e3e9ef),
	.w5(32'hba84b307),
	.w6(32'hb9df2d60),
	.w7(32'hba9e682f),
	.w8(32'hbac2b224),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97591bf),
	.w1(32'h3855dff8),
	.w2(32'h389a8011),
	.w3(32'hba7afc86),
	.w4(32'hba840125),
	.w5(32'h398ca25d),
	.w6(32'hb9cea086),
	.w7(32'hba60d885),
	.w8(32'hb93c337b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf50f92),
	.w1(32'hbaef0810),
	.w2(32'hba05f6d1),
	.w3(32'hbb84cf19),
	.w4(32'hb9c86fc6),
	.w5(32'hbb1da3c7),
	.w6(32'hbbcd9125),
	.w7(32'hbb6f13ef),
	.w8(32'hb8655665),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a882d92),
	.w1(32'h3a10d917),
	.w2(32'h3a4e3d40),
	.w3(32'h3a6677b8),
	.w4(32'h3a87ec84),
	.w5(32'h38bcf1aa),
	.w6(32'h398b1431),
	.w7(32'h3a2d26df),
	.w8(32'h39d86f95),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb590f63),
	.w1(32'hba342e92),
	.w2(32'hb900bc98),
	.w3(32'hbb18cec0),
	.w4(32'hbb7bdf9d),
	.w5(32'h3a4d9a82),
	.w6(32'hbac5358c),
	.w7(32'hb8db16d5),
	.w8(32'hba60c57c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule