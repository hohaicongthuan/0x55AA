module layer_10_featuremap_348(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07275),
	.w1(32'hbb9fecdb),
	.w2(32'hbb8b6022),
	.w3(32'hbb4ee40f),
	.w4(32'hbb87e056),
	.w5(32'hbb4cd090),
	.w6(32'hbb79175a),
	.w7(32'hbb9da5bf),
	.w8(32'hbb0109c3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0b512),
	.w1(32'hb98965af),
	.w2(32'hba773de7),
	.w3(32'h3a6f231f),
	.w4(32'h3ac0ad5a),
	.w5(32'h3aab4c95),
	.w6(32'h3ae82b5d),
	.w7(32'hba8e4c83),
	.w8(32'h3a279c4c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f49dd),
	.w1(32'h3a43ba14),
	.w2(32'hbb093a25),
	.w3(32'h3ad03c04),
	.w4(32'hb9ac5b05),
	.w5(32'h3b019040),
	.w6(32'hbb7d6f43),
	.w7(32'hb9588b1b),
	.w8(32'h3ae05398),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fbe72),
	.w1(32'h3b96674e),
	.w2(32'h3b7168ce),
	.w3(32'h3b4d8a82),
	.w4(32'h3b27a070),
	.w5(32'hbb2f9e73),
	.w6(32'h3b454370),
	.w7(32'h3b2b674e),
	.w8(32'h3aa70d26),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa353a),
	.w1(32'hbb8a2af3),
	.w2(32'hbbea1cce),
	.w3(32'hbbaa18d3),
	.w4(32'hbbccb6bf),
	.w5(32'h3a62d86b),
	.w6(32'hba82bdf8),
	.w7(32'hbb59415e),
	.w8(32'hb9f03cb7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a094949),
	.w1(32'hb95b73df),
	.w2(32'hba05a686),
	.w3(32'h3a2807ce),
	.w4(32'h3a5170b4),
	.w5(32'hb989f05d),
	.w6(32'h3a351c9b),
	.w7(32'h3a289b4d),
	.w8(32'h37f755a3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b232836),
	.w1(32'h3abd7c81),
	.w2(32'hb97972d4),
	.w3(32'h3a74251a),
	.w4(32'h3ac5c40f),
	.w5(32'h3b4145d3),
	.w6(32'h3aae63ab),
	.w7(32'h39eb014a),
	.w8(32'h3a83a362),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e99bf),
	.w1(32'h3ab8b7fa),
	.w2(32'h3bb3e193),
	.w3(32'h3b706046),
	.w4(32'h3ad2d2e9),
	.w5(32'h3b2824a3),
	.w6(32'h3b7a4fd0),
	.w7(32'h3b42824e),
	.w8(32'h3aac844d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e2f01),
	.w1(32'h3a190c13),
	.w2(32'h3862a9a2),
	.w3(32'h3b47ae57),
	.w4(32'h3b280c00),
	.w5(32'h3a9eacf3),
	.w6(32'h3af66cbc),
	.w7(32'h3ae632ce),
	.w8(32'h3a0340ae),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b677c20),
	.w1(32'h3aa52996),
	.w2(32'h3a89cf1a),
	.w3(32'h3b3fa1af),
	.w4(32'h3b22b524),
	.w5(32'h3b69796b),
	.w6(32'h3b07ed34),
	.w7(32'h3ab6ee9e),
	.w8(32'h3a33be13),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4d76c),
	.w1(32'hb90afa6b),
	.w2(32'hbb1d6a56),
	.w3(32'h3aa94d0c),
	.w4(32'h390ef53c),
	.w5(32'h3ba10775),
	.w6(32'h3a8dc8dd),
	.w7(32'hba5a8584),
	.w8(32'h3b8866bd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1bdf3),
	.w1(32'hb9765f5c),
	.w2(32'hbb0b0c8c),
	.w3(32'h3bd5648e),
	.w4(32'h3a1d573a),
	.w5(32'hba9a34e0),
	.w6(32'hba4f0556),
	.w7(32'hbad1dd2c),
	.w8(32'hba9f48bc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97244bd),
	.w1(32'hb9528ca9),
	.w2(32'hbab71edc),
	.w3(32'hba200d73),
	.w4(32'hba541ae4),
	.w5(32'hb9876113),
	.w6(32'h3a723a4e),
	.w7(32'h364842d6),
	.w8(32'hba5a2514),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9425717),
	.w1(32'h3ad82b22),
	.w2(32'hb9103758),
	.w3(32'hb9af1b65),
	.w4(32'hb90b9dba),
	.w5(32'h3ba60a5e),
	.w6(32'hb9c35db4),
	.w7(32'hbac25f24),
	.w8(32'h3b259dab),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858700b),
	.w1(32'h39912137),
	.w2(32'hb5af1a57),
	.w3(32'h3b4cd177),
	.w4(32'hb94dc616),
	.w5(32'hbb02f21d),
	.w6(32'h3ad8be73),
	.w7(32'h3ab51d09),
	.w8(32'hbb4967a0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1bd7f),
	.w1(32'hba3610b3),
	.w2(32'hb9b62131),
	.w3(32'hba14837c),
	.w4(32'hb9e455f0),
	.w5(32'hb8a244a7),
	.w6(32'hba59d6e9),
	.w7(32'hb9e2354d),
	.w8(32'hbaaa69a6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9ebb6),
	.w1(32'hbaa32bfc),
	.w2(32'hbab44870),
	.w3(32'h3a0b6a15),
	.w4(32'h3a9d084f),
	.w5(32'h39b4da64),
	.w6(32'h3a48588c),
	.w7(32'h39e572db),
	.w8(32'hb9de70e4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa1064),
	.w1(32'h3b2841b0),
	.w2(32'h3b00e4b5),
	.w3(32'h3b505a73),
	.w4(32'h3a89db2e),
	.w5(32'h3b8d52c4),
	.w6(32'h3b47a667),
	.w7(32'h3aa0a5c0),
	.w8(32'h3b70b741),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86813a),
	.w1(32'h39b74835),
	.w2(32'h3b3d1a76),
	.w3(32'hb9b3b1cd),
	.w4(32'h3a43d060),
	.w5(32'hbaaee470),
	.w6(32'h3bb72ef5),
	.w7(32'h3b6f2446),
	.w8(32'hba6036e9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437002),
	.w1(32'hba762afe),
	.w2(32'hbaad19f2),
	.w3(32'hbb2fdbba),
	.w4(32'hbadbdc91),
	.w5(32'h3a05f4a1),
	.w6(32'hbb3e008c),
	.w7(32'hbb5dd0c2),
	.w8(32'hb9beb093),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef07a3),
	.w1(32'hb9afdb14),
	.w2(32'h3a3a058c),
	.w3(32'hba29d011),
	.w4(32'h3a188212),
	.w5(32'h3afa9822),
	.w6(32'hb8bff4ee),
	.w7(32'hb8cfbcc8),
	.w8(32'h3b594027),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29efc1),
	.w1(32'h3b497f76),
	.w2(32'h3b581109),
	.w3(32'h39f7bf6c),
	.w4(32'h3ad948e7),
	.w5(32'h3b051c66),
	.w6(32'h3b0f7d47),
	.w7(32'h3b55826e),
	.w8(32'h399c05de),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78107),
	.w1(32'h3b981104),
	.w2(32'h3b550337),
	.w3(32'h3b8a541e),
	.w4(32'h3b864029),
	.w5(32'h3bb9fbcc),
	.w6(32'h3b3d9a04),
	.w7(32'h3b917215),
	.w8(32'h3b6cd08f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac97cb7),
	.w1(32'h3b480100),
	.w2(32'h3b73b125),
	.w3(32'h3ace3ea6),
	.w4(32'h3b7bbbbc),
	.w5(32'hbadb3c2d),
	.w6(32'h3a4f1fa6),
	.w7(32'h3b384f62),
	.w8(32'hbae43fff),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075982),
	.w1(32'hbaac11ef),
	.w2(32'hbae90ae8),
	.w3(32'hbaa981fc),
	.w4(32'hbadd7885),
	.w5(32'h3a7f4a47),
	.w6(32'hbb40a56a),
	.w7(32'hbab5be29),
	.w8(32'h3a0d97b9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68bea6),
	.w1(32'h3b02a2cb),
	.w2(32'h3ab90c37),
	.w3(32'h3b44f7de),
	.w4(32'h3a9f919e),
	.w5(32'h39d6bd8a),
	.w6(32'h3b4c6cfe),
	.w7(32'h3b4e9141),
	.w8(32'h3b0c3cec),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadcf65),
	.w1(32'h3ae83d9d),
	.w2(32'h3b074d7d),
	.w3(32'h3ab2cd83),
	.w4(32'h3ab6cd5f),
	.w5(32'hbaea13de),
	.w6(32'h3b9a3a99),
	.w7(32'h3b88efca),
	.w8(32'hbb0d8e65),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d347c),
	.w1(32'hbb8b2caf),
	.w2(32'hbb6047c9),
	.w3(32'hbaf19a7b),
	.w4(32'hbab14593),
	.w5(32'hbac46d69),
	.w6(32'hbaf1b570),
	.w7(32'hbacdf31c),
	.w8(32'h39eac22a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1e55),
	.w1(32'h394267b8),
	.w2(32'hbb12180f),
	.w3(32'hbac96715),
	.w4(32'hbb316b32),
	.w5(32'hbb0fb29d),
	.w6(32'hbaa6f264),
	.w7(32'hbafb2551),
	.w8(32'hbb7993d8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3fd31),
	.w1(32'h3a2b7835),
	.w2(32'hba42da8f),
	.w3(32'h3b254629),
	.w4(32'h39be9ff5),
	.w5(32'hbb06730d),
	.w6(32'hb8a83cfe),
	.w7(32'hb9476848),
	.w8(32'hbb2255b5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d9eb5),
	.w1(32'hbb8a85ad),
	.w2(32'hbabe614a),
	.w3(32'hbbb7e3e7),
	.w4(32'hbb87c486),
	.w5(32'h3b6c4b71),
	.w6(32'hbb8d3b24),
	.w7(32'hbb8709c8),
	.w8(32'h385cd042),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35497),
	.w1(32'hbad64d87),
	.w2(32'hbac15590),
	.w3(32'h3b413f66),
	.w4(32'h3b5ef10d),
	.w5(32'hbbd713d8),
	.w6(32'hbbb2ee4b),
	.w7(32'h3a9935c8),
	.w8(32'hbb69268a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34ddb6),
	.w1(32'hba6125ca),
	.w2(32'h3ba02239),
	.w3(32'hbb5c2ca9),
	.w4(32'h399a9a58),
	.w5(32'hbad843ba),
	.w6(32'h3b93df57),
	.w7(32'h3b8d5bed),
	.w8(32'hba34ad0a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8accf3),
	.w1(32'hbb0bab34),
	.w2(32'h375a4f80),
	.w3(32'h3add876c),
	.w4(32'h3ae7e35d),
	.w5(32'hbb148e21),
	.w6(32'h3a2e080f),
	.w7(32'h3b07b5e7),
	.w8(32'h3a98e79c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88fb95),
	.w1(32'h3b271ac2),
	.w2(32'h3acd42d8),
	.w3(32'hb9c775e3),
	.w4(32'h3a4a605b),
	.w5(32'hb9e164d7),
	.w6(32'hbafd650f),
	.w7(32'hb8ed34cb),
	.w8(32'hbb17a761),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ca539),
	.w1(32'hbb8b9ddb),
	.w2(32'hbb747a77),
	.w3(32'hba2e33b8),
	.w4(32'hba29083f),
	.w5(32'hbb8145ff),
	.w6(32'hba3768ef),
	.w7(32'hbb3df27e),
	.w8(32'h3b4c9e21),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5da60),
	.w1(32'h3b23dce9),
	.w2(32'h3ba7c9fe),
	.w3(32'hbaba682e),
	.w4(32'hba61b207),
	.w5(32'h3a4e6f4a),
	.w6(32'h3bc4871f),
	.w7(32'h3bc750aa),
	.w8(32'hbb13c9a4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe213),
	.w1(32'hbb884710),
	.w2(32'hbbb80c17),
	.w3(32'h380a6ac1),
	.w4(32'hba5b2eb3),
	.w5(32'hbbb91457),
	.w6(32'h3a32c307),
	.w7(32'hbaeab499),
	.w8(32'hbbb8be29),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2513e),
	.w1(32'hbc08465d),
	.w2(32'hbbfc7092),
	.w3(32'hbb837e65),
	.w4(32'hbb816d19),
	.w5(32'hbbd0a83e),
	.w6(32'hbbd6e502),
	.w7(32'hbb718db0),
	.w8(32'hbb62cec3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39822a7f),
	.w1(32'hbae430c5),
	.w2(32'hbaf7ca0d),
	.w3(32'hbbad137b),
	.w4(32'hbb67de7c),
	.w5(32'hba346dab),
	.w6(32'hbb8b2331),
	.w7(32'hbb1737c5),
	.w8(32'h3b01a91e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ac27c),
	.w1(32'h3a5c0af3),
	.w2(32'hbaddcba8),
	.w3(32'h39212ca8),
	.w4(32'hbb061460),
	.w5(32'h3b408c64),
	.w6(32'hb98b2474),
	.w7(32'hbabcc586),
	.w8(32'h3b3d49c4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45b57d),
	.w1(32'h3b68e92e),
	.w2(32'h3a9bb0f4),
	.w3(32'h3b6b2b57),
	.w4(32'h3afab9b3),
	.w5(32'h39abd2c5),
	.w6(32'h3b6ff63c),
	.w7(32'h3b6acb67),
	.w8(32'hbad4ff26),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9902c59),
	.w1(32'hba8bde1e),
	.w2(32'hb911fa40),
	.w3(32'h3b5791ef),
	.w4(32'h3b17455b),
	.w5(32'h3a8f1c09),
	.w6(32'h3a68f61e),
	.w7(32'h3a22cfbe),
	.w8(32'hbaed39d7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d7ece),
	.w1(32'hb96ebe28),
	.w2(32'hb9fb3a4f),
	.w3(32'h3bd1c100),
	.w4(32'h3b7df7e3),
	.w5(32'h3bd9425e),
	.w6(32'h3bc0ba47),
	.w7(32'hbad14f46),
	.w8(32'h3c268d1b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c220d35),
	.w1(32'h3c44fcf6),
	.w2(32'h3c2b1cf9),
	.w3(32'h3c28b534),
	.w4(32'h3c113a28),
	.w5(32'h3a7bff9f),
	.w6(32'h3c6b1822),
	.w7(32'h3c583d8c),
	.w8(32'h3a93b663),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c2e9),
	.w1(32'h3a7fc95f),
	.w2(32'h3b0eb780),
	.w3(32'h3a32a259),
	.w4(32'h3aa032ce),
	.w5(32'h3aa8dbb8),
	.w6(32'h3a93aeee),
	.w7(32'h3af98916),
	.w8(32'h3b2e452e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585533),
	.w1(32'h3ac27447),
	.w2(32'h3a840517),
	.w3(32'h3ad9f72f),
	.w4(32'h397d2bfd),
	.w5(32'h3b0e3c2b),
	.w6(32'h3b0d6140),
	.w7(32'h3b74a95e),
	.w8(32'h3b0f7fd3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8d889),
	.w1(32'h3baca851),
	.w2(32'h3b8e0b4c),
	.w3(32'h3bbc5dc8),
	.w4(32'h3bd2a928),
	.w5(32'h3b507cab),
	.w6(32'h3ba0b2d9),
	.w7(32'h3ba6e8ea),
	.w8(32'h3ac92158),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb247204),
	.w1(32'hbb085be2),
	.w2(32'hba8c35f4),
	.w3(32'hb6ca1017),
	.w4(32'h38b033c2),
	.w5(32'h3b007376),
	.w6(32'hbaca5cbc),
	.w7(32'hba001883),
	.w8(32'h3b600333),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180a88),
	.w1(32'h3b512804),
	.w2(32'h3b3e59c7),
	.w3(32'h3a3d4e4c),
	.w4(32'h3a8e2a89),
	.w5(32'h3ae85a02),
	.w6(32'h3ad99e80),
	.w7(32'h3b50cd68),
	.w8(32'hb96efa74),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf6c87),
	.w1(32'h39a62480),
	.w2(32'hbb192a76),
	.w3(32'hba838de4),
	.w4(32'hb9ffea1d),
	.w5(32'h3b132e5c),
	.w6(32'h3acce43f),
	.w7(32'hba140657),
	.w8(32'h3b803432),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c0c1),
	.w1(32'h3b62fbaf),
	.w2(32'h3b99f56c),
	.w3(32'h3bf1316c),
	.w4(32'h3b7521b9),
	.w5(32'h3b722327),
	.w6(32'h3c04cba4),
	.w7(32'h3a8c1cca),
	.w8(32'h3a9b9f44),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1008),
	.w1(32'h3acc952a),
	.w2(32'h3a2d6e9b),
	.w3(32'h3b12f3bc),
	.w4(32'hbab89ab4),
	.w5(32'hbb3efc6a),
	.w6(32'hb983510d),
	.w7(32'hba18f79a),
	.w8(32'hba3f5b18),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0af836),
	.w1(32'hb92827e3),
	.w2(32'hb98dba39),
	.w3(32'h3ac2fcac),
	.w4(32'hba0da39c),
	.w5(32'hb9117b2d),
	.w6(32'hbb136ccd),
	.w7(32'hba9555a4),
	.w8(32'hba8baad0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2492b7),
	.w1(32'hba7fb2c7),
	.w2(32'hba18a001),
	.w3(32'hbb39af1e),
	.w4(32'hb8ac080a),
	.w5(32'hbb05df8a),
	.w6(32'hbb07fb2a),
	.w7(32'hbb405842),
	.w8(32'hba64fd85),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5490fb),
	.w1(32'h3b1c26b9),
	.w2(32'hb9e34a93),
	.w3(32'hb9d06475),
	.w4(32'h3b70aa31),
	.w5(32'hbaac89a9),
	.w6(32'hba8c2b4d),
	.w7(32'hba1270db),
	.w8(32'hba3be7cc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af854b),
	.w1(32'h38ea0ad6),
	.w2(32'hba402fb7),
	.w3(32'hbb15f1ef),
	.w4(32'hba3a9b25),
	.w5(32'hbae8fa26),
	.w6(32'hbb0bbafc),
	.w7(32'hba528fd7),
	.w8(32'hbb186810),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f4e0),
	.w1(32'hbad4ae4a),
	.w2(32'hbb89e0e0),
	.w3(32'hba35d9a8),
	.w4(32'hb9cdaeef),
	.w5(32'h3b20e403),
	.w6(32'hbb0da9de),
	.w7(32'hbb88d03a),
	.w8(32'h3b351b83),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff8795),
	.w1(32'h3b2a5c64),
	.w2(32'h3a8b1b25),
	.w3(32'h3b1713ed),
	.w4(32'h3ac74e72),
	.w5(32'hba15e3f5),
	.w6(32'h3ac71ba4),
	.w7(32'h3b1ec984),
	.w8(32'hbb8180b3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e08b6),
	.w1(32'hbaef8b91),
	.w2(32'h3a178826),
	.w3(32'hbae5a656),
	.w4(32'h3aacb598),
	.w5(32'hba1bb2de),
	.w6(32'hbb1c7d9f),
	.w7(32'h399bcefb),
	.w8(32'hbad35b68),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6038),
	.w1(32'hbb3b7194),
	.w2(32'hba9ad1f1),
	.w3(32'hb82d9cc8),
	.w4(32'hb9fa1941),
	.w5(32'h3b7aa2c8),
	.w6(32'hbad64844),
	.w7(32'hbab49194),
	.w8(32'h3b1397dd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c6e46),
	.w1(32'h3aeb3496),
	.w2(32'h3a75e787),
	.w3(32'h3ab95911),
	.w4(32'h3ae83215),
	.w5(32'hbaef19cb),
	.w6(32'h3b6d14a2),
	.w7(32'h3ad1074a),
	.w8(32'h3b10adbe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0b98f),
	.w1(32'hb933780b),
	.w2(32'h384b8dc9),
	.w3(32'hbb2a58d6),
	.w4(32'hba283ff0),
	.w5(32'hb9f5a1a7),
	.w6(32'h3a2df6c9),
	.w7(32'h3a7c87aa),
	.w8(32'h3b081207),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7c170),
	.w1(32'h3a69ccec),
	.w2(32'hba9358b8),
	.w3(32'hba106073),
	.w4(32'hb9cbd3d8),
	.w5(32'hbb42c882),
	.w6(32'hba5d1b83),
	.w7(32'h3917d5b3),
	.w8(32'hbadef047),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37817468),
	.w1(32'h3a31b9c7),
	.w2(32'hb98d2399),
	.w3(32'hba680ab2),
	.w4(32'h3b1863fb),
	.w5(32'hbafbeec6),
	.w6(32'hbb395279),
	.w7(32'hbad74d7d),
	.w8(32'hbb231e46),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa50d7b),
	.w1(32'hbaa8f381),
	.w2(32'hb9af3de9),
	.w3(32'hba4b5361),
	.w4(32'hba55031d),
	.w5(32'h3b4f187a),
	.w6(32'hbb22667d),
	.w7(32'hbb25f43d),
	.w8(32'h3b6b9a8e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae94568),
	.w1(32'hba23d6f3),
	.w2(32'hb9898e67),
	.w3(32'h3b20d0d5),
	.w4(32'hba1c6549),
	.w5(32'h3b2ab697),
	.w6(32'h3ad61d5e),
	.w7(32'hba79382f),
	.w8(32'hba4445d7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80be00e),
	.w1(32'hba0601ba),
	.w2(32'hba6b6f50),
	.w3(32'hb86cc1d6),
	.w4(32'hbab3bf26),
	.w5(32'hbb51eb50),
	.w6(32'hb95a80ec),
	.w7(32'hb9f6fee8),
	.w8(32'hbb92c5ba),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccbe32),
	.w1(32'h3a871156),
	.w2(32'hba48382d),
	.w3(32'h3a5347fd),
	.w4(32'h3aa194a7),
	.w5(32'h3ae441cf),
	.w6(32'h3aceca2b),
	.w7(32'h39059047),
	.w8(32'h39570860),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb267c1d),
	.w1(32'hbb94aa22),
	.w2(32'hbbea5d67),
	.w3(32'h3b76f904),
	.w4(32'hbaadb8d9),
	.w5(32'hbabc8841),
	.w6(32'h3b3dd43d),
	.w7(32'hbb31cf39),
	.w8(32'h3ad55844),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b429eb2),
	.w1(32'h3b968711),
	.w2(32'h3bcb5d67),
	.w3(32'h3b944426),
	.w4(32'h3b1b2bc2),
	.w5(32'h3aa8d749),
	.w6(32'h3c148669),
	.w7(32'h3bb5b779),
	.w8(32'h3a6c000d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8cb8),
	.w1(32'hb9ac9611),
	.w2(32'h3a7aa11e),
	.w3(32'hb9f77521),
	.w4(32'hba4fbd94),
	.w5(32'h3a95ecf2),
	.w6(32'hba08ee16),
	.w7(32'hba0218d3),
	.w8(32'hbb12dbc8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0be366),
	.w1(32'hba4b86eb),
	.w2(32'hb8baf15a),
	.w3(32'h3908076b),
	.w4(32'h39c8808d),
	.w5(32'hbb9b44a5),
	.w6(32'hbb39a792),
	.w7(32'hbb478204),
	.w8(32'hbba1ddf9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c77e),
	.w1(32'hbb865d51),
	.w2(32'hbb2469d9),
	.w3(32'h3a3db62b),
	.w4(32'hba6c3583),
	.w5(32'h3ac70351),
	.w6(32'hba99f96c),
	.w7(32'h394ede6f),
	.w8(32'h3a4cd88c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77554ce),
	.w1(32'hbb30db8d),
	.w2(32'hbb592b33),
	.w3(32'hb8c3e765),
	.w4(32'hbab46f36),
	.w5(32'hbaf06f8a),
	.w6(32'hbb123ad0),
	.w7(32'hbb5c2391),
	.w8(32'hbb906b53),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74f504),
	.w1(32'hbb01e252),
	.w2(32'hbaab578c),
	.w3(32'hba31d91d),
	.w4(32'hba047196),
	.w5(32'h3b35ac1f),
	.w6(32'hba763730),
	.w7(32'hba9c35ae),
	.w8(32'h3a5a245c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75b936),
	.w1(32'h3b10d31e),
	.w2(32'h3b27d371),
	.w3(32'h3b221708),
	.w4(32'h3a98c52b),
	.w5(32'h3b5d62f7),
	.w6(32'h3b39cd97),
	.w7(32'h3b42f67f),
	.w8(32'h3ba18059),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35b67e),
	.w1(32'h3b2ff6d6),
	.w2(32'h3a539325),
	.w3(32'h3b8ce56b),
	.w4(32'h39c3ed0f),
	.w5(32'h3af36195),
	.w6(32'h3bda7591),
	.w7(32'hb8e7c890),
	.w8(32'hbb10b2e6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383bd503),
	.w1(32'hbb61fa6e),
	.w2(32'h3a19255a),
	.w3(32'hb98e95ad),
	.w4(32'hba2d5a43),
	.w5(32'h3a919716),
	.w6(32'hbb87f707),
	.w7(32'hbb05ab20),
	.w8(32'h3a7d45b1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0066),
	.w1(32'hba5d3193),
	.w2(32'h36b5e4a5),
	.w3(32'hb9fb0b9d),
	.w4(32'h390156dc),
	.w5(32'h3b978274),
	.w6(32'hb9069c92),
	.w7(32'h3958b00f),
	.w8(32'h3b02adeb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86c2c0),
	.w1(32'h3a9dc166),
	.w2(32'h3b1476ce),
	.w3(32'h3a73c97b),
	.w4(32'hb919bd45),
	.w5(32'hbb113511),
	.w6(32'hba8adc02),
	.w7(32'hba92dd91),
	.w8(32'hbb5c646f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a0a0),
	.w1(32'hbb597827),
	.w2(32'hbb501b89),
	.w3(32'hb8f04485),
	.w4(32'hba310961),
	.w5(32'h3a168fd3),
	.w6(32'hbab51a8e),
	.w7(32'h38ab8053),
	.w8(32'hbafc1ec7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafac6bd),
	.w1(32'hbae7e39b),
	.w2(32'hbb1d1fd9),
	.w3(32'hbb30d15f),
	.w4(32'hba210443),
	.w5(32'h395db848),
	.w6(32'hba8ffc86),
	.w7(32'hba5bf254),
	.w8(32'h396e2c4b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a033592),
	.w1(32'hbb5ad837),
	.w2(32'hbb8c965a),
	.w3(32'hbb2702f3),
	.w4(32'hbb8f6394),
	.w5(32'h3a3e2743),
	.w6(32'hbb4f72c4),
	.w7(32'hbb8de005),
	.w8(32'h39abf1cc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e5edc),
	.w1(32'hba9cd650),
	.w2(32'hbacc7f28),
	.w3(32'hbab06e1a),
	.w4(32'hb96515c6),
	.w5(32'h3a281b82),
	.w6(32'h3a776472),
	.w7(32'h394a4c3e),
	.w8(32'hb97dbdcc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad762cc),
	.w1(32'hbb3766b3),
	.w2(32'hbaf4f29e),
	.w3(32'hbb38d7af),
	.w4(32'hbb2765a1),
	.w5(32'h3b01b974),
	.w6(32'hbb0c2f46),
	.w7(32'hbaf6fcaf),
	.w8(32'h3b0d460d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a7dd6),
	.w1(32'hbaadf1f6),
	.w2(32'hbb1c8ac5),
	.w3(32'h3b4e8dd8),
	.w4(32'hba6d7767),
	.w5(32'hb9e8e312),
	.w6(32'h3a204c4c),
	.w7(32'h39bb8c3a),
	.w8(32'hb9ee6e7f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94fead),
	.w1(32'hbaa22c61),
	.w2(32'hba97db5d),
	.w3(32'hba3bf4d9),
	.w4(32'hba55ff91),
	.w5(32'hbacf98eb),
	.w6(32'hba425dc3),
	.w7(32'hb9fc82d0),
	.w8(32'hbad46b8c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8d327),
	.w1(32'hb98672d3),
	.w2(32'hb91ad314),
	.w3(32'h39e73257),
	.w4(32'h39c55af8),
	.w5(32'h3a84510f),
	.w6(32'h3aab3343),
	.w7(32'h3a3faf59),
	.w8(32'h3a0c535f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147b6f),
	.w1(32'h3b8be6d1),
	.w2(32'h3b5ad476),
	.w3(32'h3b24c40d),
	.w4(32'h3a65c786),
	.w5(32'h3b60a628),
	.w6(32'h3b03daeb),
	.w7(32'h3b3f856e),
	.w8(32'h3b9a477e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f700cb),
	.w1(32'hbac2f69e),
	.w2(32'hbb052d9f),
	.w3(32'hba8c921b),
	.w4(32'h3af37e58),
	.w5(32'hba6f1848),
	.w6(32'hba9092f0),
	.w7(32'hb8c66d81),
	.w8(32'hbb6ef689),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b9721),
	.w1(32'h3b81a613),
	.w2(32'hbb1796b2),
	.w3(32'h3b83b63b),
	.w4(32'h3a9a8899),
	.w5(32'h3ad3e0ac),
	.w6(32'h3b9686dd),
	.w7(32'h39ce17a3),
	.w8(32'h3b8314e4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff1d8b),
	.w1(32'h3a93952d),
	.w2(32'hbb5115f7),
	.w3(32'h3afc32f2),
	.w4(32'h3b3d19be),
	.w5(32'hbb61fe03),
	.w6(32'h3a5d3910),
	.w7(32'h3b817f18),
	.w8(32'h3974f54d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc0757),
	.w1(32'h3ba4073a),
	.w2(32'h3a32a35d),
	.w3(32'h3b654b4c),
	.w4(32'h3a450064),
	.w5(32'h397ea4f7),
	.w6(32'h3ba3c811),
	.w7(32'h3b2efd58),
	.w8(32'hbad49462),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a689ff),
	.w1(32'hba761472),
	.w2(32'h39e4ca44),
	.w3(32'hb9f91118),
	.w4(32'h3a75a1ab),
	.w5(32'h3bc5fbee),
	.w6(32'hba5d81fe),
	.w7(32'hba161920),
	.w8(32'h3a7869c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199216),
	.w1(32'hba66ea73),
	.w2(32'h3a791749),
	.w3(32'h3c0f3d46),
	.w4(32'h3bc6dc32),
	.w5(32'hbb3b1f93),
	.w6(32'hba6c1ccc),
	.w7(32'h3afe6017),
	.w8(32'hbb9c4d7c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5cbe8),
	.w1(32'hbb5c6b63),
	.w2(32'hbac83160),
	.w3(32'hbbad61da),
	.w4(32'hbaaf02c7),
	.w5(32'hbb78614d),
	.w6(32'hbc0680ef),
	.w7(32'hbb3b24f8),
	.w8(32'hbba2803c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9abd4e),
	.w1(32'h3b9bf79c),
	.w2(32'h3bc36dc1),
	.w3(32'hb95c560f),
	.w4(32'h3b571b71),
	.w5(32'h3ba1399a),
	.w6(32'h3b1f592b),
	.w7(32'h3bbc883f),
	.w8(32'h3bca8141),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c752b),
	.w1(32'h3b840741),
	.w2(32'h39bc061d),
	.w3(32'h3bafe7af),
	.w4(32'h3aedd91f),
	.w5(32'hbc07a0d6),
	.w6(32'h3bd494ca),
	.w7(32'h3b1dd3ac),
	.w8(32'hbb67515e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e5c23),
	.w1(32'hba7b982e),
	.w2(32'hb9e37c5e),
	.w3(32'hbc32d26c),
	.w4(32'hbc337fc5),
	.w5(32'hba7d78a6),
	.w6(32'hbb843142),
	.w7(32'hbbba42c2),
	.w8(32'h3b2b2427),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2158e2),
	.w1(32'h3b4948fd),
	.w2(32'hbb145a87),
	.w3(32'h3b5925c2),
	.w4(32'hbb6173a8),
	.w5(32'hbb9a1b9c),
	.w6(32'h3bc8c20e),
	.w7(32'h3aa36734),
	.w8(32'hbb85da8d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9bc24),
	.w1(32'hbb4d0d04),
	.w2(32'hbae5e00b),
	.w3(32'hb93401e8),
	.w4(32'h3b0edecb),
	.w5(32'h3b5dfdf5),
	.w6(32'h3b169939),
	.w7(32'h3a423607),
	.w8(32'hbaaf5d7a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154c3b),
	.w1(32'h39788566),
	.w2(32'h3aa237bf),
	.w3(32'h3aec5375),
	.w4(32'hba87b12e),
	.w5(32'hb9f40e26),
	.w6(32'h3ab8da11),
	.w7(32'hb9cb567c),
	.w8(32'hbb8730f3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68c7a),
	.w1(32'hbbc12dec),
	.w2(32'hbb745c32),
	.w3(32'h3b119bd5),
	.w4(32'h3a05b8af),
	.w5(32'hbaca6d61),
	.w6(32'hbb80c3be),
	.w7(32'hbb3fa2ab),
	.w8(32'hbaca6d43),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ea50a),
	.w1(32'h3bcaaa00),
	.w2(32'h3b4c6046),
	.w3(32'h3af7aeca),
	.w4(32'hbb10c9ed),
	.w5(32'hbaeb6926),
	.w6(32'h3c6f4715),
	.w7(32'h3b0de969),
	.w8(32'h3ac76466),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d369c),
	.w1(32'h3acb44fe),
	.w2(32'hb8b996a0),
	.w3(32'hbb87ae6a),
	.w4(32'hbb888733),
	.w5(32'hbbee19d0),
	.w6(32'hbb6a56e9),
	.w7(32'hbb68bb0a),
	.w8(32'hbba21ba3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a41cd1),
	.w1(32'h3b9922da),
	.w2(32'hbb821224),
	.w3(32'hbbe1d40c),
	.w4(32'hbb754739),
	.w5(32'hbabaeaf7),
	.w6(32'hbbcf971a),
	.w7(32'hbbccee8a),
	.w8(32'h3af081d7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66136b),
	.w1(32'hba9c3c24),
	.w2(32'h3b1f0ec2),
	.w3(32'hbbaa9b0e),
	.w4(32'hbb0e31c8),
	.w5(32'hbb84f068),
	.w6(32'h3a169189),
	.w7(32'h3ae38d23),
	.w8(32'hbb11330a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7ca1),
	.w1(32'hbb34e825),
	.w2(32'hbb9f360b),
	.w3(32'hbb030bdb),
	.w4(32'hbb55a8c4),
	.w5(32'h3bd2f83e),
	.w6(32'h3a0e30ad),
	.w7(32'hbb73fd9c),
	.w8(32'h3be41b1c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba82a07),
	.w1(32'h3b6594bc),
	.w2(32'h3b87c6c4),
	.w3(32'h3c01405e),
	.w4(32'h3bcc5698),
	.w5(32'hbb92c759),
	.w6(32'h3ba9db32),
	.w7(32'h3c0a7b24),
	.w8(32'h3a8fb278),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818967),
	.w1(32'h3b88dcd3),
	.w2(32'hbb862dfa),
	.w3(32'hbc00615a),
	.w4(32'hbbff2dbb),
	.w5(32'h3a4322b4),
	.w6(32'h3a965c19),
	.w7(32'hbaffcaae),
	.w8(32'h3b594f89),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a84fa),
	.w1(32'hba99635b),
	.w2(32'hbb30485f),
	.w3(32'h3ab0eebc),
	.w4(32'h3aeb61a3),
	.w5(32'h3bf2e5d3),
	.w6(32'hb91f2e09),
	.w7(32'hbb54a108),
	.w8(32'h3b9e7ed3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c24d),
	.w1(32'h3a97f0bc),
	.w2(32'hbb8e2d1a),
	.w3(32'h3b448855),
	.w4(32'h3a0dfe27),
	.w5(32'h3b403df8),
	.w6(32'h3bd8211d),
	.w7(32'h3a0ed397),
	.w8(32'hbb3281d1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92db91d),
	.w1(32'hb9007713),
	.w2(32'h3a1bb4ff),
	.w3(32'h3bad1d2e),
	.w4(32'h3b1b7593),
	.w5(32'hbc131d87),
	.w6(32'h3b19d6af),
	.w7(32'hba1cb686),
	.w8(32'hbb541ced),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb78af),
	.w1(32'h3b8e2471),
	.w2(32'h3bda43a0),
	.w3(32'hbb394794),
	.w4(32'h3b864644),
	.w5(32'hba3f5aac),
	.w6(32'hbaf5986e),
	.w7(32'h3b73fc00),
	.w8(32'h3b259599),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f563e),
	.w1(32'hbb09f355),
	.w2(32'hbb5f536e),
	.w3(32'h3921905b),
	.w4(32'hba9b4217),
	.w5(32'h3bfe6015),
	.w6(32'h3a9b05c2),
	.w7(32'hbb5ea156),
	.w8(32'h3b0e4411),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f0be6),
	.w1(32'h3a654c84),
	.w2(32'h3b107e18),
	.w3(32'h3c22f44c),
	.w4(32'h3bdb83c8),
	.w5(32'hbb9b9d13),
	.w6(32'h3b461c95),
	.w7(32'h3bcc18a5),
	.w8(32'hbb80ad25),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f12f8c),
	.w1(32'h3b2e4fd7),
	.w2(32'h3be8a0d8),
	.w3(32'hbbe9e5e9),
	.w4(32'h3a579859),
	.w5(32'h3ad6da63),
	.w6(32'h3a7cbbe2),
	.w7(32'hbb9b7114),
	.w8(32'hbb076679),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092faa),
	.w1(32'h3934e24e),
	.w2(32'hb905f7ad),
	.w3(32'h3a1eab87),
	.w4(32'hbb1e0821),
	.w5(32'h3c252a4d),
	.w6(32'hbacc0c5e),
	.w7(32'hbba68823),
	.w8(32'h3be97f8f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38871323),
	.w1(32'h3c209705),
	.w2(32'h3bd6a5a6),
	.w3(32'h3c735e93),
	.w4(32'h3c033fde),
	.w5(32'hbb256e46),
	.w6(32'h3c51188f),
	.w7(32'h3bf6090e),
	.w8(32'hbb4db3f8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb150),
	.w1(32'hbb831732),
	.w2(32'hbb88609b),
	.w3(32'h3b0da0c7),
	.w4(32'h3b5d32c3),
	.w5(32'hbb8ecd0e),
	.w6(32'h3b5fd9d4),
	.w7(32'h3a56e4a3),
	.w8(32'hbad6aba6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820678),
	.w1(32'h3b163359),
	.w2(32'hbad30e13),
	.w3(32'hbbf8e428),
	.w4(32'hbb9acb90),
	.w5(32'hbac3e32b),
	.w6(32'hba8e5a22),
	.w7(32'hbbd8fb56),
	.w8(32'hbbbf3fe8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14aa8f),
	.w1(32'hbbeba613),
	.w2(32'hbba6b369),
	.w3(32'h3c01060c),
	.w4(32'h3bf341a2),
	.w5(32'h3a5e1ecd),
	.w6(32'h3b707e0a),
	.w7(32'h3a38f73e),
	.w8(32'h3b2abc85),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e021),
	.w1(32'h3b472cdd),
	.w2(32'h3b1443d6),
	.w3(32'hbab87f00),
	.w4(32'h3b2d3ed8),
	.w5(32'h3a93ef0d),
	.w6(32'h3b0c528c),
	.w7(32'h3b81b90f),
	.w8(32'hbac78cb7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0d0f),
	.w1(32'hbba8f544),
	.w2(32'hbb6d1637),
	.w3(32'h3be2876c),
	.w4(32'h3bbf9ce5),
	.w5(32'h3a895acf),
	.w6(32'h3c1fce3a),
	.w7(32'h3bf0ba72),
	.w8(32'hbb08d7b7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a919608),
	.w1(32'hbb5ec87d),
	.w2(32'hbb91ead6),
	.w3(32'hba1db864),
	.w4(32'h3ab3944e),
	.w5(32'hbb8f2f16),
	.w6(32'hbb22db4f),
	.w7(32'hbb90485e),
	.w8(32'h3b4bae04),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0921),
	.w1(32'h3aa854fe),
	.w2(32'h3b0da6e2),
	.w3(32'hbb9f523e),
	.w4(32'hba888545),
	.w5(32'hbb93cca7),
	.w6(32'h3a0257eb),
	.w7(32'h3a801f86),
	.w8(32'hbb9ef553),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f427f),
	.w1(32'h3908c446),
	.w2(32'h3b1c6592),
	.w3(32'h3a0721e0),
	.w4(32'h3b07f91e),
	.w5(32'h3ba0d90b),
	.w6(32'hbb139932),
	.w7(32'h3b17c48c),
	.w8(32'h3bbb209c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dee65),
	.w1(32'h3b75cd03),
	.w2(32'h3b24b53b),
	.w3(32'h3b9a26f8),
	.w4(32'h3b0c444f),
	.w5(32'hba276828),
	.w6(32'h3c3b07c5),
	.w7(32'h3b6b805f),
	.w8(32'hbb49c296),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e7fb9),
	.w1(32'h3b1680a0),
	.w2(32'h3accc01f),
	.w3(32'h3865eb3a),
	.w4(32'h3b4ee2ad),
	.w5(32'hba8ab43c),
	.w6(32'h3b00e966),
	.w7(32'hbaa1f199),
	.w8(32'h3a900fa5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec638d),
	.w1(32'h3b514f9b),
	.w2(32'hbb09a277),
	.w3(32'h3a1792bb),
	.w4(32'hbb9bcbd4),
	.w5(32'hb9efb73c),
	.w6(32'hba894310),
	.w7(32'hbb920064),
	.w8(32'hbb8359e2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6c47a),
	.w1(32'hbb84954a),
	.w2(32'hbb167e3d),
	.w3(32'h3a31af22),
	.w4(32'h3b4eb971),
	.w5(32'h3911333c),
	.w6(32'hbb71f695),
	.w7(32'hbb3ec22a),
	.w8(32'h39da536b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4e6cb),
	.w1(32'hbb73bbcf),
	.w2(32'hbb991f5e),
	.w3(32'h3ae7f84a),
	.w4(32'hbb08344f),
	.w5(32'h3984d1db),
	.w6(32'h3b0d803e),
	.w7(32'h3b8179df),
	.w8(32'hb96bff77),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c6904),
	.w1(32'hbaf036ce),
	.w2(32'hb9dabaac),
	.w3(32'h3ac95ed8),
	.w4(32'h3ad4bbed),
	.w5(32'h3a3b2d4a),
	.w6(32'h3af15946),
	.w7(32'h3a9abca7),
	.w8(32'hbb340312),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaffe8),
	.w1(32'h3a1246b1),
	.w2(32'hbaf8685e),
	.w3(32'h3b4ef4f7),
	.w4(32'h3b0d63b7),
	.w5(32'h3b9a0c4a),
	.w6(32'h3b80f9da),
	.w7(32'h3a602b68),
	.w8(32'h3bb09db5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a132724),
	.w1(32'h3b0a9677),
	.w2(32'h3b10febb),
	.w3(32'hbac2d4af),
	.w4(32'hbbe905f4),
	.w5(32'h3b9729ed),
	.w6(32'h3a3dd338),
	.w7(32'hbb1d2aa7),
	.w8(32'h3b8167aa),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07e25f),
	.w1(32'h3b38ca71),
	.w2(32'hb94fc21b),
	.w3(32'h3bafe686),
	.w4(32'h3b9f15a4),
	.w5(32'hb9b9443a),
	.w6(32'h3b97be15),
	.w7(32'h3bd9e42a),
	.w8(32'hba571d1b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba317cc2),
	.w1(32'hbaae6854),
	.w2(32'hb93182a7),
	.w3(32'h3b0e43d8),
	.w4(32'h3b457db1),
	.w5(32'h39245994),
	.w6(32'h3ac2c2da),
	.w7(32'h3b0de0d5),
	.w8(32'hbb41161d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869285),
	.w1(32'hbb0ca050),
	.w2(32'hbb485f60),
	.w3(32'hba6f8631),
	.w4(32'h39c31d3f),
	.w5(32'h3a833839),
	.w6(32'hbb159c05),
	.w7(32'hbb2e930c),
	.w8(32'hbb8b2b02),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9780),
	.w1(32'h3baa19ee),
	.w2(32'h38db2435),
	.w3(32'h3ba815ab),
	.w4(32'h3aa3970f),
	.w5(32'hbaae8c48),
	.w6(32'hbafa6b3c),
	.w7(32'hbac4b438),
	.w8(32'h39dffbc6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c3bf),
	.w1(32'hbbe5aa9b),
	.w2(32'h3929aa75),
	.w3(32'hbbbdd168),
	.w4(32'hbb85c1be),
	.w5(32'hbbd58b5a),
	.w6(32'h3a98668a),
	.w7(32'h390022e0),
	.w8(32'hba9af9a5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4637cf),
	.w1(32'hbbbb0c43),
	.w2(32'hbb9e5e6b),
	.w3(32'hbbad2b92),
	.w4(32'hb9bc72c3),
	.w5(32'hbbe92af2),
	.w6(32'hbc08f276),
	.w7(32'hbbdef002),
	.w8(32'hbba7842d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9544ec),
	.w1(32'hba203595),
	.w2(32'hbbab2da7),
	.w3(32'hbba2c05b),
	.w4(32'hbb971f8f),
	.w5(32'hbb247a6e),
	.w6(32'hbb21db85),
	.w7(32'hbb88f529),
	.w8(32'hbbbaf4e9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9370f),
	.w1(32'hba0c28d5),
	.w2(32'hbb94f580),
	.w3(32'hbb19b4c5),
	.w4(32'hba57f4d1),
	.w5(32'hba311c49),
	.w6(32'hbaf333ea),
	.w7(32'hbaee0a14),
	.w8(32'h3b03a606),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6811a4),
	.w1(32'hb9d8e40c),
	.w2(32'h3b6c141d),
	.w3(32'h39ba22d8),
	.w4(32'h3a973a74),
	.w5(32'hbb8dee7e),
	.w6(32'h3ba6e698),
	.w7(32'h3b087bcb),
	.w8(32'hbb5ded15),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee2dc5),
	.w1(32'hbb312480),
	.w2(32'hbafecbd2),
	.w3(32'hbba7e34f),
	.w4(32'hbba4077c),
	.w5(32'hba5eb8cf),
	.w6(32'hbb632cb1),
	.w7(32'hbb6669dc),
	.w8(32'h3a9e01d7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8554b3),
	.w1(32'h39075608),
	.w2(32'hbb9cd72f),
	.w3(32'hba917223),
	.w4(32'h3aa5a56e),
	.w5(32'hba991e80),
	.w6(32'h3b8ec0b6),
	.w7(32'hbb0d48cf),
	.w8(32'hb7c6e18b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075d3a),
	.w1(32'h39cf791a),
	.w2(32'hba4d17c1),
	.w3(32'hbb049e0d),
	.w4(32'hba982fca),
	.w5(32'hbb22ea5b),
	.w6(32'hba71cb44),
	.w7(32'hbb8e7888),
	.w8(32'hbb88c53e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3429b5),
	.w1(32'hba8105e4),
	.w2(32'h39c05415),
	.w3(32'hbb15584c),
	.w4(32'h3a953a74),
	.w5(32'h3bcb16fa),
	.w6(32'hbb96e4f1),
	.w7(32'hbad36b8f),
	.w8(32'h3b28721b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af39264),
	.w1(32'h3a8a1ff4),
	.w2(32'h3b611826),
	.w3(32'h3c107bfe),
	.w4(32'h3b82a427),
	.w5(32'h3b9ec838),
	.w6(32'h3b932f87),
	.w7(32'h3b3466ca),
	.w8(32'hbb2f2b1f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c98f8),
	.w1(32'hba345482),
	.w2(32'h3affa89c),
	.w3(32'hb96a409b),
	.w4(32'hbb582725),
	.w5(32'hbbe85a0a),
	.w6(32'hbb5ff6d5),
	.w7(32'hbab54743),
	.w8(32'hbc0eea2a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940c88),
	.w1(32'hbb2fa3bb),
	.w2(32'hba8f44d5),
	.w3(32'hbb828d2f),
	.w4(32'hbb264647),
	.w5(32'hba521c15),
	.w6(32'hbb4c1291),
	.w7(32'hbaf1b7d3),
	.w8(32'h39deee46),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb586183),
	.w1(32'hbb48624a),
	.w2(32'hbb4dde64),
	.w3(32'h3aa9183c),
	.w4(32'h399994b6),
	.w5(32'hbb758918),
	.w6(32'h3b7b83e1),
	.w7(32'hb91104d4),
	.w8(32'hb9f4faac),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b4dc7),
	.w1(32'hb994fd44),
	.w2(32'hbb8c932d),
	.w3(32'hbbc14405),
	.w4(32'hbbb48f61),
	.w5(32'hbb828efb),
	.w6(32'h3a376eec),
	.w7(32'h39a998d7),
	.w8(32'hbb6df301),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1a06),
	.w1(32'hbac0cd81),
	.w2(32'hbb8592b2),
	.w3(32'hbab70538),
	.w4(32'hbb8c4eac),
	.w5(32'h3bcb9377),
	.w6(32'h39fe944c),
	.w7(32'hbaef8123),
	.w8(32'h3c00f8ad),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde62a3),
	.w1(32'h3b975d3c),
	.w2(32'h3b56d1fb),
	.w3(32'h3c0e8cb1),
	.w4(32'h3bc0e167),
	.w5(32'h3a9735d9),
	.w6(32'h3bf67c67),
	.w7(32'h3c2422a4),
	.w8(32'h3b46352e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c4714),
	.w1(32'h3b422257),
	.w2(32'hba5cb5b1),
	.w3(32'h3ad8d49d),
	.w4(32'h3b6d812f),
	.w5(32'hbad77e62),
	.w6(32'h3a4803ee),
	.w7(32'hba0407e6),
	.w8(32'h3aeb9076),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ffe3b),
	.w1(32'h3af49b87),
	.w2(32'h3b8612ed),
	.w3(32'hbb6fb7a6),
	.w4(32'hba04d3be),
	.w5(32'hbae0b71f),
	.w6(32'h39427713),
	.w7(32'hbb053631),
	.w8(32'h3b64c724),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054092),
	.w1(32'h3c1e4445),
	.w2(32'h3bd79173),
	.w3(32'hbbf2117a),
	.w4(32'hbb53d13a),
	.w5(32'h3b95dbb4),
	.w6(32'hba0f3ce6),
	.w7(32'h3be73a26),
	.w8(32'hbae08490),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cc826),
	.w1(32'hbb088f59),
	.w2(32'h3b47c6ee),
	.w3(32'h3c437f63),
	.w4(32'h3c347f2a),
	.w5(32'hbbf798af),
	.w6(32'hbb302131),
	.w7(32'h3b3e373a),
	.w8(32'h3a8a795f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc3be),
	.w1(32'hba9e6ba4),
	.w2(32'hbb7979e6),
	.w3(32'hbb6ac5cf),
	.w4(32'h3b2be584),
	.w5(32'hbbb65496),
	.w6(32'h3b0c9573),
	.w7(32'h3b6c366d),
	.w8(32'hbb2acae1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19186f),
	.w1(32'hbb2bb879),
	.w2(32'h3a9e3957),
	.w3(32'hbc023d5b),
	.w4(32'hbbb3e04b),
	.w5(32'h3b3029ae),
	.w6(32'hbb3817f3),
	.w7(32'hbb1a2056),
	.w8(32'hba156e80),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e38088),
	.w1(32'hbb3ee6a9),
	.w2(32'hba89b139),
	.w3(32'h3919d07c),
	.w4(32'hbb627ea0),
	.w5(32'hbc090b11),
	.w6(32'h3ac44361),
	.w7(32'hb9d79ad9),
	.w8(32'hbb4f736b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbc197),
	.w1(32'hbb4b04e0),
	.w2(32'hbbb5a5f4),
	.w3(32'hbc08ce7f),
	.w4(32'hbc0fce55),
	.w5(32'h3ac8f0ec),
	.w6(32'hbbf2456b),
	.w7(32'hbc0352a8),
	.w8(32'h3bce1ef1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7587b8),
	.w1(32'h3b07cb52),
	.w2(32'hbb44b3a1),
	.w3(32'hbbbce89a),
	.w4(32'hbb3832e3),
	.w5(32'h3baef3e8),
	.w6(32'h3c707b04),
	.w7(32'h3c096b4b),
	.w8(32'h3b687dc0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb501cf1),
	.w1(32'h3c044a0a),
	.w2(32'h3b29c119),
	.w3(32'h3c07304a),
	.w4(32'h3bf812d1),
	.w5(32'h3ae743ad),
	.w6(32'h3c47a01d),
	.w7(32'h3b8fe9b5),
	.w8(32'hba6ff9a0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68ac94),
	.w1(32'hbba55068),
	.w2(32'hbb917a47),
	.w3(32'h3adcc925),
	.w4(32'h3990f1b8),
	.w5(32'hba89504f),
	.w6(32'h3aaa7481),
	.w7(32'hb9cee30f),
	.w8(32'hbba2bba8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65f3d3),
	.w1(32'hb99e3946),
	.w2(32'hbb29f097),
	.w3(32'h3ac86fb5),
	.w4(32'hbbb840ba),
	.w5(32'hbacb099c),
	.w6(32'hbbb30104),
	.w7(32'hbbc23089),
	.w8(32'hbb30b327),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117550),
	.w1(32'h3b33a77c),
	.w2(32'h396e18ff),
	.w3(32'h3b231dae),
	.w4(32'h3b0c0345),
	.w5(32'hbb12b3e6),
	.w6(32'h3a14abd0),
	.w7(32'hba201040),
	.w8(32'h3b3c7818),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabff28e),
	.w1(32'h3a753203),
	.w2(32'hb99e104b),
	.w3(32'hbba1dbc4),
	.w4(32'hbb9a1faa),
	.w5(32'h3c852ff0),
	.w6(32'h3ad6d8da),
	.w7(32'h39e52a2d),
	.w8(32'h3c171afd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eab28),
	.w1(32'h3bec993d),
	.w2(32'hba9dbc8d),
	.w3(32'h3c4a0d85),
	.w4(32'h3c7aaf6b),
	.w5(32'hbc6742dc),
	.w6(32'h3c45cbe4),
	.w7(32'h3c2b4076),
	.w8(32'hbbcd2f67),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900811),
	.w1(32'h3ad71026),
	.w2(32'h38d36154),
	.w3(32'hbc2d3284),
	.w4(32'hbc08c765),
	.w5(32'hbb14da82),
	.w6(32'hbbd0f87f),
	.w7(32'hbc20154f),
	.w8(32'hbab50dd9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54a308),
	.w1(32'h3b39737a),
	.w2(32'h3b89344b),
	.w3(32'h3bda7159),
	.w4(32'h3ba89f0e),
	.w5(32'h3b6d7245),
	.w6(32'h3bd5b423),
	.w7(32'h3b9f8928),
	.w8(32'h3c4a6108),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c406d5e),
	.w1(32'hbab593b5),
	.w2(32'h3b6d92bb),
	.w3(32'hb90c2e4d),
	.w4(32'hbb79eeea),
	.w5(32'hbbc04386),
	.w6(32'h3a52db9b),
	.w7(32'h3b2db05f),
	.w8(32'h3b06e475),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ba952),
	.w1(32'h3c185dbd),
	.w2(32'h3c0ea3a4),
	.w3(32'hbbabae1a),
	.w4(32'hbba2e665),
	.w5(32'h3c164a2a),
	.w6(32'hba1d2efa),
	.w7(32'hba38b54c),
	.w8(32'h3b8ef4c6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad562c7),
	.w1(32'hba46e98a),
	.w2(32'hba2de3de),
	.w3(32'h3c25b090),
	.w4(32'h3c0b9c8e),
	.w5(32'hbb2184d0),
	.w6(32'h3bdd2b9a),
	.w7(32'h3bc6bbc0),
	.w8(32'hba63fb79),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb179ffd),
	.w1(32'hbba4af2b),
	.w2(32'hba2c1e46),
	.w3(32'hb9a93a32),
	.w4(32'h3b0a2adc),
	.w5(32'h3bb660df),
	.w6(32'hba737320),
	.w7(32'h3b309f12),
	.w8(32'h3af13b86),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973edd),
	.w1(32'hba0b1c1b),
	.w2(32'hbb348fc9),
	.w3(32'h3bb8e4a4),
	.w4(32'h38851f25),
	.w5(32'hba9435aa),
	.w6(32'h3bccd831),
	.w7(32'h39c4a731),
	.w8(32'h3b882a62),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20709e),
	.w1(32'hb840aa70),
	.w2(32'hbbc33b23),
	.w3(32'h3a48f504),
	.w4(32'hbaba5848),
	.w5(32'hbb95db6b),
	.w6(32'h3b95005f),
	.w7(32'hb9fe3051),
	.w8(32'hbbc94a6c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818b38),
	.w1(32'h3b7f9ad1),
	.w2(32'h3bb73581),
	.w3(32'hb9a25b63),
	.w4(32'h3b22e62f),
	.w5(32'hbb618fa0),
	.w6(32'hbbf99063),
	.w7(32'hbbc6d2f4),
	.w8(32'hbbb24751),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf66bce),
	.w1(32'hbb58a882),
	.w2(32'hbbeadb61),
	.w3(32'hba9534d3),
	.w4(32'h3a5c3bc0),
	.w5(32'hbbd4125f),
	.w6(32'hbaca2129),
	.w7(32'hbb88adfb),
	.w8(32'hba15491a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1bd9),
	.w1(32'h3b52ef83),
	.w2(32'h3ae99e78),
	.w3(32'hbc2b2baf),
	.w4(32'hbc648d55),
	.w5(32'hbacc84f9),
	.w6(32'h3a829b62),
	.w7(32'hbbcde35d),
	.w8(32'hbb52cada),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474fb3),
	.w1(32'h3a1d75b8),
	.w2(32'h3b0c4146),
	.w3(32'hb9d78860),
	.w4(32'hba284066),
	.w5(32'hbb7cf9be),
	.w6(32'hba196423),
	.w7(32'hbb07b858),
	.w8(32'hbaa8ec45),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78e44b),
	.w1(32'hbaefe357),
	.w2(32'hba6592cd),
	.w3(32'hbaa4196b),
	.w4(32'hbad4f467),
	.w5(32'h3a14038c),
	.w6(32'hba077520),
	.w7(32'h3b0c3f6b),
	.w8(32'hb86ade5f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d358bf),
	.w1(32'hbb19ce47),
	.w2(32'hbadcd8b1),
	.w3(32'h3a8f06fa),
	.w4(32'h39e4e74a),
	.w5(32'hba737160),
	.w6(32'hbacd55b2),
	.w7(32'h3af91ce7),
	.w8(32'h3b468fae),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5054),
	.w1(32'h3afd266e),
	.w2(32'h3a1038cc),
	.w3(32'hbb5ab4ca),
	.w4(32'hbb8ff7ff),
	.w5(32'h3b59fd36),
	.w6(32'h3ae75ec3),
	.w7(32'hbbbb7f23),
	.w8(32'hb9692d13),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f7bd),
	.w1(32'h3b2849f7),
	.w2(32'hbb341ab5),
	.w3(32'h3bdd03c5),
	.w4(32'h3ae4fa88),
	.w5(32'h3c1f1109),
	.w6(32'h3bda2398),
	.w7(32'h3b8619f6),
	.w8(32'h3bf0d460),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8338),
	.w1(32'hbb9fe36a),
	.w2(32'h3b66e40c),
	.w3(32'h3c925068),
	.w4(32'h3bc8b983),
	.w5(32'h3aaa0416),
	.w6(32'h3c4bf775),
	.w7(32'h3be6fb49),
	.w8(32'h3aebf377),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3597a0),
	.w1(32'hbaf84adc),
	.w2(32'hbb65bcdc),
	.w3(32'hbb4d91ae),
	.w4(32'hbb5bd556),
	.w5(32'hbb8850a5),
	.w6(32'h38d8635b),
	.w7(32'hba4b2f8d),
	.w8(32'h3aa4a9e6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83dcc1),
	.w1(32'hb98e236f),
	.w2(32'hba87adfe),
	.w3(32'hbc0a4d5e),
	.w4(32'hbbd05897),
	.w5(32'hbae97ad0),
	.w6(32'h3a479f69),
	.w7(32'hba2811ac),
	.w8(32'hbba1427f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41bd18),
	.w1(32'hbbbb6331),
	.w2(32'hbb3f9a30),
	.w3(32'hba018250),
	.w4(32'hba5c24a5),
	.w5(32'hbb36289f),
	.w6(32'h3b704a74),
	.w7(32'h3b71107a),
	.w8(32'hbaf3fbfe),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99270c7),
	.w1(32'hbb1f20a2),
	.w2(32'hbabbf42e),
	.w3(32'hbba6eb00),
	.w4(32'hbbb69225),
	.w5(32'h3abbf1e9),
	.w6(32'hbb7174c2),
	.w7(32'hbb5d51f4),
	.w8(32'hba95e2bb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fecab),
	.w1(32'hbb649924),
	.w2(32'hbac47cea),
	.w3(32'hbafb5086),
	.w4(32'hbb4ac86c),
	.w5(32'h3a174fb1),
	.w6(32'hbb375c52),
	.w7(32'hbabde916),
	.w8(32'hbbb6ead6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d97b7),
	.w1(32'hbab581ae),
	.w2(32'h38ccaf2a),
	.w3(32'h3b1fbeed),
	.w4(32'h3ab31815),
	.w5(32'hb94bfa48),
	.w6(32'h3b114270),
	.w7(32'h3a31b7a6),
	.w8(32'h3b28e4e9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575e59),
	.w1(32'hb9ca2415),
	.w2(32'hbaf8c81b),
	.w3(32'hbb34eead),
	.w4(32'hbbebe5c6),
	.w5(32'hba988f24),
	.w6(32'h3b10c5a3),
	.w7(32'hbb9e2915),
	.w8(32'h3a935f78),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f278),
	.w1(32'hbb070e08),
	.w2(32'hbb840492),
	.w3(32'h3af37e9a),
	.w4(32'h3b95c19e),
	.w5(32'hbb9f5775),
	.w6(32'hb841bdce),
	.w7(32'h3b78efaf),
	.w8(32'hbb2a6ef7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba281aaa),
	.w1(32'hba75d2a8),
	.w2(32'hbb6cfc24),
	.w3(32'hbb160bdc),
	.w4(32'hbbc1e2a6),
	.w5(32'hbbf7984e),
	.w6(32'hbb3d4e1a),
	.w7(32'hbba14ed3),
	.w8(32'h3a82c405),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a264),
	.w1(32'h3b35f0a1),
	.w2(32'h3afafbfe),
	.w3(32'hbc0c3bc9),
	.w4(32'hbbcf53e0),
	.w5(32'h3be62d3a),
	.w6(32'hbae8d010),
	.w7(32'hbb9bfd01),
	.w8(32'h3ba7f135),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb423067),
	.w1(32'h3a0371ba),
	.w2(32'hbb6a6f9b),
	.w3(32'h3c186c1c),
	.w4(32'h3c0a1f7d),
	.w5(32'hba9fe2da),
	.w6(32'h3c355a39),
	.w7(32'h3bbf7fd9),
	.w8(32'h3a21ff30),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967196d),
	.w1(32'hbb7911d0),
	.w2(32'hbb80c0ae),
	.w3(32'hbbd3af43),
	.w4(32'hbb860fdc),
	.w5(32'h3bbba452),
	.w6(32'hbbc2c5db),
	.w7(32'hbbdb1d45),
	.w8(32'h388012c6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ff025),
	.w1(32'hba0ec71a),
	.w2(32'hbafea5d8),
	.w3(32'h3bfbc891),
	.w4(32'h3bbe337c),
	.w5(32'hb9e7ddf0),
	.w6(32'h3b854d1c),
	.w7(32'h3b3db2ea),
	.w8(32'h3aa68a8c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3948),
	.w1(32'h3baba77c),
	.w2(32'h3b96a1e9),
	.w3(32'hbb6b894f),
	.w4(32'hb9d3f117),
	.w5(32'h3a6f8021),
	.w6(32'h3b1f733c),
	.w7(32'h3b546c2f),
	.w8(32'h397661f5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db226),
	.w1(32'h3b13f4da),
	.w2(32'hbb8e508c),
	.w3(32'h3a6a74f8),
	.w4(32'hbaae2fd0),
	.w5(32'hba54ec72),
	.w6(32'h3b818c66),
	.w7(32'hbb6784df),
	.w8(32'hbb029046),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa33937),
	.w1(32'hbb9af4d4),
	.w2(32'hb90d8b30),
	.w3(32'hba1feda3),
	.w4(32'h3b0ce260),
	.w5(32'h3aad3bd2),
	.w6(32'hbbccb036),
	.w7(32'h3a789280),
	.w8(32'hbb4a85b4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06fca9),
	.w1(32'hbaf93875),
	.w2(32'hbb5e2b37),
	.w3(32'h3934247c),
	.w4(32'hbb2cbeea),
	.w5(32'hbc123175),
	.w6(32'h3aa5429c),
	.w7(32'hbaa0f160),
	.w8(32'hbc117979),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96090a),
	.w1(32'hbb7b69d0),
	.w2(32'hbaaab4f7),
	.w3(32'hbbb15b1e),
	.w4(32'hbb9434de),
	.w5(32'h39a8d962),
	.w6(32'hbbfbf6d9),
	.w7(32'hbbf8ba91),
	.w8(32'h3abf6bb0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca4e8d),
	.w1(32'hbae4feaf),
	.w2(32'hbb64f7b4),
	.w3(32'hbb4c49c4),
	.w4(32'hbbbd7698),
	.w5(32'hbb0e05c6),
	.w6(32'hbb2c9e68),
	.w7(32'hbba2b231),
	.w8(32'h3ad43222),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d767c),
	.w1(32'hbaff02c4),
	.w2(32'hba43708d),
	.w3(32'hbaf18ae9),
	.w4(32'hbb1752dc),
	.w5(32'h3bd4af29),
	.w6(32'h3b1b434f),
	.w7(32'h38b3f611),
	.w8(32'h3b0201e4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2117),
	.w1(32'h39f83754),
	.w2(32'h3a765d3c),
	.w3(32'h3bc0189e),
	.w4(32'h3b17ec22),
	.w5(32'hba7086fa),
	.w6(32'hbb5e0eed),
	.w7(32'hbb613d19),
	.w8(32'hbaaf1376),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b0a0b),
	.w1(32'hbae34e30),
	.w2(32'hbb1c7c99),
	.w3(32'hbb552555),
	.w4(32'hbb0b95e0),
	.w5(32'h3b8844cb),
	.w6(32'hba95612d),
	.w7(32'hba0e0336),
	.w8(32'hbabb8a97),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cf7f),
	.w1(32'hbab645f7),
	.w2(32'hba8c7f03),
	.w3(32'h3afd7c82),
	.w4(32'hbadba10d),
	.w5(32'hbc13ed4d),
	.w6(32'hbb4b6970),
	.w7(32'hbbc6c431),
	.w8(32'hbc33f22b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bd5ff),
	.w1(32'hbc0d6ae0),
	.w2(32'hbc02a703),
	.w3(32'hbb55f94f),
	.w4(32'hbad9b808),
	.w5(32'h3b48ea68),
	.w6(32'hbbd4e36b),
	.w7(32'hbbfc51c6),
	.w8(32'hbb6a3265),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93c9f8),
	.w1(32'h3a314c33),
	.w2(32'h3b025ed1),
	.w3(32'h3ba9f339),
	.w4(32'h3b85807d),
	.w5(32'h3ae668cb),
	.w6(32'h39cc3204),
	.w7(32'h3ae86d1f),
	.w8(32'h3ab246be),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7564),
	.w1(32'hbb7e004a),
	.w2(32'h3814e0b8),
	.w3(32'hba8edd9b),
	.w4(32'hbb82fbd2),
	.w5(32'hbbcaafcd),
	.w6(32'h39839f1b),
	.w7(32'h3ae962a0),
	.w8(32'hb9bcf95e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39331fc7),
	.w1(32'h3c0c4989),
	.w2(32'h386d2d03),
	.w3(32'hbbb82006),
	.w4(32'hbc4a4402),
	.w5(32'h3b67d195),
	.w6(32'hbb1e7bd7),
	.w7(32'hbbbf059f),
	.w8(32'h39e94d13),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a892458),
	.w1(32'hba63ac42),
	.w2(32'hb95ba312),
	.w3(32'h392b8e07),
	.w4(32'hba0482b7),
	.w5(32'h3a462d41),
	.w6(32'h3bb87425),
	.w7(32'h3b3fb4c6),
	.w8(32'hb9fff993),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e28bc),
	.w1(32'hbac5af57),
	.w2(32'hbb1948cd),
	.w3(32'h3a1ad5c8),
	.w4(32'hb9963338),
	.w5(32'hbc08d663),
	.w6(32'h3b8034ca),
	.w7(32'h38cfb34e),
	.w8(32'hba475f9a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22ec25),
	.w1(32'h3aa3bf9e),
	.w2(32'h3ae4f4d1),
	.w3(32'hbbdf3cd8),
	.w4(32'h3adf1dee),
	.w5(32'hbb22dbb1),
	.w6(32'hbbcfd095),
	.w7(32'h3853d054),
	.w8(32'hbb86f67e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10dbe),
	.w1(32'h3bab2e9a),
	.w2(32'h3abfe367),
	.w3(32'hbb232a3e),
	.w4(32'h39716739),
	.w5(32'hbc0a7b6b),
	.w6(32'h3b538826),
	.w7(32'hb926f2c4),
	.w8(32'hbb228291),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea2c8),
	.w1(32'hbae44fd7),
	.w2(32'h3a5e4c96),
	.w3(32'hbb9e52a7),
	.w4(32'hbb549ffe),
	.w5(32'hbbebb509),
	.w6(32'hbb7f97f0),
	.w7(32'hbb37119b),
	.w8(32'hbb223d2b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92997),
	.w1(32'h3b6cc562),
	.w2(32'hb9871c9e),
	.w3(32'hbb5eb0a0),
	.w4(32'hbb8c6899),
	.w5(32'hbb0a7b8d),
	.w6(32'h3a325b0f),
	.w7(32'h3a49dab1),
	.w8(32'hbb0f9f88),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2afcc7),
	.w1(32'h397afee5),
	.w2(32'h3a7b6246),
	.w3(32'h3a7dcbd3),
	.w4(32'hb9755c53),
	.w5(32'h399362b2),
	.w6(32'h3a4c8be0),
	.w7(32'hbb17b6f2),
	.w8(32'h3b79083d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63c84),
	.w1(32'h3bf1d132),
	.w2(32'h3b53c098),
	.w3(32'h3aad46bc),
	.w4(32'h3b9d7e79),
	.w5(32'h3b70c0e9),
	.w6(32'h3b5480bc),
	.w7(32'h3ba4a053),
	.w8(32'h3af5982b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d750),
	.w1(32'h3be56fa4),
	.w2(32'hbb01cee4),
	.w3(32'h3c06c7ca),
	.w4(32'h3bdcd058),
	.w5(32'h3aac6f01),
	.w6(32'hbaab7f9e),
	.w7(32'h3a28b15f),
	.w8(32'hbba0d18b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da877),
	.w1(32'hbb57f03b),
	.w2(32'hbb1fac8b),
	.w3(32'h3bb3ff38),
	.w4(32'h3986c8ad),
	.w5(32'hbb8cdd1e),
	.w6(32'hba7af874),
	.w7(32'h394819b3),
	.w8(32'hbba7bcbe),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87bd4b),
	.w1(32'hb8dbb9e4),
	.w2(32'hb9f721e1),
	.w3(32'hbb234412),
	.w4(32'h3abaadbe),
	.w5(32'hba892cd9),
	.w6(32'hbb3b96f3),
	.w7(32'h3a4df217),
	.w8(32'hbbe8eb6e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275808),
	.w1(32'hbb5217ab),
	.w2(32'h3ba4e0fe),
	.w3(32'h3a78a3dc),
	.w4(32'h3ae2de89),
	.w5(32'h3bf21358),
	.w6(32'hbba088a0),
	.w7(32'h3ae2e7c8),
	.w8(32'h3c14c1dd),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0f157),
	.w1(32'hbb6a6b51),
	.w2(32'hbbc9bf93),
	.w3(32'h3b94e878),
	.w4(32'hbbd4bc88),
	.w5(32'h3bec4ef5),
	.w6(32'h3b7fd017),
	.w7(32'hbc2a0911),
	.w8(32'hb8b70c7b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfab3d),
	.w1(32'hbc41ec66),
	.w2(32'hbc4551e8),
	.w3(32'hbb24f523),
	.w4(32'hba8c3174),
	.w5(32'hbc22a040),
	.w6(32'h3a789551),
	.w7(32'hbc7d24b4),
	.w8(32'hbc13ba6a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e849),
	.w1(32'h3b5d7ca6),
	.w2(32'h3b9ff335),
	.w3(32'hba4d81fc),
	.w4(32'hbb15a249),
	.w5(32'h3b83782f),
	.w6(32'hbc179cb7),
	.w7(32'hbb331107),
	.w8(32'hbb1720ca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48c3bf),
	.w1(32'h3b477699),
	.w2(32'h3b21d0c3),
	.w3(32'hba81b388),
	.w4(32'h3b4f056e),
	.w5(32'h3c43d13e),
	.w6(32'h3a1a3486),
	.w7(32'hba604fc6),
	.w8(32'h3b4216bd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0376),
	.w1(32'h3c358374),
	.w2(32'h3ab3adab),
	.w3(32'h3c8d85ed),
	.w4(32'h3b5813b3),
	.w5(32'h39c93c0e),
	.w6(32'h3bafc152),
	.w7(32'h3ca7434b),
	.w8(32'h3c2bb479),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1836c8),
	.w1(32'hbb6474fd),
	.w2(32'h3aa4f3d2),
	.w3(32'h3c912a8f),
	.w4(32'h3bbc868a),
	.w5(32'h3b884245),
	.w6(32'h3c7f43fd),
	.w7(32'hbc112350),
	.w8(32'h3a5a6147),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a744),
	.w1(32'hbac2473b),
	.w2(32'hbb123547),
	.w3(32'h3b865ead),
	.w4(32'h3b82a56e),
	.w5(32'hbc29fc4e),
	.w6(32'h38d75b75),
	.w7(32'hba8d030e),
	.w8(32'hbbb9d616),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724346),
	.w1(32'h3bb5802c),
	.w2(32'h3b524bf0),
	.w3(32'h3aaa545d),
	.w4(32'h3ae7afee),
	.w5(32'h3a749de6),
	.w6(32'h3cf4db81),
	.w7(32'h3b950dd2),
	.w8(32'hba3135bb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e292),
	.w1(32'hbbcdf6a3),
	.w2(32'hbb50b561),
	.w3(32'hbb7c0e02),
	.w4(32'hbb2ad36d),
	.w5(32'h3b729d40),
	.w6(32'h3b5ffc12),
	.w7(32'hbbfb424a),
	.w8(32'hbba07ce2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb7dc),
	.w1(32'hbbaada4c),
	.w2(32'h3b6051cd),
	.w3(32'h3b3ede9a),
	.w4(32'h3b122b00),
	.w5(32'h3abf83c4),
	.w6(32'hbc107dc9),
	.w7(32'h39088a64),
	.w8(32'h3b381ef6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac08f75),
	.w1(32'hbaef1b6e),
	.w2(32'hbb03bd56),
	.w3(32'h399a85c9),
	.w4(32'hbb087161),
	.w5(32'h3bcfec68),
	.w6(32'h3b742790),
	.w7(32'hbb67e3b9),
	.w8(32'h3bf6a860),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b678f43),
	.w1(32'h39ae20da),
	.w2(32'h3c572843),
	.w3(32'h3c7c410e),
	.w4(32'h3c6b40ec),
	.w5(32'hbae146b3),
	.w6(32'h3cb34549),
	.w7(32'h3c4fca7f),
	.w8(32'hbc070f44),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62a997),
	.w1(32'h3b95c72c),
	.w2(32'hb9dcb93e),
	.w3(32'hbb96856e),
	.w4(32'h39b50952),
	.w5(32'hbc7ce8df),
	.w6(32'hbbc0aa30),
	.w7(32'h3b2d2e0d),
	.w8(32'hbc67cab2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f2a1),
	.w1(32'hbc38963c),
	.w2(32'hbbffe490),
	.w3(32'hbbb08098),
	.w4(32'hbba361c2),
	.w5(32'h3a96a9cc),
	.w6(32'hbb971af5),
	.w7(32'hbbe63f9b),
	.w8(32'hbb1b66b4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf525b8),
	.w1(32'h3a528713),
	.w2(32'h35d3e90f),
	.w3(32'hbac50dd9),
	.w4(32'hbab03fc5),
	.w5(32'hbae5675d),
	.w6(32'hbb64ac0a),
	.w7(32'h3b85d78b),
	.w8(32'hb9b3ff73),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc5a7),
	.w1(32'hbc09766d),
	.w2(32'hbc04cb8e),
	.w3(32'hbbb4132e),
	.w4(32'hbbbd6491),
	.w5(32'h3a0b579c),
	.w6(32'hbb8c2f97),
	.w7(32'hbc60d22c),
	.w8(32'hbbed9810),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5407c5),
	.w1(32'h397a1b95),
	.w2(32'hbb91c6e1),
	.w3(32'hbb2a7b3d),
	.w4(32'hb73879e7),
	.w5(32'hbb9a602b),
	.w6(32'hbc770390),
	.w7(32'h3ad55b79),
	.w8(32'hbbe098d7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc384f6),
	.w1(32'hbb9cf30d),
	.w2(32'hbb5bc07e),
	.w3(32'hbbb7d5c6),
	.w4(32'hbbab79cc),
	.w5(32'hbc72306b),
	.w6(32'hbc0038fe),
	.w7(32'hbb66494f),
	.w8(32'hbb9b0d1f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ae10),
	.w1(32'hbc21803f),
	.w2(32'hbc08552e),
	.w3(32'hbc399b9b),
	.w4(32'hbbde9820),
	.w5(32'h3b343ae8),
	.w6(32'hbcbe6d13),
	.w7(32'hbcb5ca87),
	.w8(32'hbbd4bfaf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab39f2d),
	.w1(32'h3b65f463),
	.w2(32'h3bf92e02),
	.w3(32'h3b09027b),
	.w4(32'h3868d683),
	.w5(32'h3c570881),
	.w6(32'hbba1c425),
	.w7(32'hbb13e52f),
	.w8(32'hbbddbd92),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f74b03),
	.w1(32'h3b4bf4ae),
	.w2(32'h3c934e23),
	.w3(32'h3b7fb99d),
	.w4(32'h3c354ddd),
	.w5(32'h3bd131d0),
	.w6(32'hbce4fea9),
	.w7(32'h3c331602),
	.w8(32'h3c08878d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2cb5),
	.w1(32'h3c7cd018),
	.w2(32'h3beea38f),
	.w3(32'hbb421934),
	.w4(32'h3c22e524),
	.w5(32'hba9eafb5),
	.w6(32'hbcb43e3e),
	.w7(32'h3c80b7b1),
	.w8(32'hbbfcae6d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a957a60),
	.w1(32'h3bb40699),
	.w2(32'hba96dd97),
	.w3(32'hbb84dc9f),
	.w4(32'h3b2b4886),
	.w5(32'hbc145edd),
	.w6(32'h3ac71f73),
	.w7(32'h3b79a9d5),
	.w8(32'h3807f083),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452709),
	.w1(32'h3b043b34),
	.w2(32'hbaffe423),
	.w3(32'hbbb04314),
	.w4(32'h3a94baf9),
	.w5(32'hbae9550d),
	.w6(32'h3ba4e3e7),
	.w7(32'hbb3d1a7a),
	.w8(32'hbb82c374),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa38a59),
	.w1(32'hbb19290f),
	.w2(32'hbaa10aa9),
	.w3(32'hbbd62ccd),
	.w4(32'hbc09f708),
	.w5(32'hbb886759),
	.w6(32'hbaa2c10a),
	.w7(32'hbbd11d38),
	.w8(32'h3a4a2bb8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f9457),
	.w1(32'h3b06dd9f),
	.w2(32'hbb91287e),
	.w3(32'hbb985241),
	.w4(32'hbabc8137),
	.w5(32'hbb118d00),
	.w6(32'h3bca8e20),
	.w7(32'hbacc0ad5),
	.w8(32'hbb16c660),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bf808),
	.w1(32'hba858134),
	.w2(32'h3b57dcab),
	.w3(32'h3aa0f80f),
	.w4(32'hbb1afed9),
	.w5(32'h3a9f0bc1),
	.w6(32'hb9af1cdb),
	.w7(32'h3afd9977),
	.w8(32'h3bb7f005),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9572ae),
	.w1(32'h3acdbeaf),
	.w2(32'h3b1f0cd0),
	.w3(32'h3b230c27),
	.w4(32'h3b76f95d),
	.w5(32'h3be279f2),
	.w6(32'h3c0a2ade),
	.w7(32'hba93f794),
	.w8(32'hbb0dbc30),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb264f3),
	.w1(32'hbc066ddc),
	.w2(32'hbb0c836f),
	.w3(32'hbaec798a),
	.w4(32'hbb708821),
	.w5(32'hbb37d4c1),
	.w6(32'hbb09e2a5),
	.w7(32'hba39f230),
	.w8(32'h3ae46311),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule