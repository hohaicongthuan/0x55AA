module layer_10_featuremap_305(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36888308),
	.w1(32'h37a065a8),
	.w2(32'h37cb7ff4),
	.w3(32'h36ce4239),
	.w4(32'h3827ef21),
	.w5(32'h381735e1),
	.w6(32'h36e9e57e),
	.w7(32'h3793625a),
	.w8(32'h37961ed5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbda0a),
	.w1(32'hbb7bfa76),
	.w2(32'hbb096492),
	.w3(32'hbb53e7fd),
	.w4(32'hbb6a0861),
	.w5(32'hbaea8091),
	.w6(32'hbab7cd78),
	.w7(32'hba06fc6e),
	.w8(32'hb9d28e1a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ba5b5),
	.w1(32'hb760cf61),
	.w2(32'hb790c5fa),
	.w3(32'hb6bd9bc8),
	.w4(32'hb6024b68),
	.w5(32'hb6957c73),
	.w6(32'h37952b26),
	.w7(32'h371ee504),
	.w8(32'h361f2eb1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874c20e),
	.w1(32'hba55df1a),
	.w2(32'hbad8584a),
	.w3(32'h39cc74ad),
	.w4(32'hba6d008b),
	.w5(32'h39db2cb6),
	.w6(32'hb9bbc61d),
	.w7(32'hbad168d5),
	.w8(32'hb9f96afc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb588c8cc),
	.w1(32'hb75af48f),
	.w2(32'h3738d656),
	.w3(32'h37102953),
	.w4(32'h37405b64),
	.w5(32'h3730d63a),
	.w6(32'hb83644f7),
	.w7(32'hb84b2fb2),
	.w8(32'h37045be4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3749783b),
	.w1(32'h37a29307),
	.w2(32'h36249bba),
	.w3(32'h36d42124),
	.w4(32'hb6f33329),
	.w5(32'hb7b2506f),
	.w6(32'h378eeba3),
	.w7(32'hb77ec162),
	.w8(32'hb75a4a56),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5271),
	.w1(32'hbc0a170d),
	.w2(32'hb972882f),
	.w3(32'hbb87bdbe),
	.w4(32'hbaafb746),
	.w5(32'h3bef450c),
	.w6(32'hbb3f99a9),
	.w7(32'h3bbd3c5b),
	.w8(32'h3c56732a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85a8dd),
	.w1(32'h3c302ee3),
	.w2(32'hb8df982e),
	.w3(32'h3c2dc91c),
	.w4(32'h3c266c07),
	.w5(32'h3c01e90f),
	.w6(32'h3c80622d),
	.w7(32'h3bfcadf7),
	.w8(32'hbbe6dec9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a07bc),
	.w1(32'h39212020),
	.w2(32'h38dab1bd),
	.w3(32'h398e0991),
	.w4(32'h38a41771),
	.w5(32'h3782e893),
	.w6(32'h391e133e),
	.w7(32'hb379322e),
	.w8(32'h38912160),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d3e3c),
	.w1(32'h3a136a1f),
	.w2(32'h3a3c89d7),
	.w3(32'h3ac250bd),
	.w4(32'h3acc6239),
	.w5(32'h3b3ceb2f),
	.w6(32'hbae0f67c),
	.w7(32'h3af0fec7),
	.w8(32'h39a8ccf1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1c193),
	.w1(32'h386490c2),
	.w2(32'h3900e920),
	.w3(32'h381c8992),
	.w4(32'h3530fec2),
	.w5(32'h388dfb11),
	.w6(32'hb7a251df),
	.w7(32'hb6e4e6f0),
	.w8(32'h38d5357e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a688d),
	.w1(32'hbc0a5022),
	.w2(32'hbad5e9fd),
	.w3(32'hbb8b4206),
	.w4(32'hbbf3d124),
	.w5(32'h3bfcda18),
	.w6(32'hbaf5e9f0),
	.w7(32'h3ab31e46),
	.w8(32'h3c44a947),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9d7be),
	.w1(32'h3bab4487),
	.w2(32'h3b87b7e3),
	.w3(32'h3bd98366),
	.w4(32'h3bedaf06),
	.w5(32'h3bba6201),
	.w6(32'h3b3010a3),
	.w7(32'h3ba98705),
	.w8(32'h3ad3a5e1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0da7b1),
	.w1(32'h3b901c12),
	.w2(32'h3b47421f),
	.w3(32'h3a12e876),
	.w4(32'h3b939b59),
	.w5(32'hba3bbdf7),
	.w6(32'h3aad0dfc),
	.w7(32'h3b72213a),
	.w8(32'h39cc1464),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65bbe2),
	.w1(32'hbb30ffbd),
	.w2(32'h38cc3fa8),
	.w3(32'hbb33c6f9),
	.w4(32'hbb7f05b0),
	.w5(32'hbb33522e),
	.w6(32'hbabb22c9),
	.w7(32'hbac28589),
	.w8(32'hb9b8581b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab170de),
	.w1(32'h39c6d85b),
	.w2(32'hba15c8da),
	.w3(32'h3af8da99),
	.w4(32'h3a64c79c),
	.w5(32'hbb42ca17),
	.w6(32'hbaa67a66),
	.w7(32'h3aab3c8d),
	.w8(32'hbafa66fd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7a029),
	.w1(32'hb8ad4287),
	.w2(32'h381b1a9f),
	.w3(32'hb8417aec),
	.w4(32'hb893a09d),
	.w5(32'hb7a9ada1),
	.w6(32'hb9162e8e),
	.w7(32'hb88544cb),
	.w8(32'h38b04463),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cd689),
	.w1(32'h3ae2b668),
	.w2(32'hb9957673),
	.w3(32'h3bb093e2),
	.w4(32'h3c37b03d),
	.w5(32'h3c05322d),
	.w6(32'hbb5476d0),
	.w7(32'h3b0d22e8),
	.w8(32'hbaa12639),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc38e8),
	.w1(32'h3b4d866d),
	.w2(32'h3aeb7464),
	.w3(32'h3b879b9e),
	.w4(32'h3bbfdffc),
	.w5(32'h3b9ebb37),
	.w6(32'hb9f03ab2),
	.w7(32'h3b336b9e),
	.w8(32'h3a3038f4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9014150),
	.w1(32'hb96a95e3),
	.w2(32'hb8fdb873),
	.w3(32'hb8bfad23),
	.w4(32'hb99e0671),
	.w5(32'hb89112a5),
	.w6(32'hb7e28df0),
	.w7(32'hb8b6970f),
	.w8(32'h38dc1a3b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36414938),
	.w1(32'h38bd2b77),
	.w2(32'h38b949d7),
	.w3(32'hb67b1c9c),
	.w4(32'hb7ffce74),
	.w5(32'h387cdfb3),
	.w6(32'hb7de8f82),
	.w7(32'hb73a3f7f),
	.w8(32'hb8a67495),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c01cf),
	.w1(32'h3904eef1),
	.w2(32'h39b53adc),
	.w3(32'hba234da7),
	.w4(32'hba9d9553),
	.w5(32'hba4bafe7),
	.w6(32'hb9484e92),
	.w7(32'hb9353548),
	.w8(32'hb9d28a67),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59975),
	.w1(32'h39c2a2f5),
	.w2(32'h3bb2ec1f),
	.w3(32'h3b8d48ba),
	.w4(32'hbb93f8c9),
	.w5(32'h3b730e22),
	.w6(32'hbc04b0a9),
	.w7(32'hbbd97c9e),
	.w8(32'h3a0c845d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb832f34),
	.w1(32'hbb19f884),
	.w2(32'hba29477b),
	.w3(32'hbb76888f),
	.w4(32'hbb37090c),
	.w5(32'hbb340045),
	.w6(32'hbbd4e444),
	.w7(32'hbba16512),
	.w8(32'hbb86046f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe38a04),
	.w1(32'hbbc202c3),
	.w2(32'hbaf0590f),
	.w3(32'hbc0113a0),
	.w4(32'hbc20f3a2),
	.w5(32'hbc012b19),
	.w6(32'hbb28b026),
	.w7(32'hbb85d293),
	.w8(32'hbbd30816),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a007d3),
	.w1(32'hb91a581f),
	.w2(32'hb8d9503f),
	.w3(32'h39025430),
	.w4(32'hb730ef1a),
	.w5(32'hb8a63b94),
	.w6(32'h381e2264),
	.w7(32'hb83170aa),
	.w8(32'h38055d2e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351fb013),
	.w1(32'hb8441a5d),
	.w2(32'hb8a15fe1),
	.w3(32'hb8a4c991),
	.w4(32'hb9182e6a),
	.w5(32'hb9147ba1),
	.w6(32'hb7995fef),
	.w7(32'hb88b9723),
	.w8(32'hb8da22d4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b498423),
	.w1(32'hbb3d0480),
	.w2(32'h3accec58),
	.w3(32'h3b0ce1d4),
	.w4(32'hbbc1ceab),
	.w5(32'hbb9eac81),
	.w6(32'h3bf02117),
	.w7(32'h3b00eac1),
	.w8(32'hbb7f2168),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a719805),
	.w1(32'h3a740a06),
	.w2(32'h393b2851),
	.w3(32'h38f06b46),
	.w4(32'hb676de36),
	.w5(32'h38b70146),
	.w6(32'hb91d949e),
	.w7(32'hb9986d88),
	.w8(32'hb9a4af0c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd689e8),
	.w1(32'hbbd59d14),
	.w2(32'hbb050613),
	.w3(32'hbaec92cb),
	.w4(32'hbbc2a632),
	.w5(32'hbbefbbfa),
	.w6(32'hbaf288ea),
	.w7(32'hbb178070),
	.w8(32'hbb9e3b98),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780c1d0),
	.w1(32'h36803177),
	.w2(32'hb72f1ee8),
	.w3(32'h3793139b),
	.w4(32'h3615bf81),
	.w5(32'hb82cb15f),
	.w6(32'hb8176971),
	.w7(32'hb831a853),
	.w8(32'h36246f84),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f6f18b),
	.w1(32'hb895966a),
	.w2(32'hb85f7194),
	.w3(32'hb826e1e8),
	.w4(32'hb898bbc4),
	.w5(32'hb51346ca),
	.w6(32'h37eaafd9),
	.w7(32'hb73d2605),
	.w8(32'hb577585f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab439ba),
	.w1(32'hbac73f48),
	.w2(32'hba8ac144),
	.w3(32'hba979f6c),
	.w4(32'h3974af43),
	.w5(32'h3aa173f0),
	.w6(32'hbb1c06ef),
	.w7(32'hba3218eb),
	.w8(32'hb933a959),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f51fa),
	.w1(32'hb9287bc9),
	.w2(32'h3a3478d1),
	.w3(32'hba8eb398),
	.w4(32'hbacd89f2),
	.w5(32'hba0c9c0c),
	.w6(32'hb9c2e9f2),
	.w7(32'hba76b714),
	.w8(32'hba5c4d20),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba838f8d),
	.w1(32'hba878870),
	.w2(32'hba86e24c),
	.w3(32'h392ab9ce),
	.w4(32'hba2065bb),
	.w5(32'hba228a84),
	.w6(32'h3a3f7994),
	.w7(32'h3b074adb),
	.w8(32'h3ac74e56),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbdf2f),
	.w1(32'hbadde285),
	.w2(32'hb951f516),
	.w3(32'hb9ae88b5),
	.w4(32'hb90e2d71),
	.w5(32'h3b9a784d),
	.w6(32'hb9fe9eb2),
	.w7(32'hba450ae9),
	.w8(32'h3ab2b107),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22557d),
	.w1(32'hbb6df0bf),
	.w2(32'h3c0eabd3),
	.w3(32'h3aa99620),
	.w4(32'hbcb3c42a),
	.w5(32'h3bf91211),
	.w6(32'hbb15dcd3),
	.w7(32'hbc74537e),
	.w8(32'h3cb1925d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f73b),
	.w1(32'hbb97e9c5),
	.w2(32'hbadd5984),
	.w3(32'hbbad6ed4),
	.w4(32'hbc63c743),
	.w5(32'hbc66a670),
	.w6(32'hba0fec21),
	.w7(32'hbb9ab17b),
	.w8(32'hbc2fdb07),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4a86),
	.w1(32'h39837c8d),
	.w2(32'h3bbae69a),
	.w3(32'hb92d1ef8),
	.w4(32'hbba9652f),
	.w5(32'hbb33890d),
	.w6(32'hba830e99),
	.w7(32'h3ab3fa8c),
	.w8(32'hbafaf3b7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e94e),
	.w1(32'hbafbabf2),
	.w2(32'hbaabba76),
	.w3(32'hbb15d839),
	.w4(32'hbb6c87ac),
	.w5(32'hbb1a1c5b),
	.w6(32'hba47d8ec),
	.w7(32'hbacc0c51),
	.w8(32'hba88b24b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3820bf0d),
	.w1(32'h3734637b),
	.w2(32'h3423fab0),
	.w3(32'h380f1ba2),
	.w4(32'hb7a7bb5c),
	.w5(32'hb801af80),
	.w6(32'h38795c23),
	.w7(32'h381c8a14),
	.w8(32'h384f5252),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d37e1f),
	.w1(32'hb89da0d5),
	.w2(32'hb8933585),
	.w3(32'hb803dfb6),
	.w4(32'hb94094bc),
	.w5(32'hb94dbe80),
	.w6(32'h3872e5f6),
	.w7(32'hb84323c5),
	.w8(32'hb902075e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397eeb4a),
	.w1(32'h3919ee81),
	.w2(32'h3a03dde2),
	.w3(32'hb70c3be9),
	.w4(32'hb8899481),
	.w5(32'h3a409cb1),
	.w6(32'h39af097e),
	.w7(32'h387ed1aa),
	.w8(32'h39fe9a4e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10bccd),
	.w1(32'h3b8cf5cf),
	.w2(32'h3af35c98),
	.w3(32'h3bcd3b25),
	.w4(32'h3bba3e2a),
	.w5(32'h3a0d8bf0),
	.w6(32'hbafeb9a5),
	.w7(32'h3b44d0bd),
	.w8(32'hbba6563d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf0a4),
	.w1(32'hbb9d3603),
	.w2(32'hbaf63aaf),
	.w3(32'hbb6fb949),
	.w4(32'hbbe682ee),
	.w5(32'hbbb6146e),
	.w6(32'hbb993d0b),
	.w7(32'hbbdb391f),
	.w8(32'hbbd54cf5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a89d),
	.w1(32'hbaa8ff09),
	.w2(32'hbab849ae),
	.w3(32'hbb825f0e),
	.w4(32'hbbd7d338),
	.w5(32'hbb5eb628),
	.w6(32'hbbee3450),
	.w7(32'hbbf70e84),
	.w8(32'hbbe5ab71),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33aba4),
	.w1(32'hbb4b748a),
	.w2(32'hbb2b1c6c),
	.w3(32'hbb1e05d5),
	.w4(32'hbb9e2c04),
	.w5(32'hbbb1b7af),
	.w6(32'hbb3f58d4),
	.w7(32'hbb8faae3),
	.w8(32'hbbbd1308),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45e395),
	.w1(32'h3bb48808),
	.w2(32'h3ba4f133),
	.w3(32'h3c1044b2),
	.w4(32'h3c543fe7),
	.w5(32'h3c78a620),
	.w6(32'hba25dc9d),
	.w7(32'h3b75deda),
	.w8(32'h3bb0cc25),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3819fbe1),
	.w1(32'hb5798965),
	.w2(32'h389bd0a7),
	.w3(32'h380d0f2a),
	.w4(32'hb73779a5),
	.w5(32'h388d7672),
	.w6(32'h386bb56a),
	.w7(32'h37c583b3),
	.w8(32'h39041219),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5fe36),
	.w1(32'hb913aa4a),
	.w2(32'h371ead26),
	.w3(32'hb8db32ac),
	.w4(32'hb99ec372),
	.w5(32'hb8953fa6),
	.w6(32'hb89518aa),
	.w7(32'hb949a1d3),
	.w8(32'hb835c3f2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7aa01),
	.w1(32'hb89f7cff),
	.w2(32'hb6a3879e),
	.w3(32'hb8b2ef40),
	.w4(32'hb851802f),
	.w5(32'hb7783522),
	.w6(32'hb805936e),
	.w7(32'hb871a9c6),
	.w8(32'hb7f277ad),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14fa8c),
	.w1(32'h3b147519),
	.w2(32'h3aa11dfd),
	.w3(32'h3ab9488e),
	.w4(32'h39a0b81f),
	.w5(32'hba812555),
	.w6(32'hb9b3ad97),
	.w7(32'h39a9bd04),
	.w8(32'hb9a7840f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb049c),
	.w1(32'hba271fbf),
	.w2(32'hba8f1b2f),
	.w3(32'h3a24dd79),
	.w4(32'hba061898),
	.w5(32'h39c18439),
	.w6(32'h3a0bbf80),
	.w7(32'hbaa59d6d),
	.w8(32'hba8ab328),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8b395),
	.w1(32'hba2db3ed),
	.w2(32'hbb7f4b6a),
	.w3(32'h3b770df1),
	.w4(32'h3bae5683),
	.w5(32'h3b82c649),
	.w6(32'hbb6312f8),
	.w7(32'h3abd1888),
	.w8(32'hbb48ff2b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1230b8),
	.w1(32'h3a7a3cae),
	.w2(32'h3aa153a0),
	.w3(32'h3a94461e),
	.w4(32'hb8fda1f0),
	.w5(32'hba1e8ea4),
	.w6(32'h39dfcca2),
	.w7(32'hbaa1b7e7),
	.w8(32'hbb84e538),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16e0e6),
	.w1(32'hb9a71731),
	.w2(32'hb80b3d18),
	.w3(32'hb9e384d5),
	.w4(32'hb9f32f1b),
	.w5(32'hb9720b35),
	.w6(32'hb9112c26),
	.w7(32'hb8da1ff9),
	.w8(32'hb6c227c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7979b26),
	.w1(32'hb7d06b53),
	.w2(32'hb853d5f3),
	.w3(32'hb8384675),
	.w4(32'hb8dd24c7),
	.w5(32'hb8a8872d),
	.w6(32'hb60ca383),
	.w7(32'hb8b05718),
	.w8(32'hb8886966),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959a5d8),
	.w1(32'h392e63e8),
	.w2(32'h3a0f3cef),
	.w3(32'hba4a14a2),
	.w4(32'h39009864),
	.w5(32'h38beb102),
	.w6(32'hb9c0d42d),
	.w7(32'h3a1c0e95),
	.w8(32'h38d2b9a2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe0616),
	.w1(32'hb984c133),
	.w2(32'hb9192c2c),
	.w3(32'hb93322a2),
	.w4(32'hba334c8d),
	.w5(32'hb945acb7),
	.w6(32'h38c2e2d3),
	.w7(32'hb9d313eb),
	.w8(32'hb94ddc1a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9868ec1),
	.w1(32'hba04ad83),
	.w2(32'hb9723a0d),
	.w3(32'hb90b0f07),
	.w4(32'hb82014c7),
	.w5(32'h392e5bfe),
	.w6(32'hb60d7a4c),
	.w7(32'h39622541),
	.w8(32'h38c3a96f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ea9e6),
	.w1(32'h3a0b7195),
	.w2(32'hba41f402),
	.w3(32'h3b252134),
	.w4(32'h3b33cc35),
	.w5(32'h3ab7916d),
	.w6(32'hba054865),
	.w7(32'h3adba41e),
	.w8(32'hba5beaf4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d48a0),
	.w1(32'h388f3ca3),
	.w2(32'hbb1fe8eb),
	.w3(32'h3ba279cd),
	.w4(32'h3a459b57),
	.w5(32'hbbe50613),
	.w6(32'h3b51fb7c),
	.w7(32'h3b3e8d5d),
	.w8(32'hbbe003b0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37285109),
	.w1(32'hb6d6dfb4),
	.w2(32'hb577cd81),
	.w3(32'h37c22d22),
	.w4(32'hb6c1c62e),
	.w5(32'hb821040f),
	.w6(32'h35d28e91),
	.w7(32'hb687539a),
	.w8(32'hb5091ed7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce8f66),
	.w1(32'hb801d060),
	.w2(32'hb788ade6),
	.w3(32'hb70a4f85),
	.w4(32'hb7d9da7f),
	.w5(32'hb8461f08),
	.w6(32'hb401f782),
	.w7(32'h35a8df51),
	.w8(32'hb7bb4841),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e35e4),
	.w1(32'hb92691a8),
	.w2(32'hb8bfa5e7),
	.w3(32'hb9678856),
	.w4(32'hb9257293),
	.w5(32'hb8790e19),
	.w6(32'hb949c64a),
	.w7(32'hb900ab09),
	.w8(32'hb865e126),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba7ad3),
	.w1(32'h37b5ed9a),
	.w2(32'h3734a111),
	.w3(32'hb6814ae8),
	.w4(32'hb7c9a808),
	.w5(32'hb8395a78),
	.w6(32'h38324da3),
	.w7(32'hb60e921d),
	.w8(32'hb81960c0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8644),
	.w1(32'hbbd4e58f),
	.w2(32'hbc17dd34),
	.w3(32'hbb4d84c5),
	.w4(32'hbbbf2518),
	.w5(32'hbc580567),
	.w6(32'h396e7397),
	.w7(32'h3bed7996),
	.w8(32'hbbd6fe31),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202c43),
	.w1(32'hb9ba6fd3),
	.w2(32'hb95cefae),
	.w3(32'hbb470a77),
	.w4(32'hba69a8f3),
	.w5(32'h3bae0764),
	.w6(32'hbbafde77),
	.w7(32'hbb8fb544),
	.w8(32'hbbe85392),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa85b),
	.w1(32'h3ae7d5cb),
	.w2(32'hb9fbd6da),
	.w3(32'h3a9e4b8e),
	.w4(32'h3a921a50),
	.w5(32'hbb3d26fc),
	.w6(32'hbb87d29d),
	.w7(32'hbb045ea7),
	.w8(32'hbba75582),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1775de),
	.w1(32'hbbf73d09),
	.w2(32'hbae734f6),
	.w3(32'hbc3961e8),
	.w4(32'hbc8f0feb),
	.w5(32'hbc493500),
	.w6(32'hbb69e6d5),
	.w7(32'hbbe0b699),
	.w8(32'hbc16dc3f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb757f732),
	.w1(32'h378de654),
	.w2(32'h37fba86b),
	.w3(32'hb80bd6b4),
	.w4(32'hb8243aa8),
	.w5(32'h38331cd3),
	.w6(32'h36c20404),
	.w7(32'hb7c283c0),
	.w8(32'h387d0a8a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36207a15),
	.w1(32'h3591d0ec),
	.w2(32'h360d31fe),
	.w3(32'hb73a1a6c),
	.w4(32'hb8874b2e),
	.w5(32'hb8ada952),
	.w6(32'h383690ba),
	.w7(32'h36127f00),
	.w8(32'hb82a0ac7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ee938),
	.w1(32'h37c2b96b),
	.w2(32'h380d5c3d),
	.w3(32'h3895b3e3),
	.w4(32'hb75cc771),
	.w5(32'hb869696e),
	.w6(32'h38d51b2b),
	.w7(32'h3880b9fc),
	.w8(32'hb5f22270),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a1c49),
	.w1(32'h3a567434),
	.w2(32'hb9e99fbe),
	.w3(32'h3af10ded),
	.w4(32'h3b2d72ed),
	.w5(32'h3a9a1ee7),
	.w6(32'h3ab660f0),
	.w7(32'h3ace397b),
	.w8(32'hba6795c6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb697317d),
	.w1(32'hb7f74f2e),
	.w2(32'hb831fb6c),
	.w3(32'hb73c7b7e),
	.w4(32'hb83a837c),
	.w5(32'hb7a1dd92),
	.w6(32'h37d4a560),
	.w7(32'h36961fe0),
	.w8(32'h37835169),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d850),
	.w1(32'h3aa54933),
	.w2(32'hba31b580),
	.w3(32'h3ab30caa),
	.w4(32'hba0636b0),
	.w5(32'h39d17ced),
	.w6(32'hba0c9404),
	.w7(32'hbab2d637),
	.w8(32'hbab01b05),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0af35),
	.w1(32'h3b0418e4),
	.w2(32'h3a0d511e),
	.w3(32'h3b706f25),
	.w4(32'h3bb6ffb0),
	.w5(32'h3bf73973),
	.w6(32'h3ae0696d),
	.w7(32'hba58e385),
	.w8(32'h39d5987b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ba6a1),
	.w1(32'h3a890277),
	.w2(32'h3af4e3fa),
	.w3(32'h3a9cba0a),
	.w4(32'hba8271b1),
	.w5(32'hb98a34d1),
	.w6(32'h39a45110),
	.w7(32'h399bbed3),
	.w8(32'hba8590b1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964d6e8),
	.w1(32'h3a415dba),
	.w2(32'hba737a5d),
	.w3(32'hb8a3b1db),
	.w4(32'h3b13bcff),
	.w5(32'hba462252),
	.w6(32'hbb00bdfd),
	.w7(32'h3a8b8cc3),
	.w8(32'hbb11b839),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407245),
	.w1(32'hbaf5573c),
	.w2(32'hbad07aae),
	.w3(32'hbaf0995e),
	.w4(32'hbbb11e85),
	.w5(32'hbb50a616),
	.w6(32'h39bf66c9),
	.w7(32'h3b757f74),
	.w8(32'h3b6af784),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a62d4),
	.w1(32'hb9c232f0),
	.w2(32'h3a6f9e05),
	.w3(32'h395e9cac),
	.w4(32'hbb117f40),
	.w5(32'hbb293b45),
	.w6(32'h388b6e7e),
	.w7(32'hb9d01b9b),
	.w8(32'hbb3d5d52),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b533a2d),
	.w1(32'h3a64d13c),
	.w2(32'h3a9c3d6d),
	.w3(32'h3b0a73b5),
	.w4(32'h3b3688aa),
	.w5(32'h3b8307f9),
	.w6(32'hba440376),
	.w7(32'h3a9100fd),
	.w8(32'h3af1fe30),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3791d74c),
	.w1(32'h38019a51),
	.w2(32'h3785c6c5),
	.w3(32'h37b310af),
	.w4(32'h372ff20b),
	.w5(32'hb7b6232e),
	.w6(32'h381012d5),
	.w7(32'h3814dc2a),
	.w8(32'hb7da71f6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c9327),
	.w1(32'hb6291683),
	.w2(32'h37830eff),
	.w3(32'h383553ae),
	.w4(32'hb4d6d329),
	.w5(32'hb459f38e),
	.w6(32'h38c35c10),
	.w7(32'h38877ca8),
	.w8(32'h380fd9e7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e24959),
	.w1(32'h379de968),
	.w2(32'hb868b59f),
	.w3(32'hb8016eb9),
	.w4(32'hb757af2d),
	.w5(32'hb83bd2de),
	.w6(32'hb8726332),
	.w7(32'hb77e7fe4),
	.w8(32'hb8869c1b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba018cbe),
	.w1(32'h39227883),
	.w2(32'h3812941f),
	.w3(32'h391145c7),
	.w4(32'h3a4f7ceb),
	.w5(32'h39adf294),
	.w6(32'h38bfb0ba),
	.w7(32'h3a4272a8),
	.w8(32'h399dc2f3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53efd4),
	.w1(32'hbb19ec8c),
	.w2(32'h39995e38),
	.w3(32'hbb93451e),
	.w4(32'hbc1307f0),
	.w5(32'hbba09b38),
	.w6(32'hbb17e5e6),
	.w7(32'hbb8fae9f),
	.w8(32'hbb15eb48),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d66ec),
	.w1(32'h395add37),
	.w2(32'hb7a5b6ae),
	.w3(32'h39c98fae),
	.w4(32'hb8fbe51f),
	.w5(32'h3994ac07),
	.w6(32'h39b15fd5),
	.w7(32'hb8c13175),
	.w8(32'hb8eea406),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337dfd),
	.w1(32'hbb79baf5),
	.w2(32'hbb5119b1),
	.w3(32'hbb9a464c),
	.w4(32'hbbb27fbb),
	.w5(32'hbb165c96),
	.w6(32'hbb9de5c8),
	.w7(32'hbbcd4af6),
	.w8(32'hbb897a20),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1867a),
	.w1(32'h3b59d8e0),
	.w2(32'h3adc49d3),
	.w3(32'h3b85a9ac),
	.w4(32'h3bfee555),
	.w5(32'h3c0288be),
	.w6(32'hbb33efb9),
	.w7(32'h3ae5caa4),
	.w8(32'h3b0a4605),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e6ef3),
	.w1(32'hb9474fc4),
	.w2(32'h3b3e9a90),
	.w3(32'h3a84fb67),
	.w4(32'hba9aa3aa),
	.w5(32'h39df32bf),
	.w6(32'hb918ffd2),
	.w7(32'hbaa1a0e7),
	.w8(32'hbacc31cc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d086d),
	.w1(32'hbb8f4689),
	.w2(32'h3b16b94e),
	.w3(32'hbb903506),
	.w4(32'hbc2b2ee7),
	.w5(32'hbae46a1e),
	.w6(32'hbb4ac09a),
	.w7(32'hbbb065d1),
	.w8(32'h3bba7648),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab569c3),
	.w1(32'hb9b586d5),
	.w2(32'h3a010f98),
	.w3(32'hbb21fb06),
	.w4(32'hba4ea92b),
	.w5(32'hba128a0d),
	.w6(32'hba815bd8),
	.w7(32'hba404068),
	.w8(32'hbb4e9373),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd2754),
	.w1(32'h3a947d4e),
	.w2(32'hbb28eaae),
	.w3(32'hbb0dc0e3),
	.w4(32'hb984c628),
	.w5(32'hbb85913e),
	.w6(32'hbc012e26),
	.w7(32'hba9469a0),
	.w8(32'hbbaec5d0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd49eb1),
	.w1(32'hbba9aa0c),
	.w2(32'hbad4341d),
	.w3(32'hbbfb3269),
	.w4(32'hbbf07382),
	.w5(32'hbb8cc1e9),
	.w6(32'hbb6e7e3b),
	.w7(32'hbb86cdbc),
	.w8(32'hbb1a3574),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f9702),
	.w1(32'hbb840ca5),
	.w2(32'hbaf87146),
	.w3(32'h3a50de75),
	.w4(32'hbb29d92c),
	.w5(32'hbb649566),
	.w6(32'h3998b619),
	.w7(32'hb981d61f),
	.w8(32'hba92e06e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860f7c4),
	.w1(32'h3897c5a7),
	.w2(32'h393d3f93),
	.w3(32'h370fcc2a),
	.w4(32'h39196e36),
	.w5(32'h39895f57),
	.w6(32'h392b83e0),
	.w7(32'h3989bbfa),
	.w8(32'h39142195),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b198bbd),
	.w1(32'hbad07f7a),
	.w2(32'hbb07048b),
	.w3(32'h3a8fc690),
	.w4(32'h3b752d2f),
	.w5(32'h3ba335cc),
	.w6(32'hbb80d7c7),
	.w7(32'hba02793d),
	.w8(32'hba8a937c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15047b),
	.w1(32'hbb12c184),
	.w2(32'h3be76a4c),
	.w3(32'hba023b43),
	.w4(32'hbb14ae7f),
	.w5(32'hbc9ead28),
	.w6(32'hb980102c),
	.w7(32'h3c23bf0d),
	.w8(32'hbc0f7b9f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e21d8),
	.w1(32'hba990a4e),
	.w2(32'h3c1c2828),
	.w3(32'h3bb89f4e),
	.w4(32'hbc948c99),
	.w5(32'h3bc93f12),
	.w6(32'h3b64a71d),
	.w7(32'hbc72f3a5),
	.w8(32'h3a0e14ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc824315),
	.w1(32'hbbdd7edc),
	.w2(32'h3bc1d4b8),
	.w3(32'hbb8b8efc),
	.w4(32'hbc5c6574),
	.w5(32'hbc6334eb),
	.w6(32'hbbff2345),
	.w7(32'h3bb117b2),
	.w8(32'hbb395989),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5df57),
	.w1(32'hbbe5cd52),
	.w2(32'h3950b4f2),
	.w3(32'hbc540c2f),
	.w4(32'hbc6f54fb),
	.w5(32'hbc498a6c),
	.w6(32'hbc2502ff),
	.w7(32'hbc8c0f98),
	.w8(32'hbc4773fc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60541a),
	.w1(32'hbc1e0a19),
	.w2(32'h3a5a96ef),
	.w3(32'hbb62d0c6),
	.w4(32'hbc9a1712),
	.w5(32'hbb34302d),
	.w6(32'hbc0809b3),
	.w7(32'hbc90de46),
	.w8(32'h3b65b0d6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb702306),
	.w1(32'hbc1c9ab2),
	.w2(32'hbc0a9d36),
	.w3(32'hbba760eb),
	.w4(32'hbc1713e6),
	.w5(32'h3b8a123b),
	.w6(32'hbabfa80c),
	.w7(32'hbb869864),
	.w8(32'hbb4ff25b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00011c),
	.w1(32'h3c5b5241),
	.w2(32'h3c0bb519),
	.w3(32'h3c51930b),
	.w4(32'hbc0bb86f),
	.w5(32'h3c1eb8b5),
	.w6(32'hbbd5804c),
	.w7(32'hbc12f193),
	.w8(32'h3c8d3ce5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5353fa),
	.w1(32'h3b839964),
	.w2(32'h3b3b2a83),
	.w3(32'hba9682da),
	.w4(32'hba6140f1),
	.w5(32'hbb9427ce),
	.w6(32'h3ab44f11),
	.w7(32'hbadb02c1),
	.w8(32'hbc21eea7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371174),
	.w1(32'hbb5cbbc1),
	.w2(32'h3b1ac3c0),
	.w3(32'hbc0db1c4),
	.w4(32'hbb95c677),
	.w5(32'hbb6403d8),
	.w6(32'hbc02ee4a),
	.w7(32'hba08a86b),
	.w8(32'hbc184622),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1a14),
	.w1(32'hba856aa3),
	.w2(32'hb92a1b92),
	.w3(32'hbac57e62),
	.w4(32'hbbcf651f),
	.w5(32'h3aeb9a72),
	.w6(32'h3bd6ecb7),
	.w7(32'h3b5ace82),
	.w8(32'h3a6e9586),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0115d),
	.w1(32'h3c1706dd),
	.w2(32'h3c9462d3),
	.w3(32'h3c00dace),
	.w4(32'h3ca04939),
	.w5(32'h3cd57f6e),
	.w6(32'h3ba5e4d1),
	.w7(32'h3cb4171f),
	.w8(32'h3cce3b5b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f590e),
	.w1(32'h3c9a2e7f),
	.w2(32'hbbc628cd),
	.w3(32'h3c5e158b),
	.w4(32'hbc56cf41),
	.w5(32'hbbfebdcf),
	.w6(32'h3bec5456),
	.w7(32'hbc0cc12a),
	.w8(32'h3b021b98),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2295d),
	.w1(32'h3b8e427e),
	.w2(32'h3c487d30),
	.w3(32'h39663bb4),
	.w4(32'hbb82d53d),
	.w5(32'h3b2f8404),
	.w6(32'hbb5d66fe),
	.w7(32'hbb7e7fec),
	.w8(32'h3b0be869),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0f38a),
	.w1(32'hbbe7a26d),
	.w2(32'h3bea12c6),
	.w3(32'hbb9e9a44),
	.w4(32'hbb64ecb4),
	.w5(32'h3c202038),
	.w6(32'hbc0a29ed),
	.w7(32'hb7017273),
	.w8(32'h3c494e1f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dd7a2),
	.w1(32'hbb96eec5),
	.w2(32'hbbb5cb6f),
	.w3(32'hbb2d2724),
	.w4(32'hbae0a475),
	.w5(32'h399b0eaf),
	.w6(32'hbc828fd5),
	.w7(32'hbc5a8193),
	.w8(32'hbbf3934d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019f88),
	.w1(32'h3b3fe9c0),
	.w2(32'hbb1717e4),
	.w3(32'h3b140024),
	.w4(32'h3b8fd5f5),
	.w5(32'hbab2f273),
	.w6(32'h3b8de94c),
	.w7(32'h3c2efb84),
	.w8(32'h3afd33b6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa7310),
	.w1(32'hbb5065a3),
	.w2(32'hbb555c3e),
	.w3(32'hbc29f166),
	.w4(32'h3c24bcb5),
	.w5(32'hba8c16a9),
	.w6(32'hbbb015a2),
	.w7(32'h3c5c6f0c),
	.w8(32'h3ab79133),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65c5a0),
	.w1(32'hbbfb5e18),
	.w2(32'h3bee7b61),
	.w3(32'h3a8e1105),
	.w4(32'h3ae08b2c),
	.w5(32'h3bcc2971),
	.w6(32'hbb541522),
	.w7(32'hbb339b0b),
	.w8(32'hbba3c87e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc90fe6),
	.w1(32'h3c2f8e19),
	.w2(32'h3be7d3df),
	.w3(32'h3c51cc97),
	.w4(32'h3c158bcd),
	.w5(32'hbb542483),
	.w6(32'h3c433f18),
	.w7(32'h3c1b9fe7),
	.w8(32'hbc51b13a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4045b),
	.w1(32'hbc5a02ad),
	.w2(32'hbbb8de3a),
	.w3(32'hbbf47da4),
	.w4(32'hbc0f471e),
	.w5(32'hbbaf03f5),
	.w6(32'hbc61b448),
	.w7(32'hbc0b21d5),
	.w8(32'hbc43ca07),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19a7f5),
	.w1(32'hbac049f2),
	.w2(32'hbbb618f2),
	.w3(32'h3b4a72c4),
	.w4(32'hbb200203),
	.w5(32'h3a29cfb5),
	.w6(32'h3ac7c4be),
	.w7(32'h3b23783e),
	.w8(32'h3c19438c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42ee44),
	.w1(32'h3a621b22),
	.w2(32'h3b8310b4),
	.w3(32'h3bc6082a),
	.w4(32'h3c0552f2),
	.w5(32'hbb9a55e4),
	.w6(32'h3c482da5),
	.w7(32'h3c5b328e),
	.w8(32'hbb87089e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42937e),
	.w1(32'hbb2ddbdc),
	.w2(32'hbab37bd5),
	.w3(32'h3c4994f9),
	.w4(32'hb9e28142),
	.w5(32'h3c0b4f60),
	.w6(32'h3bc14db9),
	.w7(32'hbb9fd8e7),
	.w8(32'h3bf942b6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa62a),
	.w1(32'h3c3383e2),
	.w2(32'hb9ad68d1),
	.w3(32'h3b4a72cd),
	.w4(32'hbc13d79f),
	.w5(32'h3bd716ed),
	.w6(32'h3c88263b),
	.w7(32'hbcccbd31),
	.w8(32'h3c9f3a79),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a558),
	.w1(32'hbbbaeec9),
	.w2(32'hbbeb7c0a),
	.w3(32'hbae976a9),
	.w4(32'h3b968a1c),
	.w5(32'hbb35405a),
	.w6(32'hbbf2da62),
	.w7(32'hbc753b47),
	.w8(32'h3b8fc94a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3572ff),
	.w1(32'h3bbc14d9),
	.w2(32'hbba4c7e3),
	.w3(32'hbc058af5),
	.w4(32'hbb169a78),
	.w5(32'hbc2be2fd),
	.w6(32'hbc2d2c18),
	.w7(32'hbca80c08),
	.w8(32'h3c8244dd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb543),
	.w1(32'h39e84906),
	.w2(32'hba1331f5),
	.w3(32'hbb3a44f2),
	.w4(32'hba863786),
	.w5(32'h3b49260b),
	.w6(32'hbc09db3c),
	.w7(32'hbc273050),
	.w8(32'h3b9b62e3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a094dc8),
	.w1(32'hbadc0b31),
	.w2(32'hbbdab7a6),
	.w3(32'hbc31d52c),
	.w4(32'hb9527b5d),
	.w5(32'h3bbf7de9),
	.w6(32'hbb3dd186),
	.w7(32'hbb848d0f),
	.w8(32'h3ba1eb24),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab006c),
	.w1(32'hb944bd51),
	.w2(32'hbb401525),
	.w3(32'h3b094473),
	.w4(32'h3c0b9c9d),
	.w5(32'hbb657756),
	.w6(32'h3b459c1c),
	.w7(32'h3b656406),
	.w8(32'h3b975aa8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10830),
	.w1(32'h3b95a7c6),
	.w2(32'h3bf4ca53),
	.w3(32'hbbbeddc2),
	.w4(32'h3bf22a03),
	.w5(32'h3cc82c6a),
	.w6(32'hbbfbfecf),
	.w7(32'h3b974a0c),
	.w8(32'h3cb08839),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f1a0e),
	.w1(32'h3c8fff06),
	.w2(32'hbba26df3),
	.w3(32'h3c94fc1d),
	.w4(32'hbbc031c8),
	.w5(32'hbb98b381),
	.w6(32'h3a06771b),
	.w7(32'hbc718e5b),
	.w8(32'hbb176612),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3493),
	.w1(32'hbb4eba2b),
	.w2(32'hbc312ed1),
	.w3(32'hbc22fbcb),
	.w4(32'h3bdb26f5),
	.w5(32'hbba93636),
	.w6(32'hbc2c6c1e),
	.w7(32'hbc103ab7),
	.w8(32'hbc246b4e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac35431),
	.w1(32'hbb2dc470),
	.w2(32'hbbbea6ac),
	.w3(32'hba839d69),
	.w4(32'h3c0652d0),
	.w5(32'hbb354e6f),
	.w6(32'h3963fef9),
	.w7(32'hbbe55a26),
	.w8(32'hbc129428),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08d5e8),
	.w1(32'h3a9860e8),
	.w2(32'h3ad233ae),
	.w3(32'h3ab92614),
	.w4(32'h3b0d8f18),
	.w5(32'hbb2bdd8b),
	.w6(32'h3abdcc23),
	.w7(32'h3baee313),
	.w8(32'h38919c4b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81cc12),
	.w1(32'h3c334c99),
	.w2(32'hbb708870),
	.w3(32'h3b86ddbb),
	.w4(32'h3b9b742f),
	.w5(32'h3bbb0d8f),
	.w6(32'h3c0f0dd2),
	.w7(32'hbbd5eca4),
	.w8(32'h3ba3646f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c245327),
	.w1(32'h3ba52ca1),
	.w2(32'hb9926495),
	.w3(32'h3b36ad38),
	.w4(32'hbc012bd3),
	.w5(32'hbb083fb0),
	.w6(32'hbb5017d3),
	.w7(32'hbb953a15),
	.w8(32'h3bb26f8a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1caf24),
	.w1(32'h3b73e628),
	.w2(32'hbb877e1d),
	.w3(32'h3b50a3f0),
	.w4(32'h3c0dfec1),
	.w5(32'h3c027b1c),
	.w6(32'hbbb90388),
	.w7(32'h3bc8101e),
	.w8(32'h3b1dcf4c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a6924),
	.w1(32'h3c13b43b),
	.w2(32'h3b9aef64),
	.w3(32'h3b66929f),
	.w4(32'h3b320bce),
	.w5(32'h3a2fc970),
	.w6(32'h3c75e285),
	.w7(32'h3b8effa1),
	.w8(32'hbae9f50f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05fa01),
	.w1(32'h3c120f1f),
	.w2(32'hba5402ed),
	.w3(32'h3c06bbc9),
	.w4(32'hba101310),
	.w5(32'h3c1fb60f),
	.w6(32'h3957fbcf),
	.w7(32'hbbb3240a),
	.w8(32'h3c3655a0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c763526),
	.w1(32'h3a52e7e5),
	.w2(32'hbc0400f7),
	.w3(32'hbac9c588),
	.w4(32'hbc0265d6),
	.w5(32'h3bbabf74),
	.w6(32'hbc5958a8),
	.w7(32'hbc768a60),
	.w8(32'hba58f673),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0610),
	.w1(32'hbb2a51d7),
	.w2(32'hbba68d5f),
	.w3(32'hbbbc211f),
	.w4(32'hbc21359b),
	.w5(32'hbbfe7736),
	.w6(32'hbbe6129b),
	.w7(32'hbc956cc6),
	.w8(32'hbc0d3e35),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37c19),
	.w1(32'hbbbb8cdd),
	.w2(32'hbb9f0307),
	.w3(32'hbc24cc52),
	.w4(32'hbab1a7a1),
	.w5(32'h3c0d6137),
	.w6(32'h3af63eac),
	.w7(32'hbb78c6a9),
	.w8(32'h3bc926f5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968a1a),
	.w1(32'hbbf3a96f),
	.w2(32'hbab7c165),
	.w3(32'hbc52b2e1),
	.w4(32'hbc6476ff),
	.w5(32'hba4e48ac),
	.w6(32'hbbfee9bc),
	.w7(32'hbc3996c5),
	.w8(32'h3ba42d5d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25448),
	.w1(32'hbbd1361c),
	.w2(32'h3b83ec96),
	.w3(32'hbc08d1d0),
	.w4(32'h3acf0309),
	.w5(32'hbc3eff76),
	.w6(32'hbc358118),
	.w7(32'hbb0a50e3),
	.w8(32'hbb1f70c8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e57b),
	.w1(32'hbc23c8a4),
	.w2(32'hbb948a56),
	.w3(32'hbc1f652d),
	.w4(32'hbc1fe8d5),
	.w5(32'hbaa881e5),
	.w6(32'hbc5601ac),
	.w7(32'hbc0dcd8c),
	.w8(32'h3a708aa6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ce43c),
	.w1(32'h3b408217),
	.w2(32'h3b4c8336),
	.w3(32'h391b4181),
	.w4(32'h3af14bed),
	.w5(32'h3b8d0bfc),
	.w6(32'hbc23a029),
	.w7(32'hbc031f3d),
	.w8(32'h3ba34044),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8f6a9),
	.w1(32'h3c190e05),
	.w2(32'hbbec8590),
	.w3(32'hbb2763c9),
	.w4(32'hbc07b279),
	.w5(32'hbb1b73cc),
	.w6(32'h3bd8cbd8),
	.w7(32'h3a822bb6),
	.w8(32'h3a8d003d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1cf1),
	.w1(32'h3b90d5cc),
	.w2(32'hba30c8f4),
	.w3(32'hbb547b09),
	.w4(32'hbb1a14bc),
	.w5(32'hbb2f0916),
	.w6(32'h3ad092d4),
	.w7(32'hbbda7541),
	.w8(32'hbb3879d0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfb1ec),
	.w1(32'hbbb8f969),
	.w2(32'hba7c5ef3),
	.w3(32'hbc09088d),
	.w4(32'hbc6158c0),
	.w5(32'hbb9aacd7),
	.w6(32'hbbaf3f23),
	.w7(32'hbc16d228),
	.w8(32'hbb6d7bdb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8821d6),
	.w1(32'h3be36957),
	.w2(32'h3b417e57),
	.w3(32'hba7582ef),
	.w4(32'h3c846408),
	.w5(32'h3c4b990b),
	.w6(32'h3b3b899e),
	.w7(32'h3bea9f04),
	.w8(32'h3bb5e057),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3f949),
	.w1(32'h3b2184b3),
	.w2(32'hbc286f9f),
	.w3(32'h38edb7b0),
	.w4(32'hbbc7c17d),
	.w5(32'h3b5cdcac),
	.w6(32'h3c353f25),
	.w7(32'hbc906bb6),
	.w8(32'hba399aa9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761048),
	.w1(32'h3bb8726d),
	.w2(32'h3a97ed2e),
	.w3(32'h3c1fe9c4),
	.w4(32'h3b8f20e3),
	.w5(32'hbb29a54d),
	.w6(32'h3c448c64),
	.w7(32'h3c1b5c0a),
	.w8(32'hbbdd6c1d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2616a6),
	.w1(32'hbb231bf7),
	.w2(32'hbb3cf284),
	.w3(32'hba188339),
	.w4(32'hbb25195c),
	.w5(32'h3baba907),
	.w6(32'hb87bdcd5),
	.w7(32'hbac77f4b),
	.w8(32'h3c5ec1dc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5c89e),
	.w1(32'hbb2ebe55),
	.w2(32'h3b1dfa5a),
	.w3(32'hbc775940),
	.w4(32'hbc3ebc4d),
	.w5(32'h3b79cead),
	.w6(32'hbca0bc62),
	.w7(32'hbc6d2e22),
	.w8(32'h3b4586cd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e96c),
	.w1(32'hbbe32c3f),
	.w2(32'h3aa12fe8),
	.w3(32'h3b0ec769),
	.w4(32'hbc15e124),
	.w5(32'hbc619087),
	.w6(32'h3bb1c6e7),
	.w7(32'hbb32064c),
	.w8(32'hbc2278dd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7447),
	.w1(32'hbba40f28),
	.w2(32'h3ae2f5df),
	.w3(32'hbc0fcdcd),
	.w4(32'hbc703f4c),
	.w5(32'hbb0b0404),
	.w6(32'hbc52054b),
	.w7(32'h3a14132a),
	.w8(32'hbba344e9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6df1f7),
	.w1(32'hb9fc0ae9),
	.w2(32'h3c121b34),
	.w3(32'h3b3f7f08),
	.w4(32'h3c3cb3ef),
	.w5(32'h3c80119b),
	.w6(32'hba909a1c),
	.w7(32'h3c7aab22),
	.w8(32'h3c971a90),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01996c),
	.w1(32'h3caa0e2f),
	.w2(32'hbb67b05d),
	.w3(32'h3c8224e3),
	.w4(32'hbb964d17),
	.w5(32'hb9e96087),
	.w6(32'h3bb89ffa),
	.w7(32'hbc55dc1a),
	.w8(32'hbb9420ea),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc09f),
	.w1(32'hbb12aded),
	.w2(32'hbb9f66b5),
	.w3(32'hbc5638be),
	.w4(32'hbb4f9f9b),
	.w5(32'hbae55a0c),
	.w6(32'hbb9648e5),
	.w7(32'hbbd4e923),
	.w8(32'h3a5404e4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e4678),
	.w1(32'h3bcc31ef),
	.w2(32'h3b41c368),
	.w3(32'h3b006d34),
	.w4(32'h3b04629c),
	.w5(32'hbc165ddc),
	.w6(32'h3bec52dd),
	.w7(32'hbc0c6e17),
	.w8(32'h3b2e410d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38083e42),
	.w1(32'h3bdc43e7),
	.w2(32'h3b851ddf),
	.w3(32'hba885800),
	.w4(32'hbc18b81b),
	.w5(32'hb91fd346),
	.w6(32'hbbe5baaf),
	.w7(32'hbc86bccb),
	.w8(32'hba0333ee),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0febd),
	.w1(32'h3b9f6b04),
	.w2(32'hbb476be5),
	.w3(32'h3b62096e),
	.w4(32'h3b1d7dd0),
	.w5(32'hb9bbc833),
	.w6(32'h3b603dd6),
	.w7(32'h3bced86c),
	.w8(32'h3aed9cad),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedca1d),
	.w1(32'hbba57178),
	.w2(32'h3b856199),
	.w3(32'h3a108d69),
	.w4(32'hbb89ece7),
	.w5(32'hbb3eda3f),
	.w6(32'hbbebe430),
	.w7(32'h3c188921),
	.w8(32'hb9cb84bd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc559ad),
	.w1(32'h3afeda33),
	.w2(32'hbb994784),
	.w3(32'hbbf05fed),
	.w4(32'hbbdd0932),
	.w5(32'h3bb9b354),
	.w6(32'hbb92de9e),
	.w7(32'hbc1d0605),
	.w8(32'hbb7ddb79),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c701b),
	.w1(32'hba2f42a4),
	.w2(32'hbbaf13ae),
	.w3(32'h3b21b448),
	.w4(32'h3b3e0d62),
	.w5(32'hbc50b418),
	.w6(32'h3b3d5067),
	.w7(32'hbc1c87e4),
	.w8(32'hbc53d1e9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f45db),
	.w1(32'hbb850195),
	.w2(32'hbb5ba68a),
	.w3(32'h3b141cfb),
	.w4(32'hbbd05540),
	.w5(32'hbb2c8b90),
	.w6(32'h3b7d75f0),
	.w7(32'hbba1f904),
	.w8(32'hbbd05a90),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50e97),
	.w1(32'hbb84267f),
	.w2(32'h3bba9767),
	.w3(32'hbb09d9b3),
	.w4(32'hbb0d8f78),
	.w5(32'h3c07c1e8),
	.w6(32'hbbc20453),
	.w7(32'hba5408bd),
	.w8(32'h3c343faa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f74d),
	.w1(32'hbc423016),
	.w2(32'hbaa5fa0f),
	.w3(32'hbc076b2a),
	.w4(32'hbab473a6),
	.w5(32'hba0e6349),
	.w6(32'hbceea2ea),
	.w7(32'hbbbcee28),
	.w8(32'h3c74a057),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28915),
	.w1(32'hbb062897),
	.w2(32'hb9f372a2),
	.w3(32'hbb95bdf6),
	.w4(32'h3b0376b7),
	.w5(32'h3b870e1b),
	.w6(32'h3ba7f79f),
	.w7(32'hbbe0a481),
	.w8(32'hba324106),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd19509),
	.w1(32'hbc7d93ab),
	.w2(32'hbb5efabc),
	.w3(32'hbc4a3705),
	.w4(32'hbc749159),
	.w5(32'hbac303d3),
	.w6(32'hbc2a8b44),
	.w7(32'hbb38421c),
	.w8(32'hbb449a32),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab18c3f),
	.w1(32'h3b507ade),
	.w2(32'h3bc4d65b),
	.w3(32'hb9847293),
	.w4(32'h3b145994),
	.w5(32'h3a542a41),
	.w6(32'h3aa192fb),
	.w7(32'h3a85de57),
	.w8(32'hbbc66c47),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18b286),
	.w1(32'hbb29cbb8),
	.w2(32'hba5a9fab),
	.w3(32'hbad71ae3),
	.w4(32'h39161245),
	.w5(32'hba8faa7b),
	.w6(32'h3ac1acd0),
	.w7(32'h3c1ab869),
	.w8(32'h3b41c6ad),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc630de),
	.w1(32'hbb09d625),
	.w2(32'h3bbabcf4),
	.w3(32'h3adb8d06),
	.w4(32'h3c09f11d),
	.w5(32'hbbe127b0),
	.w6(32'hbb884b48),
	.w7(32'hbae65d83),
	.w8(32'h3b0134b9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf868d),
	.w1(32'h3b944c30),
	.w2(32'h3c04825b),
	.w3(32'h3b5701e2),
	.w4(32'h3bc9bfbf),
	.w5(32'hbb7dd99e),
	.w6(32'h3bd262cf),
	.w7(32'h3b80caad),
	.w8(32'hbb57783e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16dc15),
	.w1(32'h3c4a2598),
	.w2(32'h3c0a6c38),
	.w3(32'h3bc83065),
	.w4(32'h3bf2e2d7),
	.w5(32'hbb2a554f),
	.w6(32'h3b3919c6),
	.w7(32'h3c76e51d),
	.w8(32'h3b57d464),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914b4b),
	.w1(32'hbb77361b),
	.w2(32'hbc0ec50c),
	.w3(32'h3c2784f5),
	.w4(32'h3ae4f6b6),
	.w5(32'hbbafc8a7),
	.w6(32'h3c9dc050),
	.w7(32'h3c0b7008),
	.w8(32'hbbd7ab43),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8833f5),
	.w1(32'hbc33705d),
	.w2(32'hbbc0702c),
	.w3(32'hbab6a50a),
	.w4(32'hbb6032c2),
	.w5(32'h3c4542e9),
	.w6(32'hbbd550a6),
	.w7(32'h3a56efc8),
	.w8(32'h3bf796ac),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5bdb6),
	.w1(32'h3b968a0d),
	.w2(32'hbbbd5e61),
	.w3(32'h3b86f3a5),
	.w4(32'hbb57d5af),
	.w5(32'hbbf54e4a),
	.w6(32'h3b06a29a),
	.w7(32'hbb615765),
	.w8(32'h3b93d529),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe8983),
	.w1(32'hbbc5256f),
	.w2(32'hbb45c222),
	.w3(32'hbba0ddad),
	.w4(32'hbc6f0e79),
	.w5(32'h3a51766a),
	.w6(32'hbbe1f930),
	.w7(32'hbc8eefca),
	.w8(32'h3bac932a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44cd01),
	.w1(32'h3b959613),
	.w2(32'h3b666464),
	.w3(32'h3b9b0bf8),
	.w4(32'h3baab78f),
	.w5(32'hbb4a3310),
	.w6(32'h3a00a88a),
	.w7(32'h3bb0fd70),
	.w8(32'hbb6fd2cc),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0ae5),
	.w1(32'h39b65e38),
	.w2(32'h3c15b5b5),
	.w3(32'h3aa402e4),
	.w4(32'hbb516ed7),
	.w5(32'hbb3b4950),
	.w6(32'h3b813cd9),
	.w7(32'h3971f3c8),
	.w8(32'hbb046b6a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbf564),
	.w1(32'hbbed0d53),
	.w2(32'hbbacbd27),
	.w3(32'hbbb522c6),
	.w4(32'hbb195854),
	.w5(32'hbbfc8d08),
	.w6(32'hbb059b72),
	.w7(32'h3920ca00),
	.w8(32'hbb4b36da),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5df36),
	.w1(32'hbb97a3fc),
	.w2(32'h3b70c37b),
	.w3(32'h3bd4940b),
	.w4(32'hbb285471),
	.w5(32'hbc0bceab),
	.w6(32'h3a044bc7),
	.w7(32'hbb5fa7be),
	.w8(32'hbc630916),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72ca1b),
	.w1(32'hbc646475),
	.w2(32'hbc00bcbc),
	.w3(32'hbc20e626),
	.w4(32'hbbd72d9f),
	.w5(32'h3b4e9e4a),
	.w6(32'hbb7318e6),
	.w7(32'hbc5db902),
	.w8(32'h3a9904bc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e849c),
	.w1(32'h3a229c99),
	.w2(32'hbb35db0d),
	.w3(32'hbb8263c8),
	.w4(32'h3bf9e05e),
	.w5(32'hbbea1bd6),
	.w6(32'hba3cf424),
	.w7(32'h3b3fd3d4),
	.w8(32'hbb226d99),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0449c6),
	.w1(32'h395364bc),
	.w2(32'hbb352fee),
	.w3(32'hbc0af380),
	.w4(32'h3c01a7ac),
	.w5(32'hbb58fb91),
	.w6(32'hbb9b2caa),
	.w7(32'hbb470072),
	.w8(32'hbbc9fd95),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e624),
	.w1(32'h39a3f556),
	.w2(32'hba52d19a),
	.w3(32'hbb1e7ac7),
	.w4(32'h3a93e806),
	.w5(32'hb9eece0d),
	.w6(32'hbb4a1d6f),
	.w7(32'h3c2c5aef),
	.w8(32'hba4397bc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfbb77),
	.w1(32'hbc55863b),
	.w2(32'h3aff0bca),
	.w3(32'hbc102a93),
	.w4(32'hbba4cce8),
	.w5(32'h3bcdd1e7),
	.w6(32'hbaf41d35),
	.w7(32'hbbca330d),
	.w8(32'h3c2faf4c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38cc3a),
	.w1(32'h3bfe5a5b),
	.w2(32'h3addfc74),
	.w3(32'h3bcf7794),
	.w4(32'h3b70a5fd),
	.w5(32'hbc652cfa),
	.w6(32'hbaf67965),
	.w7(32'h3a9002f0),
	.w8(32'hbce40160),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc585b34),
	.w1(32'h3b7f2026),
	.w2(32'h3bd85ff8),
	.w3(32'h3c95eca3),
	.w4(32'h3cdacd4b),
	.w5(32'h3b35b960),
	.w6(32'h3c9e0d90),
	.w7(32'h3d50ceb3),
	.w8(32'h3c0d06c5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e445),
	.w1(32'hbbe0d7f2),
	.w2(32'h3b7969e6),
	.w3(32'hbbb2e80c),
	.w4(32'hbc5edd1d),
	.w5(32'hbc306401),
	.w6(32'h3ba009f0),
	.w7(32'hbc03d6e6),
	.w8(32'h3ac6b4cb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a7e9b),
	.w1(32'hbb400183),
	.w2(32'hb9f794ad),
	.w3(32'hbbee63ed),
	.w4(32'hbaf61d59),
	.w5(32'h3be4465f),
	.w6(32'hbb8b5724),
	.w7(32'hb793fb54),
	.w8(32'h3c1e4958),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc7b6),
	.w1(32'h3953145e),
	.w2(32'hbb75a9d7),
	.w3(32'h3b198ebb),
	.w4(32'h3b89f1d7),
	.w5(32'hbaaace55),
	.w6(32'h3b69cd9d),
	.w7(32'hbb9816a1),
	.w8(32'hba643b30),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8dfd),
	.w1(32'hba506fdb),
	.w2(32'hbb8543bb),
	.w3(32'hbbdcf10f),
	.w4(32'hbb91db5c),
	.w5(32'h3b07d152),
	.w6(32'hba117f94),
	.w7(32'hbbce653b),
	.w8(32'h3a16ec15),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab9183),
	.w1(32'h3b206830),
	.w2(32'hba7a6bf9),
	.w3(32'hbb7cd967),
	.w4(32'h3c69b5b9),
	.w5(32'hb93bf99d),
	.w6(32'hbbbc3e47),
	.w7(32'hbb8b9a30),
	.w8(32'h3b9060cd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ee785),
	.w1(32'hbc0db37e),
	.w2(32'hbbb1bf72),
	.w3(32'h3b4ff3cf),
	.w4(32'h3b074cf3),
	.w5(32'h3bb08de7),
	.w6(32'h39c23ab3),
	.w7(32'hbb9ad572),
	.w8(32'h3c065e47),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcd5ac),
	.w1(32'hbbd5e668),
	.w2(32'hbbc77c57),
	.w3(32'hba92b3ce),
	.w4(32'h3ac3f81a),
	.w5(32'hba3d2eef),
	.w6(32'hb93c188b),
	.w7(32'hbc334396),
	.w8(32'h3b2325d6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedabd3),
	.w1(32'hbc09b9bb),
	.w2(32'hbb8976a9),
	.w3(32'hbb993b89),
	.w4(32'hbc1d4afe),
	.w5(32'hbbb07291),
	.w6(32'hbb21dc3e),
	.w7(32'hbb4b390c),
	.w8(32'hbb702bb3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241e14),
	.w1(32'hbaf50a2d),
	.w2(32'h3bdb01be),
	.w3(32'hbc0ac7d3),
	.w4(32'h3b16657f),
	.w5(32'hbc27f68a),
	.w6(32'hbbe3121f),
	.w7(32'h3bebcf22),
	.w8(32'hbbb6adea),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf5f7),
	.w1(32'h3ab60cca),
	.w2(32'hb9ced9ad),
	.w3(32'h3be2ab22),
	.w4(32'h3ba0e707),
	.w5(32'h3b17668d),
	.w6(32'h3c02cd7f),
	.w7(32'h3b927435),
	.w8(32'hbbc686a7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c515),
	.w1(32'h3b9ba87b),
	.w2(32'h3c2f1be3),
	.w3(32'h3bb32613),
	.w4(32'h3b8d1f40),
	.w5(32'h3aa37e5f),
	.w6(32'h3bacb7ce),
	.w7(32'h3c1e64e7),
	.w8(32'h3b91facb),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86759),
	.w1(32'hbbdc17d1),
	.w2(32'hbc50d7b0),
	.w3(32'h3ba9d0ed),
	.w4(32'hbc9bebf1),
	.w5(32'h3c34210b),
	.w6(32'h3bd5ebac),
	.w7(32'hbc9c2168),
	.w8(32'h3bf0f493),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e745c),
	.w1(32'h3c2c5264),
	.w2(32'h3bc0787e),
	.w3(32'h3c81243a),
	.w4(32'h3ab61a07),
	.w5(32'h3be21dd0),
	.w6(32'hbbcac5dc),
	.w7(32'hbbb58e92),
	.w8(32'hbaff86f0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8133),
	.w1(32'h3b2b2232),
	.w2(32'h378ec067),
	.w3(32'hbb8705a7),
	.w4(32'hb95ecaf0),
	.w5(32'h3c1b4854),
	.w6(32'h3baf9dc9),
	.w7(32'hbbfa76e8),
	.w8(32'h3c6bd390),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c553a35),
	.w1(32'hbb8e53e9),
	.w2(32'h3b0f33b7),
	.w3(32'hbc02acba),
	.w4(32'h3c08db42),
	.w5(32'h3c3fc2a8),
	.w6(32'hbc7d7163),
	.w7(32'h3b750438),
	.w8(32'h3c4e7dab),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e77a1),
	.w1(32'h3adb9efe),
	.w2(32'h3baa1c60),
	.w3(32'hbb97f762),
	.w4(32'hbc48ce9b),
	.w5(32'hbbaa24fb),
	.w6(32'h3b937b7f),
	.w7(32'hba658a88),
	.w8(32'hbbd2e279),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1adf1),
	.w1(32'hbb2a6fd2),
	.w2(32'h3b6fddb0),
	.w3(32'h3acb9dcc),
	.w4(32'hbb97b1b8),
	.w5(32'hbc1fbb26),
	.w6(32'h3a4d0027),
	.w7(32'hb9dd60d9),
	.w8(32'hbc2afe04),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9e912),
	.w1(32'hbbd28de6),
	.w2(32'hbbf8625f),
	.w3(32'hbb46d7c6),
	.w4(32'hbbf17a87),
	.w5(32'hbb3cb109),
	.w6(32'hba8707af),
	.w7(32'hbb1b17cc),
	.w8(32'h3ab2578c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a0bd),
	.w1(32'hbbfec590),
	.w2(32'hbb1d350e),
	.w3(32'h3bc32f4a),
	.w4(32'hbc072bb6),
	.w5(32'h3b68c06e),
	.w6(32'hb9226d3c),
	.w7(32'hbc061205),
	.w8(32'h3bed4fe6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c043bfb),
	.w1(32'hb93db9ad),
	.w2(32'hbbe90a72),
	.w3(32'h3b449272),
	.w4(32'hbc23ac36),
	.w5(32'hbb8ceb28),
	.w6(32'hbb8e896e),
	.w7(32'hbc14a263),
	.w8(32'hbc8d926d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7121c),
	.w1(32'h39a863e2),
	.w2(32'h3b8c2002),
	.w3(32'h3bacbff5),
	.w4(32'h3c8c2666),
	.w5(32'h3af9a644),
	.w6(32'h3b39f82a),
	.w7(32'h3c3cc866),
	.w8(32'h3c475018),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3044),
	.w1(32'h3b5d0a2c),
	.w2(32'h3ba05f24),
	.w3(32'hbb9953b0),
	.w4(32'hbacf8263),
	.w5(32'hbb8cf4fb),
	.w6(32'h39c020d2),
	.w7(32'hbb41982a),
	.w8(32'hbbb79e91),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83d68),
	.w1(32'hbbd88d9c),
	.w2(32'h3b388307),
	.w3(32'hba8bd457),
	.w4(32'hbbc82fb0),
	.w5(32'h3a7e84f7),
	.w6(32'hbb20641b),
	.w7(32'hbbf2fe0a),
	.w8(32'hbbd85806),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c678),
	.w1(32'hba6c5281),
	.w2(32'hbb9b6a84),
	.w3(32'hbc0fda01),
	.w4(32'hbc0f1a4a),
	.w5(32'h3b5c8e9b),
	.w6(32'hbc13a340),
	.w7(32'hbc5ad727),
	.w8(32'hbbe82cef),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d117),
	.w1(32'hb9859943),
	.w2(32'hbac81468),
	.w3(32'hb89ddc7b),
	.w4(32'hbac8cf97),
	.w5(32'h3b47d028),
	.w6(32'hbb8c2988),
	.w7(32'hbbe8198c),
	.w8(32'h3a415bcf),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac1eb),
	.w1(32'h3a024394),
	.w2(32'h3b1ebb4d),
	.w3(32'h3ba88caa),
	.w4(32'h3b98c706),
	.w5(32'hbc3db22a),
	.w6(32'h3b7fea9d),
	.w7(32'hbb1c5e4c),
	.w8(32'hbc40bf9e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d619f),
	.w1(32'hbcdaa0d4),
	.w2(32'hbb404bb0),
	.w3(32'hbc5f2fb4),
	.w4(32'hbc0caba4),
	.w5(32'h3b47a883),
	.w6(32'hbc932242),
	.w7(32'h3bab9f79),
	.w8(32'h3c35d9b1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2417eb),
	.w1(32'h3a78ed05),
	.w2(32'hbaa8c0ee),
	.w3(32'hbb704622),
	.w4(32'h3a537348),
	.w5(32'h3b45fd06),
	.w6(32'h3bb5c81c),
	.w7(32'h3b012ca8),
	.w8(32'h3bcea22d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf500f),
	.w1(32'h3c5aa2f1),
	.w2(32'h3b0fa6b4),
	.w3(32'h3b46b9b2),
	.w4(32'hba583606),
	.w5(32'h3bb14ef7),
	.w6(32'h3b24db41),
	.w7(32'h39ae19ca),
	.w8(32'h3b5e5089),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7ec45),
	.w1(32'hbbc9d5ca),
	.w2(32'hba0b3ff8),
	.w3(32'hbc7ba994),
	.w4(32'hbc5096e7),
	.w5(32'h3cd772a4),
	.w6(32'hbcdbb004),
	.w7(32'hbc8aacb1),
	.w8(32'h3c8b3b70),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4db52c),
	.w1(32'h3a51968a),
	.w2(32'hbc34070d),
	.w3(32'h3a9001af),
	.w4(32'hbbffc8d0),
	.w5(32'h391c3419),
	.w6(32'hbc3bd67f),
	.w7(32'hbc79c87b),
	.w8(32'hbb194138),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9839e70),
	.w1(32'hbb4338db),
	.w2(32'hbb839e39),
	.w3(32'hba57a870),
	.w4(32'h3b0cd723),
	.w5(32'hbbda341e),
	.w6(32'hbb08a0a5),
	.w7(32'hbb1bff62),
	.w8(32'h3ad5a36e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d093),
	.w1(32'h3b8d2b14),
	.w2(32'hbc318444),
	.w3(32'h3b171067),
	.w4(32'hba7aaa20),
	.w5(32'hbacc8062),
	.w6(32'h3b88750a),
	.w7(32'h3b8a81fc),
	.w8(32'hbc3e6588),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33c7c6),
	.w1(32'hbc462a50),
	.w2(32'hbb66021c),
	.w3(32'h3a4ee4de),
	.w4(32'h39f3075e),
	.w5(32'h3c065470),
	.w6(32'hbb876e56),
	.w7(32'h3b820877),
	.w8(32'h3ba84fd7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39d013),
	.w1(32'h3bead6cb),
	.w2(32'hbc1cfea8),
	.w3(32'h3c0bc4e2),
	.w4(32'hbc33d53a),
	.w5(32'h3a193d98),
	.w6(32'hbbdb12e7),
	.w7(32'hbc9bf8af),
	.w8(32'h3a23f4bb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd43d),
	.w1(32'h3b285da3),
	.w2(32'hbc135286),
	.w3(32'hb95e33cb),
	.w4(32'h3c428665),
	.w5(32'hbb456690),
	.w6(32'h3ac21e9d),
	.w7(32'hbbd32cbf),
	.w8(32'hbb650e12),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecfc6d),
	.w1(32'hbbaad376),
	.w2(32'hbb314cee),
	.w3(32'h3703006f),
	.w4(32'hbb322a20),
	.w5(32'h3b219557),
	.w6(32'hbb7cd475),
	.w7(32'h3a0cfb07),
	.w8(32'hbc18387f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca200cf),
	.w1(32'h3c5d0bc7),
	.w2(32'h3c07d377),
	.w3(32'h3b7a7a6b),
	.w4(32'hbb6c4eef),
	.w5(32'h3b6bb301),
	.w6(32'h3a472fec),
	.w7(32'h3c1af727),
	.w8(32'h3a4f8b06),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f85f6c),
	.w1(32'h3a0b1f60),
	.w2(32'h3b00d899),
	.w3(32'h3a2a5536),
	.w4(32'h3b99ab1e),
	.w5(32'hbc1793e3),
	.w6(32'hbb4a24a9),
	.w7(32'h3a371c4e),
	.w8(32'hbc7aa642),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae5c98),
	.w1(32'h3bae00bc),
	.w2(32'h39d63e2a),
	.w3(32'h3ba228c2),
	.w4(32'hbb09fb5c),
	.w5(32'h3bb6ca4a),
	.w6(32'h3c02b5c4),
	.w7(32'h3becaaff),
	.w8(32'h3ad24284),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0649f),
	.w1(32'hbb58f76d),
	.w2(32'h3afee4e2),
	.w3(32'hbb97c13b),
	.w4(32'hbbaf64fa),
	.w5(32'hbb6254db),
	.w6(32'hbbce1730),
	.w7(32'hbb83ba75),
	.w8(32'hbb906c2e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabadaa9),
	.w1(32'hb95ed621),
	.w2(32'h3aa264b8),
	.w3(32'hbbffef9c),
	.w4(32'hbb4d8049),
	.w5(32'hba2c74f3),
	.w6(32'hbc228c84),
	.w7(32'h3bbec279),
	.w8(32'h3a98cefa),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c536b01),
	.w1(32'hbb802e98),
	.w2(32'hbbc844ae),
	.w3(32'h3c39ed4d),
	.w4(32'hbaa7d21f),
	.w5(32'h3b549d85),
	.w6(32'h3c33ebda),
	.w7(32'hbc25c8a9),
	.w8(32'h3b41d683),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac37a7),
	.w1(32'h3b7af340),
	.w2(32'h39945975),
	.w3(32'h3a824cea),
	.w4(32'h3a485dc2),
	.w5(32'h3bc63afc),
	.w6(32'h3c4215d4),
	.w7(32'h3c954384),
	.w8(32'h3c21f7f8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ef6f),
	.w1(32'hbbab8eff),
	.w2(32'hbb565f7f),
	.w3(32'hbaace8a9),
	.w4(32'hbaec131d),
	.w5(32'hbc974de4),
	.w6(32'h3b75eaed),
	.w7(32'h3b003f79),
	.w8(32'hbc8da550),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc309e40),
	.w1(32'h3bf964ba),
	.w2(32'h3c440dd6),
	.w3(32'hbbd1f04a),
	.w4(32'hbb0a1c91),
	.w5(32'hbaa09df4),
	.w6(32'hba07040a),
	.w7(32'h3c0c71d0),
	.w8(32'hbb8c9196),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837e1f),
	.w1(32'hbc02f6a0),
	.w2(32'h3aea9826),
	.w3(32'hbb98bc52),
	.w4(32'h3a79b6d9),
	.w5(32'hbbc5824d),
	.w6(32'hb9971136),
	.w7(32'h3c597ee7),
	.w8(32'hbc18bd1f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb639242),
	.w1(32'hbbd4a9d4),
	.w2(32'h3a369a0c),
	.w3(32'hbb3771d9),
	.w4(32'hbb848633),
	.w5(32'h3bef882c),
	.w6(32'hbc1a85e4),
	.w7(32'hba84364d),
	.w8(32'h3a911f7b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0479e4),
	.w1(32'hbad1303b),
	.w2(32'hbb3635f1),
	.w3(32'hbb5373af),
	.w4(32'h3b3482e0),
	.w5(32'h38bf2f64),
	.w6(32'hbb8c8915),
	.w7(32'h39b0f0f2),
	.w8(32'h3a99d76d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dfb77),
	.w1(32'h3b218e8d),
	.w2(32'h3b54cc4e),
	.w3(32'h3bcebc24),
	.w4(32'h3bc5112c),
	.w5(32'hbb93e038),
	.w6(32'h3b274708),
	.w7(32'h3b606f51),
	.w8(32'hbb7ee810),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307d5e),
	.w1(32'hbb999283),
	.w2(32'h3a8c50ff),
	.w3(32'hb9e09e19),
	.w4(32'h3bf2fdc2),
	.w5(32'hbb1dc684),
	.w6(32'hbbe4c579),
	.w7(32'h3b3e3dc4),
	.w8(32'h3a8fccc3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa1ad3),
	.w1(32'hbc24df8a),
	.w2(32'hbc1eda22),
	.w3(32'h3b1df989),
	.w4(32'hbb8b8a3a),
	.w5(32'hbb7cb4ae),
	.w6(32'h3c969418),
	.w7(32'hbc37f453),
	.w8(32'hbb6de77a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81a51),
	.w1(32'hbb9febc9),
	.w2(32'h3b49834c),
	.w3(32'hba2ca38c),
	.w4(32'h3b5242c0),
	.w5(32'h3b8a63fd),
	.w6(32'hbc09d663),
	.w7(32'hbbad6c6c),
	.w8(32'hbad02f6b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ae125),
	.w1(32'hba58b634),
	.w2(32'h3bb8866e),
	.w3(32'h3b42e886),
	.w4(32'hba9e192b),
	.w5(32'h3b390a4b),
	.w6(32'hbbdde0fa),
	.w7(32'hbacebbde),
	.w8(32'hbc14f970),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64213f),
	.w1(32'h3c0b4aa8),
	.w2(32'hbb66495c),
	.w3(32'h3a44c1f7),
	.w4(32'hbbf80485),
	.w5(32'hba81c88e),
	.w6(32'h3b455a10),
	.w7(32'hbbeca4ab),
	.w8(32'hbb911c47),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30679),
	.w1(32'hbb747fa6),
	.w2(32'hbc2124ca),
	.w3(32'h3b6f130c),
	.w4(32'h3b05979c),
	.w5(32'hbb9e296a),
	.w6(32'h3c875281),
	.w7(32'hba9f871e),
	.w8(32'hbb7ec49d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc45c),
	.w1(32'hbb570711),
	.w2(32'hbb69a30c),
	.w3(32'h3a4f8cb8),
	.w4(32'h3a96b48b),
	.w5(32'h3a9c6b1e),
	.w6(32'hbaac6e96),
	.w7(32'hbabf612d),
	.w8(32'h3b100d5a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb81c5),
	.w1(32'hbb50a8ef),
	.w2(32'h3b395d78),
	.w3(32'hbbb8b69e),
	.w4(32'hbba2c970),
	.w5(32'hba8df866),
	.w6(32'hbbcc21f4),
	.w7(32'h3b67e2d2),
	.w8(32'h3678ebcb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118f36),
	.w1(32'h39cacfea),
	.w2(32'hbb83d9c1),
	.w3(32'h3aa3563f),
	.w4(32'h3991dc6e),
	.w5(32'hbb0ccebd),
	.w6(32'hbab4c527),
	.w7(32'h3aba8db2),
	.w8(32'hbc4d42d9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90590),
	.w1(32'h3b48c40f),
	.w2(32'h3a76f581),
	.w3(32'hbb2659b4),
	.w4(32'hb80a3d6a),
	.w5(32'hbb530463),
	.w6(32'h3ae717cc),
	.w7(32'h3b6103f3),
	.w8(32'hbba7cf4d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cc155),
	.w1(32'h3c1a44d9),
	.w2(32'hbc51a87c),
	.w3(32'h3c3ab07d),
	.w4(32'h3b44dc94),
	.w5(32'h3ba6e5a1),
	.w6(32'h3d4e6606),
	.w7(32'hbae51e56),
	.w8(32'h3b7e2fe3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ad59),
	.w1(32'h3c23cf7f),
	.w2(32'h38c67820),
	.w3(32'h3bd5dcfc),
	.w4(32'hba6bf55b),
	.w5(32'hbb0757bd),
	.w6(32'h3c590468),
	.w7(32'hbbbb7137),
	.w8(32'hbb2845a7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a18b8),
	.w1(32'hbba37731),
	.w2(32'hbb350d84),
	.w3(32'hbb5d5bba),
	.w4(32'hbb5afb99),
	.w5(32'hba28b374),
	.w6(32'hbc2df089),
	.w7(32'hba64e91a),
	.w8(32'h393bde5f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb747b),
	.w1(32'h3acfb054),
	.w2(32'h3baaa3a2),
	.w3(32'hbb1dbcef),
	.w4(32'h3b37aca7),
	.w5(32'h3b62fd29),
	.w6(32'hbb6cbf16),
	.w7(32'h3b309507),
	.w8(32'hbb301040),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c58c7),
	.w1(32'h3a802ab4),
	.w2(32'h3b853274),
	.w3(32'hbb12c68c),
	.w4(32'h392423a7),
	.w5(32'h3c404228),
	.w6(32'hbb28539d),
	.w7(32'hba4d84f5),
	.w8(32'h3a8f8925),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afcd3),
	.w1(32'hbae6516f),
	.w2(32'hbb37e9c8),
	.w3(32'h3ad9245a),
	.w4(32'hbc07ae5b),
	.w5(32'hbc00a72f),
	.w6(32'hbc03b507),
	.w7(32'hbb95df9b),
	.w8(32'hbba5ece1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a077829),
	.w1(32'hbae24f56),
	.w2(32'hba4815fe),
	.w3(32'hbb8aaf32),
	.w4(32'h3989e372),
	.w5(32'h3acd6757),
	.w6(32'hbb379d56),
	.w7(32'h3b117dd5),
	.w8(32'h3a8ccfa1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95ae0c),
	.w1(32'hbb008a92),
	.w2(32'hbbbbc255),
	.w3(32'hbbb2ac28),
	.w4(32'hbc38e12d),
	.w5(32'hbb779d43),
	.w6(32'hbac9ddf1),
	.w7(32'hbc3b2ea5),
	.w8(32'hbc16929e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule