module layer_10_featuremap_337(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c373),
	.w1(32'h3c889757),
	.w2(32'h3c0b68c4),
	.w3(32'hbb460e63),
	.w4(32'hb9b90953),
	.w5(32'hbc0cc925),
	.w6(32'h3a6340c3),
	.w7(32'h3be25e95),
	.w8(32'hbba47a6c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244be1),
	.w1(32'hbb629a96),
	.w2(32'hbaf7682b),
	.w3(32'hbb373330),
	.w4(32'h3ad5e576),
	.w5(32'hbac167c1),
	.w6(32'hbb9d8471),
	.w7(32'h3abee11b),
	.w8(32'hbb90cd31),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d487),
	.w1(32'hba48432f),
	.w2(32'hbb9afbf8),
	.w3(32'h3bc0b3a3),
	.w4(32'h3b3bdc30),
	.w5(32'hbb30e4e0),
	.w6(32'hbb1105c7),
	.w7(32'h3b112662),
	.w8(32'hbb37c653),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dbf42),
	.w1(32'hba878c29),
	.w2(32'hbb749aba),
	.w3(32'hbb480381),
	.w4(32'hbb63657f),
	.w5(32'hbacf9314),
	.w6(32'hbb08aacf),
	.w7(32'hbb41752b),
	.w8(32'h3bc88ce7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f69792),
	.w1(32'h38cecea7),
	.w2(32'hbba73f20),
	.w3(32'hba8d6ddf),
	.w4(32'hba97cbbf),
	.w5(32'hbbaf7c33),
	.w6(32'h38ac852b),
	.w7(32'h3b802ec3),
	.w8(32'hbb7c1370),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f837e),
	.w1(32'h3ba6351a),
	.w2(32'hb9a9c43b),
	.w3(32'hba59bf98),
	.w4(32'h3ad725d0),
	.w5(32'h3b7554be),
	.w6(32'hbad7e803),
	.w7(32'hbb3dbdc3),
	.w8(32'h3bcdefd3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3352f),
	.w1(32'h3b019ad7),
	.w2(32'h3b002c7c),
	.w3(32'hbaf664aa),
	.w4(32'h3af4dcf8),
	.w5(32'hbb04c7c3),
	.w6(32'hbb3e4a0b),
	.w7(32'h3a64b80d),
	.w8(32'h3aec0674),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40345e),
	.w1(32'h3c15df44),
	.w2(32'h3ba16e88),
	.w3(32'hbbc92cd7),
	.w4(32'hbbe6f481),
	.w5(32'h3ad1c734),
	.w6(32'h3ab7298e),
	.w7(32'hba429a87),
	.w8(32'h39bce48a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0de481),
	.w1(32'h3b89ded8),
	.w2(32'h3b53c258),
	.w3(32'h3b048c1f),
	.w4(32'h3b41f02a),
	.w5(32'hbb9b2035),
	.w6(32'hb6610138),
	.w7(32'h3b5a5089),
	.w8(32'hbb83a392),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962a7f7),
	.w1(32'h3b89c3ad),
	.w2(32'h3ae51d3d),
	.w3(32'h38dcb345),
	.w4(32'h3b8759b6),
	.w5(32'hbc19aada),
	.w6(32'hba93383a),
	.w7(32'hba6e7b68),
	.w8(32'hbc0a0156),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c1a2),
	.w1(32'h3b291810),
	.w2(32'hb995ef55),
	.w3(32'hbbbaa9eb),
	.w4(32'hbb21eab1),
	.w5(32'hbb144643),
	.w6(32'hbbb060c4),
	.w7(32'hbb3aa43b),
	.w8(32'hbba5768e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1e7cb),
	.w1(32'hbb511b08),
	.w2(32'h3aa4d950),
	.w3(32'hbb0846ab),
	.w4(32'hbb3a8dc6),
	.w5(32'h3b0a0737),
	.w6(32'hbb0aebbf),
	.w7(32'hbbe71da2),
	.w8(32'h3bb93b3c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985af67),
	.w1(32'h3b88e19b),
	.w2(32'hb99a165c),
	.w3(32'h3b3be6aa),
	.w4(32'hbb463818),
	.w5(32'hbc1b007b),
	.w6(32'h3c0b961a),
	.w7(32'h3c0b1913),
	.w8(32'hbc67c240),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdea2ab),
	.w1(32'hb96c4ef0),
	.w2(32'h3bff01ca),
	.w3(32'hbb5d22a6),
	.w4(32'h3bc64bdc),
	.w5(32'hbae12b7a),
	.w6(32'hbbc904a3),
	.w7(32'h3c4857c7),
	.w8(32'hbb56e517),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6ef8),
	.w1(32'h396a95a0),
	.w2(32'hbb0a9d78),
	.w3(32'hbb79bc61),
	.w4(32'hbb06fe3d),
	.w5(32'hbc43e2b1),
	.w6(32'hb9904c79),
	.w7(32'hbaf78084),
	.w8(32'hbc5cfd1b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecfbb5),
	.w1(32'h3a78409a),
	.w2(32'hbbe363c0),
	.w3(32'hbc0e65d9),
	.w4(32'hbb82299e),
	.w5(32'hbba95090),
	.w6(32'hbb5b9e62),
	.w7(32'hbc3bc033),
	.w8(32'h3b95f848),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8db770),
	.w1(32'h3b1174df),
	.w2(32'hbb0af0be),
	.w3(32'hba6fc242),
	.w4(32'hba2d82d1),
	.w5(32'hba8cb01b),
	.w6(32'h3acef344),
	.w7(32'hbb2ecd54),
	.w8(32'hb9ea1175),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf58664),
	.w1(32'h3a9b57c3),
	.w2(32'h3b365996),
	.w3(32'h3ad47679),
	.w4(32'h3b10a022),
	.w5(32'hbb7fcb8c),
	.w6(32'h3a476fd3),
	.w7(32'h3b8958d8),
	.w8(32'hbb6e0475),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad82342),
	.w1(32'h3aa3d44e),
	.w2(32'hbb1821d5),
	.w3(32'hbb7b388b),
	.w4(32'hbae1ee8c),
	.w5(32'hba951bf8),
	.w6(32'hbb53e94f),
	.w7(32'hbb98b1ec),
	.w8(32'h3b74e8f7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb028baa),
	.w1(32'hb8d0ee86),
	.w2(32'h3accac10),
	.w3(32'hbc109e58),
	.w4(32'hbb85e982),
	.w5(32'h3b74479c),
	.w6(32'hbc334a8f),
	.w7(32'hbb4c1dec),
	.w8(32'h3aa089d8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9174a),
	.w1(32'h3b41cd9e),
	.w2(32'hb924fbd4),
	.w3(32'hbb0f4c10),
	.w4(32'h3b59a6c0),
	.w5(32'h3b7651f8),
	.w6(32'hbbd8b302),
	.w7(32'hbb3faa58),
	.w8(32'h3bd1448b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53abe9),
	.w1(32'hbb4c07e4),
	.w2(32'hbb4d4cdd),
	.w3(32'h3a9cc5ac),
	.w4(32'hba963317),
	.w5(32'hb92e8abd),
	.w6(32'h3aded4b7),
	.w7(32'hbaa2d58d),
	.w8(32'hbbcfe9c1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba905208),
	.w1(32'h3b22f3ba),
	.w2(32'h3b085fe1),
	.w3(32'h3b755ada),
	.w4(32'h39991a4b),
	.w5(32'hbc17fc2f),
	.w6(32'h3b1948e2),
	.w7(32'hbb67c87d),
	.w8(32'hbc7b83af),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab11e),
	.w1(32'hbbd35c48),
	.w2(32'hbb356bf3),
	.w3(32'hbc28fb40),
	.w4(32'hbc04507c),
	.w5(32'hbbb531e4),
	.w6(32'hbc2949bf),
	.w7(32'hbc4693e0),
	.w8(32'h39008abf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfaa8f),
	.w1(32'h3b659dc4),
	.w2(32'h3b32ae8a),
	.w3(32'h3b1b23f5),
	.w4(32'h3c2fb935),
	.w5(32'hbb709df3),
	.w6(32'h394515b5),
	.w7(32'hb793e3ff),
	.w8(32'h3a1b8db2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a958042),
	.w1(32'h3b244345),
	.w2(32'hbab89fdf),
	.w3(32'hbb822708),
	.w4(32'hba66b10c),
	.w5(32'h3a97bdc5),
	.w6(32'h3b166474),
	.w7(32'hbb8e2252),
	.w8(32'h3b51432a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b441b11),
	.w1(32'h3a0b0b88),
	.w2(32'hba309b6d),
	.w3(32'h3a0b19a7),
	.w4(32'h3a2b5336),
	.w5(32'h3b8f32e3),
	.w6(32'h3ad83467),
	.w7(32'h3a773cca),
	.w8(32'h3b41c11f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83262),
	.w1(32'h3c03d73a),
	.w2(32'h3b50e1f9),
	.w3(32'h3bf17d8f),
	.w4(32'h3b92560c),
	.w5(32'hbb82b762),
	.w6(32'h3b81a20e),
	.w7(32'h3c03a12e),
	.w8(32'hbb02cb46),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba996c1),
	.w1(32'h3bfb6f6a),
	.w2(32'h3c7d1750),
	.w3(32'h3b90eb54),
	.w4(32'h3c8cd2f6),
	.w5(32'hbbbbf75e),
	.w6(32'h3affc07e),
	.w7(32'h3c9925d3),
	.w8(32'hbb820858),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1487f0),
	.w1(32'h3ba15a70),
	.w2(32'h3ba9cee1),
	.w3(32'hbb4ec448),
	.w4(32'h3adf07cf),
	.w5(32'h3a44ef55),
	.w6(32'h3af18a70),
	.w7(32'h3c4cd983),
	.w8(32'hbbfb5d18),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45c1d1),
	.w1(32'h3bbeaec9),
	.w2(32'h3b717e95),
	.w3(32'h3a033403),
	.w4(32'hb9d1cc73),
	.w5(32'h3c0dc033),
	.w6(32'h39fda20e),
	.w7(32'h3b5ab835),
	.w8(32'h3c10ce79),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f9e41),
	.w1(32'hbb6e651f),
	.w2(32'h3ba4f4cb),
	.w3(32'h3be14231),
	.w4(32'h3bd1b1cf),
	.w5(32'h3a537469),
	.w6(32'h3b99fff8),
	.w7(32'h3b86f8a8),
	.w8(32'h3bf52da0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d60dc),
	.w1(32'h3ba34e38),
	.w2(32'h3bb46462),
	.w3(32'h3b3d0d21),
	.w4(32'h3ae8ae2f),
	.w5(32'hbbd848cb),
	.w6(32'h3bc1b6ce),
	.w7(32'h3ab8926b),
	.w8(32'hbb85a12d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdffa00),
	.w1(32'hba054596),
	.w2(32'h3b92c6a8),
	.w3(32'hb9aaefe0),
	.w4(32'h3be932ec),
	.w5(32'h3ace7cdd),
	.w6(32'hba4f3cc6),
	.w7(32'h3be01fe7),
	.w8(32'h3b855201),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be79bd4),
	.w1(32'h3c52794b),
	.w2(32'h3b7efcdc),
	.w3(32'h3b45f548),
	.w4(32'h3bde5da1),
	.w5(32'h3ba3c849),
	.w6(32'h3c01335c),
	.w7(32'hbb9e7a02),
	.w8(32'h3bc936f5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cc9d9),
	.w1(32'hbb8471aa),
	.w2(32'h3ba06dde),
	.w3(32'hbb4e0bc8),
	.w4(32'h3b85c421),
	.w5(32'hba99462e),
	.w6(32'hbc3d8840),
	.w7(32'h3aad9fe5),
	.w8(32'h3a4777cc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b9de),
	.w1(32'hbb021e3e),
	.w2(32'hbb5e4505),
	.w3(32'hbb8aab34),
	.w4(32'h3b9883ad),
	.w5(32'hbb0c3b4f),
	.w6(32'hb96bd8f8),
	.w7(32'hba03c716),
	.w8(32'hbb404f83),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70228b),
	.w1(32'h3bafa3b8),
	.w2(32'h3b26a0d3),
	.w3(32'hbafaec11),
	.w4(32'h3b2fe42f),
	.w5(32'h3b8f603c),
	.w6(32'hbb805f1d),
	.w7(32'hbb23e604),
	.w8(32'hbacdb582),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3156c7),
	.w1(32'hbb901120),
	.w2(32'hbb37b340),
	.w3(32'h3bd3b37f),
	.w4(32'h3b0ac0d9),
	.w5(32'hbc02fbfe),
	.w6(32'hbb84f3d6),
	.w7(32'h3a527b23),
	.w8(32'hbbac9207),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29073),
	.w1(32'hbaf5f67e),
	.w2(32'hbc0611a3),
	.w3(32'hbb6d8db3),
	.w4(32'hbb7f1294),
	.w5(32'hbc9a18a2),
	.w6(32'h3b84ada6),
	.w7(32'hbb9118bb),
	.w8(32'hbcd81c8e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc726f72),
	.w1(32'hbbb050ef),
	.w2(32'hbbf65b1d),
	.w3(32'hbbd5426b),
	.w4(32'hbbca7af9),
	.w5(32'hba77776b),
	.w6(32'h3ac9b1dd),
	.w7(32'hbc7feb5f),
	.w8(32'h3b12c95f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2b1b),
	.w1(32'hbaf38bfa),
	.w2(32'hbaf77c1e),
	.w3(32'hbabbcf88),
	.w4(32'hbb07d9c4),
	.w5(32'h3be0a2bd),
	.w6(32'hbb255b0f),
	.w7(32'hbb2fa8fc),
	.w8(32'hbabe7803),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0978),
	.w1(32'h3b0d47db),
	.w2(32'h3b2fb2b5),
	.w3(32'h3bc49108),
	.w4(32'h398fd143),
	.w5(32'hbbc6a2cf),
	.w6(32'hb9b64629),
	.w7(32'h3a9a19f1),
	.w8(32'hbb8b41c9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4800cf),
	.w1(32'hbafc7bd7),
	.w2(32'hbad118d6),
	.w3(32'hba60352a),
	.w4(32'hba26dab7),
	.w5(32'h38da57d8),
	.w6(32'hba93240e),
	.w7(32'h3b19a690),
	.w8(32'h3b72cd74),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2330),
	.w1(32'hbb2a7c14),
	.w2(32'h3a1fb2c4),
	.w3(32'hbaf0e243),
	.w4(32'hbad89b57),
	.w5(32'hbb032a74),
	.w6(32'hba7ff396),
	.w7(32'hbb23b630),
	.w8(32'h3a86c2be),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45bd02),
	.w1(32'h3b23a18f),
	.w2(32'hbb1f4b0c),
	.w3(32'h3bb307e4),
	.w4(32'hbae3bacb),
	.w5(32'hbb8f9a9b),
	.w6(32'h3b9c7837),
	.w7(32'hbb4665dc),
	.w8(32'hbb71f969),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9450be),
	.w1(32'hbb643bf1),
	.w2(32'hbb9217fc),
	.w3(32'hbb80d0b6),
	.w4(32'hbb3aa841),
	.w5(32'h3bc331d4),
	.w6(32'hbb100744),
	.w7(32'hbb6e95af),
	.w8(32'h3ba8ccbb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25b97),
	.w1(32'h3a259ceb),
	.w2(32'h3a99a561),
	.w3(32'h3b26100a),
	.w4(32'hb982dbf3),
	.w5(32'h3b1ca7dd),
	.w6(32'h3a8ba288),
	.w7(32'h39e63644),
	.w8(32'hbae24f9a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4b3c),
	.w1(32'h3bd2b9f3),
	.w2(32'h3bfab9bf),
	.w3(32'h3ae394ca),
	.w4(32'h3b256ca6),
	.w5(32'h3b3795c9),
	.w6(32'h3a2a5d1f),
	.w7(32'h3c38b834),
	.w8(32'h3bbd5878),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7381ab),
	.w1(32'hba32579a),
	.w2(32'hbb8c2bf4),
	.w3(32'hbae6513b),
	.w4(32'hba481da5),
	.w5(32'h39dae400),
	.w6(32'h3b1c6db1),
	.w7(32'h3b0e0d4c),
	.w8(32'h3b0928b0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c76d7),
	.w1(32'hbb85f1bb),
	.w2(32'hbae80efd),
	.w3(32'hb96798ea),
	.w4(32'h3a7fb6df),
	.w5(32'hbac3cf29),
	.w6(32'hbac2b450),
	.w7(32'h3b24671d),
	.w8(32'hbb03402c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb035dc3),
	.w1(32'hbabba71f),
	.w2(32'h39ebdf19),
	.w3(32'h39f725a8),
	.w4(32'hbb83c525),
	.w5(32'hbbb27e0e),
	.w6(32'hbb03dfc9),
	.w7(32'hbae041da),
	.w8(32'hbc21a3f0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe96336),
	.w1(32'h3b74908b),
	.w2(32'h3c8ad582),
	.w3(32'hbc04c72a),
	.w4(32'h3a91cae6),
	.w5(32'hbbb8e617),
	.w6(32'hbbfe59ca),
	.w7(32'h3c0220b4),
	.w8(32'hbb906ffa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b67b),
	.w1(32'h3b0d746a),
	.w2(32'hbb823d3d),
	.w3(32'hbb984429),
	.w4(32'hbb240635),
	.w5(32'hbb4d7e70),
	.w6(32'h3ad134f7),
	.w7(32'hbb437ac1),
	.w8(32'hbb86ee92),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4859a6),
	.w1(32'hbb9b9499),
	.w2(32'h3947b75a),
	.w3(32'hbbb4301c),
	.w4(32'hbb57eff6),
	.w5(32'hbc1800e6),
	.w6(32'hbbcb933c),
	.w7(32'hbb3f1e50),
	.w8(32'hba4fd74f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf86bc2),
	.w1(32'h3bb610ed),
	.w2(32'h399c6099),
	.w3(32'hbbc99561),
	.w4(32'h3bba9de0),
	.w5(32'hbc942421),
	.w6(32'hba9d078b),
	.w7(32'hba4adc13),
	.w8(32'hbce085ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85e7b5),
	.w1(32'hbbb82679),
	.w2(32'hbc84e441),
	.w3(32'hbbe04483),
	.w4(32'hbc7d6f9f),
	.w5(32'hbbb2b9c7),
	.w6(32'h3bc784ed),
	.w7(32'hbcd94844),
	.w8(32'hbbe857ac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01efa7),
	.w1(32'hbb034cd4),
	.w2(32'hbba898b3),
	.w3(32'hbb7970b2),
	.w4(32'hbb89985f),
	.w5(32'h3b99d77e),
	.w6(32'hbb890481),
	.w7(32'hbac5d4b2),
	.w8(32'h3beae23d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8213d0),
	.w1(32'h391be794),
	.w2(32'hbaf160a5),
	.w3(32'hbb23da91),
	.w4(32'h3a5ccaea),
	.w5(32'h3bb28ed1),
	.w6(32'h3a5b922a),
	.w7(32'h3b41fb3f),
	.w8(32'h3c8e2d7b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0439db),
	.w1(32'hbc1073c0),
	.w2(32'hbb254664),
	.w3(32'h3b0c68f1),
	.w4(32'h3ae1ee3e),
	.w5(32'h3ae5b9b6),
	.w6(32'h3ade6b05),
	.w7(32'h38ce1172),
	.w8(32'hb94988b6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ef487),
	.w1(32'h3a7843d5),
	.w2(32'h3b9a73cf),
	.w3(32'h3b23008a),
	.w4(32'h3be197ef),
	.w5(32'hbb8f9cee),
	.w6(32'h3aff8fcb),
	.w7(32'h3bfb95c0),
	.w8(32'hbac8fe67),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf025a7),
	.w1(32'h3b203c90),
	.w2(32'hbb89403e),
	.w3(32'hba17b555),
	.w4(32'h3a4410a1),
	.w5(32'h3bb316ac),
	.w6(32'h3b840f38),
	.w7(32'h3aee79fd),
	.w8(32'h3c09401b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeaeaa),
	.w1(32'h3c02a391),
	.w2(32'h3bd4d3ea),
	.w3(32'h3b3767b7),
	.w4(32'h3ae3f7c8),
	.w5(32'hbb0b2bc5),
	.w6(32'h3bc895b4),
	.w7(32'h3bd1ce38),
	.w8(32'hbbb6490e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac466e0),
	.w1(32'h3b2d1401),
	.w2(32'h3b064f6e),
	.w3(32'h3a4b9244),
	.w4(32'h3b908dd1),
	.w5(32'hbb8369f2),
	.w6(32'hbb49ce73),
	.w7(32'hb9f19248),
	.w8(32'hbb76be62),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e03e),
	.w1(32'h3b554fb2),
	.w2(32'hba29e979),
	.w3(32'hbad9aadc),
	.w4(32'hbbb45c98),
	.w5(32'h3bd38c90),
	.w6(32'h3bbe94fe),
	.w7(32'hbb254434),
	.w8(32'hbbaeceaf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a3fd8),
	.w1(32'hba8fbbf7),
	.w2(32'h3bfe7917),
	.w3(32'hbb14b19e),
	.w4(32'hbbb15428),
	.w5(32'hba794a94),
	.w6(32'hbb1593fb),
	.w7(32'hbb0644dc),
	.w8(32'hbaf073f1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67718a),
	.w1(32'h3c3abd35),
	.w2(32'h3bec0dc5),
	.w3(32'hbb81f7ff),
	.w4(32'hbbb10fd7),
	.w5(32'h396f8a46),
	.w6(32'hbb477c89),
	.w7(32'h3b84fbd4),
	.w8(32'hbb31bcd8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83bbff),
	.w1(32'hbb7c6f0b),
	.w2(32'hbb42a048),
	.w3(32'hba5f22ef),
	.w4(32'h3b359f4f),
	.w5(32'hbc4d5b2f),
	.w6(32'hbace46ff),
	.w7(32'h3b52b61e),
	.w8(32'hbc014518),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc497c0b),
	.w1(32'hbbffd29f),
	.w2(32'hbae4f109),
	.w3(32'hbc59ba18),
	.w4(32'hbb568d55),
	.w5(32'h3adcfb4c),
	.w6(32'hbbd1b86d),
	.w7(32'hbb4f21cb),
	.w8(32'h39b16395),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8056d),
	.w1(32'h3b3f4ffe),
	.w2(32'h3aeb525f),
	.w3(32'h3bc1d921),
	.w4(32'h3b208685),
	.w5(32'hb98c31b1),
	.w6(32'h3857efa0),
	.w7(32'h3bacf142),
	.w8(32'hba61dd59),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a807077),
	.w1(32'hba719d4b),
	.w2(32'hbb4db6c2),
	.w3(32'hba6c99c9),
	.w4(32'h393260f2),
	.w5(32'hbb938773),
	.w6(32'hbb4ef4b9),
	.w7(32'hbb7fcf50),
	.w8(32'hbb5bc692),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57484c),
	.w1(32'h3beb5935),
	.w2(32'hbb6d9680),
	.w3(32'h3a7b9c18),
	.w4(32'hbb348918),
	.w5(32'hbab70910),
	.w6(32'h3b7ac2f0),
	.w7(32'hbbbd25e7),
	.w8(32'hba62e4fb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38591211),
	.w1(32'hbbc714bd),
	.w2(32'hbab3e7b0),
	.w3(32'hbac8fa4e),
	.w4(32'hbba56316),
	.w5(32'hbb81c21a),
	.w6(32'h3acb84f6),
	.w7(32'h3b6ed01d),
	.w8(32'h3a0e330c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2363),
	.w1(32'h392cb900),
	.w2(32'h3abf2fc5),
	.w3(32'h3a54bea4),
	.w4(32'h3b3f4290),
	.w5(32'hbc1d6bf4),
	.w6(32'h3b8cdc8c),
	.w7(32'h3c038ddd),
	.w8(32'hbc67ef3e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddaeea),
	.w1(32'h3c003326),
	.w2(32'h3b835e14),
	.w3(32'hbb280a1e),
	.w4(32'hbaa5d93c),
	.w5(32'hbbceef5d),
	.w6(32'hbb87fee1),
	.w7(32'hba878327),
	.w8(32'hbbb6c80c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc03b4),
	.w1(32'hbb80a327),
	.w2(32'h3af420f5),
	.w3(32'h3a472501),
	.w4(32'hb8f03298),
	.w5(32'hb961279c),
	.w6(32'hba972c58),
	.w7(32'h3b80c3d0),
	.w8(32'hbc19d834),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c5cb),
	.w1(32'h3b73c3cd),
	.w2(32'h397d8153),
	.w3(32'h3b6ebd14),
	.w4(32'h38e645a9),
	.w5(32'hbb2435f3),
	.w6(32'h3bcecc57),
	.w7(32'hbb825a7d),
	.w8(32'hbab07a0e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b903),
	.w1(32'hbb632d98),
	.w2(32'hbba9a980),
	.w3(32'hbb6f1a78),
	.w4(32'hbbba3807),
	.w5(32'hbba8deb9),
	.w6(32'hbb97ada2),
	.w7(32'hbbdfa739),
	.w8(32'hbbbb0e98),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca1dc6),
	.w1(32'h3a43b1c0),
	.w2(32'hbb914ab7),
	.w3(32'hbb635e65),
	.w4(32'hbb194ebf),
	.w5(32'hbc177a3a),
	.w6(32'h38511b69),
	.w7(32'hbadc9f6c),
	.w8(32'hbba2ccb7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4603),
	.w1(32'h3ba283d2),
	.w2(32'hbacd3924),
	.w3(32'hbac1ab5a),
	.w4(32'h3a9e810a),
	.w5(32'hbaa6ca29),
	.w6(32'hbac09c4e),
	.w7(32'hba45ec27),
	.w8(32'hbb7067c3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85111),
	.w1(32'hbaa23b64),
	.w2(32'hba8d347a),
	.w3(32'hbbbcc969),
	.w4(32'hbb1d0105),
	.w5(32'hba02c4ef),
	.w6(32'hbaec0940),
	.w7(32'hb97eea36),
	.w8(32'hbb31974d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f1700),
	.w1(32'hba123a3f),
	.w2(32'h3a8c738b),
	.w3(32'h399e77b1),
	.w4(32'h3b070e4e),
	.w5(32'hbbda562d),
	.w6(32'hba8f9447),
	.w7(32'h3bb6a345),
	.w8(32'hbc1e7985),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ec713),
	.w1(32'hba21022b),
	.w2(32'hbc146ae5),
	.w3(32'hbaa88e21),
	.w4(32'h39838c0f),
	.w5(32'h3b36946e),
	.w6(32'h3a6f78d5),
	.w7(32'hbb8fbb68),
	.w8(32'h3ba0ddbf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c6714),
	.w1(32'hbbc77df5),
	.w2(32'hbc017339),
	.w3(32'hbb2dabd7),
	.w4(32'hbb746be3),
	.w5(32'h3a0d8dcf),
	.w6(32'hbb109c43),
	.w7(32'hbbd66ed6),
	.w8(32'hbb55a5a4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b97ab),
	.w1(32'h3aa26bee),
	.w2(32'hbb0cb970),
	.w3(32'h3b862ffe),
	.w4(32'h3b8274b6),
	.w5(32'hbbf27287),
	.w6(32'h3af6060b),
	.w7(32'h3a7e6e87),
	.w8(32'hbbf7528b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9353bc),
	.w1(32'h3a1c5493),
	.w2(32'h3b18ebf6),
	.w3(32'hbb90a80c),
	.w4(32'hba72a638),
	.w5(32'h3bc52487),
	.w6(32'hbb9dd563),
	.w7(32'h3aa1eee1),
	.w8(32'h3bd9f037),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4030d),
	.w1(32'h3b58e249),
	.w2(32'h3acaf48f),
	.w3(32'h3b2d4f2a),
	.w4(32'h3b9dca73),
	.w5(32'h3a40f7e8),
	.w6(32'h3af66871),
	.w7(32'h3baf405c),
	.w8(32'hbab5ec3f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eadd5),
	.w1(32'h3a384c6e),
	.w2(32'h3be32075),
	.w3(32'hbb03280d),
	.w4(32'hbb8aef40),
	.w5(32'hba10931c),
	.w6(32'hbaf480b9),
	.w7(32'h3a7acbf5),
	.w8(32'h3bca8620),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b75ff),
	.w1(32'h3b2d928c),
	.w2(32'h3af23b6f),
	.w3(32'hbaf289b8),
	.w4(32'h3b0d3724),
	.w5(32'hbc3c73f5),
	.w6(32'h3a49b2e8),
	.w7(32'h3a429c7b),
	.w8(32'hbc96795d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22c22c),
	.w1(32'h3c02a386),
	.w2(32'h3c3dfa62),
	.w3(32'hbb5541c3),
	.w4(32'h3b810525),
	.w5(32'h39fd9c7d),
	.w6(32'h3b9c0d33),
	.w7(32'h3c2cef4c),
	.w8(32'h39e2963c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984c34),
	.w1(32'hb9b96781),
	.w2(32'h3af6ce59),
	.w3(32'h3b936f24),
	.w4(32'h3bb3f3bb),
	.w5(32'hbb80c3b0),
	.w6(32'hbb4d8ddc),
	.w7(32'h3c0897b1),
	.w8(32'hbbb76724),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc63d3),
	.w1(32'hbb2d363c),
	.w2(32'hbbbeb4bb),
	.w3(32'hbc0ecf3d),
	.w4(32'hbb913155),
	.w5(32'hbbdf8cad),
	.w6(32'hbbd8a9ed),
	.w7(32'hbbcf2995),
	.w8(32'hbb8f89d4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87b774),
	.w1(32'hbbcd0fd7),
	.w2(32'hbb369475),
	.w3(32'hbc0b02b9),
	.w4(32'hbba39139),
	.w5(32'hbadaf200),
	.w6(32'hbbdeaf79),
	.w7(32'hba31e7fa),
	.w8(32'h3aac913b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed6aca),
	.w1(32'hbaa2d21a),
	.w2(32'hbb2ec036),
	.w3(32'hbb060dc1),
	.w4(32'hbb01ed9b),
	.w5(32'hbb008ba4),
	.w6(32'h3a47f3ba),
	.w7(32'hba8ad62e),
	.w8(32'hbb4fbe43),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69e573),
	.w1(32'h3c2eef07),
	.w2(32'h3bf184a2),
	.w3(32'hb9912cf1),
	.w4(32'h3bad1667),
	.w5(32'h3b8fa002),
	.w6(32'h3b0293b1),
	.w7(32'h3b838d2b),
	.w8(32'h3b09f88c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de3f7),
	.w1(32'h3b1a0e7c),
	.w2(32'h3ae729af),
	.w3(32'h3b91031a),
	.w4(32'h3a3df438),
	.w5(32'hbb8343b2),
	.w6(32'hba079e60),
	.w7(32'hbb6bb877),
	.w8(32'hbb4f7032),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb179945),
	.w1(32'hbb91e471),
	.w2(32'hbbc4c0be),
	.w3(32'hbb482fcf),
	.w4(32'hbba7f84a),
	.w5(32'hbca93558),
	.w6(32'hba338001),
	.w7(32'hbbbd27ba),
	.w8(32'hbcb81f2b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b64d),
	.w1(32'hbba3dc82),
	.w2(32'hbc5b0232),
	.w3(32'hbc2d42be),
	.w4(32'hbc58e542),
	.w5(32'h3ba41f3b),
	.w6(32'hbb4dc710),
	.w7(32'hbc6ea708),
	.w8(32'h3bcac96d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cb2b3),
	.w1(32'hbaafba6f),
	.w2(32'h3aa2cd0b),
	.w3(32'hb940d20f),
	.w4(32'h3b48fef6),
	.w5(32'h3b52ed4a),
	.w6(32'h3b2829da),
	.w7(32'h3b09d02b),
	.w8(32'hba205640),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6b4d),
	.w1(32'hbc019236),
	.w2(32'hbb91f8b9),
	.w3(32'hbad4c951),
	.w4(32'hb87c5d73),
	.w5(32'hbb53a9b3),
	.w6(32'hbb9f26af),
	.w7(32'hbbaa4ece),
	.w8(32'hba9cf867),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5c4d9),
	.w1(32'h39f5538e),
	.w2(32'hba8a88a4),
	.w3(32'h3ad054b4),
	.w4(32'hb89ea77c),
	.w5(32'hbb31ac6c),
	.w6(32'h3b2c30fb),
	.w7(32'h3aeb6539),
	.w8(32'hbc1e1998),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2314ad),
	.w1(32'hbc34995d),
	.w2(32'hbbfeb970),
	.w3(32'hbb5edbda),
	.w4(32'hbabd0303),
	.w5(32'hbb1c7cf6),
	.w6(32'hbc26dd73),
	.w7(32'hbbeaf29f),
	.w8(32'hbb0dbcd5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb439bd3),
	.w1(32'hbc067477),
	.w2(32'hbba1d5b7),
	.w3(32'hbbfcc58a),
	.w4(32'hbb87f5cd),
	.w5(32'hbc472992),
	.w6(32'hbbf8c895),
	.w7(32'hbba9d75d),
	.w8(32'hbc364ff5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c29e4),
	.w1(32'hbc3907a5),
	.w2(32'hbc3a60b9),
	.w3(32'hbc23a7a8),
	.w4(32'hbc2aab96),
	.w5(32'hbb9d5e24),
	.w6(32'hbc1af708),
	.w7(32'hbc565237),
	.w8(32'hbbc89b3c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478330),
	.w1(32'hbbf6eb5c),
	.w2(32'hbbdc9637),
	.w3(32'hbb8904e0),
	.w4(32'hbab1f2eb),
	.w5(32'hbc8b93a9),
	.w6(32'hbbe92c2a),
	.w7(32'hbc096eea),
	.w8(32'hbc896d3c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc826df3),
	.w1(32'hbc7241e6),
	.w2(32'hbc625d81),
	.w3(32'hbc8de90c),
	.w4(32'hbc8d751b),
	.w5(32'h3b356bda),
	.w6(32'hbc78ec95),
	.w7(32'hbc620937),
	.w8(32'h3a0170ae),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd60fb0),
	.w1(32'h3b7e6f72),
	.w2(32'h3c127018),
	.w3(32'hbbf11b5c),
	.w4(32'h3b79ed34),
	.w5(32'hbbf7ad5c),
	.w6(32'hbbb6fbca),
	.w7(32'h3b9286eb),
	.w8(32'hbba549b9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba76f0f),
	.w1(32'hbc231eee),
	.w2(32'hbbe53779),
	.w3(32'hbc1ddf42),
	.w4(32'hbbd439e2),
	.w5(32'h3b92194e),
	.w6(32'hbc0dfef4),
	.w7(32'hbbde74f5),
	.w8(32'h3b6936e4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b557831),
	.w1(32'hbbc71e50),
	.w2(32'hbb0bf24a),
	.w3(32'hbb86a495),
	.w4(32'hb82956cb),
	.w5(32'hbb8c1555),
	.w6(32'hbb76c488),
	.w7(32'hbb1478bf),
	.w8(32'hbb0575ad),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf5f8),
	.w1(32'hba26745c),
	.w2(32'h3a8836f3),
	.w3(32'hbac15985),
	.w4(32'h3974c57b),
	.w5(32'hbb0f2612),
	.w6(32'h3aa932c2),
	.w7(32'h3ab9551b),
	.w8(32'hbc16a135),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc599c35),
	.w1(32'hbc5a663f),
	.w2(32'hbc0f81c2),
	.w3(32'hbc03e67c),
	.w4(32'hbbf2868a),
	.w5(32'h3aed5175),
	.w6(32'hbc228285),
	.w7(32'hbc0bad07),
	.w8(32'hb9925beb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae04dad),
	.w1(32'hbb064ee8),
	.w2(32'hbbd89c41),
	.w3(32'h3afcc4fa),
	.w4(32'hba25c81c),
	.w5(32'hbb22a609),
	.w6(32'h3abe446b),
	.w7(32'hbb1f9aa8),
	.w8(32'hbb7d9d8d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ecacb),
	.w1(32'h3b81ee3e),
	.w2(32'h3b803641),
	.w3(32'h3915292d),
	.w4(32'h3a794130),
	.w5(32'h3b7baeb9),
	.w6(32'hb8a40b00),
	.w7(32'h39be443f),
	.w8(32'h3b41f792),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb086b45),
	.w1(32'hbad0e46e),
	.w2(32'hbab4e45f),
	.w3(32'h3b9c2672),
	.w4(32'h3ab8f6ac),
	.w5(32'hbbcbedf0),
	.w6(32'h3b1c8778),
	.w7(32'h3b8a020c),
	.w8(32'hbb9a3264),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b678a),
	.w1(32'h39a0b111),
	.w2(32'hbb25d9af),
	.w3(32'hbbed7e12),
	.w4(32'hbbc19638),
	.w5(32'h3baa8d1c),
	.w6(32'hba8f419e),
	.w7(32'hbbb0d085),
	.w8(32'h3a37de57),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089583),
	.w1(32'hbaee1568),
	.w2(32'hbb9baf90),
	.w3(32'h3bd69cca),
	.w4(32'h3b9a096e),
	.w5(32'h3c1058da),
	.w6(32'h3b0cbe23),
	.w7(32'h39ae1363),
	.w8(32'h3b94a58a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ace5),
	.w1(32'h3bafb274),
	.w2(32'h3baad8cd),
	.w3(32'h3c11635b),
	.w4(32'h3bd7903a),
	.w5(32'hbb868d61),
	.w6(32'h3b8607bc),
	.w7(32'h3b7379c1),
	.w8(32'hbb4d6bf9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e99dfa),
	.w1(32'hbc01479c),
	.w2(32'hbb61baa0),
	.w3(32'hbbb92e68),
	.w4(32'h3bcf0f34),
	.w5(32'hbb090642),
	.w6(32'hbb82e7e4),
	.w7(32'h3ba8952e),
	.w8(32'hbbb380db),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f66f),
	.w1(32'hbc4d8d44),
	.w2(32'hbb8aa103),
	.w3(32'hbc3cbc84),
	.w4(32'hbb4cbaf9),
	.w5(32'h3cd3c004),
	.w6(32'hbc79adc3),
	.w7(32'hbc170bea),
	.w8(32'h3d0320fa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe02cd),
	.w1(32'h3cef3ffd),
	.w2(32'h3caef50d),
	.w3(32'h3cf992c5),
	.w4(32'h3cba4d89),
	.w5(32'h3a97d8b4),
	.w6(32'h3d2c3b80),
	.w7(32'h3cd5999d),
	.w8(32'h399d1ef0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39f36),
	.w1(32'h3b2f25c2),
	.w2(32'hbb494ea9),
	.w3(32'h3b137184),
	.w4(32'hb9e919e8),
	.w5(32'h3b9c784a),
	.w6(32'h3b782488),
	.w7(32'h39dd304f),
	.w8(32'h3b99590f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894bec),
	.w1(32'h3c2e6f53),
	.w2(32'h3afddac9),
	.w3(32'h3c176391),
	.w4(32'h3bade528),
	.w5(32'hbb85df76),
	.w6(32'h3c285b05),
	.w7(32'h3a0f36e6),
	.w8(32'hbbb49211),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c72ac3),
	.w1(32'hbba5e33f),
	.w2(32'hbadfe718),
	.w3(32'hbb8600ae),
	.w4(32'hb67eb032),
	.w5(32'h3a16ee23),
	.w6(32'hbba077a2),
	.w7(32'h39049bfa),
	.w8(32'h3ab4545c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986e452),
	.w1(32'h3a9ad160),
	.w2(32'h3ac49e24),
	.w3(32'hbab478c2),
	.w4(32'h3ad5e8c5),
	.w5(32'hba8d422c),
	.w6(32'hbb03e1cc),
	.w7(32'h3a4985e7),
	.w8(32'hbb53c652),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb014c6),
	.w1(32'hbbd7d862),
	.w2(32'h3917a201),
	.w3(32'hbb1b7947),
	.w4(32'h3a671876),
	.w5(32'hbaa9492c),
	.w6(32'hb98ad9fb),
	.w7(32'h3bb8f3a0),
	.w8(32'hbad63c57),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e1fda),
	.w1(32'hbaa126a9),
	.w2(32'hbaddf4ac),
	.w3(32'hbb08a145),
	.w4(32'hbb6975db),
	.w5(32'hbc07a9da),
	.w6(32'hbba797ae),
	.w7(32'hbba6624a),
	.w8(32'hbb25fe68),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0e4d),
	.w1(32'hbc18137b),
	.w2(32'hbbfcf2ec),
	.w3(32'hbc1ac27a),
	.w4(32'hbb36aa0c),
	.w5(32'hbbabcde2),
	.w6(32'hbb95af30),
	.w7(32'hbb1fae26),
	.w8(32'hbbae5fe8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3f2b),
	.w1(32'h3a28dc96),
	.w2(32'hbbb42a2b),
	.w3(32'hba989669),
	.w4(32'hbc1320f1),
	.w5(32'hbb468625),
	.w6(32'h3a202992),
	.w7(32'hbbeea8c1),
	.w8(32'hb98f9c1d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7df5),
	.w1(32'h3ba499a7),
	.w2(32'h3c2f2900),
	.w3(32'h3abaf983),
	.w4(32'h3bf7efa5),
	.w5(32'hbc39d285),
	.w6(32'h3c12290b),
	.w7(32'h3c391f21),
	.w8(32'hbc0247b6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987c40),
	.w1(32'hbc2eda4d),
	.w2(32'hbc228dc3),
	.w3(32'hbc56c0cb),
	.w4(32'hbbe8ed7b),
	.w5(32'hbbd38a67),
	.w6(32'hbc64ca3c),
	.w7(32'hbc15e484),
	.w8(32'hbba54d66),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6088f8),
	.w1(32'hbc62ebdc),
	.w2(32'hbc5788bc),
	.w3(32'hbc00375a),
	.w4(32'hbbe4d74b),
	.w5(32'hbba7bb2e),
	.w6(32'hbc087708),
	.w7(32'hbbfa16a8),
	.w8(32'hbbe9a060),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38c85),
	.w1(32'hbbfe6f04),
	.w2(32'hbc0b1bc9),
	.w3(32'hbba0a885),
	.w4(32'hbb6055a2),
	.w5(32'hbb9f4978),
	.w6(32'hbbc99c2f),
	.w7(32'hbbac9119),
	.w8(32'hbb2d7dfb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bc43c),
	.w1(32'h3ae3b7ec),
	.w2(32'hbb616db9),
	.w3(32'hbadfb87f),
	.w4(32'hbb8f86aa),
	.w5(32'hbb094f24),
	.w6(32'hba269f4f),
	.w7(32'hbbb5ed6f),
	.w8(32'hbb039835),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cd892),
	.w1(32'hbabce868),
	.w2(32'hbaab71a6),
	.w3(32'h3aa2ad36),
	.w4(32'h3b06859f),
	.w5(32'hba6ad7dd),
	.w6(32'h3b36a2cd),
	.w7(32'h3aa9e59f),
	.w8(32'h39ec3f9e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2b244),
	.w1(32'h3b58855d),
	.w2(32'h3a17337d),
	.w3(32'h3bb510fb),
	.w4(32'h3bb119ad),
	.w5(32'h3c0224f3),
	.w6(32'h3c03a25e),
	.w7(32'h3bb54ce5),
	.w8(32'h3b916881),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab105ff),
	.w1(32'h3b9634cf),
	.w2(32'h3b5019a6),
	.w3(32'h3bf95a51),
	.w4(32'h3ba5f86a),
	.w5(32'hba114797),
	.w6(32'h3be6c5ba),
	.w7(32'h3b98b029),
	.w8(32'hbb1e687f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2de3c2),
	.w1(32'h3b7eb422),
	.w2(32'h3ba60e69),
	.w3(32'h3b634929),
	.w4(32'h3b9f1b95),
	.w5(32'hbbdf41bd),
	.w6(32'h3b465783),
	.w7(32'h3b8942a4),
	.w8(32'hbbc0ecbb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf795c),
	.w1(32'hbbcf3052),
	.w2(32'hbb9f80a3),
	.w3(32'hbb94808d),
	.w4(32'hbac493b3),
	.w5(32'hbbaf003c),
	.w6(32'hbb2af531),
	.w7(32'hbb56e5e1),
	.w8(32'hbbbeed4f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe91ba5),
	.w1(32'hbb792f70),
	.w2(32'hbb60af35),
	.w3(32'hbaf29d55),
	.w4(32'hba2e9740),
	.w5(32'hbb76a2ff),
	.w6(32'hba2b69de),
	.w7(32'hba9be202),
	.w8(32'hbac2d8f0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d82a),
	.w1(32'hbc43c2e3),
	.w2(32'hbc601307),
	.w3(32'hbbee694a),
	.w4(32'hbbf3753c),
	.w5(32'hbc03e587),
	.w6(32'hbbbdcd73),
	.w7(32'hbbc1f12b),
	.w8(32'hbc0d9d63),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb040f6),
	.w1(32'hbac523fc),
	.w2(32'hbbd083e5),
	.w3(32'hbbf16f0a),
	.w4(32'hbc4fe240),
	.w5(32'h3b04dd5d),
	.w6(32'hbbc6e8f1),
	.w7(32'hbc0e6ff2),
	.w8(32'hb980ef56),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c4d6e),
	.w1(32'hbb9aa4b8),
	.w2(32'hbb9302de),
	.w3(32'hbb6709ef),
	.w4(32'hbb08eac5),
	.w5(32'hbbbaa64f),
	.w6(32'hbba26ee9),
	.w7(32'hbb877a7c),
	.w8(32'hbc016c6e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3978a6),
	.w1(32'hbc0cba54),
	.w2(32'hbc07699f),
	.w3(32'hbbcc5872),
	.w4(32'hbc0e8cd3),
	.w5(32'hbc24cb78),
	.w6(32'hbb9284e7),
	.w7(32'hbbc61b20),
	.w8(32'hbc4bd258),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6469),
	.w1(32'hbbf01f32),
	.w2(32'hbbf45f93),
	.w3(32'hbbb88d4a),
	.w4(32'hbbb1e010),
	.w5(32'hbb889a47),
	.w6(32'hbbfde981),
	.w7(32'hbbf839f0),
	.w8(32'hbb65739e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7931db),
	.w1(32'hbbdfc599),
	.w2(32'hbbc1af10),
	.w3(32'hbb307874),
	.w4(32'hbb8dd7d5),
	.w5(32'hbbe96aa8),
	.w6(32'hbb85bd3c),
	.w7(32'hbb6a6a2e),
	.w8(32'hbc0d5b94),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00dd4),
	.w1(32'hbc0be0df),
	.w2(32'hbb87f1de),
	.w3(32'hbc15565d),
	.w4(32'hbba292fa),
	.w5(32'h3aae0418),
	.w6(32'hbc057887),
	.w7(32'hbbbee3ea),
	.w8(32'hbb62283e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee77a),
	.w1(32'hbbd93cf4),
	.w2(32'hbb21aa14),
	.w3(32'h3af2eca8),
	.w4(32'h3bb68c1d),
	.w5(32'hbb2684aa),
	.w6(32'hb8c9a6a3),
	.w7(32'hbb0e925a),
	.w8(32'h3aa95bca),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f11d),
	.w1(32'hb95347ca),
	.w2(32'h3a8de5d0),
	.w3(32'hbb61e60f),
	.w4(32'hbadf5b19),
	.w5(32'hbb874a10),
	.w6(32'hbb1e6172),
	.w7(32'hba502d13),
	.w8(32'hbbddf11e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc768d6),
	.w1(32'hbb16a9db),
	.w2(32'hbb0c6b39),
	.w3(32'h3b1e0a18),
	.w4(32'h395e3fe3),
	.w5(32'h3c0f655c),
	.w6(32'hb989a9bc),
	.w7(32'hbad6f2f8),
	.w8(32'h3bb24ba1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75f885),
	.w1(32'h3a949c4b),
	.w2(32'hba071f5b),
	.w3(32'h3bb009e3),
	.w4(32'h3b3b8a66),
	.w5(32'h3af92b11),
	.w6(32'h3a9d0b18),
	.w7(32'hb8f02091),
	.w8(32'h3b132151),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1ca7),
	.w1(32'hbaf77192),
	.w2(32'hbb3b0268),
	.w3(32'h3a1bc353),
	.w4(32'h3a0250a4),
	.w5(32'hbb53c612),
	.w6(32'h3a9c27d4),
	.w7(32'h3a18207d),
	.w8(32'hbc2542ad),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcff06),
	.w1(32'hba211cda),
	.w2(32'h3a0e094b),
	.w3(32'h3ae61ebf),
	.w4(32'h39b19f93),
	.w5(32'h3b832fcc),
	.w6(32'h3b5156af),
	.w7(32'hb98a84f2),
	.w8(32'h3b4ed54b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef6c1b),
	.w1(32'hbb257c05),
	.w2(32'hba03912e),
	.w3(32'h3b7cf062),
	.w4(32'h3bce7f3a),
	.w5(32'hbbc06372),
	.w6(32'hb9b11a1c),
	.w7(32'h3b23c389),
	.w8(32'hbbbbe054),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1af6d0),
	.w1(32'hbc0c3603),
	.w2(32'hbc17b67e),
	.w3(32'hbb75fcef),
	.w4(32'hbc0d4d9d),
	.w5(32'h3b19308c),
	.w6(32'hbb1ecebe),
	.w7(32'hbbdbdab8),
	.w8(32'hbaf2aa33),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb033278),
	.w1(32'hbbb6895f),
	.w2(32'hbbb527fe),
	.w3(32'hba351579),
	.w4(32'hbb77339f),
	.w5(32'hbb3af08f),
	.w6(32'hbbdfbe6b),
	.w7(32'hbbccab43),
	.w8(32'h3a819fc1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b1fab),
	.w1(32'h3b643376),
	.w2(32'h3bfc738f),
	.w3(32'h3aa0da26),
	.w4(32'h3b9ff77b),
	.w5(32'h3aafc0e7),
	.w6(32'h3bc897f4),
	.w7(32'h3bf9b8d0),
	.w8(32'h3b3b1ac5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad52934),
	.w1(32'h38264b00),
	.w2(32'hba7e796b),
	.w3(32'hba3a3979),
	.w4(32'h3ba7544a),
	.w5(32'hba7920de),
	.w6(32'hbae226b7),
	.w7(32'hbb1dbde1),
	.w8(32'hb9b062ba),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b239088),
	.w1(32'h3b048d1e),
	.w2(32'hbaa066b3),
	.w3(32'h3b284a9a),
	.w4(32'h3b3e48e0),
	.w5(32'hbb79aa6e),
	.w6(32'h3ae1be00),
	.w7(32'hbafa6b17),
	.w8(32'hbb6cc81f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84d973),
	.w1(32'hbc17e1a0),
	.w2(32'hbb671016),
	.w3(32'hbc31d06c),
	.w4(32'hbb9de884),
	.w5(32'hbb77982d),
	.w6(32'hbc28255f),
	.w7(32'hbbf656d5),
	.w8(32'hbbc3ab1a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3876da),
	.w1(32'hbc29dbe6),
	.w2(32'hbbf57c4c),
	.w3(32'hbc309466),
	.w4(32'hbbf6b2cf),
	.w5(32'hbbf3239b),
	.w6(32'hbbe19a08),
	.w7(32'hbba105aa),
	.w8(32'hbc1a3652),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23cea2),
	.w1(32'hbb9d6412),
	.w2(32'hbc4b6ad0),
	.w3(32'h394541ac),
	.w4(32'hbb4bf969),
	.w5(32'hbc312ea6),
	.w6(32'h3aab3570),
	.w7(32'hbc3a75e7),
	.w8(32'hbc507fc1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc381336),
	.w1(32'hbc4dec71),
	.w2(32'hbc2375d1),
	.w3(32'hbc5c7992),
	.w4(32'hbbf97603),
	.w5(32'hbb2b1fd0),
	.w6(32'hbc5145b6),
	.w7(32'hbc303b2b),
	.w8(32'hb94dd4a9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866f01),
	.w1(32'hbb9de24a),
	.w2(32'hbbbec451),
	.w3(32'hbb30ad84),
	.w4(32'hbb53fd68),
	.w5(32'hba7efd5a),
	.w6(32'hba75403c),
	.w7(32'hbb98037e),
	.w8(32'hbbd0b2fc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaf3c2),
	.w1(32'hbc073722),
	.w2(32'hbc0bae6a),
	.w3(32'hbb213940),
	.w4(32'hbb49bc3d),
	.w5(32'hbc16482a),
	.w6(32'hbbd5dd8d),
	.w7(32'hbbd95bbb),
	.w8(32'hbb3c110c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4ab0),
	.w1(32'hbbbe3de1),
	.w2(32'hbba87495),
	.w3(32'hbc1045c9),
	.w4(32'hbbca1d04),
	.w5(32'hbc009817),
	.w6(32'hbad94695),
	.w7(32'hbaeac4e2),
	.w8(32'hbbfe1a55),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ca53),
	.w1(32'hbad24e6a),
	.w2(32'hbc172c44),
	.w3(32'h3a2ff10a),
	.w4(32'hbba6ea1a),
	.w5(32'h3a15e8de),
	.w6(32'h3a7b79cb),
	.w7(32'hbc048e19),
	.w8(32'h3afb49cf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f6173),
	.w1(32'h369a179a),
	.w2(32'h3b34c845),
	.w3(32'hbba91232),
	.w4(32'h3b437a56),
	.w5(32'h3c1ded02),
	.w6(32'hb99f486a),
	.w7(32'h3b8890ed),
	.w8(32'h3c31622a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7b600),
	.w1(32'hb9bb13ac),
	.w2(32'hbbe4fdfb),
	.w3(32'h3bad244b),
	.w4(32'h3aadb16e),
	.w5(32'h3b82e385),
	.w6(32'hba39d674),
	.w7(32'hbbdb46d0),
	.w8(32'h3bb590f8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b862bcb),
	.w1(32'h3b663ed5),
	.w2(32'h3af2bc76),
	.w3(32'hb9a3da14),
	.w4(32'h3996a3cb),
	.w5(32'hbc000640),
	.w6(32'h3ac6f2ae),
	.w7(32'hbaf814c7),
	.w8(32'hbb40904b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe98ebe),
	.w1(32'hbbe801c9),
	.w2(32'hbc1e6067),
	.w3(32'hbbabacc0),
	.w4(32'hbbfa62a6),
	.w5(32'hbb67e74b),
	.w6(32'h39ec62f8),
	.w7(32'hbb84f196),
	.w8(32'hbbc98eea),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63f7a9),
	.w1(32'hba73c554),
	.w2(32'hbaf5790e),
	.w3(32'hbaccf055),
	.w4(32'hba5085b7),
	.w5(32'hbbf65c04),
	.w6(32'hb9f4a9bf),
	.w7(32'hbb0cfbd0),
	.w8(32'hbc6ba6d1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bd377),
	.w1(32'hbca9679c),
	.w2(32'hbc6cbdcf),
	.w3(32'hbc82ad1c),
	.w4(32'hbc2643df),
	.w5(32'hbaac9a36),
	.w6(32'hbcc799a9),
	.w7(32'hbc8b2906),
	.w8(32'h3b1370ec),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d2846),
	.w1(32'h3bb0ae6a),
	.w2(32'hba489946),
	.w3(32'h3bf9b0eb),
	.w4(32'h3b68aca3),
	.w5(32'hbab3b587),
	.w6(32'h3c568738),
	.w7(32'h3b2817a7),
	.w8(32'h3b1104e9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af92b68),
	.w1(32'hbb373055),
	.w2(32'hb9224db0),
	.w3(32'hbb927de8),
	.w4(32'h3b0610fe),
	.w5(32'h3b8f9599),
	.w6(32'hbad35d05),
	.w7(32'h3b296c73),
	.w8(32'h3bbd24b7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7d325),
	.w1(32'hba717788),
	.w2(32'h3a972532),
	.w3(32'h3b87ee62),
	.w4(32'h3ba1fe28),
	.w5(32'h3bb593a0),
	.w6(32'h3b19064a),
	.w7(32'h3b1c4802),
	.w8(32'h3b836afd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e21e),
	.w1(32'h3b3b15f4),
	.w2(32'hb9912788),
	.w3(32'h3b300321),
	.w4(32'hba08ac38),
	.w5(32'hbc5ec8b5),
	.w6(32'h389f89f9),
	.w7(32'hba3ca86f),
	.w8(32'hbc56f49a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc546725),
	.w1(32'hbc1bef53),
	.w2(32'hbbfeef69),
	.w3(32'hbc4a8235),
	.w4(32'hbc4917bc),
	.w5(32'h3b2b7bbf),
	.w6(32'hbbd7870f),
	.w7(32'hbbedf640),
	.w8(32'h3a5687f2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2afef0),
	.w1(32'hbb638ec5),
	.w2(32'hbbe3554b),
	.w3(32'h3ab6076c),
	.w4(32'hbb76adae),
	.w5(32'h3b5967ec),
	.w6(32'hb99eecf9),
	.w7(32'hbb98f568),
	.w8(32'hb953a8ca),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dccc1),
	.w1(32'hbc17ef8c),
	.w2(32'hbafd2cc0),
	.w3(32'hbbc233fa),
	.w4(32'hbb872244),
	.w5(32'h3a6d7ab1),
	.w6(32'hbbf83993),
	.w7(32'hbb29dd7b),
	.w8(32'h3b6e490d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c156f82),
	.w1(32'h3b241f75),
	.w2(32'h3bd72dc5),
	.w3(32'hba83c533),
	.w4(32'h3bc97d75),
	.w5(32'h3a3d4940),
	.w6(32'h3b84f719),
	.w7(32'h3bd6904d),
	.w8(32'hb9abf0e6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec06e6),
	.w1(32'h3b40020a),
	.w2(32'h3b0818f7),
	.w3(32'h3b5f42f2),
	.w4(32'h37b35b33),
	.w5(32'hbb3bc44d),
	.w6(32'h3b65760a),
	.w7(32'h3a98a826),
	.w8(32'h3b0bb26d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61339c),
	.w1(32'hbb0a2af8),
	.w2(32'hbc3635a2),
	.w3(32'hbb343c8e),
	.w4(32'hbc209814),
	.w5(32'hb9d0d345),
	.w6(32'h3ad1004c),
	.w7(32'hbc508b4f),
	.w8(32'h3aeb1b3d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01512),
	.w1(32'h3b5a0585),
	.w2(32'h3b324bcc),
	.w3(32'hbb069ad4),
	.w4(32'hbb2f79fa),
	.w5(32'hbbb61451),
	.w6(32'h396e4d41),
	.w7(32'hba990842),
	.w8(32'hbbfd1485),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4eeda),
	.w1(32'hbc12c0fe),
	.w2(32'hbaee55ea),
	.w3(32'hbbdaf1b2),
	.w4(32'h3a8b84f9),
	.w5(32'h3b17c2a1),
	.w6(32'hbc1613bb),
	.w7(32'hbb8f6972),
	.w8(32'h3ac453fb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9401a7),
	.w1(32'h3ae9a689),
	.w2(32'h3b297a8e),
	.w3(32'hb89e17a0),
	.w4(32'hba07e152),
	.w5(32'hba0b928e),
	.w6(32'hbaaff12c),
	.w7(32'hbb15ca9a),
	.w8(32'hbb13e974),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9783),
	.w1(32'hbb9f553e),
	.w2(32'hbb58f310),
	.w3(32'hbb99c7eb),
	.w4(32'h38d15ca2),
	.w5(32'h39dc4d12),
	.w6(32'hbbcc5d65),
	.w7(32'hbbdad11a),
	.w8(32'hb8fb44ea),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37b2bf),
	.w1(32'hbaae02e0),
	.w2(32'hbb71787f),
	.w3(32'h3b19fbe1),
	.w4(32'hbb1aa772),
	.w5(32'h3c61b259),
	.w6(32'h3b53d262),
	.w7(32'hbaa70186),
	.w8(32'h3c2757e1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308d99),
	.w1(32'h3b968e4c),
	.w2(32'h3c4c6d31),
	.w3(32'h3b8be57a),
	.w4(32'h3c0b847f),
	.w5(32'hbaf32c01),
	.w6(32'hbaffe080),
	.w7(32'h3c2bdc7a),
	.w8(32'hbb657860),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae00c6),
	.w1(32'hbb853861),
	.w2(32'hba34a7c2),
	.w3(32'hbbdb27a8),
	.w4(32'hbb3ecb8d),
	.w5(32'hbbc18fd0),
	.w6(32'hbb8f5a13),
	.w7(32'hba914d79),
	.w8(32'hbb56f1e7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf33900),
	.w1(32'hbc52579d),
	.w2(32'hbc113df1),
	.w3(32'hbbe2a460),
	.w4(32'hbb630db6),
	.w5(32'hbbfed45a),
	.w6(32'hbba9d9f3),
	.w7(32'hbb87c87d),
	.w8(32'hbbebd2f5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71eb07),
	.w1(32'hbb8ac6c0),
	.w2(32'hbb84e597),
	.w3(32'hbc19700c),
	.w4(32'hbbf61a84),
	.w5(32'h3a867e4e),
	.w6(32'hbc19907b),
	.w7(32'hbc098131),
	.w8(32'h3b57c810),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2161b),
	.w1(32'h3aa22308),
	.w2(32'h3ad45971),
	.w3(32'h3755cc02),
	.w4(32'h3a50a585),
	.w5(32'hba937dd9),
	.w6(32'h3b313d60),
	.w7(32'h3a32297d),
	.w8(32'h3a82d06e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f41cb3),
	.w1(32'hbbb4010b),
	.w2(32'hbb88ab9b),
	.w3(32'hbb860218),
	.w4(32'hba240cf2),
	.w5(32'hbaf0dbef),
	.w6(32'hbb106d02),
	.w7(32'hbb773780),
	.w8(32'hbb3593b8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebe230),
	.w1(32'hbafa3841),
	.w2(32'h3aa745b2),
	.w3(32'hbb8fb9ad),
	.w4(32'hbb073915),
	.w5(32'hbb43cd87),
	.w6(32'hbbc073d7),
	.w7(32'hbae1b6b8),
	.w8(32'hbb5784be),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb836b),
	.w1(32'hbb7664ce),
	.w2(32'hbbc627b0),
	.w3(32'hbba82c54),
	.w4(32'hbb3ca84f),
	.w5(32'hba7a6326),
	.w6(32'hbb772a9c),
	.w7(32'hbb0ba8e5),
	.w8(32'hbb99f53e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f5755),
	.w1(32'hbb706f99),
	.w2(32'hbb3436bb),
	.w3(32'hbbf7c005),
	.w4(32'hbc250c23),
	.w5(32'hbaee07cd),
	.w6(32'hbc3e8695),
	.w7(32'hbbdea8ea),
	.w8(32'hbb4401ce),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8032),
	.w1(32'hbb9aa35f),
	.w2(32'hbbcd368e),
	.w3(32'hbb8211c2),
	.w4(32'hbb95d133),
	.w5(32'hbc3ead36),
	.w6(32'hbae78cc0),
	.w7(32'hbbb42edb),
	.w8(32'hbc92dcf2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc684d0e),
	.w1(32'hbca55e03),
	.w2(32'hbc5198c7),
	.w3(32'hbca2a9fd),
	.w4(32'hbc19687c),
	.w5(32'h3a057c09),
	.w6(32'hbcac7ca0),
	.w7(32'hbc61a301),
	.w8(32'hba372c34),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2349eb),
	.w1(32'hb9611ac1),
	.w2(32'hbaeeca7e),
	.w3(32'h3b9583c5),
	.w4(32'h3b20cd77),
	.w5(32'hbaee81ef),
	.w6(32'h3b5931cb),
	.w7(32'hb920b0cf),
	.w8(32'hbb61ebb5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e3ca),
	.w1(32'h390936dd),
	.w2(32'hb9060de6),
	.w3(32'hbb9e7617),
	.w4(32'hbab2a2a4),
	.w5(32'hbb36dbe9),
	.w6(32'hbba28689),
	.w7(32'h3a96076a),
	.w8(32'hbb3705a4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba228ce6),
	.w1(32'hba09dabe),
	.w2(32'h3a98bdb6),
	.w3(32'hbba9eae8),
	.w4(32'hbb8359dc),
	.w5(32'hbc27ef91),
	.w6(32'hbb65d68f),
	.w7(32'h384de632),
	.w8(32'hbc09ccb6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2f58),
	.w1(32'hbc1bddfc),
	.w2(32'hbc0a9e6e),
	.w3(32'hbc7b77ee),
	.w4(32'hbc50bfbd),
	.w5(32'hbc2acc61),
	.w6(32'hbc122d87),
	.w7(32'hbc17326d),
	.w8(32'hbc13167e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26842b),
	.w1(32'hbbba65d2),
	.w2(32'hbc116f17),
	.w3(32'hbc17d741),
	.w4(32'hbbb93a23),
	.w5(32'hbba6e360),
	.w6(32'hbbe21289),
	.w7(32'hbc07f913),
	.w8(32'hbba61940),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b67e8),
	.w1(32'hbb0a5e19),
	.w2(32'hbabe9f0f),
	.w3(32'hbc010fd7),
	.w4(32'hbbf75821),
	.w5(32'hb97871e6),
	.w6(32'hbbb0bb51),
	.w7(32'hbb8e043e),
	.w8(32'hbb3d27ef),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901e8af),
	.w1(32'hbaa48edd),
	.w2(32'h3aaf0de4),
	.w3(32'hbb34d90e),
	.w4(32'h3aa4e18e),
	.w5(32'h3bab7f42),
	.w6(32'hbba3379c),
	.w7(32'hb89d357d),
	.w8(32'h3b20e827),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd47d3c),
	.w1(32'h3a5daec6),
	.w2(32'h3b74c0ad),
	.w3(32'h3b38a7d3),
	.w4(32'h3bc05062),
	.w5(32'hbbd885c7),
	.w6(32'hba5ca98b),
	.w7(32'h3a1a8816),
	.w8(32'hbbc1d079),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0207),
	.w1(32'hbc12c3b2),
	.w2(32'hbc2a156a),
	.w3(32'hbc04c472),
	.w4(32'hbbe38550),
	.w5(32'hbbb20066),
	.w6(32'hbbfa9e7b),
	.w7(32'hbc0876b0),
	.w8(32'hbbbd35d1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb41e8e),
	.w1(32'hbb8f4948),
	.w2(32'hbae73fa3),
	.w3(32'hbba9d9e7),
	.w4(32'hb9a043ac),
	.w5(32'hbb17d262),
	.w6(32'hbb5aa6ed),
	.w7(32'h3a5984fd),
	.w8(32'hbb9962b3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f353),
	.w1(32'hbabde2c0),
	.w2(32'hbbb41276),
	.w3(32'hbb75a485),
	.w4(32'hbbe489f6),
	.w5(32'hbc902732),
	.w6(32'hbbe61045),
	.w7(32'hbc23ab17),
	.w8(32'hbc89daad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ffc45),
	.w1(32'hbc966b42),
	.w2(32'hbc7a910f),
	.w3(32'hbc9d3046),
	.w4(32'hbc8ce8ea),
	.w5(32'h3b4c64f7),
	.w6(32'hbc733e23),
	.w7(32'hbc71b693),
	.w8(32'h3b76351b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bd6dc),
	.w1(32'hbb821cec),
	.w2(32'hbb72a711),
	.w3(32'hbab7cab1),
	.w4(32'h394a54c8),
	.w5(32'h3a79e4b6),
	.w6(32'hbac474f4),
	.w7(32'hbb235457),
	.w8(32'hbbdbc14a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39ada8),
	.w1(32'hbc1101e2),
	.w2(32'hbc26b638),
	.w3(32'hbbbd3404),
	.w4(32'hbb801372),
	.w5(32'h3ac839d3),
	.w6(32'hbc7cb693),
	.w7(32'hbc20777d),
	.w8(32'h3aed45a8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa96165),
	.w1(32'hbb54d588),
	.w2(32'hbb667a6f),
	.w3(32'hb9ca0c0d),
	.w4(32'h39f17076),
	.w5(32'hbbd198a6),
	.w6(32'hbb424adc),
	.w7(32'hbadb19a1),
	.w8(32'hbbb751b2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dba13),
	.w1(32'hbc65c961),
	.w2(32'hbba524eb),
	.w3(32'hbc1922aa),
	.w4(32'hbb298d37),
	.w5(32'hbbe05d84),
	.w6(32'hbc0b9576),
	.w7(32'hbb273a64),
	.w8(32'hbbd75c3a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc496472),
	.w1(32'hbc4465f4),
	.w2(32'hbc3b5cb4),
	.w3(32'hbbf12e43),
	.w4(32'hbc01b77e),
	.w5(32'hbb622bd3),
	.w6(32'hbbe2dbb9),
	.w7(32'hbc124c56),
	.w8(32'hbb60c27c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca1000),
	.w1(32'h3b118373),
	.w2(32'h3a9a2bf3),
	.w3(32'hbbc01365),
	.w4(32'hbbb08dc0),
	.w5(32'h3ba7e851),
	.w6(32'hbbd824ec),
	.w7(32'hbb93e32f),
	.w8(32'h3b910971),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3413c9),
	.w1(32'h3b9a1944),
	.w2(32'h3b4bad96),
	.w3(32'h3c04e42b),
	.w4(32'h3bbd0be3),
	.w5(32'hbb42bc76),
	.w6(32'h3c179908),
	.w7(32'h3bd7df89),
	.w8(32'hb973ed62),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0568c5),
	.w1(32'h3ab06308),
	.w2(32'hbb70f295),
	.w3(32'h3a62039b),
	.w4(32'hbba2f719),
	.w5(32'hbb6db64a),
	.w6(32'h3921d3cd),
	.w7(32'hbbd57e3c),
	.w8(32'hbb9931ac),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92fbab),
	.w1(32'h39bd74dd),
	.w2(32'hbb1588dc),
	.w3(32'hbb4a7056),
	.w4(32'hbb1e2c6b),
	.w5(32'h390f5b79),
	.w6(32'h3a0e8e72),
	.w7(32'hbb858524),
	.w8(32'h3a8d4767),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa47037),
	.w1(32'h3b07ce52),
	.w2(32'hbbd2ff90),
	.w3(32'h3b239cd6),
	.w4(32'hbb94bbbb),
	.w5(32'hbc01e34c),
	.w6(32'h3a774838),
	.w7(32'hbbb979ce),
	.w8(32'hbc143796),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bca67),
	.w1(32'hbc3d6d8c),
	.w2(32'hbc819c4e),
	.w3(32'hbb9cde41),
	.w4(32'hbc2a854e),
	.w5(32'h39549b1d),
	.w6(32'hbbafc878),
	.w7(32'hbc555e31),
	.w8(32'hbaff02e4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2f5e),
	.w1(32'hbc0635e6),
	.w2(32'hbc2eb989),
	.w3(32'hbb38c6e7),
	.w4(32'hbb388a27),
	.w5(32'hbc32b621),
	.w6(32'hbb9936a7),
	.w7(32'hbc0467fd),
	.w8(32'hbc4f07b9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fe410),
	.w1(32'hbb9b6159),
	.w2(32'hbc1c0d8d),
	.w3(32'hbb9006f2),
	.w4(32'hbc0a0757),
	.w5(32'hbc2c10d8),
	.w6(32'hbb9b52b7),
	.w7(32'hbc2ee08e),
	.w8(32'hbc210b36),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08114e),
	.w1(32'h3a9705ce),
	.w2(32'hbad8945e),
	.w3(32'hbc1f7063),
	.w4(32'hbc228180),
	.w5(32'hbc0d0ea0),
	.w6(32'hbb0180e3),
	.w7(32'hbbd5a25f),
	.w8(32'hbbf5e8bc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe81fc1),
	.w1(32'hbbe75fd0),
	.w2(32'hbbeb4ec5),
	.w3(32'hbc311815),
	.w4(32'hbc113754),
	.w5(32'hbc278c96),
	.w6(32'hbc191bae),
	.w7(32'hbc158b89),
	.w8(32'hbc8842dd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867898),
	.w1(32'hbc549f67),
	.w2(32'hbc44d06a),
	.w3(32'hbbeb40a9),
	.w4(32'hbc13c1fe),
	.w5(32'hba30a5e3),
	.w6(32'hbc0d7428),
	.w7(32'hbc764194),
	.w8(32'h3997daf8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a884367),
	.w1(32'hbaf62b15),
	.w2(32'hbacc52d4),
	.w3(32'hbb884c69),
	.w4(32'hbb9276b7),
	.w5(32'hbb17abe1),
	.w6(32'hbbb9897c),
	.w7(32'hbb938f8d),
	.w8(32'h3bb6c511),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb3fc),
	.w1(32'h3a1aec6b),
	.w2(32'h39a5846f),
	.w3(32'h3a7a42ac),
	.w4(32'h3b9be3a2),
	.w5(32'h3ba73036),
	.w6(32'hbb3f15bb),
	.w7(32'hbb36eca6),
	.w8(32'h3b19c5c4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22c643),
	.w1(32'hbb9f43a8),
	.w2(32'hba2f163b),
	.w3(32'hbb5a9c26),
	.w4(32'hb9fa1d86),
	.w5(32'h3af4e1ce),
	.w6(32'hbaf71d80),
	.w7(32'hbb523450),
	.w8(32'hbbb1ffbc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38cbae),
	.w1(32'hbb65bafa),
	.w2(32'hbc2753d7),
	.w3(32'hbb544993),
	.w4(32'hbbbb78a9),
	.w5(32'hbb307d40),
	.w6(32'hbab9ec9c),
	.w7(32'hbbf6e11e),
	.w8(32'hbab54106),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474b88),
	.w1(32'h39f51932),
	.w2(32'hbb80e8a6),
	.w3(32'hbb3c647b),
	.w4(32'h398aaf8a),
	.w5(32'h3aac2c4f),
	.w6(32'h3c47cd43),
	.w7(32'h3b34bc60),
	.w8(32'h3b994d9f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba68f9),
	.w1(32'h3c062bf7),
	.w2(32'h3b392a59),
	.w3(32'hbbb8bd12),
	.w4(32'hbb53b4ce),
	.w5(32'hbb07f75c),
	.w6(32'h3b3eabfc),
	.w7(32'h3c254923),
	.w8(32'hbb2ae050),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90632f2),
	.w1(32'h399de76e),
	.w2(32'hba9a1e78),
	.w3(32'h3baab0ea),
	.w4(32'hbb2f2472),
	.w5(32'h3a215c23),
	.w6(32'hbba6e0a4),
	.w7(32'hbbedae42),
	.w8(32'h3a94753e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1351),
	.w1(32'hbacd0756),
	.w2(32'h3b6bbfe8),
	.w3(32'hbb6ce27b),
	.w4(32'h3a004c94),
	.w5(32'hbb0da66d),
	.w6(32'hb9dcc040),
	.w7(32'hba1e909d),
	.w8(32'h3bf3fc4b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d70e),
	.w1(32'hbbc31f66),
	.w2(32'hbabefc3f),
	.w3(32'h3c6a3c2c),
	.w4(32'h3b93b173),
	.w5(32'h3bb09efa),
	.w6(32'h3c5e8303),
	.w7(32'hbb816d2b),
	.w8(32'h3b8f1149),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af87b68),
	.w1(32'h3ac9a234),
	.w2(32'h3942a361),
	.w3(32'h3ab2b1f9),
	.w4(32'h3b9d21a6),
	.w5(32'h3b55f095),
	.w6(32'hb8fc75a5),
	.w7(32'hba989f0f),
	.w8(32'h3a98a7e0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bcbc5),
	.w1(32'hb9320b6d),
	.w2(32'h39a7aa77),
	.w3(32'hbb4a4d88),
	.w4(32'hbb87d15c),
	.w5(32'h3a57a218),
	.w6(32'hbb748c80),
	.w7(32'hbb5af612),
	.w8(32'hbb09c259),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24da58),
	.w1(32'hbb336a06),
	.w2(32'hbaec04c3),
	.w3(32'h3b0fa6b8),
	.w4(32'h38e77d92),
	.w5(32'hb994ed7c),
	.w6(32'hbb4cc56f),
	.w7(32'hbb8254b7),
	.w8(32'h3a8cdf68),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947f994),
	.w1(32'hbb62c055),
	.w2(32'h3905d701),
	.w3(32'h3bbcc227),
	.w4(32'h3b4ce054),
	.w5(32'hbb181101),
	.w6(32'hba20bf14),
	.w7(32'hbbac0743),
	.w8(32'hba364901),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9092f40),
	.w1(32'h3b4e08da),
	.w2(32'h3b3b0959),
	.w3(32'h3adf1ad3),
	.w4(32'hba1e4adc),
	.w5(32'hba752970),
	.w6(32'h3b4214d7),
	.w7(32'hba32b31b),
	.w8(32'hbb85e199),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d437),
	.w1(32'hbae50a0b),
	.w2(32'hbb277604),
	.w3(32'h3b38126b),
	.w4(32'hbb2ffff3),
	.w5(32'hbb84e141),
	.w6(32'hb91b4c94),
	.w7(32'hbbd2afea),
	.w8(32'hb8ff851a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3612),
	.w1(32'hba8952bf),
	.w2(32'hbbcc0123),
	.w3(32'hbbce4f86),
	.w4(32'h3a230511),
	.w5(32'h3b259b4d),
	.w6(32'h3cab7e63),
	.w7(32'h3c4fb286),
	.w8(32'h3af7d9ae),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3055a),
	.w1(32'hb873cb2c),
	.w2(32'hbba6281b),
	.w3(32'h3b727114),
	.w4(32'h3bc259cf),
	.w5(32'hbb6004b7),
	.w6(32'hba130831),
	.w7(32'h3b5c7bf1),
	.w8(32'hbacdceee),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba714c4b),
	.w1(32'h3a2811dc),
	.w2(32'h39973780),
	.w3(32'h3a820281),
	.w4(32'hbb04226c),
	.w5(32'hbab0c71d),
	.w6(32'h3b336502),
	.w7(32'hbb7ee65e),
	.w8(32'hbabe01c5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ca2d2),
	.w1(32'hbaebdd87),
	.w2(32'hbb5869a5),
	.w3(32'hbb3832cb),
	.w4(32'h390e9de4),
	.w5(32'h3b3fc017),
	.w6(32'hba0508ac),
	.w7(32'hb8916abb),
	.w8(32'hbb1aebf9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cd400),
	.w1(32'hbae16a18),
	.w2(32'hbb2e6e12),
	.w3(32'h393c86b5),
	.w4(32'hbb0fa910),
	.w5(32'hba36d4b8),
	.w6(32'hbb5c0ce5),
	.w7(32'hbb59a6ff),
	.w8(32'hbb4c8205),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8241a7),
	.w1(32'hbb654f3a),
	.w2(32'hbb482c7d),
	.w3(32'hbb117b4b),
	.w4(32'h39c73bdb),
	.w5(32'hb986f810),
	.w6(32'hbb645110),
	.w7(32'hbb3b8620),
	.w8(32'hba4dec71),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ada0aa),
	.w1(32'hbaf57677),
	.w2(32'hba4751ab),
	.w3(32'hbc137eff),
	.w4(32'hbadd2cb1),
	.w5(32'h3bbbcb0a),
	.w6(32'hbbddbe45),
	.w7(32'h3a17cfd5),
	.w8(32'h3ae28e05),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8aa91),
	.w1(32'h3bc990cb),
	.w2(32'h3b4d2d70),
	.w3(32'h398a9fab),
	.w4(32'hb8cc47c4),
	.w5(32'hba85eb2e),
	.w6(32'h3c068322),
	.w7(32'h3ba8d43d),
	.w8(32'h3a8e6845),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b78e0),
	.w1(32'hbb23d251),
	.w2(32'hb985b466),
	.w3(32'h3ab56da8),
	.w4(32'hbab7435f),
	.w5(32'hbb6fd933),
	.w6(32'h3aeeb0f3),
	.w7(32'hbb858d12),
	.w8(32'hbc1452b2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda823),
	.w1(32'h39934c6d),
	.w2(32'h3b518273),
	.w3(32'h3b5953f3),
	.w4(32'hba284cde),
	.w5(32'hb997e88c),
	.w6(32'hbb2dec64),
	.w7(32'hbb86c469),
	.w8(32'h39dafc64),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ae49c),
	.w1(32'hbaf67349),
	.w2(32'h3b9c62ad),
	.w3(32'h3a85855d),
	.w4(32'hba139e54),
	.w5(32'h3835a1b1),
	.w6(32'hbb4a32f4),
	.w7(32'hb94bfb2e),
	.w8(32'hbb7c169c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c12e4),
	.w1(32'hbac8935e),
	.w2(32'hba789194),
	.w3(32'h3b46eefe),
	.w4(32'hba20c858),
	.w5(32'h3ae1d64b),
	.w6(32'hba53b972),
	.w7(32'hb7f21def),
	.w8(32'h3b942f8f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b8459),
	.w1(32'hbbab984b),
	.w2(32'hbb80f4f4),
	.w3(32'hbc2d6ba3),
	.w4(32'hbbe937d1),
	.w5(32'h3a579a21),
	.w6(32'h3b7c4b8a),
	.w7(32'h3ae168a8),
	.w8(32'hba28187d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83e039),
	.w1(32'hbb1aa80b),
	.w2(32'h3a175c95),
	.w3(32'h3b5223cc),
	.w4(32'hba37dd9d),
	.w5(32'h3aa54547),
	.w6(32'hbb3589ff),
	.w7(32'hbb4c48fa),
	.w8(32'h3b4edfca),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f989),
	.w1(32'h3b814b29),
	.w2(32'h3b419eb5),
	.w3(32'hbb0b233f),
	.w4(32'h3b20032d),
	.w5(32'h3a1d1471),
	.w6(32'h3adeec6c),
	.w7(32'h3be27085),
	.w8(32'hba03600a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule