module layer_10_featuremap_307(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb735528),
	.w1(32'hbb2d6d5d),
	.w2(32'hbbce14a1),
	.w3(32'hbbc4ec0f),
	.w4(32'hbbbd5eb9),
	.w5(32'hbb7c7d75),
	.w6(32'hbc0363a7),
	.w7(32'hbc05aced),
	.w8(32'h3a966146),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163ef6),
	.w1(32'hbbf3d258),
	.w2(32'hbb9be6a0),
	.w3(32'h3b44aa5b),
	.w4(32'hbbe894f3),
	.w5(32'h3bc777a7),
	.w6(32'h3b78eb66),
	.w7(32'hbb06caf2),
	.w8(32'hba8da30c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5168),
	.w1(32'h3b16a9c0),
	.w2(32'h3ae33365),
	.w3(32'hbb99a179),
	.w4(32'hba25edd5),
	.w5(32'h3b94d289),
	.w6(32'h3b044e68),
	.w7(32'hb5e760ed),
	.w8(32'h3b821feb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191c26),
	.w1(32'h3b3c82c7),
	.w2(32'h3b95b2f4),
	.w3(32'h3b7fc842),
	.w4(32'h3c1584b4),
	.w5(32'hbbc74e98),
	.w6(32'hba19d350),
	.w7(32'h3bfcedcd),
	.w8(32'hbcd91edb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27b2fb),
	.w1(32'h3bcdf9bf),
	.w2(32'h3b3ad60d),
	.w3(32'hbb92d844),
	.w4(32'h3b6252f2),
	.w5(32'h3b32842d),
	.w6(32'hbc7a8e47),
	.w7(32'hbca377d4),
	.w8(32'hba6d631f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68387a),
	.w1(32'hbb817e38),
	.w2(32'hbbc4d5c2),
	.w3(32'h3af4e01c),
	.w4(32'h3b5f17eb),
	.w5(32'hba6c6df5),
	.w6(32'hbb99702e),
	.w7(32'hbb1ba7f0),
	.w8(32'hbaf797f9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1c2c9),
	.w1(32'hbac9d172),
	.w2(32'hba5e3a09),
	.w3(32'h3b601d2a),
	.w4(32'hba29f49b),
	.w5(32'hbbb2360c),
	.w6(32'hbb1c6a46),
	.w7(32'h3a5d2ff2),
	.w8(32'hbaa96be1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd577a0),
	.w1(32'hbb622f0f),
	.w2(32'hbbf4a8ab),
	.w3(32'hbbdafa85),
	.w4(32'hbb53d401),
	.w5(32'h3bda8fc6),
	.w6(32'hbc260a01),
	.w7(32'hbb880086),
	.w8(32'h3b45a8c2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba726b0),
	.w1(32'hbbad1bb4),
	.w2(32'hbbb6abd0),
	.w3(32'h3b6ffcc8),
	.w4(32'h3b53d69d),
	.w5(32'h39b07a3a),
	.w6(32'hbb4225db),
	.w7(32'hb9ea5c35),
	.w8(32'hbad99dd6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3aaf4),
	.w1(32'hbb649dbf),
	.w2(32'hbb8cc1d4),
	.w3(32'hbaee4b37),
	.w4(32'h3bb0d28d),
	.w5(32'h3c4a6fa4),
	.w6(32'hbbf1843c),
	.w7(32'hbb0d7e2e),
	.w8(32'h3a8b4db1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb3631),
	.w1(32'hbb350d09),
	.w2(32'hbb962b53),
	.w3(32'h3b8e87f7),
	.w4(32'h3bd1e28b),
	.w5(32'hba853bcc),
	.w6(32'hbb84c397),
	.w7(32'hba135076),
	.w8(32'hbbf512a7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc866b),
	.w1(32'hbbb17b19),
	.w2(32'hbaa8bbe4),
	.w3(32'hbc44e796),
	.w4(32'hb8cce599),
	.w5(32'hbc54dbb0),
	.w6(32'hbc123ea1),
	.w7(32'h3ae8a950),
	.w8(32'hbc103022),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93462),
	.w1(32'h3be7ec85),
	.w2(32'hba124178),
	.w3(32'hbcf6d658),
	.w4(32'hbc704cc9),
	.w5(32'h3b81760e),
	.w6(32'hbc573eb3),
	.w7(32'hbb74e950),
	.w8(32'h3b9c1bbf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22d734),
	.w1(32'h38eeb611),
	.w2(32'hba834183),
	.w3(32'h39dcf4d0),
	.w4(32'hbb300f6a),
	.w5(32'h3b98655c),
	.w6(32'h3bb56b21),
	.w7(32'hba859417),
	.w8(32'h3c07f70f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6e2c1),
	.w1(32'hbb54ece1),
	.w2(32'hbae1ec51),
	.w3(32'h3b8cd57f),
	.w4(32'h3b597f8c),
	.w5(32'h3a8572f7),
	.w6(32'hbaf8a21a),
	.w7(32'hba5231ce),
	.w8(32'h3b563d35),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03069),
	.w1(32'hbba59750),
	.w2(32'hbb1c0421),
	.w3(32'h3b7330b0),
	.w4(32'h3aa26cd5),
	.w5(32'hbb348e22),
	.w6(32'h3b870526),
	.w7(32'h3ba7d7d8),
	.w8(32'hba611946),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a7166),
	.w1(32'hbc876688),
	.w2(32'hbc6a0323),
	.w3(32'h3a8637ba),
	.w4(32'h3b1ac214),
	.w5(32'hbc253f7f),
	.w6(32'hbb5efd16),
	.w7(32'hba7789e3),
	.w8(32'hbb30f828),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389e13),
	.w1(32'h3aa73675),
	.w2(32'hbb149b3e),
	.w3(32'hbca0c311),
	.w4(32'hbc5837d6),
	.w5(32'hba802bd0),
	.w6(32'hbc49e157),
	.w7(32'hbb0dad42),
	.w8(32'h3befa901),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47986f),
	.w1(32'hbb913628),
	.w2(32'hbba4af59),
	.w3(32'hbb466df1),
	.w4(32'hba4eb051),
	.w5(32'h3b012579),
	.w6(32'h3b33de36),
	.w7(32'h3b62ff2d),
	.w8(32'hbb9373c2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02c256),
	.w1(32'h3acbfc96),
	.w2(32'h3be5bc2f),
	.w3(32'hbb0e2710),
	.w4(32'hbabbf6c1),
	.w5(32'hbabd647f),
	.w6(32'h3c05a1ee),
	.w7(32'h3b34f423),
	.w8(32'h3a16e6e5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0387c0),
	.w1(32'h3b9072ea),
	.w2(32'h3c10486e),
	.w3(32'hbb1f98b3),
	.w4(32'hbb2a1001),
	.w5(32'h3bf8a99a),
	.w6(32'h3b12bb71),
	.w7(32'h3bd22f8d),
	.w8(32'h3a64ce64),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1977),
	.w1(32'hbb4e6015),
	.w2(32'h395564df),
	.w3(32'h3c23f1f7),
	.w4(32'h3c28e226),
	.w5(32'hbbb95fa0),
	.w6(32'hbb944501),
	.w7(32'h3b6526be),
	.w8(32'hbb93a3c9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560d46),
	.w1(32'h3b4e1018),
	.w2(32'hbbdbe1a6),
	.w3(32'hbbf99327),
	.w4(32'hbb238f27),
	.w5(32'hbc6dd8bc),
	.w6(32'hbb5c91e6),
	.w7(32'hbb00f93c),
	.w8(32'hbb0badc8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164a3c),
	.w1(32'h3c4da12a),
	.w2(32'h3b765e25),
	.w3(32'hbc855e9a),
	.w4(32'hbc05bb7f),
	.w5(32'h3c660f3f),
	.w6(32'hbb4fab0f),
	.w7(32'h3a804f3a),
	.w8(32'h3b9ba6cb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86e2245),
	.w1(32'h3b5f8e35),
	.w2(32'h3ba20d5d),
	.w3(32'hbb742a35),
	.w4(32'h3bd2c569),
	.w5(32'h3bbe54d9),
	.w6(32'h3cb374f4),
	.w7(32'h3b154929),
	.w8(32'h3c4a70c8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bc7e97),
	.w1(32'hbc7561b9),
	.w2(32'hbbc7b508),
	.w3(32'h3c2b29e0),
	.w4(32'h3c01d3b9),
	.w5(32'h3c0306ac),
	.w6(32'h3b987c7b),
	.w7(32'h39aeb5a3),
	.w8(32'h3a08cf01),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187730),
	.w1(32'hbca26850),
	.w2(32'hbc7a403f),
	.w3(32'h3c868874),
	.w4(32'h3c3b78e9),
	.w5(32'hba279c3c),
	.w6(32'hbaa571c7),
	.w7(32'hba69c91b),
	.w8(32'hbb15c21e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71650d),
	.w1(32'hbb34fc3d),
	.w2(32'hbb731377),
	.w3(32'hbbb4288a),
	.w4(32'hbba020c1),
	.w5(32'hbb65e9fc),
	.w6(32'hbbc83a01),
	.w7(32'hbc005aa5),
	.w8(32'hbbee78b5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba222047),
	.w1(32'hbaf466a1),
	.w2(32'h3aa2ec73),
	.w3(32'hbbf8cd11),
	.w4(32'hbb9ca9e5),
	.w5(32'hba9553f4),
	.w6(32'h3b5b487b),
	.w7(32'h3a951cad),
	.w8(32'hbb4b6738),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74e489),
	.w1(32'h3b4f0e89),
	.w2(32'hbb8faf6a),
	.w3(32'hbbc648df),
	.w4(32'hbbb2d9ab),
	.w5(32'h3c8ab4bb),
	.w6(32'h3b258470),
	.w7(32'h3a7c1528),
	.w8(32'h3abdabc9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b01dd),
	.w1(32'h3bab8671),
	.w2(32'h3b8eafaa),
	.w3(32'h3cb7d4b8),
	.w4(32'h3c29212d),
	.w5(32'hbc2b5c02),
	.w6(32'h3cb7ff66),
	.w7(32'h3ba22023),
	.w8(32'hbba62168),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4988f),
	.w1(32'hbbbce840),
	.w2(32'hbb9ed9a8),
	.w3(32'hbc523c91),
	.w4(32'hbc304bbc),
	.w5(32'hbb80691d),
	.w6(32'hbb6ab587),
	.w7(32'hbc5363a4),
	.w8(32'h3c4e3bce),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfec22),
	.w1(32'hbcab1eb2),
	.w2(32'hbc49f055),
	.w3(32'h3ccef83f),
	.w4(32'h3c3da252),
	.w5(32'hbbc1dc39),
	.w6(32'h3b5e18e6),
	.w7(32'h3bc8287a),
	.w8(32'h3be99016),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fa971),
	.w1(32'h3c95bf94),
	.w2(32'h3c44bc84),
	.w3(32'hbc5e5ce1),
	.w4(32'hbc3fee2f),
	.w5(32'hbb540f90),
	.w6(32'h3ba66a67),
	.w7(32'h3b0f2d07),
	.w8(32'hbb51b6bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aae5b),
	.w1(32'hbad6ee8b),
	.w2(32'hb9cddd34),
	.w3(32'hbc395c96),
	.w4(32'hbad44115),
	.w5(32'h3b2726ac),
	.w6(32'h3b1fb724),
	.w7(32'h3af78657),
	.w8(32'hbba16d80),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063fe9),
	.w1(32'h3b830937),
	.w2(32'h3b473465),
	.w3(32'hbc217263),
	.w4(32'hba0b3519),
	.w5(32'h3c41799d),
	.w6(32'h393fb0fc),
	.w7(32'h3ab0e7d6),
	.w8(32'h3b8a4ae1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba920c4e),
	.w1(32'hbb896fc1),
	.w2(32'hbb7bcc54),
	.w3(32'h3c353ec8),
	.w4(32'h3b2aee40),
	.w5(32'h3c3aecb1),
	.w6(32'h3c8b4343),
	.w7(32'h3c296e75),
	.w8(32'hba462040),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978bcb),
	.w1(32'hbc090d2c),
	.w2(32'hbbb8d302),
	.w3(32'h3ca5378c),
	.w4(32'h3c2bf7db),
	.w5(32'h3991d303),
	.w6(32'h3b6d7d40),
	.w7(32'h3a92a87e),
	.w8(32'hbc080671),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33f2b3),
	.w1(32'h3c362ae7),
	.w2(32'h3c4cf3f7),
	.w3(32'h3b4d2528),
	.w4(32'hbc11d3ca),
	.w5(32'hbb9d9f49),
	.w6(32'h3ba20bff),
	.w7(32'hbbea0571),
	.w8(32'h3a93c9e4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa6a4f),
	.w1(32'h3c2f992c),
	.w2(32'h3bd4d6d4),
	.w3(32'hbc47c5a2),
	.w4(32'hbb579cc3),
	.w5(32'hbb3a3849),
	.w6(32'hbbc2dba7),
	.w7(32'h3b6cd3f6),
	.w8(32'hbb764328),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad825),
	.w1(32'hba22758e),
	.w2(32'hba8d0568),
	.w3(32'hbc33e480),
	.w4(32'h3a5170f2),
	.w5(32'h3b62ea71),
	.w6(32'hbc03413c),
	.w7(32'h3a007400),
	.w8(32'hba8a12ad),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb6d93),
	.w1(32'hbc36f25f),
	.w2(32'hbbcba73e),
	.w3(32'h3be1025c),
	.w4(32'h3bb72f6f),
	.w5(32'h3c330f2a),
	.w6(32'hbbd5cb33),
	.w7(32'hbae70ddc),
	.w8(32'h3bf27a7b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1257),
	.w1(32'hbc144d4f),
	.w2(32'hbb24c759),
	.w3(32'h3c291033),
	.w4(32'h3b7ec5df),
	.w5(32'h3c4d487e),
	.w6(32'hba89186d),
	.w7(32'h3bff4dac),
	.w8(32'hbb62908e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb10113),
	.w1(32'hbd24a8c8),
	.w2(32'hbcc39e72),
	.w3(32'h3cf61ccc),
	.w4(32'h3c59e1d2),
	.w5(32'h3b5149c3),
	.w6(32'h3bf074cc),
	.w7(32'hbaeb0cb9),
	.w8(32'h3c0cc279),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1446),
	.w1(32'hbc4ff5cb),
	.w2(32'hbbbc3e62),
	.w3(32'h3c307180),
	.w4(32'h3b7f13b9),
	.w5(32'h3b6f9332),
	.w6(32'hbc0abb06),
	.w7(32'hbba561c0),
	.w8(32'h3a6a715f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b6e1e),
	.w1(32'h3a1d2c86),
	.w2(32'h3c0fdbb1),
	.w3(32'hbaf894b7),
	.w4(32'hbb26216e),
	.w5(32'h3c10d032),
	.w6(32'h3b3e75f2),
	.w7(32'hba6aa8a5),
	.w8(32'h3b87214e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbc883),
	.w1(32'hbbd1ffa4),
	.w2(32'h3a53110d),
	.w3(32'h3b0dfc0b),
	.w4(32'h3c19d6e7),
	.w5(32'h3bfaf57d),
	.w6(32'h3b717faa),
	.w7(32'h3b789acd),
	.w8(32'h38834500),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc608e66),
	.w1(32'hbbcc4a69),
	.w2(32'hbbcb6679),
	.w3(32'hbaf3f589),
	.w4(32'h3c120a93),
	.w5(32'h3b3af779),
	.w6(32'hbc2e0852),
	.w7(32'h3a4a99c5),
	.w8(32'h3baba6c0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbca88),
	.w1(32'h3c903699),
	.w2(32'h3c2d8f52),
	.w3(32'hbb746242),
	.w4(32'hbb3d6ce6),
	.w5(32'h3b69d776),
	.w6(32'hba779d11),
	.w7(32'h3baacbd0),
	.w8(32'hb9fc5d5f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09cc26),
	.w1(32'hbbd78723),
	.w2(32'hbb805c5f),
	.w3(32'h3c0e75ef),
	.w4(32'h3c2cb8a3),
	.w5(32'hbc384b2e),
	.w6(32'hbb921d69),
	.w7(32'h39b98c77),
	.w8(32'hbafab847),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d074),
	.w1(32'h3c20d35c),
	.w2(32'hbc04d695),
	.w3(32'hbb910239),
	.w4(32'h39c59e8f),
	.w5(32'hba452460),
	.w6(32'h3b68e25f),
	.w7(32'hbaf1652c),
	.w8(32'hbbe2086f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4673ae),
	.w1(32'hbc293380),
	.w2(32'hbb740324),
	.w3(32'hba1f1f86),
	.w4(32'hb91277fa),
	.w5(32'h3c034a04),
	.w6(32'hbc178b2d),
	.w7(32'h3a81090a),
	.w8(32'h3af1b4a1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d0f40),
	.w1(32'h3ae76609),
	.w2(32'hbc04355e),
	.w3(32'hbb92a9f0),
	.w4(32'hbb08b76f),
	.w5(32'h3b89ce87),
	.w6(32'h3b8f87ea),
	.w7(32'hbb74fb16),
	.w8(32'h3b12e8d5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba379c85),
	.w1(32'hbc278e94),
	.w2(32'hbc2758c0),
	.w3(32'h3c1d2794),
	.w4(32'hbc264439),
	.w5(32'hbb0cb524),
	.w6(32'h3b78404c),
	.w7(32'h3c002a3a),
	.w8(32'hba84a9de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae049ae),
	.w1(32'h3b659707),
	.w2(32'h3b6f72b9),
	.w3(32'hbb280fa9),
	.w4(32'hb903970c),
	.w5(32'hbad13b9e),
	.w6(32'h3bc35518),
	.w7(32'h3ba3732a),
	.w8(32'h3a0a1086),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43c93),
	.w1(32'h3a412648),
	.w2(32'hb9ba3a06),
	.w3(32'hb9384ac2),
	.w4(32'h3bbeaeba),
	.w5(32'hbb6f4864),
	.w6(32'h3b9745f2),
	.w7(32'h39dd9c57),
	.w8(32'h39dcfae1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b074674),
	.w1(32'h398e9e61),
	.w2(32'hbb6d2764),
	.w3(32'hbb749ea4),
	.w4(32'h3befd7d3),
	.w5(32'h3c10bf9b),
	.w6(32'hbb89b7ae),
	.w7(32'hb815b85b),
	.w8(32'h3b5f2c2f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdea61b),
	.w1(32'hbba3fc04),
	.w2(32'h3a32c03e),
	.w3(32'h3c1b963c),
	.w4(32'hbbc9234f),
	.w5(32'h3896de85),
	.w6(32'h3b866730),
	.w7(32'hba450af8),
	.w8(32'hbabbd2ff),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53c0ac),
	.w1(32'hbc1d8fde),
	.w2(32'hbbfbb696),
	.w3(32'h3ba95f49),
	.w4(32'h3be318b6),
	.w5(32'h3c227cda),
	.w6(32'hbb899b4f),
	.w7(32'hbaf9b203),
	.w8(32'hbbe2b861),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7c1f8),
	.w1(32'hbc09e8e6),
	.w2(32'hbb69787d),
	.w3(32'h3bc7228c),
	.w4(32'h3c3bd2c6),
	.w5(32'hbbc8bd01),
	.w6(32'hbb4f5e48),
	.w7(32'hbb87a7eb),
	.w8(32'hbbe31bd4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94122),
	.w1(32'hbb3d6225),
	.w2(32'hbb398eb0),
	.w3(32'hbb9217a1),
	.w4(32'h3a9a8b76),
	.w5(32'hbad095a9),
	.w6(32'hbb7ba3e9),
	.w7(32'hbb0f3a4e),
	.w8(32'hba3b37a6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac10a2),
	.w1(32'hbb8d29d5),
	.w2(32'hbb9070b0),
	.w3(32'h3bf777e1),
	.w4(32'h3b802595),
	.w5(32'h39c85381),
	.w6(32'hbb38e472),
	.w7(32'hbb9f50c2),
	.w8(32'hbc0b467c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e7c4),
	.w1(32'h39b54f1d),
	.w2(32'hbaaac1a5),
	.w3(32'hbb333c64),
	.w4(32'hbb872592),
	.w5(32'hbb81e3b6),
	.w6(32'h3c4965c8),
	.w7(32'hbbbcfec9),
	.w8(32'hbb0005a5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c58c),
	.w1(32'h3bbd7cea),
	.w2(32'h3b8e547c),
	.w3(32'hbc23a2f4),
	.w4(32'h3ad8e11b),
	.w5(32'h3a1a520f),
	.w6(32'hba6d6d54),
	.w7(32'h3b1f8494),
	.w8(32'hbc218e9d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a625),
	.w1(32'h3c2a6c8d),
	.w2(32'h3b4383c4),
	.w3(32'hbbbf8e81),
	.w4(32'hb900561f),
	.w5(32'h3ba221d9),
	.w6(32'h3b77ae05),
	.w7(32'h3b982b58),
	.w8(32'h3a5b3f3a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cda4e),
	.w1(32'h3b8de247),
	.w2(32'hbb00365a),
	.w3(32'h3b973624),
	.w4(32'h3b4aa2a1),
	.w5(32'hba75bc3e),
	.w6(32'h3c4b5b6d),
	.w7(32'hbaa2c3f0),
	.w8(32'hbb850536),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8048fe),
	.w1(32'h3b085a74),
	.w2(32'hbb9f0852),
	.w3(32'hbbad5939),
	.w4(32'hbaa8e193),
	.w5(32'h3bdcec99),
	.w6(32'hbbab2eb9),
	.w7(32'hbbe1cff3),
	.w8(32'h3b151f92),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d6b2f),
	.w1(32'hbc50ac46),
	.w2(32'hbc0c0d31),
	.w3(32'h3b66f451),
	.w4(32'h3c12ca67),
	.w5(32'hbc2ea903),
	.w6(32'hbb558502),
	.w7(32'h3a04f3a7),
	.w8(32'hba9ea002),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de8f5f),
	.w1(32'h3b25d57e),
	.w2(32'hbc050905),
	.w3(32'hbc337166),
	.w4(32'hbb4caedb),
	.w5(32'h3c8502dc),
	.w6(32'hbb37215a),
	.w7(32'h3b70fdab),
	.w8(32'h3bcbb9c6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e19d8),
	.w1(32'hbc8c3508),
	.w2(32'hbb54f5af),
	.w3(32'h3cbfb0a4),
	.w4(32'h3c257b71),
	.w5(32'h3ca2ee1e),
	.w6(32'hbc1dcfac),
	.w7(32'h3b2432b4),
	.w8(32'h3beb126a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5829b4),
	.w1(32'hbc3871c4),
	.w2(32'hbbf2e4fa),
	.w3(32'h3cacbc62),
	.w4(32'h3c8e1b06),
	.w5(32'hbbb6b1a5),
	.w6(32'h3b65b818),
	.w7(32'h3c30b764),
	.w8(32'hbb00e2c6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88e752),
	.w1(32'h3bfe8c40),
	.w2(32'h3be80225),
	.w3(32'hbadb7992),
	.w4(32'hbb900ab2),
	.w5(32'h3b8e5df8),
	.w6(32'h3c0b2950),
	.w7(32'hba9becb0),
	.w8(32'hbaa75300),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b678178),
	.w1(32'h3bd9d036),
	.w2(32'h3bc019cb),
	.w3(32'h3b4b66dd),
	.w4(32'h3b30d3a2),
	.w5(32'hbb88a515),
	.w6(32'h3b199248),
	.w7(32'hba791ed0),
	.w8(32'h3b8f884f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85ac69),
	.w1(32'h3c52bb39),
	.w2(32'h3bb99749),
	.w3(32'hbc4efd88),
	.w4(32'hbc4e21cd),
	.w5(32'h3aac368b),
	.w6(32'h3ba26844),
	.w7(32'hbb3fb9bf),
	.w8(32'h39f4146f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd73f6),
	.w1(32'hbb9d95fd),
	.w2(32'hbc1d024a),
	.w3(32'h3a35bd12),
	.w4(32'h3af6ba5f),
	.w5(32'hbc6d50d5),
	.w6(32'h3a90814b),
	.w7(32'h39e864e3),
	.w8(32'hbaa8aa5d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12bf00),
	.w1(32'h3cb3235e),
	.w2(32'h3c00c772),
	.w3(32'hbd030546),
	.w4(32'hbca1fd11),
	.w5(32'h3b2c7fdc),
	.w6(32'hbbac6104),
	.w7(32'hbb7ed705),
	.w8(32'h3b91f174),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d7f51),
	.w1(32'hb9eb1e98),
	.w2(32'hbb040afc),
	.w3(32'hbc8561b2),
	.w4(32'hbb00116f),
	.w5(32'hbb760c47),
	.w6(32'hba2be3b1),
	.w7(32'h39096662),
	.w8(32'hb8097a5f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afa6a),
	.w1(32'hbb1d2c45),
	.w2(32'h3aefdbec),
	.w3(32'hba1351b6),
	.w4(32'hbac35f51),
	.w5(32'hbc042b94),
	.w6(32'hbb878955),
	.w7(32'hba94caed),
	.w8(32'h3bd9d155),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111832),
	.w1(32'h3c9e73ed),
	.w2(32'h3be0295e),
	.w3(32'hbcbec3e9),
	.w4(32'hbc1b7911),
	.w5(32'h3b410818),
	.w6(32'hbb214de3),
	.w7(32'h3bfaf65b),
	.w8(32'hb95971a6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c299a),
	.w1(32'hbae407e9),
	.w2(32'hbb5b8161),
	.w3(32'h39936dd6),
	.w4(32'hba9781f7),
	.w5(32'hbc5354af),
	.w6(32'hbbb4cce8),
	.w7(32'hbbcd220e),
	.w8(32'hbae6b34e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2517e3),
	.w1(32'h3c6d9c35),
	.w2(32'hbb5cab43),
	.w3(32'hbc7c6577),
	.w4(32'hbc0e2ef5),
	.w5(32'hba418889),
	.w6(32'hbae7f55a),
	.w7(32'hba5fb4ac),
	.w8(32'h3ba6b4d3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6f8a2),
	.w1(32'h3ca36690),
	.w2(32'h3bb36620),
	.w3(32'hbc2e396c),
	.w4(32'hbbf18ef7),
	.w5(32'h3a7440eb),
	.w6(32'hbb8691ba),
	.w7(32'hbb15e5e7),
	.w8(32'hbafc94f2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdb9ec),
	.w1(32'h3bf4ecf4),
	.w2(32'hbc2e5eae),
	.w3(32'hbbc16cb5),
	.w4(32'hbba229a2),
	.w5(32'h3be63989),
	.w6(32'h3c08de65),
	.w7(32'hbb9ccbb0),
	.w8(32'hba00fb7d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37676d),
	.w1(32'h3be6ece4),
	.w2(32'h3b610a63),
	.w3(32'hbbd0eea3),
	.w4(32'h3b1c0b05),
	.w5(32'hba2adfca),
	.w6(32'hbbda1ecb),
	.w7(32'hbaed3b11),
	.w8(32'h3b2d118d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a965b83),
	.w1(32'h3b431b18),
	.w2(32'hbb9aec0f),
	.w3(32'hbb0e9f9d),
	.w4(32'hba8ce9e1),
	.w5(32'hbba8d339),
	.w6(32'h3c428cfb),
	.w7(32'h3a32100f),
	.w8(32'hbc130d12),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995246b),
	.w1(32'h3b8a3313),
	.w2(32'hbbcc6a37),
	.w3(32'hb9e7a2a2),
	.w4(32'hbb802c29),
	.w5(32'h3bae1277),
	.w6(32'hbb1325d5),
	.w7(32'hbc40260f),
	.w8(32'h3b3b64a2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41fb4d),
	.w1(32'hbc7c940e),
	.w2(32'hbc3c8bd5),
	.w3(32'h3c8c00fe),
	.w4(32'hbad8208b),
	.w5(32'hbb1d18a6),
	.w6(32'h3a3c2d1f),
	.w7(32'hba91777f),
	.w8(32'h3b2d5032),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975abb5),
	.w1(32'h3b15a420),
	.w2(32'h3bd84b85),
	.w3(32'hbb481439),
	.w4(32'hbbd79cca),
	.w5(32'hb9effdd1),
	.w6(32'h3c959063),
	.w7(32'h3b3d3ef9),
	.w8(32'hb947f72e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1f9e),
	.w1(32'hbc1212ca),
	.w2(32'hbbff4c30),
	.w3(32'h3bfa8f48),
	.w4(32'h3bb85adc),
	.w5(32'hbc18138d),
	.w6(32'hbb961981),
	.w7(32'hbb072d89),
	.w8(32'h3bb569ed),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96089),
	.w1(32'h3c16be21),
	.w2(32'hbb2ee1a3),
	.w3(32'hbc700d80),
	.w4(32'h3a8003bb),
	.w5(32'hbbc04f0f),
	.w6(32'hbb70edcc),
	.w7(32'h39b4fa39),
	.w8(32'hba86418c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90c462),
	.w1(32'h3c697cc8),
	.w2(32'h3b9d53be),
	.w3(32'hbbdc0d29),
	.w4(32'hbc4e8e83),
	.w5(32'hba80588a),
	.w6(32'h3af86d9c),
	.w7(32'h3870fe2b),
	.w8(32'h3ac5d8b0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38494c1b),
	.w1(32'hbbb7125c),
	.w2(32'hbb05c891),
	.w3(32'h3b8073c8),
	.w4(32'h3bb02c8f),
	.w5(32'hbb909258),
	.w6(32'h3a709892),
	.w7(32'hbb571c3e),
	.w8(32'hba54ed4f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012c54),
	.w1(32'hbc8b817f),
	.w2(32'hbc6da7dc),
	.w3(32'h3c6455a5),
	.w4(32'h3ae97969),
	.w5(32'hbbc1da1a),
	.w6(32'h3b2ca5bf),
	.w7(32'hbbae5cc3),
	.w8(32'hbbb943b4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af65d9d),
	.w1(32'h3bbed767),
	.w2(32'h3bbae328),
	.w3(32'h3a320d9a),
	.w4(32'hbaa2ee29),
	.w5(32'hba9db987),
	.w6(32'h3a58f785),
	.w7(32'h3ac5dca4),
	.w8(32'h3b382471),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb299a),
	.w1(32'hbbb2d16e),
	.w2(32'hbb56d4ee),
	.w3(32'h3bbceacb),
	.w4(32'h3c04ccfe),
	.w5(32'h3bb5b75f),
	.w6(32'hbb15c84e),
	.w7(32'h3a3cbfd2),
	.w8(32'hbc84f011),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cefda),
	.w1(32'hbd02c87f),
	.w2(32'hbc96b23d),
	.w3(32'h3bcaac5c),
	.w4(32'hba96ba5c),
	.w5(32'hbc3da3c4),
	.w6(32'hbcae8df6),
	.w7(32'hbc75dbed),
	.w8(32'h3b9b50d5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c17e4),
	.w1(32'h3cd36c8b),
	.w2(32'h3c83dd97),
	.w3(32'hbcf1c614),
	.w4(32'hbc95d4a5),
	.w5(32'hbb97fcde),
	.w6(32'h3b367c9a),
	.w7(32'hb9beea21),
	.w8(32'h3c0a74bc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5017af),
	.w1(32'hbbe5e206),
	.w2(32'hbc713872),
	.w3(32'h3c922343),
	.w4(32'h3bba2d95),
	.w5(32'h3bc269d6),
	.w6(32'h3bf9d5f0),
	.w7(32'hbb81a739),
	.w8(32'h3b34cca4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade5850),
	.w1(32'hbb1e1427),
	.w2(32'h3694d660),
	.w3(32'hb96e0990),
	.w4(32'h3b352e2f),
	.w5(32'h3a77057b),
	.w6(32'hbb8e9126),
	.w7(32'hba810528),
	.w8(32'hbab30f5d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0067f9),
	.w1(32'hbb033ce7),
	.w2(32'h3a9900fa),
	.w3(32'hbc20184c),
	.w4(32'hba2f7276),
	.w5(32'h3a86fbfb),
	.w6(32'hbc3619a5),
	.w7(32'hb85b43d3),
	.w8(32'h3b7bbb36),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39076),
	.w1(32'h3b78ba05),
	.w2(32'h3bdee805),
	.w3(32'h3c328f83),
	.w4(32'hbac6eb4a),
	.w5(32'h3ba87b85),
	.w6(32'h3c1e69c7),
	.w7(32'hbb31f5a0),
	.w8(32'hba76782b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c7b6c),
	.w1(32'h3bb8e4f9),
	.w2(32'h3bd11fe3),
	.w3(32'h3b505737),
	.w4(32'h3c0a1bdc),
	.w5(32'h3b56e5f7),
	.w6(32'hbac6654d),
	.w7(32'hb9a1caf2),
	.w8(32'h3a715623),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d1f73),
	.w1(32'hba912ad6),
	.w2(32'hbb168649),
	.w3(32'h39d9c23d),
	.w4(32'h39b8d805),
	.w5(32'h3a859bb0),
	.w6(32'hb9c43448),
	.w7(32'hba7a74ae),
	.w8(32'h3abb537c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a295cc),
	.w1(32'h393a5787),
	.w2(32'h3ae5b103),
	.w3(32'h39a0d9cc),
	.w4(32'hba06378a),
	.w5(32'h3b68b108),
	.w6(32'h3ab097ed),
	.w7(32'hba365071),
	.w8(32'h3b2dac66),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063649),
	.w1(32'hbb40b076),
	.w2(32'hbb4ba155),
	.w3(32'hbbc5545d),
	.w4(32'h39e9b708),
	.w5(32'hbb110131),
	.w6(32'hbbdf822d),
	.w7(32'h3b0543c2),
	.w8(32'hbae80ce9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012674),
	.w1(32'hbb9850b0),
	.w2(32'h3698f152),
	.w3(32'hbc18fcad),
	.w4(32'hbb87e56b),
	.w5(32'h3b84b98f),
	.w6(32'hbc1a2260),
	.w7(32'hbb6f2f32),
	.w8(32'h3b67dda8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b784382),
	.w1(32'hbad51f16),
	.w2(32'h3b759fbd),
	.w3(32'h3b50713f),
	.w4(32'h3b216f22),
	.w5(32'h3b26d930),
	.w6(32'hbb23903f),
	.w7(32'h39592466),
	.w8(32'h3aed7e45),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a206f98),
	.w1(32'hb8d22305),
	.w2(32'h3a881558),
	.w3(32'h3b4a2507),
	.w4(32'h3a3696d3),
	.w5(32'h3bbb6a12),
	.w6(32'h3af33500),
	.w7(32'h3b0a57b0),
	.w8(32'h3b0f0372),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1e23),
	.w1(32'hba546b9d),
	.w2(32'h3b8285de),
	.w3(32'hba0c7154),
	.w4(32'h3ba33ccf),
	.w5(32'h3c6b05dc),
	.w6(32'hbb555e82),
	.w7(32'h3aa92e20),
	.w8(32'h3c290385),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29769f),
	.w1(32'h3b8db3df),
	.w2(32'h3b39124d),
	.w3(32'h3be63b34),
	.w4(32'h3bfb24ec),
	.w5(32'hb99ad287),
	.w6(32'h3b3a6a29),
	.w7(32'h38d21264),
	.w8(32'hba337ccd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09db5a),
	.w1(32'hbb693d83),
	.w2(32'hb99f55df),
	.w3(32'hb9a73fe8),
	.w4(32'hbb4fc903),
	.w5(32'hb9a4c9b2),
	.w6(32'hbbabdabe),
	.w7(32'hbaeca431),
	.w8(32'h391df094),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b66a),
	.w1(32'h3b0a67bb),
	.w2(32'h3a83ce98),
	.w3(32'h3af36b28),
	.w4(32'hb9fe70f7),
	.w5(32'h3a7419a8),
	.w6(32'h3b2b8357),
	.w7(32'h3a2e4abe),
	.w8(32'h39aee661),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7000b7),
	.w1(32'hba8bf78a),
	.w2(32'hbb0ecf26),
	.w3(32'hbb3d7cb5),
	.w4(32'hbb033809),
	.w5(32'h3ab5a572),
	.w6(32'hbbc38d9d),
	.w7(32'hbbb4acae),
	.w8(32'h3a012f67),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4533a3),
	.w1(32'hbb271e19),
	.w2(32'hbb31239b),
	.w3(32'hbaac6819),
	.w4(32'hba99dfca),
	.w5(32'h3aa135bd),
	.w6(32'hba923696),
	.w7(32'hbb02901b),
	.w8(32'hbb10edce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0252),
	.w1(32'hbb39fb8c),
	.w2(32'hbb2a26ff),
	.w3(32'h3896524d),
	.w4(32'hbb0d72fe),
	.w5(32'h3a4d31d7),
	.w6(32'hbaa50c44),
	.w7(32'hbb260350),
	.w8(32'h3aa66b43),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f2db7),
	.w1(32'h3b67ae9d),
	.w2(32'h3b890dbd),
	.w3(32'h3abe605b),
	.w4(32'h3b40cc95),
	.w5(32'hba134db9),
	.w6(32'h3b11ff65),
	.w7(32'h3aa23321),
	.w8(32'hbac730d1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26c81),
	.w1(32'h3afc2b0b),
	.w2(32'h3abed3d2),
	.w3(32'h3a3787aa),
	.w4(32'h3b20d26a),
	.w5(32'hba78d195),
	.w6(32'h3adde96c),
	.w7(32'h3b8c4948),
	.w8(32'h3b731316),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710665),
	.w1(32'hbad926b0),
	.w2(32'hba93259f),
	.w3(32'hbb160635),
	.w4(32'hb7a6b283),
	.w5(32'hbb67d0b4),
	.w6(32'h3b85bf37),
	.w7(32'h3ae98790),
	.w8(32'hbba6519b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac85ded),
	.w1(32'hbb4e136f),
	.w2(32'hbc00b2b4),
	.w3(32'hbb84c129),
	.w4(32'hbbe01247),
	.w5(32'h3c32030c),
	.w6(32'hbbb59ce6),
	.w7(32'hbc04b9e5),
	.w8(32'h3ba27823),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d78d2),
	.w1(32'h3a62f3fe),
	.w2(32'h3a8f79e6),
	.w3(32'h3bcc6fe4),
	.w4(32'h3bda5ed1),
	.w5(32'hb993b57c),
	.w6(32'h3b4b63f8),
	.w7(32'h3ab4cd23),
	.w8(32'hb903d5ba),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae23952),
	.w1(32'hbb0ebf6d),
	.w2(32'hbb37fd2b),
	.w3(32'hbad9cdec),
	.w4(32'hba63a86b),
	.w5(32'h3a654e5f),
	.w6(32'h3a335e2e),
	.w7(32'hbab04489),
	.w8(32'h3a9aaf80),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3d962),
	.w1(32'h3b2283c4),
	.w2(32'h3a13a635),
	.w3(32'hbb1d930e),
	.w4(32'hba0437f1),
	.w5(32'h3931b1bf),
	.w6(32'hbb01bbc4),
	.w7(32'hba6870a8),
	.w8(32'h3adfac71),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee19fc),
	.w1(32'h3b5ef459),
	.w2(32'h3bac0a50),
	.w3(32'hbb9b8f76),
	.w4(32'hb9bf8229),
	.w5(32'h3933b5b9),
	.w6(32'hbbab964b),
	.w7(32'hbb6988d9),
	.w8(32'hbb771358),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77265c),
	.w1(32'hbbac4cf4),
	.w2(32'hbb7aa38b),
	.w3(32'hbb9a8a80),
	.w4(32'hbb3ddbf3),
	.w5(32'hbad838cc),
	.w6(32'hbbf6c3a7),
	.w7(32'hbba28e83),
	.w8(32'h3b2901b0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a49f50),
	.w1(32'hba17e35f),
	.w2(32'h3993c416),
	.w3(32'hbacbb7f5),
	.w4(32'h3aa54fd7),
	.w5(32'h3a810c98),
	.w6(32'hb9da26c4),
	.w7(32'hbaf66f9a),
	.w8(32'h349354f3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f9110),
	.w1(32'hbacf368a),
	.w2(32'hbab1b5ca),
	.w3(32'hb9fef0a2),
	.w4(32'hbb4624ec),
	.w5(32'h3bc0ed37),
	.w6(32'hbafd9fc0),
	.w7(32'hbb168db9),
	.w8(32'h3b9861b5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f229a),
	.w1(32'h39ba2d3c),
	.w2(32'hba84b9c9),
	.w3(32'h3b064f9c),
	.w4(32'h3b2fa271),
	.w5(32'h3b1e1072),
	.w6(32'h3aec9b4a),
	.w7(32'h3ac341c8),
	.w8(32'h3a655946),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16c813),
	.w1(32'hba3c32cf),
	.w2(32'hbb4dbc11),
	.w3(32'h3a4016c9),
	.w4(32'h39b113bf),
	.w5(32'h3bcf6515),
	.w6(32'hbad21a9d),
	.w7(32'hb9a14d48),
	.w8(32'h3ba5f433),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8c467),
	.w1(32'h3b9706cf),
	.w2(32'hb65b0b16),
	.w3(32'h3b8a671e),
	.w4(32'h3bc461ee),
	.w5(32'hbb16b4d6),
	.w6(32'h3b866ed5),
	.w7(32'hb85ca93f),
	.w8(32'hb9825144),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad14331),
	.w1(32'hba9eed88),
	.w2(32'hbb81c63d),
	.w3(32'hbabfa501),
	.w4(32'hbb278c51),
	.w5(32'hbb841272),
	.w6(32'h3aba0a70),
	.w7(32'hba684a88),
	.w8(32'hba932db8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad99298),
	.w1(32'hb9a1c49a),
	.w2(32'h3a78ea1c),
	.w3(32'hbb5e1ac1),
	.w4(32'h3a458510),
	.w5(32'hbabd9398),
	.w6(32'h3a96583f),
	.w7(32'h39898526),
	.w8(32'hbae9e4ff),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bb8f6),
	.w1(32'hbb7423a9),
	.w2(32'hbb81b7db),
	.w3(32'hbb5681f1),
	.w4(32'hbb13d0bf),
	.w5(32'h3b502c7d),
	.w6(32'hbb89a1eb),
	.w7(32'hbb4ecef0),
	.w8(32'hbb317ba9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdafc7a),
	.w1(32'h3bdce77a),
	.w2(32'h3bcdd1a1),
	.w3(32'hba434b29),
	.w4(32'h3b399baf),
	.w5(32'h3bd18a4a),
	.w6(32'hbbed0d2d),
	.w7(32'hbb927189),
	.w8(32'h3bb77cf0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba0361),
	.w1(32'h3bbef08f),
	.w2(32'h3b2117d5),
	.w3(32'h3badf72d),
	.w4(32'h3ba36f68),
	.w5(32'h3b2ee3eb),
	.w6(32'h3aaa50b7),
	.w7(32'h3980935a),
	.w8(32'h3a908aef),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f0958),
	.w1(32'h3af773f5),
	.w2(32'hbaf55349),
	.w3(32'h38f18e57),
	.w4(32'h3b71d787),
	.w5(32'h3a9fe530),
	.w6(32'hb9c67340),
	.w7(32'h3b79ecd5),
	.w8(32'hba4ac585),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b7051),
	.w1(32'h3bea9997),
	.w2(32'h3b3276c5),
	.w3(32'h3af65dd3),
	.w4(32'h3b61bf70),
	.w5(32'h3a58ab83),
	.w6(32'hb9af6de6),
	.w7(32'h3ab4d360),
	.w8(32'hbb41c387),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37907e),
	.w1(32'hbaa3f63e),
	.w2(32'hba33c2a5),
	.w3(32'hbb60465c),
	.w4(32'hbaba46dc),
	.w5(32'h3c13b11b),
	.w6(32'hbbf5ecd6),
	.w7(32'hbb602828),
	.w8(32'h3bbba3e3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96f057),
	.w1(32'h3b7490f7),
	.w2(32'hbab98af6),
	.w3(32'h3ba06be8),
	.w4(32'h3bc5f659),
	.w5(32'h39d5f769),
	.w6(32'h3a8c0d62),
	.w7(32'h3acdf66f),
	.w8(32'h3aa8c433),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5ef9b),
	.w1(32'h3ae6f87e),
	.w2(32'h3a81943f),
	.w3(32'hbb0ae2c6),
	.w4(32'hb9182334),
	.w5(32'h3b8d4b9d),
	.w6(32'hbb04a163),
	.w7(32'hbad2583a),
	.w8(32'h3b749cb3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba225de),
	.w1(32'h3a5f95cf),
	.w2(32'h3b0e160c),
	.w3(32'h3b3ad9fb),
	.w4(32'h3a7f18aa),
	.w5(32'hbaf32fbd),
	.w6(32'h3b009d87),
	.w7(32'hba34cbf5),
	.w8(32'hbb6ac27a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa4d04),
	.w1(32'hbafca7dc),
	.w2(32'hba4e01ab),
	.w3(32'hbb908d61),
	.w4(32'hbb241e36),
	.w5(32'hbaad5e0a),
	.w6(32'hbbf729de),
	.w7(32'hbb6c1705),
	.w8(32'hbb1cb153),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b9fb),
	.w1(32'h39e22456),
	.w2(32'h3b5ab6ba),
	.w3(32'hbac7d13a),
	.w4(32'hbb457c4f),
	.w5(32'h3a99452e),
	.w6(32'hb98342bf),
	.w7(32'hbaa7178f),
	.w8(32'hbaa7fc37),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7986),
	.w1(32'hbb4bc396),
	.w2(32'hbb0a8f4d),
	.w3(32'hbb472bc7),
	.w4(32'hbaf0028a),
	.w5(32'h3a7c0e95),
	.w6(32'hbbd14537),
	.w7(32'hbb00e495),
	.w8(32'h3b9d14f6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfe834),
	.w1(32'h3b8a58e3),
	.w2(32'hbad66f8a),
	.w3(32'h38e9814c),
	.w4(32'h3a4ac666),
	.w5(32'h3b53da33),
	.w6(32'h3af9068f),
	.w7(32'hbb0d2379),
	.w8(32'h39226fea),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fccd4),
	.w1(32'h3a1fe163),
	.w2(32'h3ab21aec),
	.w3(32'h3b3a9b78),
	.w4(32'h3ae48cc0),
	.w5(32'hbaaecad9),
	.w6(32'h398dbbe3),
	.w7(32'h3aac2987),
	.w8(32'hbb0245a8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b54fb),
	.w1(32'h3aa86d70),
	.w2(32'h3b4618f1),
	.w3(32'hbb3afb94),
	.w4(32'hbae7247f),
	.w5(32'hb965b506),
	.w6(32'hbb0ba9bb),
	.w7(32'hba5c31d1),
	.w8(32'h3b611d9f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5105e),
	.w1(32'hbace626d),
	.w2(32'h3afe717e),
	.w3(32'hbb3a33af),
	.w4(32'hbaec793b),
	.w5(32'h3b63b41b),
	.w6(32'h3976b4ba),
	.w7(32'h3b0ed042),
	.w8(32'h3b938041),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fd8ed),
	.w1(32'h3aa97a7b),
	.w2(32'h3a92fc41),
	.w3(32'hbb25802e),
	.w4(32'hba987c0d),
	.w5(32'h3b8fe6c4),
	.w6(32'hbb401762),
	.w7(32'hb931e068),
	.w8(32'h3bce4cc5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66bbe3),
	.w1(32'h3a7ad076),
	.w2(32'hbb17b396),
	.w3(32'hbb26b9ff),
	.w4(32'hbb0d7be7),
	.w5(32'h3bb93944),
	.w6(32'h39efe729),
	.w7(32'hbb5dda76),
	.w8(32'h3b9f29dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c5ca3),
	.w1(32'h3b8823e7),
	.w2(32'h3b0a7969),
	.w3(32'h3bcfa213),
	.w4(32'h3c0bc6d0),
	.w5(32'h3b898ff8),
	.w6(32'h3bbafb96),
	.w7(32'h3bc8d04a),
	.w8(32'h3b4f6ef4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37fd67),
	.w1(32'h3a98b00f),
	.w2(32'h388de795),
	.w3(32'h3b02e81f),
	.w4(32'h3ab96799),
	.w5(32'h39f1a419),
	.w6(32'h3a8b89b7),
	.w7(32'hbaea1d8c),
	.w8(32'h3b87311d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a098f),
	.w1(32'h3b2f2127),
	.w2(32'hbb8c3255),
	.w3(32'hbaa31967),
	.w4(32'h3a050e65),
	.w5(32'h3aa02469),
	.w6(32'hbabb85a7),
	.w7(32'hbb74fde8),
	.w8(32'h3b855e13),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42b948),
	.w1(32'h3ae02047),
	.w2(32'h3aa8c14f),
	.w3(32'hb8f0eaf4),
	.w4(32'hb9154c50),
	.w5(32'h3b05390d),
	.w6(32'h3b2c16a5),
	.w7(32'h3a2f3ee1),
	.w8(32'h3a86e6ef),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fe7b1),
	.w1(32'h3af61be3),
	.w2(32'h3aeb8b14),
	.w3(32'h3b54011d),
	.w4(32'h38b29e91),
	.w5(32'h3b72ac84),
	.w6(32'h3a21524f),
	.w7(32'h3b3e0268),
	.w8(32'h3b652b44),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30c476),
	.w1(32'h3b3239eb),
	.w2(32'h3b602026),
	.w3(32'h3ad128be),
	.w4(32'h3b0afcdb),
	.w5(32'h3bfbae9d),
	.w6(32'h3b787e34),
	.w7(32'h3b8fea7d),
	.w8(32'h3b790e0e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175bc6),
	.w1(32'h3b5377ab),
	.w2(32'h3ac8ea3f),
	.w3(32'h3bb1c412),
	.w4(32'h3b8d13f6),
	.w5(32'hbad26196),
	.w6(32'h3aab5635),
	.w7(32'hbaed5836),
	.w8(32'hba816d75),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5df866),
	.w1(32'h3a50ff1c),
	.w2(32'h3a3af799),
	.w3(32'h39804829),
	.w4(32'hbb64b1d1),
	.w5(32'h3a5be366),
	.w6(32'h3af600b8),
	.w7(32'hba3dc87a),
	.w8(32'h3ad8e966),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69484e),
	.w1(32'h3b320a62),
	.w2(32'h3a9138ff),
	.w3(32'hb9bf6f54),
	.w4(32'hba1c0a8a),
	.w5(32'h3abb8728),
	.w6(32'h3a981f01),
	.w7(32'hba8007f7),
	.w8(32'h3b96907c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5512fc),
	.w1(32'h3c29a87b),
	.w2(32'h3c143bca),
	.w3(32'h3b63d71f),
	.w4(32'h3ba8e293),
	.w5(32'h393b0fb7),
	.w6(32'h3b2baab0),
	.w7(32'h3bab3cb6),
	.w8(32'h3a7d2551),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbb0d),
	.w1(32'h3ab07227),
	.w2(32'h3b0b5ba5),
	.w3(32'h3b466ee4),
	.w4(32'h3b3a5fc7),
	.w5(32'h3bc5c147),
	.w6(32'h3b9a0204),
	.w7(32'h3b153286),
	.w8(32'h3b7d0227),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03fecf),
	.w1(32'h3bba4770),
	.w2(32'h3bd2309b),
	.w3(32'h3b81e635),
	.w4(32'h3c0102b8),
	.w5(32'hbb926582),
	.w6(32'hbabf14a1),
	.w7(32'h3c06fa3d),
	.w8(32'hbb9cc73f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c6475),
	.w1(32'hbb284a76),
	.w2(32'hbac39f85),
	.w3(32'hbb110e99),
	.w4(32'hbb0ad882),
	.w5(32'h3afb5904),
	.w6(32'hbb6d6a8e),
	.w7(32'hbafd72fc),
	.w8(32'h3b23af1c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b0b95),
	.w1(32'hb9d9909c),
	.w2(32'hbb124494),
	.w3(32'h3a0ca135),
	.w4(32'hbb60a95a),
	.w5(32'hbbb295d4),
	.w6(32'h3b3e2ad2),
	.w7(32'h3a2ed611),
	.w8(32'hbbb40cb0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061fd8),
	.w1(32'hba634a95),
	.w2(32'hba8e0fa9),
	.w3(32'hbb9c8d41),
	.w4(32'hbabc1d3d),
	.w5(32'h3aed7e5b),
	.w6(32'hbb5c38b5),
	.w7(32'hbabcae30),
	.w8(32'h3a916426),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13b2d3),
	.w1(32'h3b9d7c3a),
	.w2(32'h3b80acbd),
	.w3(32'h398d2687),
	.w4(32'h3a9ce3e9),
	.w5(32'h3bd071c7),
	.w6(32'h3b10b887),
	.w7(32'h3b3ff41f),
	.w8(32'h3c2a3129),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57d89e),
	.w1(32'h3bb49cf3),
	.w2(32'h3af656c4),
	.w3(32'h3b9edb0d),
	.w4(32'h3b21071c),
	.w5(32'hbadf34e3),
	.w6(32'h3c1759af),
	.w7(32'h3b06cda2),
	.w8(32'hbac07b9b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad111d),
	.w1(32'hba39348a),
	.w2(32'hba8df6b9),
	.w3(32'h3a414081),
	.w4(32'h3b055d33),
	.w5(32'hb8bf1df0),
	.w6(32'hbb135363),
	.w7(32'hbae8b775),
	.w8(32'h3aea6646),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f68e1),
	.w1(32'hba8e9866),
	.w2(32'hb9e0fb95),
	.w3(32'h3ba90f51),
	.w4(32'h39d1ff7f),
	.w5(32'hba54c68a),
	.w6(32'h3bddd477),
	.w7(32'h3b09424c),
	.w8(32'hbb06364f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b7ea7),
	.w1(32'hbb8bcdf9),
	.w2(32'hbb7129e5),
	.w3(32'hb8e83b1e),
	.w4(32'hba81f51f),
	.w5(32'h3ba98d73),
	.w6(32'hbb22ce71),
	.w7(32'hbb63a8df),
	.w8(32'h3a947751),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77560ca),
	.w1(32'h3a0c79dc),
	.w2(32'hba38afe2),
	.w3(32'h3b658295),
	.w4(32'h3b20311c),
	.w5(32'h3af8c136),
	.w6(32'h3b2f6eec),
	.w7(32'h3b39b8ab),
	.w8(32'h3b7fb7ee),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8ff12),
	.w1(32'h3a9a32e1),
	.w2(32'h3af37690),
	.w3(32'h3a505654),
	.w4(32'h3a288f40),
	.w5(32'hba19c455),
	.w6(32'h3af1747b),
	.w7(32'hba6ac257),
	.w8(32'h3ad4cb35),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824e6c),
	.w1(32'h3b166f93),
	.w2(32'h3a79a975),
	.w3(32'h39252e91),
	.w4(32'h3b1f9ee0),
	.w5(32'hbb03945e),
	.w6(32'h3aaab14c),
	.w7(32'h3b657ec9),
	.w8(32'hbb637377),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc636b2d),
	.w1(32'hbbd8716c),
	.w2(32'hbc1d0e98),
	.w3(32'hbb93685a),
	.w4(32'hb9eb5faa),
	.w5(32'h3bd92a73),
	.w6(32'hbb40c4be),
	.w7(32'hba515a70),
	.w8(32'h3bab62a8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393388ac),
	.w1(32'hbad6a4b0),
	.w2(32'h3b36ba40),
	.w3(32'h3a4505da),
	.w4(32'h3ac42873),
	.w5(32'h3b9ac060),
	.w6(32'hbad852c1),
	.w7(32'h3b586776),
	.w8(32'h3b2fc53d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1b278),
	.w1(32'hba4c7bd5),
	.w2(32'h3ae59d23),
	.w3(32'h3b82d00c),
	.w4(32'h3b89c2d8),
	.w5(32'h3b933bcb),
	.w6(32'hba4db429),
	.w7(32'h3b393811),
	.w8(32'h3b0e00f0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153ce4),
	.w1(32'h3a75cb2e),
	.w2(32'h39d6e335),
	.w3(32'h3b075637),
	.w4(32'h3b2a8ff6),
	.w5(32'hbb7c418a),
	.w6(32'hb919a000),
	.w7(32'h37d59605),
	.w8(32'hbb2f5b41),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b450d),
	.w1(32'hbb4db556),
	.w2(32'hbb99b71a),
	.w3(32'hbb42afd8),
	.w4(32'hbb002229),
	.w5(32'h3bdb646b),
	.w6(32'hbb433e44),
	.w7(32'hbb607ae3),
	.w8(32'h3b912bc9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb85a37),
	.w1(32'h3bb0b24e),
	.w2(32'h3b18dbec),
	.w3(32'h3bd02ebc),
	.w4(32'h3bd2178e),
	.w5(32'h3b39914b),
	.w6(32'h3bf76315),
	.w7(32'h3ba79ec0),
	.w8(32'hbac0d634),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb8e32),
	.w1(32'h39c0a734),
	.w2(32'h3b9b0bc8),
	.w3(32'h3b0e8c8a),
	.w4(32'h3b45ab67),
	.w5(32'hbb43c5f8),
	.w6(32'hbba77837),
	.w7(32'hb902fb2a),
	.w8(32'hba016c8f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4664),
	.w1(32'hbac7e6c7),
	.w2(32'hbb0f7ec4),
	.w3(32'hbad9b389),
	.w4(32'hbb358d8f),
	.w5(32'hbb68bf52),
	.w6(32'h3aa3563e),
	.w7(32'hba8cccf0),
	.w8(32'hba5eb834),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6911c59),
	.w1(32'h3a524fe8),
	.w2(32'h3a8a315c),
	.w3(32'hbb4da140),
	.w4(32'h3b1f7eca),
	.w5(32'h3a39fcf7),
	.w6(32'hb84939ce),
	.w7(32'h3afe362d),
	.w8(32'h3a8511ef),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5c87),
	.w1(32'hbb073b02),
	.w2(32'h3a3dfa1a),
	.w3(32'h3a2bce52),
	.w4(32'hbb80d3fa),
	.w5(32'h3b626bcb),
	.w6(32'h3aac8738),
	.w7(32'hbb3a439d),
	.w8(32'h3b5b7faf),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ea91a),
	.w1(32'h3af58c65),
	.w2(32'h3ad05ac6),
	.w3(32'h3afead85),
	.w4(32'hba0599fd),
	.w5(32'hba200b0e),
	.w6(32'h3abad699),
	.w7(32'h39a45917),
	.w8(32'h3a9bd4b0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2a4bd),
	.w1(32'hba56a560),
	.w2(32'hbb371e7c),
	.w3(32'hbb84dbc9),
	.w4(32'hbb8e00aa),
	.w5(32'h3a49453f),
	.w6(32'hba9d2bc1),
	.w7(32'hbb23d72f),
	.w8(32'hbabc738c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17f1f0),
	.w1(32'hbb16f7e2),
	.w2(32'hbab8bd2e),
	.w3(32'hbb30a99d),
	.w4(32'hbae0e1fa),
	.w5(32'h3ac943e3),
	.w6(32'hbb436198),
	.w7(32'hbb1701cd),
	.w8(32'h3b23bea9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6553fc),
	.w1(32'h3b09f18f),
	.w2(32'hb9bd903d),
	.w3(32'h39df3dc2),
	.w4(32'hb9d1159c),
	.w5(32'h3bb2b465),
	.w6(32'h3b249192),
	.w7(32'hbac999bf),
	.w8(32'h3b16141a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b481d10),
	.w1(32'h3bb1b067),
	.w2(32'h3ae864cb),
	.w3(32'h3bb62970),
	.w4(32'h3baf6c0a),
	.w5(32'h3b166249),
	.w6(32'h3bae2b5f),
	.w7(32'h3b917ebb),
	.w8(32'hba3ef7b5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93e575),
	.w1(32'hba96e0a6),
	.w2(32'h3b9ad1a2),
	.w3(32'hbc102527),
	.w4(32'h3c0bafc5),
	.w5(32'h3be3b69b),
	.w6(32'hbbc44548),
	.w7(32'h3c1a4a63),
	.w8(32'h3bd35fb6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c8b0),
	.w1(32'hb8cf97b5),
	.w2(32'h3ac86748),
	.w3(32'h3b72fcc8),
	.w4(32'h38b5178c),
	.w5(32'h3b77d171),
	.w6(32'hba6406a5),
	.w7(32'hbb127721),
	.w8(32'hb8ffa5b2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4ffd7),
	.w1(32'h38b222b4),
	.w2(32'h3a36ceec),
	.w3(32'hb8a400d7),
	.w4(32'h3a94c297),
	.w5(32'h3b5ca07b),
	.w6(32'hbb36bc14),
	.w7(32'h3ad1c625),
	.w8(32'h3b1e7efa),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf97cf),
	.w1(32'h3b26ca86),
	.w2(32'h3b040d3a),
	.w3(32'h3b32e171),
	.w4(32'h3b2ae053),
	.w5(32'h3a503c6f),
	.w6(32'h3aa10298),
	.w7(32'h3a67ef7c),
	.w8(32'hb9cdf925),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38894274),
	.w1(32'hb9b16265),
	.w2(32'hbabdba58),
	.w3(32'h377f6156),
	.w4(32'hbafd4a6e),
	.w5(32'h396651e2),
	.w6(32'hb8830201),
	.w7(32'hbae01d43),
	.w8(32'hba13802d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877bb0),
	.w1(32'hbb423ed7),
	.w2(32'hbb95e228),
	.w3(32'hbb3114d3),
	.w4(32'hbb8575ae),
	.w5(32'h3b078548),
	.w6(32'hbb49ce4b),
	.w7(32'hbb88f521),
	.w8(32'h3b234820),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1ead1),
	.w1(32'h3a8e695f),
	.w2(32'h3a213647),
	.w3(32'h3b302de3),
	.w4(32'h3a8e9918),
	.w5(32'h3af35f40),
	.w6(32'h3aa49a3b),
	.w7(32'hba842b5a),
	.w8(32'h3ae514ff),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4e1d1),
	.w1(32'h3b4bb1ea),
	.w2(32'hba278b64),
	.w3(32'hb98e8216),
	.w4(32'hbae8929e),
	.w5(32'hba92c641),
	.w6(32'hbaaba249),
	.w7(32'hbb46f4d9),
	.w8(32'hbb97c46c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5740e8),
	.w1(32'hbb98d0f4),
	.w2(32'hbb9986dc),
	.w3(32'hbbc4d58c),
	.w4(32'hbab511e8),
	.w5(32'h3badda6f),
	.w6(32'hbc22d9b8),
	.w7(32'hbba8f1b3),
	.w8(32'h3b97f108),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23925a),
	.w1(32'h3b7b0675),
	.w2(32'hb7173119),
	.w3(32'hb97ed112),
	.w4(32'h39b63eb4),
	.w5(32'hbb912074),
	.w6(32'h3b0cd2e0),
	.w7(32'h3a4e592a),
	.w8(32'hbbeba60f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb400a2),
	.w1(32'hbb6b6e09),
	.w2(32'hbb083e1a),
	.w3(32'hbb9531d2),
	.w4(32'hbacf4ebf),
	.w5(32'h3b34435a),
	.w6(32'hbbe1c2b5),
	.w7(32'hbb8d8c71),
	.w8(32'h3b0a2fba),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799ad8),
	.w1(32'hbaa68c65),
	.w2(32'hba88d696),
	.w3(32'hbb8943f1),
	.w4(32'hba8ea19b),
	.w5(32'h3b43b232),
	.w6(32'hba4b4732),
	.w7(32'h3a21a5c1),
	.w8(32'h3b9222af),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb1cd),
	.w1(32'h3b716ba3),
	.w2(32'h3a130210),
	.w3(32'h3b8abfc6),
	.w4(32'h3bccabcc),
	.w5(32'h3a5b5b86),
	.w6(32'h3ba52fd1),
	.w7(32'h3b91ba8e),
	.w8(32'h3b2aad13),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a35b6),
	.w1(32'h3aa7905e),
	.w2(32'hbb128612),
	.w3(32'h3acf9548),
	.w4(32'h3b098bb3),
	.w5(32'hbb51de6f),
	.w6(32'h3b8466b3),
	.w7(32'h3b203497),
	.w8(32'hbb432cd2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad365),
	.w1(32'hba0454ae),
	.w2(32'hba580674),
	.w3(32'hb824fd44),
	.w4(32'h3a14bfbf),
	.w5(32'h3b4d7f0c),
	.w6(32'hbaa7e288),
	.w7(32'hb90ac339),
	.w8(32'h3b80e018),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a4d2),
	.w1(32'h3a9fbf8e),
	.w2(32'h39bc13d1),
	.w3(32'hbbe36367),
	.w4(32'hbb49f9ba),
	.w5(32'hbab626e4),
	.w6(32'hbbbcd6da),
	.w7(32'hba9fc369),
	.w8(32'hba9ad585),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaced5f7),
	.w1(32'hbb613722),
	.w2(32'h3adbce44),
	.w3(32'hbb55efdd),
	.w4(32'hbb770b79),
	.w5(32'h3b21a892),
	.w6(32'hbba6ee98),
	.w7(32'hbb8ec5eb),
	.w8(32'h3a80d101),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9cf9),
	.w1(32'h37c86183),
	.w2(32'hb8137266),
	.w3(32'h3ad2716e),
	.w4(32'h3a356cfb),
	.w5(32'hba030f73),
	.w6(32'h3aded2f8),
	.w7(32'hbaa99dcc),
	.w8(32'hbb67c434),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf788),
	.w1(32'hbae43b56),
	.w2(32'hbb0925c0),
	.w3(32'hbafd98ae),
	.w4(32'hbb41d74d),
	.w5(32'hbad373d7),
	.w6(32'hbb78e9f4),
	.w7(32'hbb950d2e),
	.w8(32'hbb124dcb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48fd92),
	.w1(32'hbb0863ed),
	.w2(32'h3a804973),
	.w3(32'hbb608907),
	.w4(32'hbae451f6),
	.w5(32'h3b0d4cfd),
	.w6(32'hbb873a07),
	.w7(32'hbb033cee),
	.w8(32'hba2d944e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b305),
	.w1(32'hbaf3cf30),
	.w2(32'hba4e8790),
	.w3(32'hbb4f8eae),
	.w4(32'hb6fde11a),
	.w5(32'hbb30d1e5),
	.w6(32'hbbe7a855),
	.w7(32'hbb6c8f43),
	.w8(32'hbb1f11ee),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2111e2),
	.w1(32'hbb7314c1),
	.w2(32'hbb3a2d84),
	.w3(32'hbc3562ad),
	.w4(32'h3a9e4112),
	.w5(32'h3b9bce34),
	.w6(32'hbc22605b),
	.w7(32'hbb1f73e3),
	.w8(32'h3b0bcbc8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a944f),
	.w1(32'hba9560da),
	.w2(32'hba63bc3d),
	.w3(32'hbab1ff27),
	.w4(32'hbac29bc2),
	.w5(32'hbae5edc9),
	.w6(32'hba9ac10d),
	.w7(32'hbaeabae7),
	.w8(32'h3a77e386),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b2d1),
	.w1(32'h3b142630),
	.w2(32'h3af8a46c),
	.w3(32'hb8886fca),
	.w4(32'h3b6dc48d),
	.w5(32'hbb0c8cad),
	.w6(32'h3b14048a),
	.w7(32'h3b1b4869),
	.w8(32'h39a61152),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba3658),
	.w1(32'hbae79d08),
	.w2(32'hbaa32d1a),
	.w3(32'hbbbc68ed),
	.w4(32'hbb941676),
	.w5(32'hba8b22f5),
	.w6(32'hbbb9d4b6),
	.w7(32'hbba76873),
	.w8(32'h397b3446),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ce6bc),
	.w1(32'h39a64a4b),
	.w2(32'hbaaf3ff1),
	.w3(32'hbb7d74f3),
	.w4(32'hbaa5ebd4),
	.w5(32'h3b464c09),
	.w6(32'hbb182f18),
	.w7(32'hbb3139bd),
	.w8(32'h3b75492b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83764bb),
	.w1(32'h3ac27b37),
	.w2(32'h3bc1e242),
	.w3(32'hb891558f),
	.w4(32'h3bdf2a19),
	.w5(32'h3bc1a29b),
	.w6(32'hbab9907f),
	.w7(32'h3b98e196),
	.w8(32'h3b708aa6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbabe34),
	.w1(32'h3a00476e),
	.w2(32'h3b882b27),
	.w3(32'h3b84ded6),
	.w4(32'h3abd0a64),
	.w5(32'h3b3d16f5),
	.w6(32'h3b501715),
	.w7(32'h3aaba677),
	.w8(32'h3a5f2f41),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360fa1b8),
	.w1(32'hba13c30a),
	.w2(32'hb955f9e9),
	.w3(32'h3b298029),
	.w4(32'hba05a641),
	.w5(32'h3b648bcb),
	.w6(32'hb9b04513),
	.w7(32'hbafa56b4),
	.w8(32'hb9a4031e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afea13a),
	.w1(32'h3b108188),
	.w2(32'h3abf8035),
	.w3(32'h3b1fe833),
	.w4(32'h3b277a9c),
	.w5(32'hb9e5f39f),
	.w6(32'hb92e79b0),
	.w7(32'h3b042276),
	.w8(32'hb90cfab5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f30e3),
	.w1(32'h3adc2cfc),
	.w2(32'h3aad3fbd),
	.w3(32'hbb193078),
	.w4(32'h3abc6acd),
	.w5(32'hba0ae0b0),
	.w6(32'hbb371a7b),
	.w7(32'hbac4a7ac),
	.w8(32'h3aab6671),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb911b2),
	.w1(32'hb99c1a50),
	.w2(32'hbb7d1693),
	.w3(32'hbbeeef1f),
	.w4(32'h3b227383),
	.w5(32'h3bcbf4a9),
	.w6(32'hbbeff2fe),
	.w7(32'h3b1d0f2f),
	.w8(32'h3bcfaaf1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0d8a),
	.w1(32'h3a453f42),
	.w2(32'h3a89379b),
	.w3(32'hbbc51983),
	.w4(32'h3a8ffcdd),
	.w5(32'h3ab72825),
	.w6(32'hbbc076f6),
	.w7(32'h3acaacc8),
	.w8(32'hba8b2a3a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64dc35),
	.w1(32'h3bb9cdbc),
	.w2(32'h3a6cd789),
	.w3(32'h3a0b228d),
	.w4(32'hba0b860b),
	.w5(32'hbb2da2f4),
	.w6(32'h3ae693a4),
	.w7(32'hba4fc687),
	.w8(32'hba3a0150),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac03f08),
	.w1(32'h3ad77cff),
	.w2(32'hbbde512f),
	.w3(32'hbaa025c7),
	.w4(32'hbc00f27c),
	.w5(32'h3bb611d3),
	.w6(32'h3b6db97c),
	.w7(32'hbbc2ce0b),
	.w8(32'h3c14ed94),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be031ff),
	.w1(32'h3c233dfc),
	.w2(32'h3b1790ac),
	.w3(32'h3bafe9c5),
	.w4(32'h3ba9dd12),
	.w5(32'h395048cc),
	.w6(32'h3c138dc2),
	.w7(32'h3b71162e),
	.w8(32'h3b1a1bc1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b634e55),
	.w1(32'h3bc7b29e),
	.w2(32'h3bb1c188),
	.w3(32'h3aafaf41),
	.w4(32'h3af54592),
	.w5(32'hbb448cdc),
	.w6(32'h3b6cbd7b),
	.w7(32'h3925b45a),
	.w8(32'hbb001278),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83c3c0),
	.w1(32'hbb6a27f3),
	.w2(32'hbb1aa94a),
	.w3(32'hbb10f353),
	.w4(32'hbacce3bb),
	.w5(32'h3b944c33),
	.w6(32'hbb7d8e3f),
	.w7(32'hbb50ae77),
	.w8(32'h3b4592ba),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa84c97),
	.w1(32'h3b8a6190),
	.w2(32'h3b8eb69e),
	.w3(32'h3afe532f),
	.w4(32'h3b31612e),
	.w5(32'h3aefeb43),
	.w6(32'h3a2f9ebd),
	.w7(32'h3bdc7bb7),
	.w8(32'h3a46b01d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc4a53),
	.w1(32'h3b6b47ad),
	.w2(32'h3bad1b3e),
	.w3(32'h3afc890a),
	.w4(32'h3bddded9),
	.w5(32'hbbb2f81a),
	.w6(32'h3bac9689),
	.w7(32'h3bee71f7),
	.w8(32'hbb979b94),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe86087),
	.w1(32'hbc46e662),
	.w2(32'hbc0d3803),
	.w3(32'hbc0f53c0),
	.w4(32'hbbf0d95e),
	.w5(32'hbba8abbd),
	.w6(32'hbbfc1af8),
	.w7(32'hbbd986e4),
	.w8(32'hbb381b82),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3beb32),
	.w1(32'h3b5159f4),
	.w2(32'hbb6e46e2),
	.w3(32'h3b6b5d41),
	.w4(32'hbb9b8f26),
	.w5(32'hba6e7cb5),
	.w6(32'h3c462280),
	.w7(32'h3a450fe9),
	.w8(32'h3a8c2696),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a9de),
	.w1(32'h3ae03b6c),
	.w2(32'h3b2ade90),
	.w3(32'h3b84383f),
	.w4(32'h3c0c2a9c),
	.w5(32'hbb6203a4),
	.w6(32'h3b09760e),
	.w7(32'h3b1cb45b),
	.w8(32'hbbbf469c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa6c96),
	.w1(32'h385fc2cf),
	.w2(32'hbbea39d1),
	.w3(32'hbbe6bba0),
	.w4(32'h3b058fe6),
	.w5(32'h3b4a2041),
	.w6(32'hbbe60898),
	.w7(32'hbad08fb9),
	.w8(32'hbb96fcc8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93aa6),
	.w1(32'hbc394de5),
	.w2(32'hbbafcef4),
	.w3(32'hbc0913b8),
	.w4(32'hbaf711fc),
	.w5(32'h3b1268a0),
	.w6(32'hbc5f6e61),
	.w7(32'hbc277088),
	.w8(32'hbb940ed6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a98c2),
	.w1(32'hbb1915c0),
	.w2(32'hbc1dceda),
	.w3(32'h3bd570cb),
	.w4(32'hbbd21fc2),
	.w5(32'hbc0d9291),
	.w6(32'h3b6486ef),
	.w7(32'hbc0b0c7a),
	.w8(32'hbb74c6f0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc347e0e),
	.w1(32'hbb9c0ebd),
	.w2(32'hbbbf012c),
	.w3(32'hbbed7703),
	.w4(32'hbbf4ce30),
	.w5(32'hbb678d28),
	.w6(32'h3b38bfa3),
	.w7(32'hbb6446cc),
	.w8(32'hbc0bf517),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc007772),
	.w1(32'hbaf84cf6),
	.w2(32'hbaca40ea),
	.w3(32'hbc5fb88a),
	.w4(32'hba0b85f6),
	.w5(32'hb9287c0c),
	.w6(32'hbb7c16b6),
	.w7(32'h3b6713cd),
	.w8(32'h3b16afef),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec369b),
	.w1(32'h3b07e8ec),
	.w2(32'hba19a922),
	.w3(32'h3a1f4313),
	.w4(32'hbb3bc504),
	.w5(32'hbba82639),
	.w6(32'h3c001333),
	.w7(32'h3b90abcd),
	.w8(32'hbc2d7bc2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902a2f),
	.w1(32'hbc00d243),
	.w2(32'h3bc2df87),
	.w3(32'hbc42a334),
	.w4(32'h3b47bc7f),
	.w5(32'h3c142466),
	.w6(32'hbc44908a),
	.w7(32'h3a90b967),
	.w8(32'h3c0cc91a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc6b68),
	.w1(32'h3c7199d1),
	.w2(32'h3ac19810),
	.w3(32'h3c8b7b58),
	.w4(32'h3b829e11),
	.w5(32'hbc54460a),
	.w6(32'h3cda83fa),
	.w7(32'h3c195c48),
	.w8(32'hbc0c2473),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1087e8),
	.w1(32'hbb614b2e),
	.w2(32'hbc2c2f36),
	.w3(32'hbb49154a),
	.w4(32'hbbc27f98),
	.w5(32'h3aed804b),
	.w6(32'h3bde8dee),
	.w7(32'hbbaddfb3),
	.w8(32'h3a88c57f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71d211),
	.w1(32'hbb5d6f31),
	.w2(32'hbc161072),
	.w3(32'h3b25243f),
	.w4(32'h3c040fb1),
	.w5(32'h3b816359),
	.w6(32'hba7c3f55),
	.w7(32'hbb0ab72f),
	.w8(32'h3bd2bf96),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969a90),
	.w1(32'h3c1cafa4),
	.w2(32'h3b69bf32),
	.w3(32'h3c1f1ce5),
	.w4(32'h3bf62102),
	.w5(32'h3b6cd759),
	.w6(32'h3c8890c7),
	.w7(32'h3c511c13),
	.w8(32'h3be16c8d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c3b18),
	.w1(32'h3bb6861f),
	.w2(32'h3b617dad),
	.w3(32'hbb4de99a),
	.w4(32'h39b8688d),
	.w5(32'h3b02d078),
	.w6(32'hbb258af8),
	.w7(32'hba509192),
	.w8(32'h3bf00697),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5a75c),
	.w1(32'h3a3616c8),
	.w2(32'hbb34a13d),
	.w3(32'hbc332e2e),
	.w4(32'hb9d4ac8a),
	.w5(32'hbb911779),
	.w6(32'hbaf02890),
	.w7(32'hbb4bc138),
	.w8(32'hbb2ff451),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9198ac),
	.w1(32'hba2db188),
	.w2(32'hbb3cda27),
	.w3(32'hba9c5e6e),
	.w4(32'h3b99050a),
	.w5(32'hbc20610b),
	.w6(32'h3ade719e),
	.w7(32'h3b08e9c3),
	.w8(32'hbc2e4e3d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49d997),
	.w1(32'hbc1628a8),
	.w2(32'hbbd49382),
	.w3(32'hbc295845),
	.w4(32'hbc00896a),
	.w5(32'hbc08feff),
	.w6(32'hbc340028),
	.w7(32'hbbda6506),
	.w8(32'hbc890eae),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbff0f8),
	.w1(32'hbc423878),
	.w2(32'hbc261919),
	.w3(32'hbb3102c3),
	.w4(32'hbb64e0f0),
	.w5(32'h391c02e9),
	.w6(32'hbc348082),
	.w7(32'hbc13f421),
	.w8(32'h39521589),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d9c28),
	.w1(32'h3bcee9ce),
	.w2(32'h3a33a9bb),
	.w3(32'h3b1d0cc1),
	.w4(32'hba55748a),
	.w5(32'h3b64a350),
	.w6(32'h3a5ea6e9),
	.w7(32'hba01fa29),
	.w8(32'hbac216a9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03ebb2),
	.w1(32'hbb9f92a3),
	.w2(32'h3b296674),
	.w3(32'hbb57aeb1),
	.w4(32'h3b5c6d83),
	.w5(32'h3bb77490),
	.w6(32'hbb2c8b00),
	.w7(32'h3aa5efd3),
	.w8(32'h3bf1755c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c261248),
	.w1(32'h3b6a09bc),
	.w2(32'h3b3c7cf3),
	.w3(32'h3b1ae3da),
	.w4(32'h3bf08791),
	.w5(32'hbbfd3e0c),
	.w6(32'h3b340c64),
	.w7(32'h3bb41dff),
	.w8(32'hbbca95e0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902127),
	.w1(32'hbbd01d4e),
	.w2(32'hbbdfb069),
	.w3(32'hbc09eedf),
	.w4(32'hbc299fd0),
	.w5(32'hbbb65a84),
	.w6(32'hbc2f56bb),
	.w7(32'hbc062591),
	.w8(32'hbbb0aed9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d5f95),
	.w1(32'hbc37637c),
	.w2(32'hbc70572b),
	.w3(32'hbc595e14),
	.w4(32'hbbbdbc3a),
	.w5(32'hbbd2dc93),
	.w6(32'h37725b97),
	.w7(32'h3b333f4d),
	.w8(32'hbc41a469),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d124),
	.w1(32'hbbfcad5e),
	.w2(32'h3b1cec1b),
	.w3(32'hbc08db4a),
	.w4(32'hbc5b8628),
	.w5(32'hbbd59b7f),
	.w6(32'hba838801),
	.w7(32'hbbb479e3),
	.w8(32'hbb9592df),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebf016),
	.w1(32'h3b5b6455),
	.w2(32'hbbbced6c),
	.w3(32'hbbda7fd0),
	.w4(32'hbb8c838f),
	.w5(32'h3b05059c),
	.w6(32'hbc2d7bff),
	.w7(32'hb9f2471e),
	.w8(32'h3b926482),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c9dd4),
	.w1(32'hba9df600),
	.w2(32'hba64263a),
	.w3(32'hbb8ee3b7),
	.w4(32'hbaaca0d8),
	.w5(32'hbb06cd93),
	.w6(32'hbbfe4742),
	.w7(32'hbbaf86e6),
	.w8(32'h3bc95421),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc7df4),
	.w1(32'h3bb09d4c),
	.w2(32'hba5ae9cc),
	.w3(32'hbb8a5394),
	.w4(32'hbbfe64a1),
	.w5(32'hbab98329),
	.w6(32'h3c8680b9),
	.w7(32'h3b0dac42),
	.w8(32'h3b1dda5a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096c51),
	.w1(32'h3ae92346),
	.w2(32'h3b74aca5),
	.w3(32'hbb26f12f),
	.w4(32'h388e345a),
	.w5(32'h3b3c9b96),
	.w6(32'hbbe16871),
	.w7(32'hbb21221a),
	.w8(32'h3b54b883),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule