module layer_8_featuremap_123(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7bda),
	.w1(32'hb9dceb93),
	.w2(32'hba118062),
	.w3(32'hbb40702e),
	.w4(32'hba6d1b30),
	.w5(32'hbc2377c7),
	.w6(32'hba8f3469),
	.w7(32'hbb0d5fe2),
	.w8(32'hbbf57a1d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5a46e),
	.w1(32'hbb4ae71f),
	.w2(32'h3b6466da),
	.w3(32'hbb3dcbf8),
	.w4(32'h3ba60c2f),
	.w5(32'h3c74c5e0),
	.w6(32'hbb3ce82c),
	.w7(32'h3bab377a),
	.w8(32'h3c6e2e9e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79c2f4),
	.w1(32'h3c1401ed),
	.w2(32'hbb66d994),
	.w3(32'h3bb47900),
	.w4(32'hbb7703ac),
	.w5(32'hbabd916a),
	.w6(32'h3b4388e7),
	.w7(32'hbb74b751),
	.w8(32'hb953b068),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7a776),
	.w1(32'hbc04ac32),
	.w2(32'hbbf0954c),
	.w3(32'hbc0be08c),
	.w4(32'hbb6ea7ea),
	.w5(32'h3c0c62d0),
	.w6(32'hbbbb5f77),
	.w7(32'hbb9a027e),
	.w8(32'h3bc5385a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dca26),
	.w1(32'hb9885372),
	.w2(32'hbc0f113d),
	.w3(32'hba89fe73),
	.w4(32'hbab2da07),
	.w5(32'h3b9f362b),
	.w6(32'h3ab8159c),
	.w7(32'h3b880c26),
	.w8(32'h3b68f78a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99d1eb),
	.w1(32'hbaf06b5e),
	.w2(32'hbc4fa654),
	.w3(32'h3ba50c9b),
	.w4(32'hbbd71c4a),
	.w5(32'hb9353102),
	.w6(32'h3ab4c542),
	.w7(32'hbc0c31fc),
	.w8(32'hbb469274),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb687c2a),
	.w1(32'hbb8eb605),
	.w2(32'h3b890da5),
	.w3(32'hbb5f60df),
	.w4(32'hbb5ae080),
	.w5(32'hbad5b764),
	.w6(32'hbb34d9a1),
	.w7(32'h3ad7701b),
	.w8(32'hba8f4dce),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5836ba),
	.w1(32'h3b6ac834),
	.w2(32'hba61c567),
	.w3(32'h3b929a07),
	.w4(32'h3ad2f8e1),
	.w5(32'hbaa09288),
	.w6(32'h3b94271c),
	.w7(32'hbb8d10d4),
	.w8(32'hbb983353),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace003f),
	.w1(32'hbb5a5e78),
	.w2(32'hbbaeae41),
	.w3(32'hbb9abe1c),
	.w4(32'hbba0fe81),
	.w5(32'hbbc7936d),
	.w6(32'hbc1ef5f9),
	.w7(32'h3989992c),
	.w8(32'hbbd2269f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06cf35),
	.w1(32'h3a0c5ad1),
	.w2(32'hbc18f90f),
	.w3(32'h39639635),
	.w4(32'hbbca8a28),
	.w5(32'h3ac9487c),
	.w6(32'h3b0ffa87),
	.w7(32'hbb640006),
	.w8(32'hba9792cf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44ff45),
	.w1(32'hbc0fbd90),
	.w2(32'hbc0afac3),
	.w3(32'hbbc9cbbe),
	.w4(32'hbbf38c00),
	.w5(32'h3b2b1b1f),
	.w6(32'hbb230fac),
	.w7(32'hbb96c5b2),
	.w8(32'h3c5fb880),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba907c7),
	.w1(32'h3ac767b6),
	.w2(32'h3bd528f3),
	.w3(32'h3c17e075),
	.w4(32'h3baa264c),
	.w5(32'h3ad6ab39),
	.w6(32'h3bb9e42a),
	.w7(32'h3b7cf668),
	.w8(32'hbb6c1e16),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf9283),
	.w1(32'h3b279149),
	.w2(32'h38831259),
	.w3(32'h3a6e8845),
	.w4(32'h390ed4c5),
	.w5(32'h38e8e1a6),
	.w6(32'h3b811473),
	.w7(32'h3931f8e6),
	.w8(32'h3951673a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37038ecf),
	.w1(32'hb5ac32f6),
	.w2(32'hb66ba8dd),
	.w3(32'h3716eac6),
	.w4(32'hb5d42c35),
	.w5(32'hb4b50dd9),
	.w6(32'h36fe2a64),
	.w7(32'hb6321875),
	.w8(32'hb5f3b1a0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c56131),
	.w1(32'h3670ca9a),
	.w2(32'h364c24e0),
	.w3(32'h36d3dfe7),
	.w4(32'h367cd185),
	.w5(32'h3651e3df),
	.w6(32'h366af453),
	.w7(32'h35bb5bd3),
	.w8(32'h35e22ba8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368eac18),
	.w1(32'h361bc68a),
	.w2(32'h35a01cdc),
	.w3(32'h3687cd82),
	.w4(32'h360815e7),
	.w5(32'h35288267),
	.w6(32'h366d5c2c),
	.w7(32'hb4921a82),
	.w8(32'hb5a2534f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886966f),
	.w1(32'h39164d2d),
	.w2(32'h395f90bd),
	.w3(32'h38dd89af),
	.w4(32'h39948e36),
	.w5(32'h3955e056),
	.w6(32'h392f2527),
	.w7(32'h38c301cf),
	.w8(32'h391d6276),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954152d),
	.w1(32'hb9171752),
	.w2(32'hb8ad92e5),
	.w3(32'hb987bbd9),
	.w4(32'hb7a74f20),
	.w5(32'h3886bea5),
	.w6(32'hb8b1ec3d),
	.w7(32'h385ca013),
	.w8(32'h38a3a81e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3d77b),
	.w1(32'h3ab94680),
	.w2(32'hb9210f3f),
	.w3(32'h3a879c32),
	.w4(32'h39002556),
	.w5(32'hb9f71887),
	.w6(32'h3a6af039),
	.w7(32'h3a3fed30),
	.w8(32'h39ec7b91),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f901aa),
	.w1(32'hb884a75b),
	.w2(32'hba1db9e9),
	.w3(32'h3671c8ad),
	.w4(32'hb93f6924),
	.w5(32'hba0b3e2a),
	.w6(32'h394921f4),
	.w7(32'h3929901a),
	.w8(32'hb9e8917f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1fc86),
	.w1(32'hb975ad16),
	.w2(32'hb7bf5880),
	.w3(32'hb9026c47),
	.w4(32'hb907d1da),
	.w5(32'hb988fd53),
	.w6(32'h3981dd1d),
	.w7(32'h38bc7f34),
	.w8(32'hb76cf3cb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904b74f),
	.w1(32'hb6364efa),
	.w2(32'h38435d3e),
	.w3(32'hb9a1b049),
	.w4(32'hb8d89ebe),
	.w5(32'hb8a0ed8f),
	.w6(32'hb90f2f4b),
	.w7(32'h381e4f8f),
	.w8(32'h37ac1ff2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20e36c),
	.w1(32'h3b3d9164),
	.w2(32'h3b277973),
	.w3(32'h3b020404),
	.w4(32'h3b042a26),
	.w5(32'h3afc80ba),
	.w6(32'h3af0bf77),
	.w7(32'h3b23280c),
	.w8(32'h3b2e116f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9315be6),
	.w1(32'hb966ee61),
	.w2(32'hb9adb98a),
	.w3(32'hb87a0aa4),
	.w4(32'hb816f948),
	.w5(32'hb8bb49be),
	.w6(32'h39003e69),
	.w7(32'h388aae6e),
	.w8(32'hb8f9a4b9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3631f5b7),
	.w1(32'hb68c8219),
	.w2(32'h3791e768),
	.w3(32'h37ac3d96),
	.w4(32'h37abdf8e),
	.w5(32'h37e107ed),
	.w6(32'h37aa6a88),
	.w7(32'h3748dee3),
	.w8(32'h3795a7af),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a655365),
	.w1(32'h3a54563c),
	.w2(32'h39eb2d58),
	.w3(32'h3a17959b),
	.w4(32'h397f8fca),
	.w5(32'h379a7eb1),
	.w6(32'h3a06e205),
	.w7(32'h39eeabd2),
	.w8(32'h39579914),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb450317e),
	.w1(32'hb5132a72),
	.w2(32'hb3ac7c99),
	.w3(32'hb56d5db6),
	.w4(32'h351c0a08),
	.w5(32'h3600de3d),
	.w6(32'h34bee12f),
	.w7(32'h33cec99b),
	.w8(32'h34e6eccb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4e21),
	.w1(32'h3c19cad1),
	.w2(32'h3bd73271),
	.w3(32'h3bd854a6),
	.w4(32'h3c22f02f),
	.w5(32'h37023f20),
	.w6(32'h3c125a45),
	.w7(32'h3c254a4f),
	.w8(32'h3bc0104d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e9784),
	.w1(32'h3a317300),
	.w2(32'h39e868b9),
	.w3(32'h39af46e2),
	.w4(32'h39c1b17e),
	.w5(32'h39892b88),
	.w6(32'h3989d34b),
	.w7(32'h39d6b433),
	.w8(32'h39d8b747),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38006474),
	.w1(32'h38ab90f6),
	.w2(32'h381f9b25),
	.w3(32'h38322586),
	.w4(32'h38634279),
	.w5(32'h38042aa2),
	.w6(32'h38dc6482),
	.w7(32'h3911eb6a),
	.w8(32'h38c689f9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b6d40c),
	.w1(32'hb66350d7),
	.w2(32'hb6ff4a4f),
	.w3(32'h37df8115),
	.w4(32'hb5f2ee33),
	.w5(32'hb699ae2b),
	.w6(32'h362b78bd),
	.w7(32'h3778ee82),
	.w8(32'h384d5a45),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9456a9b),
	.w1(32'hb9600edd),
	.w2(32'hb92f296c),
	.w3(32'hb81578b7),
	.w4(32'hb8a2f70c),
	.w5(32'hb959128b),
	.w6(32'h386ac866),
	.w7(32'hb6e175dc),
	.w8(32'hb95f71e9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ee46f0),
	.w1(32'h3556f151),
	.w2(32'h3424c5a6),
	.w3(32'h36f668b8),
	.w4(32'h35775390),
	.w5(32'h35e62ca6),
	.w6(32'h3680b7ba),
	.w7(32'hb609c4da),
	.w8(32'hb5a075e9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac7ae8),
	.w1(32'hb32dd7a8),
	.w2(32'hb548907f),
	.w3(32'h36d57f9b),
	.w4(32'hb43ff29d),
	.w5(32'hb528b1ea),
	.w6(32'h3659caab),
	.w7(32'hb600b49f),
	.w8(32'hb641aa95),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93738f3),
	.w1(32'hb8ebff6d),
	.w2(32'hb92831eb),
	.w3(32'hb876f57f),
	.w4(32'h386adf6e),
	.w5(32'hb8660201),
	.w6(32'h3828ebc7),
	.w7(32'h393fc25c),
	.w8(32'h38a974ca),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fc5f6),
	.w1(32'h38e3d381),
	.w2(32'hb961d518),
	.w3(32'hb7aa072a),
	.w4(32'hb9c5b298),
	.w5(32'hb9cdf36a),
	.w6(32'hb88ae370),
	.w7(32'hb93e3a55),
	.w8(32'hb9abafbd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34959251),
	.w1(32'hb5d338f1),
	.w2(32'hb573b519),
	.w3(32'h360e0481),
	.w4(32'hb6084601),
	.w5(32'hb57ece86),
	.w6(32'h35a05203),
	.w7(32'hb5cef9b5),
	.w8(32'hb679162d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0c9c2),
	.w1(32'h38e8f390),
	.w2(32'h393ad397),
	.w3(32'hb9131317),
	.w4(32'h36776491),
	.w5(32'h38be9851),
	.w6(32'hb90546ff),
	.w7(32'h385b5b79),
	.w8(32'h3916a3e9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c0e340),
	.w1(32'hb654dfa7),
	.w2(32'hb65d48bc),
	.w3(32'h36a1175d),
	.w4(32'h35a1ae67),
	.w5(32'hb5aa34c3),
	.w6(32'h35894d4b),
	.w7(32'hb6851362),
	.w8(32'hb6a0b86d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789ba65),
	.w1(32'hb60a9544),
	.w2(32'h3553e8ef),
	.w3(32'h37b5fae9),
	.w4(32'h373c2de7),
	.w5(32'h365fece9),
	.w6(32'h37748738),
	.w7(32'hb6b92798),
	.w8(32'hb6fd3802),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945d12),
	.w1(32'h38f011a5),
	.w2(32'hb8c7ed39),
	.w3(32'hb5dca29e),
	.w4(32'h38d3baba),
	.w5(32'h39a29af6),
	.w6(32'h3a0633ce),
	.w7(32'h3a5c2b45),
	.w8(32'h3a23bf53),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd5c32),
	.w1(32'hb8cd401e),
	.w2(32'hb884689f),
	.w3(32'hb93ad41a),
	.w4(32'hb90d9a3d),
	.w5(32'hb8f35490),
	.w6(32'hb8f85e5f),
	.w7(32'hb8da2b16),
	.w8(32'hb8b1c7d8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358d3334),
	.w1(32'h36850608),
	.w2(32'h36ca2240),
	.w3(32'h36f7e220),
	.w4(32'h373d3790),
	.w5(32'h370870ea),
	.w6(32'h368819f2),
	.w7(32'hb60e05f9),
	.w8(32'hb5e2b824),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d68991),
	.w1(32'h3904f7ba),
	.w2(32'h38e5a1c5),
	.w3(32'h38b3bb14),
	.w4(32'h38cf2070),
	.w5(32'h38c5a16d),
	.w6(32'h38adc172),
	.w7(32'h390cf477),
	.w8(32'h38e7e2b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81213e),
	.w1(32'h3a859359),
	.w2(32'h39e411ae),
	.w3(32'h3a34d334),
	.w4(32'h39cde4f4),
	.w5(32'h38ed811f),
	.w6(32'h39f11651),
	.w7(32'h3a133ee0),
	.w8(32'h39f172ba),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bfb3f),
	.w1(32'h396bd83d),
	.w2(32'h39125867),
	.w3(32'h39153914),
	.w4(32'h3932881f),
	.w5(32'h3914316e),
	.w6(32'h39325edb),
	.w7(32'h393679c2),
	.w8(32'h393e25b7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a6371c),
	.w1(32'hb493bd24),
	.w2(32'hb5139776),
	.w3(32'h36122c43),
	.w4(32'hb4282cff),
	.w5(32'h3463d9cb),
	.w6(32'h352344b4),
	.w7(32'hb5feadca),
	.w8(32'hb594341a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05dff1),
	.w1(32'h3a0512cb),
	.w2(32'h39048027),
	.w3(32'h39f29122),
	.w4(32'h395b4ee1),
	.w5(32'h37f97d2c),
	.w6(32'h39af8c9c),
	.w7(32'h395bd11b),
	.w8(32'h392002dc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388950cc),
	.w1(32'h398838dd),
	.w2(32'h39944d9b),
	.w3(32'hb64d11aa),
	.w4(32'h397a5353),
	.w5(32'h398518b1),
	.w6(32'h37f7bb70),
	.w7(32'h3985cb85),
	.w8(32'h39bd3dd4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d00d6),
	.w1(32'h3a183a6b),
	.w2(32'h3949dcd3),
	.w3(32'h3a0b752f),
	.w4(32'h39eac79c),
	.w5(32'h397c28a5),
	.w6(32'h3a1c0872),
	.w7(32'h3a2b82b4),
	.w8(32'h3a0196a2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37034766),
	.w1(32'h36fb9107),
	.w2(32'h373f3584),
	.w3(32'hb8cd71e4),
	.w4(32'hb8f4066f),
	.w5(32'hb89d858f),
	.w6(32'hb8502517),
	.w7(32'hb82d122a),
	.w8(32'hb7438730),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e8780),
	.w1(32'h3b822838),
	.w2(32'h3af1febb),
	.w3(32'h3b5f06b4),
	.w4(32'h3b2f1c7e),
	.w5(32'h3adc417f),
	.w6(32'h3b24e942),
	.w7(32'h3b4d441b),
	.w8(32'h3b487909),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042bf2),
	.w1(32'h39e49e02),
	.w2(32'hb8646547),
	.w3(32'h3a02c43f),
	.w4(32'h394a3959),
	.w5(32'hb8ee6ae9),
	.w6(32'h39f3ac5b),
	.w7(32'h396d77fd),
	.w8(32'hb8767dad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79ee6c4),
	.w1(32'hb713560b),
	.w2(32'hb8877130),
	.w3(32'hb89dc5f6),
	.w4(32'hb8ecf5c0),
	.w5(32'hb873b8b7),
	.w6(32'hb7675246),
	.w7(32'hb8713f61),
	.w8(32'hb85e4da0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364d6d2f),
	.w1(32'hb6107ec3),
	.w2(32'hb54d53b0),
	.w3(32'h352e83e4),
	.w4(32'hb6d424d5),
	.w5(32'hb69563bf),
	.w6(32'hb6308cc4),
	.w7(32'hb7176833),
	.w8(32'hb6e6dfbf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a29e6),
	.w1(32'h3a946d90),
	.w2(32'h3a4cbe36),
	.w3(32'h3a1608ce),
	.w4(32'h3a0a3f3e),
	.w5(32'h399b0c3c),
	.w6(32'h3a52a258),
	.w7(32'h3a30bd60),
	.w8(32'h3a310284),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986971a),
	.w1(32'hb8dfc69d),
	.w2(32'hb7a90b7c),
	.w3(32'hb8c81c2d),
	.w4(32'h38e3b8a3),
	.w5(32'h389b055e),
	.w6(32'h3909a8c1),
	.w7(32'h391f8a12),
	.w8(32'h392d7f3a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c8dec),
	.w1(32'h3a23e9cd),
	.w2(32'h39c5cdba),
	.w3(32'h39471511),
	.w4(32'h3990ad5f),
	.w5(32'h3a028b53),
	.w6(32'hb5a96762),
	.w7(32'h39cf8794),
	.w8(32'h3a2105b9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b56250),
	.w1(32'h3a46f4d6),
	.w2(32'h3a2e6d01),
	.w3(32'h39c3fd0b),
	.w4(32'h3a0f5282),
	.w5(32'h39cf0a58),
	.w6(32'h39bc2bf4),
	.w7(32'h3a164ff7),
	.w8(32'h3a11fbe2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39083682),
	.w1(32'h394112db),
	.w2(32'h392d6c92),
	.w3(32'h38afaa90),
	.w4(32'h392c7a43),
	.w5(32'h38e30db1),
	.w6(32'h387438d6),
	.w7(32'h38d83617),
	.w8(32'h38cc71f6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37438347),
	.w1(32'h3696ccea),
	.w2(32'h3612c32b),
	.w3(32'h3728185e),
	.w4(32'h351571d5),
	.w5(32'hb5e4bfe4),
	.w6(32'h36aa690c),
	.w7(32'hb69ddcd2),
	.w8(32'hb684d070),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34fe2bc8),
	.w1(32'h3840ff5d),
	.w2(32'h386b4ed0),
	.w3(32'h384b7650),
	.w4(32'h3850805c),
	.w5(32'h381d7cb1),
	.w6(32'h37cff993),
	.w7(32'h3806aff6),
	.w8(32'h38408e79),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f1a38),
	.w1(32'h3988577c),
	.w2(32'h38f4573c),
	.w3(32'hb7d4f461),
	.w4(32'h3964bd23),
	.w5(32'h38e91c04),
	.w6(32'h39174f4f),
	.w7(32'h398f8d0d),
	.w8(32'h394ad99f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da5e3e),
	.w1(32'hb888cf29),
	.w2(32'hb93e5c2c),
	.w3(32'h3917f5ae),
	.w4(32'h38fb81cb),
	.w5(32'h3871202c),
	.w6(32'h38f0cb46),
	.w7(32'h38ee892e),
	.w8(32'h38c510ca),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a9250),
	.w1(32'hb84c34d5),
	.w2(32'hb8aaf5a6),
	.w3(32'h38a535cb),
	.w4(32'h37e4e9ca),
	.w5(32'hb85b57ec),
	.w6(32'h36f3d0ba),
	.w7(32'hb90616d6),
	.w8(32'hb89e936e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ef609),
	.w1(32'h39c34179),
	.w2(32'h39914ba4),
	.w3(32'h38da6f2d),
	.w4(32'h395d8f87),
	.w5(32'h39815e47),
	.w6(32'h399ef75d),
	.w7(32'h3a0a2920),
	.w8(32'h39eaf684),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b07343),
	.w1(32'h398352ff),
	.w2(32'h3931fc0c),
	.w3(32'h38fd1e18),
	.w4(32'h3981d528),
	.w5(32'h397ed9f0),
	.w6(32'h3935bf58),
	.w7(32'h39b97e4f),
	.w8(32'h39952672),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ba51e),
	.w1(32'h390ec045),
	.w2(32'h37146365),
	.w3(32'h38aa6dec),
	.w4(32'h37fd02da),
	.w5(32'h3685ab98),
	.w6(32'h392d420a),
	.w7(32'h392d2767),
	.w8(32'h38a345fc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36542eb2),
	.w1(32'h3670e0dd),
	.w2(32'h3657aa36),
	.w3(32'h36e11c5c),
	.w4(32'h36095ee5),
	.w5(32'h35e66dc5),
	.w6(32'h36948a71),
	.w7(32'h36448e41),
	.w8(32'hb59ddc64),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e3ef),
	.w1(32'h3a78ef5d),
	.w2(32'h39f724a9),
	.w3(32'h39f55c8c),
	.w4(32'h39851809),
	.w5(32'hb966ed2b),
	.w6(32'h39c19fc6),
	.w7(32'h39c95cde),
	.w8(32'h395bc594),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb501e705),
	.w1(32'hb62201b4),
	.w2(32'hb5fdfcff),
	.w3(32'h3581ef24),
	.w4(32'hb5781224),
	.w5(32'hb5a88c91),
	.w6(32'h35382014),
	.w7(32'hb59adc15),
	.w8(32'hb5843637),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b296),
	.w1(32'hb9dfcc27),
	.w2(32'hb9e16c56),
	.w3(32'hb99b9d04),
	.w4(32'hb8d11357),
	.w5(32'hb9caa4a0),
	.w6(32'hb8ba0a56),
	.w7(32'h3707d508),
	.w8(32'hb9d16c49),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6587875),
	.w1(32'hb531c9cc),
	.w2(32'hb71cefe9),
	.w3(32'h34edd16c),
	.w4(32'hb4d78d54),
	.w5(32'hb73fa317),
	.w6(32'hb5b138ea),
	.w7(32'hb68f1ef2),
	.w8(32'hb7669e14),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d2dab),
	.w1(32'h38c4d886),
	.w2(32'h388016b3),
	.w3(32'hb8925b69),
	.w4(32'hb6bbb9c5),
	.w5(32'hb690d185),
	.w6(32'hb70085b4),
	.w7(32'h38e51921),
	.w8(32'h382d807d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c72734),
	.w1(32'h3687661f),
	.w2(32'h36599b62),
	.w3(32'h36bdf4cf),
	.w4(32'h368a1d52),
	.w5(32'h35fb7744),
	.w6(32'h36a370db),
	.w7(32'h35f3bd21),
	.w8(32'h364bd1f9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d9fe3),
	.w1(32'h3aa6b731),
	.w2(32'h3a5213cf),
	.w3(32'h3a1d9b62),
	.w4(32'h3a6c74ef),
	.w5(32'h3a4249ee),
	.w6(32'h3a62f815),
	.w7(32'h3a9c7265),
	.w8(32'h3a8cfd29),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3563f3d1),
	.w1(32'hb524ad9e),
	.w2(32'hbba80579),
	.w3(32'hb630e830),
	.w4(32'hba37d644),
	.w5(32'hbbe33a4d),
	.w6(32'hb6380a05),
	.w7(32'hbb8ead20),
	.w8(32'h3ab0af9b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd674a),
	.w1(32'hb9362416),
	.w2(32'h3b940134),
	.w3(32'h3b93275b),
	.w4(32'h3b0add7f),
	.w5(32'h3ad9c610),
	.w6(32'h3b75097e),
	.w7(32'hbacb28c5),
	.w8(32'h3bbc2417),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc579bb),
	.w1(32'h3b5932b2),
	.w2(32'h39f11e4a),
	.w3(32'h3bcd1aec),
	.w4(32'h3bbf6d2d),
	.w5(32'h3bf5db13),
	.w6(32'hbab6335f),
	.w7(32'hbaf727e1),
	.w8(32'h3bdba7dd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb2c3a),
	.w1(32'h3b4367e8),
	.w2(32'hbc312f22),
	.w3(32'h3b9353b1),
	.w4(32'hb8d489e8),
	.w5(32'hbaae9887),
	.w6(32'hba7a98f3),
	.w7(32'hbaa3a882),
	.w8(32'hbce58ccc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878a22),
	.w1(32'hbc3046ce),
	.w2(32'h3a92e49d),
	.w3(32'hbbb56423),
	.w4(32'hbbae15f2),
	.w5(32'hbb1adeac),
	.w6(32'h3c2f1720),
	.w7(32'hbb434641),
	.w8(32'h3b9138c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140db7),
	.w1(32'h3b1ef5f7),
	.w2(32'hbb9ba018),
	.w3(32'h3c6685cf),
	.w4(32'h3c2bc1e1),
	.w5(32'hbc147dad),
	.w6(32'h3a1c62d1),
	.w7(32'hbb874319),
	.w8(32'h3d3fa779),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c3cb7),
	.w1(32'h3ca75652),
	.w2(32'hbc1625d7),
	.w3(32'hbbb07d2d),
	.w4(32'hbb5409d2),
	.w5(32'hbc948f84),
	.w6(32'hbcc85058),
	.w7(32'hbbb03331),
	.w8(32'hbc8daa0b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c9f5),
	.w1(32'hbc1b4a73),
	.w2(32'h3c761381),
	.w3(32'hbabbe039),
	.w4(32'hbc00f3b2),
	.w5(32'h3becc269),
	.w6(32'h3c00bb4a),
	.w7(32'hbb68d5e2),
	.w8(32'hba125689),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cfd08),
	.w1(32'h3b163494),
	.w2(32'h3c2fe54d),
	.w3(32'hba845312),
	.w4(32'hbc2603a3),
	.w5(32'h3c880622),
	.w6(32'hbb7f82ae),
	.w7(32'hba9c5a46),
	.w8(32'h3c10c9cb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90dcc8),
	.w1(32'h3a5c5922),
	.w2(32'h3c0baa8b),
	.w3(32'hbca2ebc2),
	.w4(32'hbbd666b8),
	.w5(32'h3bd9bf87),
	.w6(32'hbbbeb36f),
	.w7(32'h3c85db7f),
	.w8(32'hbc425834),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd4539),
	.w1(32'hbb0b4a2a),
	.w2(32'h3acddccf),
	.w3(32'hbc0e3932),
	.w4(32'h3cb838f9),
	.w5(32'h3ca92dd2),
	.w6(32'hbb504900),
	.w7(32'h3c71a9a8),
	.w8(32'hbc7f3e03),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ced2),
	.w1(32'h3c81b67a),
	.w2(32'hba8b2b62),
	.w3(32'hbc043188),
	.w4(32'h3c40ebbe),
	.w5(32'h3c170eea),
	.w6(32'h3bc8dd34),
	.w7(32'h3c14b437),
	.w8(32'h3b2aeb0d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eec9e),
	.w1(32'hbbb0740f),
	.w2(32'hbb2e2281),
	.w3(32'hba47df0c),
	.w4(32'h3aee11aa),
	.w5(32'hba872100),
	.w6(32'hbac42494),
	.w7(32'hbb0bab56),
	.w8(32'h3b3d88c0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbd2d1),
	.w1(32'hbb300189),
	.w2(32'h3c769417),
	.w3(32'hbc3f2d39),
	.w4(32'hbbdbbf54),
	.w5(32'h3d68e6f4),
	.w6(32'hbc5d6162),
	.w7(32'h3c730bbd),
	.w8(32'h3c560441),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c0d57),
	.w1(32'h3ccefa57),
	.w2(32'h3baf6396),
	.w3(32'hbd1c589e),
	.w4(32'h3c06e8f9),
	.w5(32'hbc16099f),
	.w6(32'hbd56b6b0),
	.w7(32'hbbd430e0),
	.w8(32'h3c929e09),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10bdc7),
	.w1(32'hba8ee151),
	.w2(32'h3b9fcf74),
	.w3(32'h3cb7b1d5),
	.w4(32'hbc935449),
	.w5(32'h3cc20a83),
	.w6(32'hbb79c0e9),
	.w7(32'hbca2ff05),
	.w8(32'h3cea7e3d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ae75),
	.w1(32'hbc4e089c),
	.w2(32'hbc160af0),
	.w3(32'h3ae01e45),
	.w4(32'h382ba069),
	.w5(32'h3caad0ff),
	.w6(32'hbca4a13d),
	.w7(32'h3c4141c7),
	.w8(32'hbc4e1a8f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25c2c),
	.w1(32'h3bc92b9a),
	.w2(32'hbcb9a776),
	.w3(32'hbbe2e229),
	.w4(32'hbc1ac300),
	.w5(32'hbd058557),
	.w6(32'hbba7214b),
	.w7(32'hbb6a13ec),
	.w8(32'h3c093ec1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc15916),
	.w1(32'h3af64c32),
	.w2(32'h3b09fc11),
	.w3(32'h3c0b1100),
	.w4(32'hb9b07c22),
	.w5(32'h3a08b2d8),
	.w6(32'h3b517f4e),
	.w7(32'hb9fce06b),
	.w8(32'hbb70c885),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ffd3),
	.w1(32'h3a55bb26),
	.w2(32'h3b49c43a),
	.w3(32'h39aefe1f),
	.w4(32'hbc1076ce),
	.w5(32'h3c55d3c6),
	.w6(32'hba91dbb4),
	.w7(32'h3b1f2085),
	.w8(32'hbc59540a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f378d),
	.w1(32'hbc579544),
	.w2(32'hbc97e62a),
	.w3(32'h3a2eb8e4),
	.w4(32'h3c1ccc56),
	.w5(32'hbcde6dcf),
	.w6(32'h3b5d3f68),
	.w7(32'h3af558f3),
	.w8(32'hba4d9e6c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc441519),
	.w1(32'h3ca27f7f),
	.w2(32'h3bbd0f89),
	.w3(32'h3c22be9e),
	.w4(32'hbc1a2a69),
	.w5(32'hbd1b071b),
	.w6(32'h3b7b19de),
	.w7(32'hbb125ede),
	.w8(32'h3d338a13),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aced883),
	.w1(32'hbb698f35),
	.w2(32'h3c02054f),
	.w3(32'h3c1a1ea5),
	.w4(32'hb9a2e2bc),
	.w5(32'hbb586f2d),
	.w6(32'hbc9b4dcb),
	.w7(32'h3bc3fcdf),
	.w8(32'hbbe7d633),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf48ecc),
	.w1(32'h3bae88e1),
	.w2(32'hbc07d273),
	.w3(32'h3b71ffa2),
	.w4(32'h3c5b892f),
	.w5(32'hbb2044fc),
	.w6(32'h3a08f126),
	.w7(32'h3c4d03ab),
	.w8(32'hbb8a8e52),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e8f46),
	.w1(32'h3bf4cb15),
	.w2(32'h3c19db2b),
	.w3(32'h3b281a05),
	.w4(32'hbbb3b352),
	.w5(32'h3c12b9a6),
	.w6(32'h3ca2f3ac),
	.w7(32'h3c14ac28),
	.w8(32'hbb46d60e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc182ddc),
	.w1(32'h3b8d2648),
	.w2(32'hbbcd9e43),
	.w3(32'h3c48a9c3),
	.w4(32'h3a1e36ab),
	.w5(32'hbc5a5070),
	.w6(32'hbbd1f17d),
	.w7(32'hbb96092e),
	.w8(32'hbc159b4a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54030),
	.w1(32'hbc31f122),
	.w2(32'hbc4b006e),
	.w3(32'h3c1395af),
	.w4(32'hbc33f9fe),
	.w5(32'h3bf97a94),
	.w6(32'hbc0ae641),
	.w7(32'h3b203031),
	.w8(32'hbcc778ea),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f73ef),
	.w1(32'h3b28af9b),
	.w2(32'h3b03ecc1),
	.w3(32'hbc525aec),
	.w4(32'h3bd3ee0d),
	.w5(32'h3a2f4421),
	.w6(32'hbb67b5f5),
	.w7(32'h3b9dc1c2),
	.w8(32'hbc78c483),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd646),
	.w1(32'h3a53ffec),
	.w2(32'h3ba74551),
	.w3(32'hbb91878a),
	.w4(32'hbba87159),
	.w5(32'hbccf0d3b),
	.w6(32'h3bec79c6),
	.w7(32'hbc8558e8),
	.w8(32'hbbc71c04),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a46fe),
	.w1(32'h3bad67d9),
	.w2(32'h3a917931),
	.w3(32'h3c17709d),
	.w4(32'h3be9ee2a),
	.w5(32'hbbea08ec),
	.w6(32'h3940f3c8),
	.w7(32'hbb7d4b87),
	.w8(32'h3cb4d93e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf8593),
	.w1(32'hb9808c79),
	.w2(32'hbcb30bf6),
	.w3(32'h3c237d6e),
	.w4(32'h3b2b0b5a),
	.w5(32'h3bb6f85e),
	.w6(32'h3aa8b1e6),
	.w7(32'h3cde5756),
	.w8(32'hbd861e58),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c385ef2),
	.w1(32'h3bc76a64),
	.w2(32'hbb9bcc6e),
	.w3(32'hbaa85054),
	.w4(32'hba962d70),
	.w5(32'hbc274224),
	.w6(32'h3d11ce7e),
	.w7(32'hbbca0f95),
	.w8(32'h3aae69ae),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6a71f),
	.w1(32'h3a542d99),
	.w2(32'hbcc4698d),
	.w3(32'h3bc84734),
	.w4(32'hbba52320),
	.w5(32'h3c278e02),
	.w6(32'h3bbc30cf),
	.w7(32'h3a68ef68),
	.w8(32'hbbaac547),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af876),
	.w1(32'h39547943),
	.w2(32'hbbc135e2),
	.w3(32'hbc70e2ac),
	.w4(32'h3c0217ad),
	.w5(32'h3c5f65df),
	.w6(32'hbc27ca5f),
	.w7(32'h3cd1c4a7),
	.w8(32'hbdb2a420),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46f9db),
	.w1(32'h3c0bf5b8),
	.w2(32'hbc221769),
	.w3(32'hbc9095ab),
	.w4(32'h3ae9decc),
	.w5(32'h3c892f89),
	.w6(32'h3cf7e25c),
	.w7(32'h3cbe3440),
	.w8(32'hbc6ac3f6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc824b8e),
	.w1(32'h3c4f7f7d),
	.w2(32'hb9faf3c5),
	.w3(32'hbc7450cd),
	.w4(32'h3be43f5f),
	.w5(32'hbb5a9682),
	.w6(32'h3a8f24bd),
	.w7(32'h3c57a501),
	.w8(32'hbc3fa9a3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff25bb),
	.w1(32'hbb148dca),
	.w2(32'hbbdf9ccb),
	.w3(32'h3c48bd3c),
	.w4(32'hbadad9ad),
	.w5(32'hbc9a33cb),
	.w6(32'hba5bf321),
	.w7(32'hbcdff053),
	.w8(32'h3d53d60c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76a53b),
	.w1(32'h3c07a788),
	.w2(32'hbc94ca93),
	.w3(32'hbbf5e57c),
	.w4(32'hbcd16f6b),
	.w5(32'hbc58becf),
	.w6(32'hbca479af),
	.w7(32'hbcc8b1ac),
	.w8(32'h3b81bce8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f199a),
	.w1(32'hbcc0f04d),
	.w2(32'hbc29d531),
	.w3(32'hbbbf86f3),
	.w4(32'hbc0089c8),
	.w5(32'h3bf336b1),
	.w6(32'hbc0123a8),
	.w7(32'hbc9e9aaa),
	.w8(32'h3d0cddf8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c592c84),
	.w1(32'hbc9f9079),
	.w2(32'h3c85d759),
	.w3(32'h3b2dea00),
	.w4(32'hbcb32b9e),
	.w5(32'h3cc7b231),
	.w6(32'hbbc9587b),
	.w7(32'h3c84d337),
	.w8(32'hbb3478c5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca00e),
	.w1(32'hbc04242d),
	.w2(32'h3a78b1ee),
	.w3(32'h3bb261eb),
	.w4(32'hbc5e9361),
	.w5(32'hbc2abdfc),
	.w6(32'h3b808009),
	.w7(32'hbca56f09),
	.w8(32'h3c8fa69e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b59d6),
	.w1(32'hbb89b980),
	.w2(32'hb9fa8b1a),
	.w3(32'h3c44233f),
	.w4(32'hbb8124ca),
	.w5(32'hbba1a097),
	.w6(32'hbd050d1c),
	.w7(32'hbb83830e),
	.w8(32'h3b238eb7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38917dde),
	.w1(32'h3a6a7437),
	.w2(32'hbc50fec3),
	.w3(32'h3b91fe13),
	.w4(32'hbbf01d46),
	.w5(32'hbc87fe29),
	.w6(32'h3b336216),
	.w7(32'h3beaca36),
	.w8(32'hbc862b59),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2f229),
	.w1(32'hbbc1eb84),
	.w2(32'hbb19db52),
	.w3(32'hbc1b8d58),
	.w4(32'hbc178ccf),
	.w5(32'hbbaadacb),
	.w6(32'h3b11fc62),
	.w7(32'hbcc1a66d),
	.w8(32'h3baeecb6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaad3fb),
	.w1(32'hbc0c2899),
	.w2(32'h3ba0ccbb),
	.w3(32'h3c120903),
	.w4(32'h3b75c73a),
	.w5(32'h3be36135),
	.w6(32'h3b58fe16),
	.w7(32'hbab4c1e6),
	.w8(32'h3c3f206f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092a58),
	.w1(32'hbbe6efb6),
	.w2(32'hbc641384),
	.w3(32'h3b85dabe),
	.w4(32'hbab9e66a),
	.w5(32'h3cac4399),
	.w6(32'hbbd2dc92),
	.w7(32'hba896de1),
	.w8(32'h3b26a91a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4c7eb),
	.w1(32'hbc1411f6),
	.w2(32'hbb2af324),
	.w3(32'h3b04ab2d),
	.w4(32'hbb0a5563),
	.w5(32'hbc08e183),
	.w6(32'h3c081ed2),
	.w7(32'hbbbbec14),
	.w8(32'h3acc765a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52cbf7),
	.w1(32'h3a072f0e),
	.w2(32'h3c95e947),
	.w3(32'h3bc2e6b8),
	.w4(32'hbc3a8d42),
	.w5(32'h3d5e8a07),
	.w6(32'h3b867d4a),
	.w7(32'h3ce84f9a),
	.w8(32'hbcf7aebe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd38da63),
	.w1(32'h3c86df34),
	.w2(32'hbc70de9f),
	.w3(32'hbd1c3e0b),
	.w4(32'hbb9ac9cf),
	.w5(32'hbc9066eb),
	.w6(32'h3c2d9ec7),
	.w7(32'hbd2331e5),
	.w8(32'h3c95ccab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca03d7),
	.w1(32'hbc52696c),
	.w2(32'hbb8bffd4),
	.w3(32'h3b5864fa),
	.w4(32'h3b09de23),
	.w5(32'h3c1a88e5),
	.w6(32'hbc587171),
	.w7(32'hba3397f3),
	.w8(32'hbb13fd6e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b618),
	.w1(32'h3b87887e),
	.w2(32'h3c025812),
	.w3(32'h3b96770c),
	.w4(32'hbbcfc16f),
	.w5(32'hbc625c62),
	.w6(32'hbb04f9a0),
	.w7(32'h3c0d083b),
	.w8(32'hbba2cd91),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49b826),
	.w1(32'h3b4c7300),
	.w2(32'h3abbe996),
	.w3(32'h3c152089),
	.w4(32'h3ac591c9),
	.w5(32'h3baf23ae),
	.w6(32'h39c921cd),
	.w7(32'h3b835cb8),
	.w8(32'hbc1f5f68),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule