module layer_10_featuremap_495(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01ff2e),
	.w1(32'hbb12f634),
	.w2(32'hbbeb2934),
	.w3(32'hbbd34400),
	.w4(32'hbb49d5d2),
	.w5(32'hbbcffa68),
	.w6(32'hbb2560e4),
	.w7(32'hbb439697),
	.w8(32'hbbb35763),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47a778),
	.w1(32'h3b210aaf),
	.w2(32'hbaa5795c),
	.w3(32'hbb73f1a9),
	.w4(32'hbb188e04),
	.w5(32'h3b855b68),
	.w6(32'hbbcd2dc0),
	.w7(32'h3b3a83f7),
	.w8(32'h3a48840e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a385000),
	.w1(32'hbbccddca),
	.w2(32'hbb96bf5b),
	.w3(32'h3be8a761),
	.w4(32'hba660b10),
	.w5(32'h3b1201b7),
	.w6(32'h3b95ee50),
	.w7(32'hbb5d5a7f),
	.w8(32'h3b68a9a4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4231),
	.w1(32'h3a9b7eae),
	.w2(32'h3ba99042),
	.w3(32'hbb56d59f),
	.w4(32'hba30beb0),
	.w5(32'h3c098fcf),
	.w6(32'hbabda54f),
	.w7(32'hba1692f3),
	.w8(32'h3b9efa61),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71019),
	.w1(32'h3a8b6d00),
	.w2(32'h37a7982a),
	.w3(32'h3bcb221d),
	.w4(32'h3a80b032),
	.w5(32'h3a92e545),
	.w6(32'h3b8f91d8),
	.w7(32'h3aab199a),
	.w8(32'hb9c05903),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dd6f7),
	.w1(32'h3bd0758b),
	.w2(32'h3b73a271),
	.w3(32'hbaaaa018),
	.w4(32'h39944e6e),
	.w5(32'h39ab4cfb),
	.w6(32'hbae90174),
	.w7(32'h3b1de4c7),
	.w8(32'h392632d1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805084),
	.w1(32'hb9867773),
	.w2(32'hbbaa544a),
	.w3(32'h3b9c2dc0),
	.w4(32'hbaf99b57),
	.w5(32'hbc0ebfce),
	.w6(32'h3b6eb28a),
	.w7(32'hbbb9bfba),
	.w8(32'hbc21e1a8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd190c8),
	.w1(32'hbb378059),
	.w2(32'hbba6b590),
	.w3(32'hbc3af0e9),
	.w4(32'h3abce843),
	.w5(32'h3b4b2f92),
	.w6(32'hbc21ff8b),
	.w7(32'h39c5040a),
	.w8(32'h3b324f91),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af468bb),
	.w1(32'hbacc1915),
	.w2(32'h3a9795a3),
	.w3(32'h3ba4119a),
	.w4(32'hbb998752),
	.w5(32'h38cb3c6e),
	.w6(32'h3b69f0f1),
	.w7(32'hbb4a7745),
	.w8(32'hbb374ab1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5931ea),
	.w1(32'hbb941d1e),
	.w2(32'hbbb78ae0),
	.w3(32'hba59f970),
	.w4(32'hb99c01e3),
	.w5(32'hbb3ee6e9),
	.w6(32'h3908e3b4),
	.w7(32'hbae26d64),
	.w8(32'hbb924df5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6091d1),
	.w1(32'hba311296),
	.w2(32'hbae8b350),
	.w3(32'hbaf859bb),
	.w4(32'hb9a9389c),
	.w5(32'hbb4ab509),
	.w6(32'hbb82bd21),
	.w7(32'hbb9e3c86),
	.w8(32'hbb23f93d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe18a8),
	.w1(32'h3b7a8f9c),
	.w2(32'hbb85c667),
	.w3(32'hbb63b894),
	.w4(32'h3b0fea46),
	.w5(32'hbb4d5be8),
	.w6(32'hb7cd1ee8),
	.w7(32'hbae252fd),
	.w8(32'hbc120130),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf23d),
	.w1(32'hbafbaa18),
	.w2(32'hbba32bbf),
	.w3(32'hbbaa06e1),
	.w4(32'hba29d09f),
	.w5(32'h3c32de6a),
	.w6(32'hbb746d55),
	.w7(32'h3b91ff04),
	.w8(32'hb9cf8b82),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd321a7),
	.w1(32'hbb8a66d4),
	.w2(32'hb97dc0f5),
	.w3(32'hbb4927f5),
	.w4(32'hbc2c0c14),
	.w5(32'h3a5be3e3),
	.w6(32'hbbcaa2f4),
	.w7(32'hba5a82a7),
	.w8(32'h3b906170),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29488),
	.w1(32'h3a836a95),
	.w2(32'hbae012b1),
	.w3(32'hbaf66ae6),
	.w4(32'hb9c1a755),
	.w5(32'h3a54458a),
	.w6(32'hbb53f7a3),
	.w7(32'hbb51dea3),
	.w8(32'hba02a492),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3c837),
	.w1(32'hb995f700),
	.w2(32'hbb1fe8ef),
	.w3(32'hbac4b353),
	.w4(32'h3aad2699),
	.w5(32'h3ae235e2),
	.w6(32'hba80624b),
	.w7(32'hba34ef7e),
	.w8(32'h3900c91a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994ec0),
	.w1(32'hbb0f320f),
	.w2(32'hbb1e0adb),
	.w3(32'hbba15f4b),
	.w4(32'h3a5f63f7),
	.w5(32'h39e7872a),
	.w6(32'hba9ce0c6),
	.w7(32'hbb0b1117),
	.w8(32'hb9e8b1bd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8796d),
	.w1(32'hbbc65fae),
	.w2(32'hbbd9cd9c),
	.w3(32'hbaf8c30f),
	.w4(32'hbb04eed8),
	.w5(32'hbb9a1083),
	.w6(32'h3a8dccf7),
	.w7(32'hbb9af940),
	.w8(32'hbb829846),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33dbe4),
	.w1(32'hba25275e),
	.w2(32'hbb9cef20),
	.w3(32'h3a1ae8c7),
	.w4(32'hbab122ce),
	.w5(32'hbaa144b3),
	.w6(32'h3a69f11c),
	.w7(32'hbb23a1a0),
	.w8(32'hbac8921c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31d148),
	.w1(32'hbb076d2a),
	.w2(32'h3b39d4f5),
	.w3(32'hb9d6f21d),
	.w4(32'hbb203b1c),
	.w5(32'h3b8f90c6),
	.w6(32'hbaa29072),
	.w7(32'hbc054874),
	.w8(32'hbaa0c085),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d44d),
	.w1(32'h3b5ed1d7),
	.w2(32'h3ab0e44a),
	.w3(32'hbb70b317),
	.w4(32'h3b16bec0),
	.w5(32'h3a86354b),
	.w6(32'hbba67e64),
	.w7(32'h3b4064f0),
	.w8(32'h3b06d7f2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ae02),
	.w1(32'h3b24d90d),
	.w2(32'h3c1a4a26),
	.w3(32'h3b0219b4),
	.w4(32'h3b95f3a9),
	.w5(32'h3c859dad),
	.w6(32'h3b876df3),
	.w7(32'h3b5afd93),
	.w8(32'h3c0dbdca),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13313f),
	.w1(32'hbb6139c4),
	.w2(32'hbbb75725),
	.w3(32'hbb6e01c7),
	.w4(32'h3b8cb9ae),
	.w5(32'hbb10ca91),
	.w6(32'hbb5993d6),
	.w7(32'hb7e5aa84),
	.w8(32'hb817f333),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9670df),
	.w1(32'hbb4030b4),
	.w2(32'h3a36dee0),
	.w3(32'hbace156a),
	.w4(32'hbad66da7),
	.w5(32'hbaafaf5a),
	.w6(32'h3b25b616),
	.w7(32'hbb4dbc65),
	.w8(32'h3a3ef4c4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7b1c0),
	.w1(32'h3bc3ed54),
	.w2(32'hb94b2093),
	.w3(32'h3b51cfa0),
	.w4(32'hbb3aa766),
	.w5(32'hbb52ea34),
	.w6(32'hba8a4e08),
	.w7(32'hbb589363),
	.w8(32'hbadd015f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e15f2b),
	.w1(32'hb92918eb),
	.w2(32'hbbc49f09),
	.w3(32'hb9bc387e),
	.w4(32'h3b163497),
	.w5(32'hbc049e56),
	.w6(32'hbb4f69b2),
	.w7(32'h3b0d6248),
	.w8(32'hbb5597e3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14e42),
	.w1(32'hbab2f2d9),
	.w2(32'hbaf48362),
	.w3(32'hbb81a900),
	.w4(32'hbabb79cd),
	.w5(32'hbb90edb5),
	.w6(32'hbb5157f5),
	.w7(32'hbae1e2b4),
	.w8(32'hbb777f87),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eda3c),
	.w1(32'h3a9c4232),
	.w2(32'hb910c55e),
	.w3(32'hbadfde82),
	.w4(32'hbb1ecc7a),
	.w5(32'hbb887faa),
	.w6(32'hbaf85bba),
	.w7(32'hbbbe6fbe),
	.w8(32'h3ae5cba2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d5e71),
	.w1(32'hb915dba6),
	.w2(32'hba635bd3),
	.w3(32'h3972308c),
	.w4(32'h3b4a32e4),
	.w5(32'h3b404508),
	.w6(32'hba293937),
	.w7(32'h3b2cc311),
	.w8(32'h398a75cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43ad6d),
	.w1(32'h3ba98def),
	.w2(32'h3b318b66),
	.w3(32'hb7cdf7c9),
	.w4(32'h3b0397d5),
	.w5(32'h3a6d06b5),
	.w6(32'h3af15248),
	.w7(32'hb9487825),
	.w8(32'hbb585e7b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f4e3),
	.w1(32'hbb4c6410),
	.w2(32'hbba352e3),
	.w3(32'hbb832eba),
	.w4(32'h3ab826f4),
	.w5(32'hba1530cd),
	.w6(32'hbaabd330),
	.w7(32'hbb8367bf),
	.w8(32'hbb85489a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4455),
	.w1(32'hba39ac70),
	.w2(32'h3ae7aaed),
	.w3(32'hbb071c22),
	.w4(32'hba490973),
	.w5(32'h3c18ff62),
	.w6(32'hbb075f4b),
	.w7(32'hbac560d4),
	.w8(32'h3a28a4e8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb1c16),
	.w1(32'hbb540736),
	.w2(32'hbb81f272),
	.w3(32'h39d96515),
	.w4(32'hb9e80505),
	.w5(32'h3af2b424),
	.w6(32'h3ad89add),
	.w7(32'hbab66513),
	.w8(32'hbba02c61),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081dea),
	.w1(32'hbb80a511),
	.w2(32'hbb59f94f),
	.w3(32'hbba56c9f),
	.w4(32'h3a0ff71a),
	.w5(32'hbae0c919),
	.w6(32'hbb9697c7),
	.w7(32'hbb5564b5),
	.w8(32'hbaf32746),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c809e),
	.w1(32'hbacfd20b),
	.w2(32'hba85ef57),
	.w3(32'hbb8f7725),
	.w4(32'hbb0f20d5),
	.w5(32'h3b1bb8f7),
	.w6(32'hbb1c1c70),
	.w7(32'h39b89409),
	.w8(32'h3b7d79da),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d53af2),
	.w1(32'hba47ba8c),
	.w2(32'hbb0f2713),
	.w3(32'h3b2903d0),
	.w4(32'hbb74ad94),
	.w5(32'hbb2f4a05),
	.w6(32'h3b874c88),
	.w7(32'hbb64cd91),
	.w8(32'hbb854d99),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d186c),
	.w1(32'h3afb8aee),
	.w2(32'hbac632cd),
	.w3(32'hbbbc7e39),
	.w4(32'h3b8784fe),
	.w5(32'h3bce3df8),
	.w6(32'hbbc9cbe9),
	.w7(32'h3b3c075a),
	.w8(32'hbbed633b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cad73),
	.w1(32'hb9b853c1),
	.w2(32'h3a59cc4c),
	.w3(32'h39ad9927),
	.w4(32'hbbe487c6),
	.w5(32'h3c3a1da4),
	.w6(32'hbaa95a4f),
	.w7(32'hbbfed258),
	.w8(32'hbb67f12c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb713294),
	.w1(32'hbb62210c),
	.w2(32'hbb828171),
	.w3(32'h3ac8e227),
	.w4(32'hbbe22888),
	.w5(32'hbbf5a6b8),
	.w6(32'h3aaff6c2),
	.w7(32'hbbef554a),
	.w8(32'hbbba0348),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f060),
	.w1(32'hbaa8fcd5),
	.w2(32'h3b1c6907),
	.w3(32'hbb57e9d9),
	.w4(32'hbb178630),
	.w5(32'h3b2be478),
	.w6(32'hbb99810a),
	.w7(32'h39fec0b0),
	.w8(32'h3b232b26),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c821c),
	.w1(32'hbad8f724),
	.w2(32'h3ae1a96e),
	.w3(32'h3af458fb),
	.w4(32'hbc0a8359),
	.w5(32'hbb2034f9),
	.w6(32'h3b5f4f32),
	.w7(32'h3ac59c35),
	.w8(32'h3b5c42c8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944c12),
	.w1(32'hba4316ed),
	.w2(32'hbb572962),
	.w3(32'h3a7c5177),
	.w4(32'hbaa4494b),
	.w5(32'h39e2054b),
	.w6(32'hbaa8c8db),
	.w7(32'hbab402ad),
	.w8(32'hb9c617b7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19ce83),
	.w1(32'hbb2d3e3d),
	.w2(32'hbaa40b71),
	.w3(32'h3a91d01d),
	.w4(32'hbbe78d86),
	.w5(32'h3c3b840e),
	.w6(32'h39307504),
	.w7(32'hbb4a70fe),
	.w8(32'h3b3d4d44),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95a73b),
	.w1(32'hbbbb45b8),
	.w2(32'hbc0684db),
	.w3(32'h398c67b2),
	.w4(32'hbb944852),
	.w5(32'hbbd253e1),
	.w6(32'h3bbaa550),
	.w7(32'hbbb4b8e4),
	.w8(32'h3b364f58),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b706f89),
	.w1(32'hbaefb478),
	.w2(32'hb944e998),
	.w3(32'h3bbdc3dc),
	.w4(32'hbb601525),
	.w5(32'h3b0fd788),
	.w6(32'h3ac05f44),
	.w7(32'hbb0f1974),
	.w8(32'h3b42066b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507bf5),
	.w1(32'hb973ec38),
	.w2(32'hb95d9244),
	.w3(32'hbaee16fc),
	.w4(32'hbaaa505a),
	.w5(32'h3b006c6f),
	.w6(32'h3a0bb783),
	.w7(32'h39351aef),
	.w8(32'hbaafbcd3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cb6ea),
	.w1(32'h393811a4),
	.w2(32'h3b15bed6),
	.w3(32'hbbb5f900),
	.w4(32'h3a15dd89),
	.w5(32'h3a1c7a30),
	.w6(32'h3ab87abc),
	.w7(32'h3b50ee0e),
	.w8(32'h3b8b10fa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a915e2f),
	.w1(32'hbb0bafe8),
	.w2(32'hbac11ea7),
	.w3(32'hbb254d7c),
	.w4(32'hbae73fdf),
	.w5(32'hb81c8051),
	.w6(32'h3b94edd0),
	.w7(32'h3b17ed7b),
	.w8(32'hba4694cf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dc833),
	.w1(32'hba4b42e4),
	.w2(32'hbb3e1e9c),
	.w3(32'h3afc0de2),
	.w4(32'hbab92946),
	.w5(32'hbbde13d0),
	.w6(32'hba8fabe2),
	.w7(32'hbb2ae1b3),
	.w8(32'hbbb0ed0e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba779bd),
	.w1(32'h3b1b0abd),
	.w2(32'h3b3fd45b),
	.w3(32'hbbb8cd25),
	.w4(32'h3b3e3d69),
	.w5(32'h38d6c2d5),
	.w6(32'hbb4d06c9),
	.w7(32'hba9ab799),
	.w8(32'h3aa3d7b0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5bbe5),
	.w1(32'h39ae0344),
	.w2(32'hbb4f64ae),
	.w3(32'h3b54400f),
	.w4(32'hb99e52c6),
	.w5(32'hbafb403c),
	.w6(32'h3baf4003),
	.w7(32'h3acdd265),
	.w8(32'hbb962982),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b53b),
	.w1(32'hbaec6515),
	.w2(32'h3a9251d3),
	.w3(32'hba2ec83e),
	.w4(32'hbb4301d9),
	.w5(32'hba57b7b7),
	.w6(32'hbb2b3fdd),
	.w7(32'hbb558fa3),
	.w8(32'h3b157376),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba717d5e),
	.w1(32'hbb070922),
	.w2(32'hbaae8f77),
	.w3(32'hbafe6caf),
	.w4(32'hbb55e35f),
	.w5(32'hbb22a09c),
	.w6(32'hbafa2e1b),
	.w7(32'hbb2e43e5),
	.w8(32'hb99fddb8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2777bf),
	.w1(32'hbbc762ca),
	.w2(32'hbbab7ca8),
	.w3(32'hba20222a),
	.w4(32'hbc0c199e),
	.w5(32'hbb2f2587),
	.w6(32'h3ab1632d),
	.w7(32'hbb06ab70),
	.w8(32'h3a16fc1c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9fdf),
	.w1(32'hba850b95),
	.w2(32'hba48f957),
	.w3(32'h3b5ef6b0),
	.w4(32'hbb3da07f),
	.w5(32'h3b05ff77),
	.w6(32'h3af45fd2),
	.w7(32'hbb282735),
	.w8(32'hbba3ae36),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b1885),
	.w1(32'hbb68c1f6),
	.w2(32'hbae04afb),
	.w3(32'hbaa8a926),
	.w4(32'hbbe8b100),
	.w5(32'h3c3f4504),
	.w6(32'hbb2986d6),
	.w7(32'h3a83c478),
	.w8(32'hbac4482c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb639d94),
	.w1(32'hb8d3959a),
	.w2(32'hbb4d4007),
	.w3(32'h3a0341f9),
	.w4(32'h3b8211d8),
	.w5(32'hbb1f5cb3),
	.w6(32'hba9fecc2),
	.w7(32'h3b0e7cfb),
	.w8(32'hbb4610cf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2199),
	.w1(32'h3b6c84e4),
	.w2(32'hb9006d6d),
	.w3(32'hbc0e7192),
	.w4(32'h3c048745),
	.w5(32'hba848ff7),
	.w6(32'hbbc6e503),
	.w7(32'h3b27f488),
	.w8(32'hbb868084),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be262),
	.w1(32'hbb74e60a),
	.w2(32'hbbd3d5d6),
	.w3(32'h3ae30b0b),
	.w4(32'hbb779b25),
	.w5(32'hbbc8d51c),
	.w6(32'hbb1a405d),
	.w7(32'hba731956),
	.w8(32'hbbca10ad),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de7df9),
	.w1(32'h3aacb943),
	.w2(32'h3abbca35),
	.w3(32'hbb5a674e),
	.w4(32'hbb1a0edb),
	.w5(32'hba82ff32),
	.w6(32'hbb5e0103),
	.w7(32'h3b4e9caf),
	.w8(32'h3a8b3952),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b720884),
	.w1(32'hbb4ab41d),
	.w2(32'hbb72d2be),
	.w3(32'hb988e02a),
	.w4(32'h3c070c4d),
	.w5(32'h395fc5ed),
	.w6(32'h398c57ec),
	.w7(32'hba492ca8),
	.w8(32'hbb78b10d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a5d7),
	.w1(32'hbb2ebbfc),
	.w2(32'h3b66fd5e),
	.w3(32'hbbfb0ffe),
	.w4(32'hbb35f429),
	.w5(32'h3bc59c01),
	.w6(32'hbb469026),
	.w7(32'hbb6adb2f),
	.w8(32'h3ba003a2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb341324),
	.w1(32'h386ddc53),
	.w2(32'hbb8588c7),
	.w3(32'hba8309d6),
	.w4(32'hbb948e7b),
	.w5(32'h3b6bdb51),
	.w6(32'h392ae6fd),
	.w7(32'hba66acf5),
	.w8(32'hbad7f69a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a756bf4),
	.w1(32'hbb37071d),
	.w2(32'hbb9ab769),
	.w3(32'hbb0814ce),
	.w4(32'hb8afc647),
	.w5(32'hbb21edb6),
	.w6(32'h3a152283),
	.w7(32'hbaa17213),
	.w8(32'hbb9ea02f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3c90),
	.w1(32'h3b72794a),
	.w2(32'h39d30f03),
	.w3(32'hbbaadd31),
	.w4(32'h3b6d9dd4),
	.w5(32'h3ac3a33a),
	.w6(32'hbc005320),
	.w7(32'h3b25c029),
	.w8(32'hba0fd63b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404a3f),
	.w1(32'hbaa53f61),
	.w2(32'hbb8adc0b),
	.w3(32'hbaa61e7c),
	.w4(32'hbb85620c),
	.w5(32'hbb884bb3),
	.w6(32'hbb19724a),
	.w7(32'hbaea1257),
	.w8(32'hbb2ce8bf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73cf5b),
	.w1(32'h3b18def8),
	.w2(32'h3b5de315),
	.w3(32'hb778172f),
	.w4(32'h3b24be38),
	.w5(32'h3c12caa0),
	.w6(32'h3a63b812),
	.w7(32'hbad1cc1a),
	.w8(32'h3a0d9b10),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9bc7),
	.w1(32'h3c312b1d),
	.w2(32'hbb6532b3),
	.w3(32'h3b1fda37),
	.w4(32'h3bb131af),
	.w5(32'hbb140199),
	.w6(32'h3a82b3a1),
	.w7(32'h3bced71b),
	.w8(32'hba89c95f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4b835),
	.w1(32'h3aae00a4),
	.w2(32'hbb108b88),
	.w3(32'h39f47398),
	.w4(32'h3ac6d939),
	.w5(32'hb9382451),
	.w6(32'h38e0fee8),
	.w7(32'h3aed083e),
	.w8(32'hba8b5f4d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45b97a),
	.w1(32'h3a94b0b8),
	.w2(32'hba57565b),
	.w3(32'hba9fb13c),
	.w4(32'hbb3c9d60),
	.w5(32'hbb1f7645),
	.w6(32'hbba2e140),
	.w7(32'hbbaea8f2),
	.w8(32'hba6e88a8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c884a),
	.w1(32'hba9c5f6e),
	.w2(32'hba8ab058),
	.w3(32'hba00b6a6),
	.w4(32'hbaa3d88b),
	.w5(32'hba91d516),
	.w6(32'h3921e5cd),
	.w7(32'hbaa68667),
	.w8(32'hba632cff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c5e5a),
	.w1(32'hb9566ff5),
	.w2(32'hb9a5dea2),
	.w3(32'hb949c1a8),
	.w4(32'hba212904),
	.w5(32'hbacaae0a),
	.w6(32'hba02cd42),
	.w7(32'h38f803b4),
	.w8(32'hba1b43bf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978354c),
	.w1(32'h3aad471b),
	.w2(32'h3a9af666),
	.w3(32'hba6083d1),
	.w4(32'h3af71124),
	.w5(32'h3a544f41),
	.w6(32'hb95e3aaa),
	.w7(32'h3b08dc27),
	.w8(32'h3b0212ce),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa33785),
	.w1(32'hb8bb92b0),
	.w2(32'hba74ad09),
	.w3(32'h3a489e48),
	.w4(32'h3a31e7b1),
	.w5(32'h38d5d4d0),
	.w6(32'h3af47764),
	.w7(32'h3a1bdf49),
	.w8(32'hba37d8a6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dd44e),
	.w1(32'hba295644),
	.w2(32'hb947754d),
	.w3(32'h39867bbb),
	.w4(32'hbaab7da3),
	.w5(32'h3a3ab80e),
	.w6(32'hb9bc0c7e),
	.w7(32'hba16f7d2),
	.w8(32'h394881f4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e5c5),
	.w1(32'hb8eebf67),
	.w2(32'hba9a0529),
	.w3(32'h3a984762),
	.w4(32'h3a08a55c),
	.w5(32'h39bf2888),
	.w6(32'hb9a6ec66),
	.w7(32'hb9163992),
	.w8(32'hbafa6c7d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64ce21),
	.w1(32'h3908b10f),
	.w2(32'hbb8320b5),
	.w3(32'hbaab6b22),
	.w4(32'h3ac79df8),
	.w5(32'h3a98c844),
	.w6(32'hbac1ad2d),
	.w7(32'h3ac90922),
	.w8(32'hbab7ef4e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38868467),
	.w1(32'h3a03f585),
	.w2(32'h3a329141),
	.w3(32'h3995e539),
	.w4(32'h39ceff28),
	.w5(32'hb98bebb9),
	.w6(32'h38aae8c5),
	.w7(32'h3a8b8d39),
	.w8(32'h3adc5f61),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933a5f),
	.w1(32'hbb0540a0),
	.w2(32'hba470b9d),
	.w3(32'h38f1f18e),
	.w4(32'hbaa3ca2a),
	.w5(32'hb8eab148),
	.w6(32'hb97b251b),
	.w7(32'hba7ef4b4),
	.w8(32'h3a08997f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48970),
	.w1(32'h396be8a7),
	.w2(32'hb98cd7c3),
	.w3(32'h3a53c04b),
	.w4(32'h3a588ac8),
	.w5(32'h3ac55333),
	.w6(32'hba970281),
	.w7(32'hbb1a96b8),
	.w8(32'hbb2f398e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbfb64),
	.w1(32'h3a33e384),
	.w2(32'h39d7f484),
	.w3(32'h3983fcdf),
	.w4(32'h3a7be494),
	.w5(32'h3a592361),
	.w6(32'h39be424e),
	.w7(32'h39a35179),
	.w8(32'h3aa7b01a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa258a5),
	.w1(32'hb9f52438),
	.w2(32'hbafca12d),
	.w3(32'h3a92d12c),
	.w4(32'hb8d2531c),
	.w5(32'hba979ee9),
	.w6(32'h3adbd090),
	.w7(32'h3a4d787b),
	.w8(32'hba98c158),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ea3db),
	.w1(32'h3a12bbb5),
	.w2(32'hb78f57c1),
	.w3(32'hb9dc72a2),
	.w4(32'h36e05240),
	.w5(32'hb97f809a),
	.w6(32'hb912697c),
	.w7(32'hb87e6d31),
	.w8(32'hb9e82119),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e136b3),
	.w1(32'h3a1a2ca0),
	.w2(32'hb90341c4),
	.w3(32'hba123e95),
	.w4(32'h39097dcd),
	.w5(32'hba7385b5),
	.w6(32'hb9a67843),
	.w7(32'hb9c1424a),
	.w8(32'h3a7ee762),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d5048),
	.w1(32'hb9da7b6e),
	.w2(32'hba43b3d0),
	.w3(32'h39c25f75),
	.w4(32'hba1671c7),
	.w5(32'hba807682),
	.w6(32'h3a54aac3),
	.w7(32'h39b2ca75),
	.w8(32'hb98da304),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939f385),
	.w1(32'h3a64f500),
	.w2(32'hb91848f8),
	.w3(32'hba6f0152),
	.w4(32'hba24506c),
	.w5(32'h3704647e),
	.w6(32'hb9ea0790),
	.w7(32'hb9cc6bd4),
	.w8(32'hba77c305),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39d2ac),
	.w1(32'h3ab03983),
	.w2(32'h3a64e0c1),
	.w3(32'hbaf2626b),
	.w4(32'hb845222d),
	.w5(32'hb81cd6a5),
	.w6(32'hbaee1837),
	.w7(32'hbab14ca2),
	.w8(32'h378c690a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f83ea6),
	.w1(32'h3a8c963f),
	.w2(32'h3a6d5873),
	.w3(32'h3a2ff251),
	.w4(32'h3a4d9226),
	.w5(32'hbac23e3f),
	.w6(32'h38e17e68),
	.w7(32'h3a75eaa4),
	.w8(32'h3a07a84c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb806f96c),
	.w1(32'hba3908bf),
	.w2(32'h37f96d71),
	.w3(32'h3893842a),
	.w4(32'hb994c6b3),
	.w5(32'h38b4493d),
	.w6(32'hbabb77a6),
	.w7(32'hbb08ca67),
	.w8(32'h3974a513),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6ed55),
	.w1(32'hb9a3749b),
	.w2(32'hb9ac24a8),
	.w3(32'hba2ec736),
	.w4(32'h3ac8ad90),
	.w5(32'h3a514aca),
	.w6(32'hb9607b4c),
	.w7(32'h39ae7b7a),
	.w8(32'hbaccf519),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ce844),
	.w1(32'hb9d06125),
	.w2(32'hba15336a),
	.w3(32'h3a2bc6ad),
	.w4(32'hbac510eb),
	.w5(32'hb9fde92c),
	.w6(32'h3a19e35d),
	.w7(32'hbabc674c),
	.w8(32'hba794cbd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad71c7f),
	.w1(32'hba1ef2e6),
	.w2(32'hbb84a6ac),
	.w3(32'h3a1b0611),
	.w4(32'h3b95bd86),
	.w5(32'hb91c1830),
	.w6(32'h3a896fef),
	.w7(32'hbaee0331),
	.w8(32'hbb1a68aa),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d9f6d),
	.w1(32'h39d946b8),
	.w2(32'h39afc654),
	.w3(32'hba069ac8),
	.w4(32'hb9b9c058),
	.w5(32'hba1fc476),
	.w6(32'hbb24bd8d),
	.w7(32'hba810a4a),
	.w8(32'hba7a5c04),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51cbca),
	.w1(32'hbb57193c),
	.w2(32'hba7006fc),
	.w3(32'hba28acdb),
	.w4(32'hb96b9eb7),
	.w5(32'h3ae865e2),
	.w6(32'hba423443),
	.w7(32'hbaa1659a),
	.w8(32'h3a6e2aba),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efd81a),
	.w1(32'hbabe4d50),
	.w2(32'hb98f310e),
	.w3(32'h393cad08),
	.w4(32'hba4891f8),
	.w5(32'h3b100a34),
	.w6(32'hb8ea4118),
	.w7(32'hba7fad6a),
	.w8(32'h3a8e3caf),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc3cc0),
	.w1(32'h39d0a996),
	.w2(32'hb99af446),
	.w3(32'hba4907c9),
	.w4(32'hba934759),
	.w5(32'h3a055408),
	.w6(32'hbaf27b07),
	.w7(32'hbace3dd3),
	.w8(32'hba10c9f6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913c080),
	.w1(32'hb9aeb04f),
	.w2(32'hb9b9aa97),
	.w3(32'hba07c2cd),
	.w4(32'hb8ae85d7),
	.w5(32'h39506191),
	.w6(32'hba56d3aa),
	.w7(32'hba453981),
	.w8(32'hba5ed456),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf8ec),
	.w1(32'hb94e1d1c),
	.w2(32'hbb13fae6),
	.w3(32'hba6b73fe),
	.w4(32'h3a1becad),
	.w5(32'hba777782),
	.w6(32'hb88b1cb3),
	.w7(32'h3a0c59ea),
	.w8(32'hbabb9566),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86dfe7),
	.w1(32'hb9ac7fde),
	.w2(32'hbafac105),
	.w3(32'h3aae824e),
	.w4(32'h3b03fb5d),
	.w5(32'h39b1b9c4),
	.w6(32'h3ab480f5),
	.w7(32'hbad913a9),
	.w8(32'hbb3dfc51),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc144b8d),
	.w1(32'h3a8f7730),
	.w2(32'hbac8f33f),
	.w3(32'hbc2c3711),
	.w4(32'h3b3c4155),
	.w5(32'h390477ae),
	.w6(32'hbbcf1207),
	.w7(32'h3b4973f5),
	.w8(32'h3a09afac),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30dd0),
	.w1(32'hba1a9165),
	.w2(32'hb76a9cba),
	.w3(32'hbbb5d40a),
	.w4(32'hbb0e44df),
	.w5(32'hba508099),
	.w6(32'hbbbe76bc),
	.w7(32'hbb75b054),
	.w8(32'h3a789692),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d27e5),
	.w1(32'h3a806ee9),
	.w2(32'hb8c44c7f),
	.w3(32'h3a228db5),
	.w4(32'h3a9d1d8b),
	.w5(32'hba9a9e36),
	.w6(32'hbb031228),
	.w7(32'hb871a81a),
	.w8(32'h3a9cbe35),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92aac7),
	.w1(32'h3b1b0ab3),
	.w2(32'h3abcf650),
	.w3(32'hbb7eda53),
	.w4(32'h3bd82256),
	.w5(32'h3a5e8220),
	.w6(32'hbac8861f),
	.w7(32'h3b692b8e),
	.w8(32'hbb7463c3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc5b3b),
	.w1(32'hb8e535e9),
	.w2(32'hbac948c0),
	.w3(32'hbaa539fa),
	.w4(32'hb9cbd417),
	.w5(32'hbae7160a),
	.w6(32'hba4e3667),
	.w7(32'hb988dbe4),
	.w8(32'h37b0b365),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3be383),
	.w1(32'hba08ecf2),
	.w2(32'hbb215107),
	.w3(32'hbc260f62),
	.w4(32'h3ac46593),
	.w5(32'h38afba9c),
	.w6(32'hbc0d3528),
	.w7(32'h3b8a400e),
	.w8(32'hbace4646),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36241e),
	.w1(32'h3a9f46e5),
	.w2(32'hbb0a1160),
	.w3(32'h3b08a70b),
	.w4(32'h39b0918e),
	.w5(32'hbb0d3a7c),
	.w6(32'h3a812f86),
	.w7(32'h3ac25adb),
	.w8(32'hbb2d7665),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39854bd0),
	.w1(32'h39c04cd3),
	.w2(32'hb9d90efd),
	.w3(32'hb6fe66d7),
	.w4(32'h398d0253),
	.w5(32'h37c926d7),
	.w6(32'h3a2065d5),
	.w7(32'h3a13925e),
	.w8(32'h3a237018),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7159309),
	.w1(32'hb9cd7675),
	.w2(32'hba65fa08),
	.w3(32'h3a00797f),
	.w4(32'h38f57e36),
	.w5(32'hb9797d5e),
	.w6(32'hba78e037),
	.w7(32'hbae6a3c8),
	.w8(32'hba051c39),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b7d4b),
	.w1(32'h3a9a69c7),
	.w2(32'hba64bb99),
	.w3(32'h3a9efd46),
	.w4(32'h3b357eee),
	.w5(32'hba8fba6c),
	.w6(32'h3ae16e50),
	.w7(32'h3adbbef0),
	.w8(32'h39041ddc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba812965),
	.w1(32'hba071fab),
	.w2(32'hbaaff1fa),
	.w3(32'hb901d405),
	.w4(32'hba2b8266),
	.w5(32'hb9ea7f39),
	.w6(32'h3a397991),
	.w7(32'hba9cd0cd),
	.w8(32'hb9d973fe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23e6cc),
	.w1(32'hbb207fb1),
	.w2(32'hbae264d5),
	.w3(32'h3a472951),
	.w4(32'hbac20fd8),
	.w5(32'hbaa82980),
	.w6(32'h3a592417),
	.w7(32'hb9ed3075),
	.w8(32'hb8c0ff1c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c7d2e),
	.w1(32'hb92d4c1f),
	.w2(32'h3a50e9c0),
	.w3(32'hbaf7bc69),
	.w4(32'hb7aae3bf),
	.w5(32'h3ab62e39),
	.w6(32'hbae3e9ce),
	.w7(32'hb89f9f03),
	.w8(32'h3a015193),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8556bc),
	.w1(32'h3baa9e9f),
	.w2(32'h3aeaf962),
	.w3(32'h39bb87da),
	.w4(32'h3b8713b8),
	.w5(32'h3adc44da),
	.w6(32'hb8a51d2b),
	.w7(32'h3b3edf37),
	.w8(32'h3aef3ace),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacce6bd),
	.w1(32'hbb1c264b),
	.w2(32'hbac2ee9a),
	.w3(32'hbac22283),
	.w4(32'hba48a757),
	.w5(32'h3b52f488),
	.w6(32'hb9163d36),
	.w7(32'hbaf1f6ab),
	.w8(32'h3b208956),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca820e),
	.w1(32'h399768d2),
	.w2(32'hba185d2c),
	.w3(32'h39496038),
	.w4(32'h3a35ee5b),
	.w5(32'hba569ab4),
	.w6(32'hb9b58ad9),
	.w7(32'h399ce8a1),
	.w8(32'hba3e3ac2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba093a3c),
	.w1(32'hb9b4f85f),
	.w2(32'hb9dacac4),
	.w3(32'hba7a77b1),
	.w4(32'hba3e3736),
	.w5(32'hba0a3d93),
	.w6(32'hba8be071),
	.w7(32'hb9f74af4),
	.w8(32'hba087ecb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba436ced),
	.w1(32'h383bc85c),
	.w2(32'hb9914d82),
	.w3(32'hba364716),
	.w4(32'h38960536),
	.w5(32'h3a49b1db),
	.w6(32'hb9be5903),
	.w7(32'h3a2d9437),
	.w8(32'h39a4eaf5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ead3b1),
	.w1(32'h39569d4d),
	.w2(32'hba10e351),
	.w3(32'h39b32a9c),
	.w4(32'h372e439b),
	.w5(32'hb9e30e22),
	.w6(32'h39f8a8a1),
	.w7(32'hba3099e5),
	.w8(32'hba50a135),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f024),
	.w1(32'h3a862cd5),
	.w2(32'h3a8e3e5d),
	.w3(32'hba611240),
	.w4(32'h3ad7828a),
	.w5(32'hb962e06e),
	.w6(32'hba2cee44),
	.w7(32'h3a8082b3),
	.w8(32'h39bcc3a3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981d001),
	.w1(32'h39a00253),
	.w2(32'h384d7631),
	.w3(32'h3aa75b01),
	.w4(32'h39cfce90),
	.w5(32'h392044b6),
	.w6(32'h3a396989),
	.w7(32'hb84f7734),
	.w8(32'h3998d3c0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f736fa),
	.w1(32'hba3c0bdb),
	.w2(32'hba84d05c),
	.w3(32'hba6a7d4d),
	.w4(32'hba2248f3),
	.w5(32'hb9926b42),
	.w6(32'hb82f55e8),
	.w7(32'hba05b301),
	.w8(32'hba3e6280),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b99c1d),
	.w1(32'hb781a548),
	.w2(32'hba6e72fc),
	.w3(32'h3a6c363c),
	.w4(32'h3b11744b),
	.w5(32'h39728d94),
	.w6(32'h39b8325f),
	.w7(32'hb9f7881c),
	.w8(32'hb9984214),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f6e1),
	.w1(32'h3ab1f69c),
	.w2(32'h3aea3ff0),
	.w3(32'h3aabada5),
	.w4(32'hbb1d1175),
	.w5(32'hb96ea67f),
	.w6(32'hbb07f586),
	.w7(32'hbb7b419c),
	.w8(32'hba890f10),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cf80c),
	.w1(32'hba2d5957),
	.w2(32'hb991118e),
	.w3(32'hb95e57aa),
	.w4(32'h38eed070),
	.w5(32'h3a382ad0),
	.w6(32'hba11c8c5),
	.w7(32'hb9866015),
	.w8(32'hb7a33acc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34c4ce),
	.w1(32'h3a31581a),
	.w2(32'hb9f3ab38),
	.w3(32'h39f563de),
	.w4(32'hb9bd224f),
	.w5(32'hbad665da),
	.w6(32'hb9bd0596),
	.w7(32'hb987de4d),
	.w8(32'hba967b1e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d1f5d),
	.w1(32'hba8da0f8),
	.w2(32'hb9e28d90),
	.w3(32'hb999cbf8),
	.w4(32'hb9faccec),
	.w5(32'hba580052),
	.w6(32'hb9f42954),
	.w7(32'hba87a9cc),
	.w8(32'hba88307c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e3e51),
	.w1(32'hbb0eabb2),
	.w2(32'hbae6c584),
	.w3(32'hba642e0c),
	.w4(32'hbb136098),
	.w5(32'hba9a1e3a),
	.w6(32'hba69d36e),
	.w7(32'hbaa84dce),
	.w8(32'hba1f8745),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4936bc),
	.w1(32'h3b68d739),
	.w2(32'hbb485701),
	.w3(32'hb9f0f699),
	.w4(32'hb9645408),
	.w5(32'hbb753dc5),
	.w6(32'h3a0ea067),
	.w7(32'hba9c6419),
	.w8(32'hba98eb73),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba567b05),
	.w1(32'hbac912b0),
	.w2(32'hbb0e8085),
	.w3(32'h3ab3ebdd),
	.w4(32'hba7a4b39),
	.w5(32'hbb0ecc05),
	.w6(32'h3a9d7f53),
	.w7(32'hbae9be54),
	.w8(32'hbaf56344),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb6bb7),
	.w1(32'hb9d77694),
	.w2(32'hb9c2c140),
	.w3(32'hb987205a),
	.w4(32'h3a536b92),
	.w5(32'h39dc80bd),
	.w6(32'h3a4339ee),
	.w7(32'h3938bb16),
	.w8(32'hb71098ff),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba554e38),
	.w1(32'h39cd1174),
	.w2(32'hba2dab70),
	.w3(32'hba503ef5),
	.w4(32'hb90c9c77),
	.w5(32'hba65ee77),
	.w6(32'hbaa47abc),
	.w7(32'hba053681),
	.w8(32'hbac15e24),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6dc79),
	.w1(32'h379c8d13),
	.w2(32'h39c5daa7),
	.w3(32'hb9b4e137),
	.w4(32'h38ad439d),
	.w5(32'h3a2a97c8),
	.w6(32'hba3c0d1a),
	.w7(32'hba50da5a),
	.w8(32'hba0264d4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70da89),
	.w1(32'hbaab387b),
	.w2(32'hba277e41),
	.w3(32'hba2e167f),
	.w4(32'h39bd37d0),
	.w5(32'h3a209be6),
	.w6(32'h3915a739),
	.w7(32'h396255e3),
	.w8(32'h3a26e899),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf7ca1),
	.w1(32'hbb37cc6d),
	.w2(32'hba355c23),
	.w3(32'hb9b616bb),
	.w4(32'hba79986c),
	.w5(32'h3af2e334),
	.w6(32'hba1854c0),
	.w7(32'hb9f655cd),
	.w8(32'h3af8c00d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06cfbd),
	.w1(32'hb88f6216),
	.w2(32'hbad6e87a),
	.w3(32'hba72a621),
	.w4(32'h3b030a6f),
	.w5(32'hbaa7115d),
	.w6(32'hb92b3b89),
	.w7(32'hb99a0e7d),
	.w8(32'hbab4c05f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934442b),
	.w1(32'h3a792f87),
	.w2(32'h3abf6f54),
	.w3(32'hba32caf0),
	.w4(32'h38aa6f85),
	.w5(32'h39983ed9),
	.w6(32'hba788a4e),
	.w7(32'hba3f136a),
	.w8(32'h39bb1dce),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa96999),
	.w1(32'hba05e901),
	.w2(32'hbb15e61d),
	.w3(32'hbaa8fe6d),
	.w4(32'h3a628c01),
	.w5(32'hba6cb4b3),
	.w6(32'hba475061),
	.w7(32'hb9f052a7),
	.w8(32'hba28407f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba644b45),
	.w1(32'hba2cad73),
	.w2(32'hbaad72c4),
	.w3(32'hba575429),
	.w4(32'h3a886539),
	.w5(32'hba4af4f7),
	.w6(32'hb95554e5),
	.w7(32'h394676e5),
	.w8(32'hbacfa615),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bc862),
	.w1(32'h3a8d06b3),
	.w2(32'h39c30f3c),
	.w3(32'hb9dc1755),
	.w4(32'h3913ee80),
	.w5(32'h3a096e0a),
	.w6(32'hba69e3d1),
	.w7(32'h3a1582d9),
	.w8(32'h3b1a412b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bc671),
	.w1(32'hb6800ccd),
	.w2(32'hb99c4047),
	.w3(32'h38ab9457),
	.w4(32'h3a82b45c),
	.w5(32'h3a39f2bd),
	.w6(32'hb9123638),
	.w7(32'h39c3f138),
	.w8(32'hba64869d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991b7a4),
	.w1(32'hb9de0489),
	.w2(32'hba78943f),
	.w3(32'hb9aaedc9),
	.w4(32'hb9d0fdea),
	.w5(32'hb9b0222d),
	.w6(32'hb732c256),
	.w7(32'hb9bc2102),
	.w8(32'hb892465b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42179),
	.w1(32'h3aaabb29),
	.w2(32'h3ae73a22),
	.w3(32'hb9518f2e),
	.w4(32'hbb368873),
	.w5(32'hbaea6e6b),
	.w6(32'hba5becff),
	.w7(32'hbb56b8b4),
	.w8(32'hbae93d2f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31ff9e),
	.w1(32'hb97602bb),
	.w2(32'hba9fa65a),
	.w3(32'hba3d3c05),
	.w4(32'hb8d8ee26),
	.w5(32'h39d7d53d),
	.w6(32'hba98d1d3),
	.w7(32'hb9784774),
	.w8(32'hb993f54b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c30588),
	.w1(32'h39abdbbb),
	.w2(32'hb96acae7),
	.w3(32'hba66c4a7),
	.w4(32'hb875cfc3),
	.w5(32'hba0fc14a),
	.w6(32'hb96d6102),
	.w7(32'hb9dd4da8),
	.w8(32'hb9eff8ef),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29d8a9),
	.w1(32'hb9d796e7),
	.w2(32'hb7c755ac),
	.w3(32'h3932be4d),
	.w4(32'hba2d25da),
	.w5(32'hb9707b3c),
	.w6(32'h398a299d),
	.w7(32'h380a40cc),
	.w8(32'hb9e43383),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae7aec),
	.w1(32'h3a2edb37),
	.w2(32'h3a5a0437),
	.w3(32'h380c09ff),
	.w4(32'h3a82fe67),
	.w5(32'h39f2dc12),
	.w6(32'hb98d587f),
	.w7(32'h39c96ab6),
	.w8(32'hb9830055),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77c7a3),
	.w1(32'hba1a8a22),
	.w2(32'hb93d4017),
	.w3(32'hbaa7dfe1),
	.w4(32'hba8757a8),
	.w5(32'h397635e1),
	.w6(32'hbb18aab9),
	.w7(32'hbb13fd55),
	.w8(32'hbad99734),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b0bc0a),
	.w1(32'hbb25bc19),
	.w2(32'hbb5d6fdb),
	.w3(32'h3a8e6f79),
	.w4(32'hba6ac7ca),
	.w5(32'hbaa5b566),
	.w6(32'h3aaf44b2),
	.w7(32'hb9a233d4),
	.w8(32'hba7fdab6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97711a9),
	.w1(32'hba02679f),
	.w2(32'hba39ec8a),
	.w3(32'h3a0de5cb),
	.w4(32'hb9bbe0bd),
	.w5(32'hb8b481f6),
	.w6(32'h3aa1dd9b),
	.w7(32'h380f5658),
	.w8(32'h39a5b5f8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee0b7f),
	.w1(32'hba3c9407),
	.w2(32'hbb541965),
	.w3(32'h394224ee),
	.w4(32'h38da4fc1),
	.w5(32'hbb0cb211),
	.w6(32'hba22f945),
	.w7(32'hba392dc7),
	.w8(32'hbada0145),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b350),
	.w1(32'hb9923f71),
	.w2(32'h3952c52c),
	.w3(32'hb81efe7c),
	.w4(32'h3a30165f),
	.w5(32'hb96cf530),
	.w6(32'h39b8f55c),
	.w7(32'hb8f78c7f),
	.w8(32'h3888cc41),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38765a25),
	.w1(32'hbaa2f66f),
	.w2(32'hbb597fbc),
	.w3(32'h3ae276fa),
	.w4(32'h3b7dba18),
	.w5(32'h3a14f4af),
	.w6(32'h39d6591b),
	.w7(32'h39f3e354),
	.w8(32'hbaee4e76),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b628),
	.w1(32'hb9abcbb5),
	.w2(32'h3a25cf1e),
	.w3(32'h3b816e5d),
	.w4(32'hba2e9d2d),
	.w5(32'hb9905a77),
	.w6(32'h3a357f4a),
	.w7(32'hbad1e28f),
	.w8(32'hba3794b0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3f238),
	.w1(32'hbb1528b3),
	.w2(32'hbb039455),
	.w3(32'hba286644),
	.w4(32'hbb1c3f8c),
	.w5(32'hba98d98f),
	.w6(32'hbab3e1fb),
	.w7(32'hbb29e8c9),
	.w8(32'hbad68ec9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada0878),
	.w1(32'h39e6d0a7),
	.w2(32'hb97212e2),
	.w3(32'hbae11ec9),
	.w4(32'h375b2a07),
	.w5(32'h3938dea3),
	.w6(32'hbaeb83a5),
	.w7(32'h396b5aba),
	.w8(32'h39f5d4ad),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9267b4a),
	.w1(32'h3ac70b28),
	.w2(32'h3b0b3d4d),
	.w3(32'h390cee3c),
	.w4(32'h3a5a9f6f),
	.w5(32'h3ac94aa4),
	.w6(32'hba07343a),
	.w7(32'h3a3b6486),
	.w8(32'h3b0b4a54),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacba2f0),
	.w1(32'hbb108725),
	.w2(32'hb991f4f7),
	.w3(32'h3669a8f8),
	.w4(32'hba75cdbc),
	.w5(32'h39f03b7b),
	.w6(32'h3a22263d),
	.w7(32'hba7e3893),
	.w8(32'h3a39ab30),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addd38f),
	.w1(32'h3a961428),
	.w2(32'h3ab935d1),
	.w3(32'h3a03299c),
	.w4(32'hb90216f6),
	.w5(32'h3a59b6bd),
	.w6(32'hb8d10b59),
	.w7(32'hb92fe4bf),
	.w8(32'h39f8e6ea),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7693da8),
	.w1(32'hba444136),
	.w2(32'hb931b2fe),
	.w3(32'h39114df3),
	.w4(32'h3a34bd04),
	.w5(32'h3a5c9a6b),
	.w6(32'h390acf10),
	.w7(32'h3a6b9e8e),
	.w8(32'h3a443c6f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d90572),
	.w1(32'h39b55cee),
	.w2(32'h3a0c375f),
	.w3(32'h3a7e499c),
	.w4(32'h398ce6c3),
	.w5(32'h39fd420e),
	.w6(32'h3a8a3481),
	.w7(32'h3a1b5c96),
	.w8(32'h3990a6b2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2794c6),
	.w1(32'h3aa731cc),
	.w2(32'hb95588e9),
	.w3(32'hb95eb658),
	.w4(32'h3ae6a753),
	.w5(32'hb918abf4),
	.w6(32'hb934e292),
	.w7(32'h3a67f596),
	.w8(32'hba2cb07c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f7976),
	.w1(32'h3997a905),
	.w2(32'hb9c469eb),
	.w3(32'h3ab1a1e4),
	.w4(32'h3a157c7a),
	.w5(32'hbac70dd8),
	.w6(32'h3a2605dd),
	.w7(32'h39c6aa47),
	.w8(32'hba2b4b20),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ab9cd),
	.w1(32'h3a3bacdc),
	.w2(32'h39ab1405),
	.w3(32'hb8612ce8),
	.w4(32'hbac0dfb0),
	.w5(32'hba6f89c1),
	.w6(32'hba2c5bab),
	.w7(32'hbaf53bb6),
	.w8(32'hb9f46ed9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5472cc),
	.w1(32'h3a5c8163),
	.w2(32'h37e36d3d),
	.w3(32'hbabb8a41),
	.w4(32'hb787b3c4),
	.w5(32'hba303182),
	.w6(32'hb9d4a95b),
	.w7(32'hb98ed104),
	.w8(32'hb9fba52c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba29b8e),
	.w1(32'h3b4e20e4),
	.w2(32'h3a4f4fe8),
	.w3(32'h3aa6f825),
	.w4(32'hbb041fe2),
	.w5(32'hbac533e4),
	.w6(32'h3a74c357),
	.w7(32'hbadc20f0),
	.w8(32'hbad04b25),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a435117),
	.w1(32'h3a0d6018),
	.w2(32'h3907368d),
	.w3(32'h3a407486),
	.w4(32'h3a0a4cfa),
	.w5(32'hb8436159),
	.w6(32'h39a64b83),
	.w7(32'h3a83b5e5),
	.w8(32'h3a41eff1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398133af),
	.w1(32'h38cc5692),
	.w2(32'hb9ad9ac3),
	.w3(32'hb9577945),
	.w4(32'h3a31dec9),
	.w5(32'h3a338883),
	.w6(32'h39d97699),
	.w7(32'h3a69f8d5),
	.w8(32'hb97e15d1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88eba64),
	.w1(32'hba30bc87),
	.w2(32'h38a337b5),
	.w3(32'hba8574cd),
	.w4(32'hba223870),
	.w5(32'h3a23832d),
	.w6(32'hba1d5003),
	.w7(32'hba6b12f6),
	.w8(32'h39ab7c47),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad1c1c),
	.w1(32'h3b14a619),
	.w2(32'hbb023397),
	.w3(32'hbb08f79d),
	.w4(32'h3adbe9fa),
	.w5(32'hb9bd2d6c),
	.w6(32'hba773efa),
	.w7(32'h3ab71a8e),
	.w8(32'hba128413),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c9a1c),
	.w1(32'h3a69fe52),
	.w2(32'h3a67ecfa),
	.w3(32'hba49aa63),
	.w4(32'h3a40a787),
	.w5(32'h3a692877),
	.w6(32'hba721142),
	.w7(32'h38ec5ed4),
	.w8(32'h393a354e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3674917f),
	.w1(32'hba492053),
	.w2(32'hb8082fdd),
	.w3(32'hba50215a),
	.w4(32'hbab445bd),
	.w5(32'hba7857f9),
	.w6(32'h39dcb843),
	.w7(32'hba5b8266),
	.w8(32'hba0dbb19),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e1feb),
	.w1(32'hb987f3ba),
	.w2(32'hb9dc8ad9),
	.w3(32'hb9270bdb),
	.w4(32'hb9b322d6),
	.w5(32'h395731d9),
	.w6(32'hba0a83a8),
	.w7(32'hba156150),
	.w8(32'hb8a53c38),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6e16),
	.w1(32'hbb6f6cad),
	.w2(32'hbb4ca093),
	.w3(32'h3a8e6b6d),
	.w4(32'hba575a7c),
	.w5(32'hba95501e),
	.w6(32'h3b0328d2),
	.w7(32'hbacef4a6),
	.w8(32'hb93b591f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab754a4),
	.w1(32'hbb016420),
	.w2(32'hba07363e),
	.w3(32'hb91fbd24),
	.w4(32'hb9f3e025),
	.w5(32'h399b8882),
	.w6(32'hb95813d8),
	.w7(32'hba47909c),
	.w8(32'h3a4a956c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27d588),
	.w1(32'hbb155224),
	.w2(32'hbb312df1),
	.w3(32'hbabf25d3),
	.w4(32'hbab5b587),
	.w5(32'hbb263400),
	.w6(32'h3a952747),
	.w7(32'hb861a092),
	.w8(32'hba346320),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d3708),
	.w1(32'h3aa8f177),
	.w2(32'h3a3b7963),
	.w3(32'hba6b33c9),
	.w4(32'h3a59ba06),
	.w5(32'h39b8b930),
	.w6(32'hba0b20df),
	.w7(32'h3a85661c),
	.w8(32'h3a92c01c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a5d51),
	.w1(32'hba809c2f),
	.w2(32'hba5eab63),
	.w3(32'hba3aed23),
	.w4(32'hba0e620f),
	.w5(32'h3a0e07bd),
	.w6(32'h3935f853),
	.w7(32'hb92c8a82),
	.w8(32'h3a96cbd0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b1906),
	.w1(32'h39db8b12),
	.w2(32'h3a2b0215),
	.w3(32'hb81c444e),
	.w4(32'hba5acc8c),
	.w5(32'hb9aaff18),
	.w6(32'hb9af33f5),
	.w7(32'h39a65997),
	.w8(32'h391aca85),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f30fb5),
	.w1(32'hb8ede758),
	.w2(32'h3a019129),
	.w3(32'h3a570d78),
	.w4(32'h3a9a4189),
	.w5(32'h39d2ce37),
	.w6(32'h3a398ba2),
	.w7(32'hb7229c81),
	.w8(32'h39448cd4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13114a),
	.w1(32'h3acfda58),
	.w2(32'hb9d11824),
	.w3(32'hba0fa303),
	.w4(32'h39f541ae),
	.w5(32'hba0ce090),
	.w6(32'hba8eef4d),
	.w7(32'h39aa0cc4),
	.w8(32'hba3d1120),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51e260),
	.w1(32'hba546bb4),
	.w2(32'h3a8408ea),
	.w3(32'hba05d476),
	.w4(32'h3a30a15d),
	.w5(32'h3ae884d5),
	.w6(32'h38202c5d),
	.w7(32'h39376ae2),
	.w8(32'h3b1374f0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf2aa3),
	.w1(32'h39be9830),
	.w2(32'h3662c4a3),
	.w3(32'h3a0e9139),
	.w4(32'h3a820573),
	.w5(32'hb9f1733a),
	.w6(32'h3782d45c),
	.w7(32'h3a87f979),
	.w8(32'h3a13a8cc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5085e1),
	.w1(32'hb982cdc3),
	.w2(32'h3a1c26a7),
	.w3(32'hb894b6b5),
	.w4(32'hba3fa197),
	.w5(32'hb981ced2),
	.w6(32'hba31a35a),
	.w7(32'hb8ac6b23),
	.w8(32'hb9c67813),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af681ab),
	.w1(32'h39da70d0),
	.w2(32'h39425d46),
	.w3(32'h3a8408c9),
	.w4(32'hba0830f5),
	.w5(32'h388f9b9f),
	.w6(32'hb93abe09),
	.w7(32'hbaa96c8d),
	.w8(32'h3b0a3347),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f0716),
	.w1(32'hba6206ad),
	.w2(32'hba9d417e),
	.w3(32'hba9d9470),
	.w4(32'h3b39c9af),
	.w5(32'h3ab0a6b9),
	.w6(32'h3a5d61c0),
	.w7(32'hba28af40),
	.w8(32'hba86df96),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec862),
	.w1(32'h3ac61036),
	.w2(32'hb712ffce),
	.w3(32'hbb90b9dc),
	.w4(32'h3aff2ff1),
	.w5(32'h3aad7983),
	.w6(32'hbba68d6a),
	.w7(32'h3af006c0),
	.w8(32'hbb2389ba),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d0021),
	.w1(32'hbaceb8a5),
	.w2(32'hb9a2bfaf),
	.w3(32'hba4ac9a9),
	.w4(32'hba6ccdf9),
	.w5(32'hba67ec1b),
	.w6(32'hba34a699),
	.w7(32'hbaa116e2),
	.w8(32'hba856d2c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978fbee),
	.w1(32'hbb0647d6),
	.w2(32'hbb551a28),
	.w3(32'h3a81dace),
	.w4(32'hbae1eb20),
	.w5(32'hbb4c24c1),
	.w6(32'h3b6239bf),
	.w7(32'hba07cf18),
	.w8(32'hbb70ad66),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cfbf8),
	.w1(32'hbb3ddfd7),
	.w2(32'hbafd6098),
	.w3(32'h3b1cf923),
	.w4(32'hbb2f0846),
	.w5(32'hba13bd55),
	.w6(32'h3a347cbf),
	.w7(32'hbb3c8221),
	.w8(32'h3a6cbf66),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3634a),
	.w1(32'h3a60a8da),
	.w2(32'hba3db351),
	.w3(32'hba8d320b),
	.w4(32'h3a8e47d9),
	.w5(32'h3a521bb1),
	.w6(32'hbac1cff1),
	.w7(32'hb9b40548),
	.w8(32'hbaeb0a18),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee9c46),
	.w1(32'hb9b28904),
	.w2(32'h374917e0),
	.w3(32'hb9e8f708),
	.w4(32'h39bbd65e),
	.w5(32'h3987d204),
	.w6(32'h3997f6cd),
	.w7(32'hba313b21),
	.w8(32'hba03f05e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900f877),
	.w1(32'hba3fefe1),
	.w2(32'h398f1c82),
	.w3(32'h38861e35),
	.w4(32'hba129f9e),
	.w5(32'h398126f1),
	.w6(32'h39107631),
	.w7(32'hb9dbe4de),
	.w8(32'h388ef561),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9793b86),
	.w1(32'h3a87f34e),
	.w2(32'h3a4ae20e),
	.w3(32'h397f4c81),
	.w4(32'h3a2064ea),
	.w5(32'h3a10fcd0),
	.w6(32'h3a1d1a1d),
	.w7(32'h3a14d0cb),
	.w8(32'h3a387883),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e8ae),
	.w1(32'h3b0953ee),
	.w2(32'hba6df2f0),
	.w3(32'h3a8d494b),
	.w4(32'h3a8f4936),
	.w5(32'hba6fc9de),
	.w6(32'h3a62460c),
	.w7(32'h394032f3),
	.w8(32'hbad0bc58),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926a577),
	.w1(32'hba2fe781),
	.w2(32'hba822809),
	.w3(32'h3a0d2bf8),
	.w4(32'h364428c0),
	.w5(32'hba13b213),
	.w6(32'h3956be8d),
	.w7(32'hb905a4fa),
	.w8(32'hba864e3f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c2aa9),
	.w1(32'hba8c7df3),
	.w2(32'h3a2bf95c),
	.w3(32'hbb0f9918),
	.w4(32'hba6da94d),
	.w5(32'h3aebee93),
	.w6(32'hbabf38ed),
	.w7(32'h39c952dc),
	.w8(32'h3b1d04dd),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fef14),
	.w1(32'h3a222edd),
	.w2(32'h3a1f1457),
	.w3(32'h3a3223d6),
	.w4(32'h3a1fe4ff),
	.w5(32'h3a8b6ad8),
	.w6(32'h3aca36f2),
	.w7(32'hb93dd70e),
	.w8(32'h3a49b615),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44bd09),
	.w1(32'hb9bade4d),
	.w2(32'hbaf694b3),
	.w3(32'h396583bb),
	.w4(32'h3a432f45),
	.w5(32'hbb14f36b),
	.w6(32'h3a293909),
	.w7(32'h39ded01e),
	.w8(32'hbb08c7e8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed0e8b),
	.w1(32'hb989fd93),
	.w2(32'hba57de2a),
	.w3(32'h399151ce),
	.w4(32'h3a4a47fb),
	.w5(32'hb9dd729d),
	.w6(32'hb9e1dce5),
	.w7(32'h3a664bb9),
	.w8(32'hb91dfd57),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c0376e),
	.w1(32'h367fcc6f),
	.w2(32'h37525c94),
	.w3(32'hb3f82e8c),
	.w4(32'h35df1828),
	.w5(32'h377ce841),
	.w6(32'hb69622dc),
	.w7(32'h36b4dfef),
	.w8(32'h3777c39f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0a27),
	.w1(32'hba77a3af),
	.w2(32'h3aa85810),
	.w3(32'hbb03e632),
	.w4(32'h39c98e77),
	.w5(32'h3adef5cf),
	.w6(32'hba387494),
	.w7(32'h39f521d2),
	.w8(32'h3ae07236),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c92b8d),
	.w1(32'hb6d361a7),
	.w2(32'h37cd4f25),
	.w3(32'hb6b2cf51),
	.w4(32'hb77d15aa),
	.w5(32'h37eae47c),
	.w6(32'h36256fca),
	.w7(32'hb7620141),
	.w8(32'h38006502),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aaca80),
	.w1(32'h3a084a8c),
	.w2(32'hba53609f),
	.w3(32'h39ea5342),
	.w4(32'h3a606494),
	.w5(32'hba5451ab),
	.w6(32'h39d70e2d),
	.w7(32'h389fef75),
	.w8(32'hba88d46e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6574d36),
	.w1(32'hb9e9ee16),
	.w2(32'hb9aeaa18),
	.w3(32'hb8c71244),
	.w4(32'hbaaec470),
	.w5(32'h39f4edce),
	.w6(32'hbae0f631),
	.w7(32'hbb123808),
	.w8(32'h3763c19d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e2dd2),
	.w1(32'h393ee51b),
	.w2(32'hb897543a),
	.w3(32'h38d5df3c),
	.w4(32'h39b15590),
	.w5(32'h38cc7434),
	.w6(32'hb91fcd63),
	.w7(32'hb9065774),
	.w8(32'h398eb3d4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a60c3f),
	.w1(32'h39a0418d),
	.w2(32'h39298f26),
	.w3(32'h38f82912),
	.w4(32'h38ba0b25),
	.w5(32'h3903e1e7),
	.w6(32'hb8458d1d),
	.w7(32'hb90f6ef3),
	.w8(32'hb90318ad),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9051adf),
	.w1(32'h38b15980),
	.w2(32'h39ef313e),
	.w3(32'h39a0833d),
	.w4(32'hb9eaef35),
	.w5(32'h3a68a1d7),
	.w6(32'hb92d5877),
	.w7(32'hba030040),
	.w8(32'h3ae92c40),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d6aae),
	.w1(32'hba8f09ad),
	.w2(32'hba274772),
	.w3(32'hb9b125a4),
	.w4(32'h383cc6db),
	.w5(32'h39a95c77),
	.w6(32'h3a104a53),
	.w7(32'h399af575),
	.w8(32'h392439aa),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeaff2),
	.w1(32'hbac1b80e),
	.w2(32'hbb31e7f9),
	.w3(32'h3a89f655),
	.w4(32'hba1770b6),
	.w5(32'hbaec5abb),
	.w6(32'h3b1e02ca),
	.w7(32'h3a586777),
	.w8(32'hba7c4bfe),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373332ea),
	.w1(32'h3768342c),
	.w2(32'h381abe9d),
	.w3(32'hb59ec762),
	.w4(32'h3722fbb0),
	.w5(32'h37901ec3),
	.w6(32'h33dfdd1e),
	.w7(32'h34d1b5c4),
	.w8(32'hb6b4cf6b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381eb1bf),
	.w1(32'h3807d607),
	.w2(32'h38b46f4b),
	.w3(32'hb79a5916),
	.w4(32'h35357781),
	.w5(32'h3838e4ef),
	.w6(32'h3893243a),
	.w7(32'hb777ddcc),
	.w8(32'h3778b037),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9ef4),
	.w1(32'h3af9d912),
	.w2(32'hbb35d111),
	.w3(32'h3aaeff06),
	.w4(32'h3ac9361b),
	.w5(32'hbb396eaf),
	.w6(32'hb9ade413),
	.w7(32'h3ae47ce1),
	.w8(32'hb9a1eb14),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c9a6),
	.w1(32'hb9b6bf14),
	.w2(32'hbaf25ff1),
	.w3(32'hbaa93437),
	.w4(32'h3a0bfcab),
	.w5(32'hba42f5eb),
	.w6(32'h390b0a4d),
	.w7(32'hb9c343ed),
	.w8(32'hba128ba5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b80d4f),
	.w1(32'h399f4eaf),
	.w2(32'h39955d23),
	.w3(32'h3a3416f0),
	.w4(32'h3a2c3967),
	.w5(32'h3a399c39),
	.w6(32'hba184378),
	.w7(32'hb94aa86d),
	.w8(32'h3a4fb430),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d9eeb),
	.w1(32'h3ba3acae),
	.w2(32'h3b03889e),
	.w3(32'h3ad96158),
	.w4(32'h3bbacf99),
	.w5(32'h3b5c3a9a),
	.w6(32'h3a18ea45),
	.w7(32'hbb491c03),
	.w8(32'hbb567153),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f90653),
	.w1(32'hb7ebd721),
	.w2(32'h38bf0a20),
	.w3(32'hb90d6950),
	.w4(32'hba0f76e2),
	.w5(32'hb870463c),
	.w6(32'hb991bcc9),
	.w7(32'hba4a580b),
	.w8(32'h38d02b8e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edc29b),
	.w1(32'hba396e85),
	.w2(32'hb937f2b6),
	.w3(32'hba14942f),
	.w4(32'hb9b748f7),
	.w5(32'h3a19d24f),
	.w6(32'hb9ff9cc2),
	.w7(32'hb9d6b593),
	.w8(32'h39be0331),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cbdb7),
	.w1(32'h3bba85bf),
	.w2(32'hbae13229),
	.w3(32'hbb41c7f7),
	.w4(32'h3b437e93),
	.w5(32'hbba1d593),
	.w6(32'hbaea4be2),
	.w7(32'h3b4a2de6),
	.w8(32'hbb654d9d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f834),
	.w1(32'hbaf1b43a),
	.w2(32'hbb41b81f),
	.w3(32'hb95ccfd4),
	.w4(32'hba213765),
	.w5(32'hbb06e603),
	.w6(32'h3ad0e2a0),
	.w7(32'hba3720f8),
	.w8(32'hbb1cc150),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d6e4),
	.w1(32'h3a6d7423),
	.w2(32'hb9fd921e),
	.w3(32'hbab4b726),
	.w4(32'h3b45f93e),
	.w5(32'h39e93373),
	.w6(32'hbaabd854),
	.w7(32'h3b5c654c),
	.w8(32'h393d32d9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1567d),
	.w1(32'h3a21ba45),
	.w2(32'h3a9352e6),
	.w3(32'hb913c250),
	.w4(32'hbaa87ae0),
	.w5(32'h395bdc1e),
	.w6(32'hba9ffe7b),
	.w7(32'hbb05eea7),
	.w8(32'hb99b6fe5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb4366),
	.w1(32'hba4fe636),
	.w2(32'h39995bbc),
	.w3(32'hb9f2ba77),
	.w4(32'hbaf30223),
	.w5(32'h39a46fe3),
	.w6(32'hba9d7238),
	.w7(32'hbb2e2961),
	.w8(32'hb905fd52),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373cd351),
	.w1(32'h370194c1),
	.w2(32'h36fa5e5a),
	.w3(32'h36b6b20e),
	.w4(32'h364709e1),
	.w5(32'h360eab9c),
	.w6(32'h36124786),
	.w7(32'hb433921f),
	.w8(32'h35bfa901),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37516129),
	.w1(32'h374992ee),
	.w2(32'h376c3609),
	.w3(32'h3704a26e),
	.w4(32'h36f0bd43),
	.w5(32'h37173be0),
	.w6(32'h37005ce5),
	.w7(32'h36c4f44d),
	.w8(32'h3702eb4d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae75e89),
	.w1(32'h3ac264df),
	.w2(32'h39b1913d),
	.w3(32'h38c48370),
	.w4(32'hb95a4395),
	.w5(32'hb991bccd),
	.w6(32'hb8b12108),
	.w7(32'hba3e9733),
	.w8(32'hba229fd5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369f8149),
	.w1(32'hb5747907),
	.w2(32'h373d98b2),
	.w3(32'h36d3542e),
	.w4(32'hb688fd82),
	.w5(32'h366c8c8a),
	.w6(32'h36690c73),
	.w7(32'hb66b4541),
	.w8(32'h360f548e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa43ba8),
	.w1(32'h3997bc2d),
	.w2(32'hbafee1b4),
	.w3(32'h396b4c43),
	.w4(32'hba2fbf3e),
	.w5(32'hbafee595),
	.w6(32'hb8b5f088),
	.w7(32'hb925501c),
	.w8(32'hbafcb457),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f865),
	.w1(32'h39dc70a1),
	.w2(32'hba93477f),
	.w3(32'hba25e771),
	.w4(32'hb97562d8),
	.w5(32'hbaa98168),
	.w6(32'h390227fc),
	.w7(32'hba498f9e),
	.w8(32'hba48a0da),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c827f),
	.w1(32'hb8e7dff1),
	.w2(32'hba021a8d),
	.w3(32'h39102a59),
	.w4(32'h39c7790b),
	.w5(32'hb95a5370),
	.w6(32'hb8836708),
	.w7(32'h39afa9c8),
	.w8(32'h387fd96a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ed932),
	.w1(32'h374f6a3b),
	.w2(32'h380a9d83),
	.w3(32'hb685fb99),
	.w4(32'h35e988b0),
	.w5(32'h37afb7df),
	.w6(32'hb7182e33),
	.w7(32'h36901595),
	.w8(32'h37d641c0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15892c),
	.w1(32'h3a048cf0),
	.w2(32'hbb1f9424),
	.w3(32'hbb85e6cf),
	.w4(32'h3b2973bd),
	.w5(32'hb8f3400d),
	.w6(32'hbb3f4d7a),
	.w7(32'h3b33bd41),
	.w8(32'hbad51954),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff510c),
	.w1(32'hb9379dee),
	.w2(32'hba518827),
	.w3(32'hba17ce7e),
	.w4(32'h38dd13d1),
	.w5(32'hb9ce352d),
	.w6(32'h3a03c3ee),
	.w7(32'hb970cbbf),
	.w8(32'hba49313f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938d1c2),
	.w1(32'hb8825ac8),
	.w2(32'h37c6331a),
	.w3(32'hb7366b92),
	.w4(32'h37f93cff),
	.w5(32'h37a56b74),
	.w6(32'hb86c92ac),
	.w7(32'hb903bc88),
	.w8(32'hb8832a71),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1ef70),
	.w1(32'hba08f293),
	.w2(32'hbabcbb0e),
	.w3(32'h3991ac2e),
	.w4(32'h39fb4ffe),
	.w5(32'hba47ad56),
	.w6(32'h39f3cb07),
	.w7(32'h3967845e),
	.w8(32'hba4af929),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffcdea),
	.w1(32'h388a25b9),
	.w2(32'h3842187a),
	.w3(32'hb6494b1c),
	.w4(32'hb8854e36),
	.w5(32'hb7caf43b),
	.w6(32'h381ccf71),
	.w7(32'hb7b8f1f8),
	.w8(32'h36890fb8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981adc0),
	.w1(32'h396b8193),
	.w2(32'hb8fc5c1a),
	.w3(32'h3901b74e),
	.w4(32'h390ae2e7),
	.w5(32'hb9b45fd4),
	.w6(32'h397b4137),
	.w7(32'h3993b0f9),
	.w8(32'h38bc5405),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c52b20),
	.w1(32'hb710d0a2),
	.w2(32'h38377462),
	.w3(32'hb7048093),
	.w4(32'h35c9b186),
	.w5(32'h3829aa75),
	.w6(32'h363289bc),
	.w7(32'h381e9f90),
	.w8(32'h37462f3a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378a002f),
	.w1(32'hb6261624),
	.w2(32'h3819bce4),
	.w3(32'h38753dfe),
	.w4(32'h37f641d8),
	.w5(32'h37eb7424),
	.w6(32'h3711b4a3),
	.w7(32'hb8494fdc),
	.w8(32'hb7bc710e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec57d0),
	.w1(32'h398abe6e),
	.w2(32'h39c81bd7),
	.w3(32'hb9cf3922),
	.w4(32'hb97a7dea),
	.w5(32'h39646233),
	.w6(32'hba93e5c8),
	.w7(32'hba10e96b),
	.w8(32'h388b5d5d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7cd26),
	.w1(32'hbb0cb865),
	.w2(32'hbb10ac71),
	.w3(32'h3aff629b),
	.w4(32'hb94d259d),
	.w5(32'hba9a173b),
	.w6(32'h3abd208f),
	.w7(32'hbb1b7fef),
	.w8(32'hba8f8172),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef464e),
	.w1(32'hbadeae90),
	.w2(32'hbadfbb8b),
	.w3(32'hb978242a),
	.w4(32'h39ab013c),
	.w5(32'hb9749565),
	.w6(32'h3a59039d),
	.w7(32'h3a1c53ba),
	.w8(32'hb97af913),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b18df),
	.w1(32'hb9df5bd4),
	.w2(32'hbaa045d4),
	.w3(32'h3a8132c9),
	.w4(32'h3a2bd957),
	.w5(32'hba0b95f6),
	.w6(32'h3acf4586),
	.w7(32'hba2e2230),
	.w8(32'hb9e4be6d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38939244),
	.w1(32'h392acc52),
	.w2(32'h3986d37c),
	.w3(32'h38d69ced),
	.w4(32'h39511ab6),
	.w5(32'h395725e9),
	.w6(32'h38a11176),
	.w7(32'h39391979),
	.w8(32'h393ab05a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3715aa0a),
	.w1(32'h383e12b2),
	.w2(32'hb8967676),
	.w3(32'hb8ca1f33),
	.w4(32'hb959b1f0),
	.w5(32'h38a3627d),
	.w6(32'hb955cba5),
	.w7(32'hb8a313bf),
	.w8(32'h38c2f0ac),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377d5a06),
	.w1(32'h380bd2ae),
	.w2(32'h37a02bfe),
	.w3(32'h37eb5227),
	.w4(32'h37fdb4df),
	.w5(32'h374641c7),
	.w6(32'h3801e5b8),
	.w7(32'h379d3154),
	.w8(32'h36f2d511),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eec3a7),
	.w1(32'hb7cf0990),
	.w2(32'hb83e5a19),
	.w3(32'h385dd13c),
	.w4(32'h381078ce),
	.w5(32'hb7386630),
	.w6(32'h383a3c54),
	.w7(32'h38038fc5),
	.w8(32'h36539ebd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09db7f),
	.w1(32'hbb206000),
	.w2(32'hbaecc769),
	.w3(32'hba47d1ff),
	.w4(32'hbaf2f7c7),
	.w5(32'hb92dcd45),
	.w6(32'hb9f4f0de),
	.w7(32'hbad915d2),
	.w8(32'hb91fa245),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38605afe),
	.w1(32'h3851e4e4),
	.w2(32'h3919b334),
	.w3(32'h36f53795),
	.w4(32'h37cef257),
	.w5(32'h38fddb57),
	.w6(32'h38718253),
	.w7(32'h38681710),
	.w8(32'h38e72da5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27378c),
	.w1(32'h38735cc5),
	.w2(32'h3998077e),
	.w3(32'h3a0ca476),
	.w4(32'h383afb1e),
	.w5(32'h39d71d51),
	.w6(32'h39da801c),
	.w7(32'hb7b9478c),
	.w8(32'h399b32ed),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aef80),
	.w1(32'hba632bb7),
	.w2(32'h399dc8e7),
	.w3(32'hba9b9eef),
	.w4(32'hb8e3d777),
	.w5(32'h3a4cec3d),
	.w6(32'hba8be4a9),
	.w7(32'hb9a49d15),
	.w8(32'h395dd01a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3652344b),
	.w1(32'h37e41b74),
	.w2(32'h389e603e),
	.w3(32'hb7a53b12),
	.w4(32'h37caf5a4),
	.w5(32'h388f4b97),
	.w6(32'hb7c28522),
	.w7(32'h37533ec3),
	.w8(32'h383cfa22),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990e278),
	.w1(32'hb8a6921b),
	.w2(32'hba2a03a7),
	.w3(32'h3a3fe2c7),
	.w4(32'h39913c6d),
	.w5(32'hb9c46d62),
	.w6(32'h3a50ab05),
	.w7(32'h39c3a5ce),
	.w8(32'hb99543cb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f895e7),
	.w1(32'hb863d691),
	.w2(32'h38e91b5d),
	.w3(32'hb8cdcdb9),
	.w4(32'hb8901969),
	.w5(32'hb8b3988a),
	.w6(32'hb88e39bf),
	.w7(32'hb8a967d2),
	.w8(32'h3303db99),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66045),
	.w1(32'hbb947741),
	.w2(32'hbb3e07b2),
	.w3(32'h3ae9d15a),
	.w4(32'hba9c86ba),
	.w5(32'h3aacb3cd),
	.w6(32'h39088d56),
	.w7(32'hbb2d5726),
	.w8(32'h3b3b50c2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39065e6f),
	.w1(32'hb86bd09e),
	.w2(32'hb9663f89),
	.w3(32'h372b5212),
	.w4(32'hb8fc85d6),
	.w5(32'hb9584c07),
	.w6(32'hb71f0de6),
	.w7(32'hb90cd551),
	.w8(32'hb90d8106),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba29f4),
	.w1(32'h3a059bd9),
	.w2(32'h39b3adde),
	.w3(32'hb8acbca7),
	.w4(32'h3ae2c719),
	.w5(32'h3ad382ff),
	.w6(32'hbb230bb4),
	.w7(32'hb9e4fd36),
	.w8(32'h3abf49f4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule