module layer_8_featuremap_26(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d073e),
	.w1(32'hba801678),
	.w2(32'hb9e64299),
	.w3(32'hba56c545),
	.w4(32'hbabe0012),
	.w5(32'hba0a5caf),
	.w6(32'h38596b4f),
	.w7(32'hb99c1a08),
	.w8(32'hb9edd036),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f284f3),
	.w1(32'hba33e611),
	.w2(32'hba164d32),
	.w3(32'hb9d01fce),
	.w4(32'hba4e7a9a),
	.w5(32'hba48121c),
	.w6(32'hb99823f9),
	.w7(32'hb9a12a91),
	.w8(32'h395433e6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398718de),
	.w1(32'hb9ad2665),
	.w2(32'hb9f86261),
	.w3(32'hb90df565),
	.w4(32'hba287d71),
	.w5(32'hba55e89c),
	.w6(32'h38ab25a3),
	.w7(32'hb7805a2d),
	.w8(32'hbb84dc78),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb962c45),
	.w1(32'h3a097ada),
	.w2(32'h3b25afc1),
	.w3(32'h3ac99a47),
	.w4(32'h3acecf6f),
	.w5(32'h39e7e9e6),
	.w6(32'hbb1810d0),
	.w7(32'hbb27bf5b),
	.w8(32'h39ae376f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944d703),
	.w1(32'hb9ec62db),
	.w2(32'hb8801e0a),
	.w3(32'h393bc738),
	.w4(32'hb9388a11),
	.w5(32'hb9873dcb),
	.w6(32'h39828946),
	.w7(32'hb97335e8),
	.w8(32'hbae465f0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60cd5d),
	.w1(32'hba5e0710),
	.w2(32'h3b18c35b),
	.w3(32'h3a94ea4b),
	.w4(32'h38cbaf05),
	.w5(32'h3b024a66),
	.w6(32'hb95ad6f2),
	.w7(32'h3a8f5f4b),
	.w8(32'h39c33aa2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fdc4c),
	.w1(32'hb8c18b9c),
	.w2(32'h38a73071),
	.w3(32'hb940dc18),
	.w4(32'hba3d2b34),
	.w5(32'hba207951),
	.w6(32'h3a0937dc),
	.w7(32'h39da6af1),
	.w8(32'h3891edd6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883fc20),
	.w1(32'hba170c0b),
	.w2(32'h39a37145),
	.w3(32'h398f4666),
	.w4(32'h3921b33b),
	.w5(32'hb8ea1b37),
	.w6(32'hb90ebff4),
	.w7(32'hb98ffe12),
	.w8(32'h38ab707b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bcd0f),
	.w1(32'h38d2050a),
	.w2(32'hb9a89c3f),
	.w3(32'h38ad9048),
	.w4(32'hb9b691b9),
	.w5(32'hba56313b),
	.w6(32'h39859a64),
	.w7(32'hb78cbe95),
	.w8(32'hbb78e20e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd86764),
	.w1(32'h3aecd60d),
	.w2(32'h3bc35e85),
	.w3(32'h3a0fd273),
	.w4(32'h3b293ae7),
	.w5(32'h3b4a270c),
	.w6(32'hbb5e1196),
	.w7(32'hbb6adb87),
	.w8(32'h3adc163b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65915d),
	.w1(32'h3a29e0fc),
	.w2(32'h390a28cd),
	.w3(32'h3a270b0f),
	.w4(32'h3a07a635),
	.w5(32'hb9b48089),
	.w6(32'h3a8cd2a8),
	.w7(32'h3a059a28),
	.w8(32'hb72f77dd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372c7d89),
	.w1(32'hb9f04013),
	.w2(32'hb9eaa0b3),
	.w3(32'hb9f8b746),
	.w4(32'hba5a1e25),
	.w5(32'hba660a41),
	.w6(32'h395076a7),
	.w7(32'h371ba087),
	.w8(32'h3a6f60d0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd5a6b),
	.w1(32'hb9301930),
	.w2(32'h373a6e55),
	.w3(32'h3949f25c),
	.w4(32'hb9bd0bb7),
	.w5(32'hba376053),
	.w6(32'h3a2f005b),
	.w7(32'h39c698d0),
	.w8(32'hbae50073),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c38c1),
	.w1(32'hba6074c2),
	.w2(32'h3b38a604),
	.w3(32'h3ad854c1),
	.w4(32'h39a51dbc),
	.w5(32'h3b29fdf3),
	.w6(32'h3775b1f0),
	.w7(32'h3ad2946a),
	.w8(32'hba6e7cc0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f81bd),
	.w1(32'hba33298b),
	.w2(32'h3a9e71bf),
	.w3(32'h39f46d2a),
	.w4(32'hba36a5d6),
	.w5(32'h3904dea4),
	.w6(32'h3984e500),
	.w7(32'h3a234d01),
	.w8(32'hba73f6c1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f162),
	.w1(32'hba625c60),
	.w2(32'h394fa32f),
	.w3(32'hba8896ba),
	.w4(32'hba820572),
	.w5(32'hb9e1dc1f),
	.w6(32'hb92d677c),
	.w7(32'hb996cc0b),
	.w8(32'h398be2b3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9369f),
	.w1(32'hba172cc2),
	.w2(32'h3ae207e9),
	.w3(32'hbb5c50ca),
	.w4(32'h3b538004),
	.w5(32'h3bd48d8b),
	.w6(32'h3b0e7dec),
	.w7(32'h3a68f4b9),
	.w8(32'h3aa18bb8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f7340),
	.w1(32'h3857ca8a),
	.w2(32'hb98260dd),
	.w3(32'h39a9d8af),
	.w4(32'hba346654),
	.w5(32'hbaa8695a),
	.w6(32'h3a374e37),
	.w7(32'h3974bd50),
	.w8(32'h3a1174b1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf0380),
	.w1(32'hbad82575),
	.w2(32'hba166c48),
	.w3(32'h39f6a7ba),
	.w4(32'h39cc979e),
	.w5(32'hbad8f07a),
	.w6(32'hb9e1a97b),
	.w7(32'hba4d3bc0),
	.w8(32'h38a2a120),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568db6),
	.w1(32'h3b0c93d3),
	.w2(32'hbbd9e2c8),
	.w3(32'h3ab4aedb),
	.w4(32'hbb8bb315),
	.w5(32'hbb24763d),
	.w6(32'h3b8c5562),
	.w7(32'hb9bbee66),
	.w8(32'h3ad97041),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2799e7),
	.w1(32'h39208c5d),
	.w2(32'hba31a623),
	.w3(32'h3a07814d),
	.w4(32'h37c6d5b7),
	.w5(32'hba655cf8),
	.w6(32'h3a6aea89),
	.w7(32'h38f64f48),
	.w8(32'h3a93a4f4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ee063),
	.w1(32'hb982afc8),
	.w2(32'hb79572e2),
	.w3(32'h395acf28),
	.w4(32'hba0f1df1),
	.w5(32'hba0bf94d),
	.w6(32'h3a68c8e2),
	.w7(32'h393beb45),
	.w8(32'h3b8159e8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef62dd),
	.w1(32'h3a624827),
	.w2(32'hba13bb84),
	.w3(32'h3ac0768a),
	.w4(32'h3af0e0bc),
	.w5(32'h3aca2b15),
	.w6(32'h3ae33ca6),
	.w7(32'h3b3c0e26),
	.w8(32'hb96f9fc1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba476462),
	.w1(32'hbabb9e27),
	.w2(32'hb98230ba),
	.w3(32'hba86c32e),
	.w4(32'hba71d0d5),
	.w5(32'hba7807a8),
	.w6(32'hbae042e3),
	.w7(32'hbae8383d),
	.w8(32'hbae6f236),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb060cc5),
	.w1(32'h3b6f6fa3),
	.w2(32'h3adea16f),
	.w3(32'hbb56e8ae),
	.w4(32'h3abeee72),
	.w5(32'h3ac2d40a),
	.w6(32'hba843d78),
	.w7(32'hbaab651b),
	.w8(32'h3b7698a4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad77912),
	.w1(32'h3a064aa6),
	.w2(32'hba2597ec),
	.w3(32'h3aad37c7),
	.w4(32'h3ab5635a),
	.w5(32'h3a9fdef6),
	.w6(32'h3acd1939),
	.w7(32'h3b1dcc12),
	.w8(32'h3b65619c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3b375),
	.w1(32'h39d3c91a),
	.w2(32'hba0a48aa),
	.w3(32'h3a8b8bb5),
	.w4(32'h3a6c12af),
	.w5(32'h3a66d6b8),
	.w6(32'h3ab19311),
	.w7(32'h3af3254b),
	.w8(32'h3acfa5e7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e6b2f),
	.w1(32'h398d9905),
	.w2(32'hba348eb6),
	.w3(32'hba15a055),
	.w4(32'h3a18facd),
	.w5(32'h39c5e1aa),
	.w6(32'h3a29f0cd),
	.w7(32'h39a5ed80),
	.w8(32'hbba01df7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f9ba3),
	.w1(32'hba93a2ce),
	.w2(32'h3b27590b),
	.w3(32'hb91c4415),
	.w4(32'h3b2e1812),
	.w5(32'h3b3662b2),
	.w6(32'hbb86bf4c),
	.w7(32'hbbac82a0),
	.w8(32'h378db892),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880e6cf),
	.w1(32'hb9b2c972),
	.w2(32'hb966c837),
	.w3(32'hb9912395),
	.w4(32'hba257f44),
	.w5(32'hba348792),
	.w6(32'h38f7b94b),
	.w7(32'hb822bf03),
	.w8(32'hbbceb884),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9246d20),
	.w1(32'h3a89367c),
	.w2(32'hba8665f8),
	.w3(32'hba9bfb83),
	.w4(32'hb9bbcbcd),
	.w5(32'h39121b9d),
	.w6(32'hbbacf533),
	.w7(32'hbbfdaa98),
	.w8(32'h39eb3a49),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1bba9),
	.w1(32'hba2c88da),
	.w2(32'hba9b2696),
	.w3(32'hbb56b82d),
	.w4(32'hbb23c091),
	.w5(32'hbb1f3220),
	.w6(32'h39f77ff5),
	.w7(32'h34d57e00),
	.w8(32'hba7124d5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b70d),
	.w1(32'hb9e78377),
	.w2(32'h3b922414),
	.w3(32'hbb87cc2d),
	.w4(32'hbb615d91),
	.w5(32'hbb10288d),
	.w6(32'h3989b088),
	.w7(32'h39400c57),
	.w8(32'hbb8570bb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ffcd0),
	.w1(32'hb9e675f1),
	.w2(32'hbb80ec0e),
	.w3(32'h3b24b17a),
	.w4(32'h3a596c22),
	.w5(32'h3b52310f),
	.w6(32'hbad15784),
	.w7(32'hbad95614),
	.w8(32'hbac8ceac),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ed16d),
	.w1(32'hba4673db),
	.w2(32'h3b239d6d),
	.w3(32'h3ac067bf),
	.w4(32'h3992666f),
	.w5(32'h3b18ad6f),
	.w6(32'h380876ef),
	.w7(32'h3ab84c38),
	.w8(32'hba1fdb5c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eefd6),
	.w1(32'hbae364ff),
	.w2(32'hba6fbe94),
	.w3(32'hba732a6d),
	.w4(32'hbaaf3468),
	.w5(32'hbaabf70c),
	.w6(32'hba7275bb),
	.w7(32'hbac8a023),
	.w8(32'h3949e9c2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8359b1),
	.w1(32'h3ac6d4a3),
	.w2(32'hb8c3133e),
	.w3(32'hbab55992),
	.w4(32'h3a43bea7),
	.w5(32'h3a8df53f),
	.w6(32'hba6a14fe),
	.w7(32'hba00695a),
	.w8(32'h38e8c9a6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397532aa),
	.w1(32'hba583517),
	.w2(32'hba269e09),
	.w3(32'hb9ce4816),
	.w4(32'hbab5a7a7),
	.w5(32'hbaaef79c),
	.w6(32'hb8414cf2),
	.w7(32'hb984ab99),
	.w8(32'hbabd108e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5d113),
	.w1(32'hba894605),
	.w2(32'h3b276ace),
	.w3(32'h3a5e5363),
	.w4(32'hbaafbdfa),
	.w5(32'hb9c1de5d),
	.w6(32'h3a5ba220),
	.w7(32'h3aa99f5b),
	.w8(32'h37e29709),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bc0d6),
	.w1(32'h3a32f0e5),
	.w2(32'hb935d295),
	.w3(32'hba3751c5),
	.w4(32'h391543e6),
	.w5(32'h390bf979),
	.w6(32'h3942055a),
	.w7(32'h398fe9e9),
	.w8(32'h3ac83e25),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a096988),
	.w1(32'h3976d1bc),
	.w2(32'hb99805d2),
	.w3(32'h39b279f4),
	.w4(32'h39f31cbe),
	.w5(32'h39def14b),
	.w6(32'h39fc3984),
	.w7(32'h3a583a8c),
	.w8(32'h3b103602),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b776c),
	.w1(32'h3a377589),
	.w2(32'hba2db01e),
	.w3(32'h39cdfa6b),
	.w4(32'h3aa3be56),
	.w5(32'h3ab075ac),
	.w6(32'h3b39979f),
	.w7(32'h3a7f9cc3),
	.w8(32'h3a65ecc1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1162),
	.w1(32'h3bfb49dd),
	.w2(32'hbc0f4af2),
	.w3(32'h39bdd597),
	.w4(32'h3bb60e02),
	.w5(32'hbae24335),
	.w6(32'h3c272df2),
	.w7(32'hbbf253a0),
	.w8(32'hbac4685a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08bdd),
	.w1(32'h3b6fbc15),
	.w2(32'h3aaa222e),
	.w3(32'hbadbfff7),
	.w4(32'h3ac419d0),
	.w5(32'h3a2de957),
	.w6(32'h3ad4b51d),
	.w7(32'h3a7a98cf),
	.w8(32'hbba09b71),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d0ea),
	.w1(32'hbb38bf42),
	.w2(32'hbb8935b7),
	.w3(32'hbb45d643),
	.w4(32'hbab94668),
	.w5(32'hbb11a29b),
	.w6(32'hbb89f5cc),
	.w7(32'hbb542554),
	.w8(32'hbb1fd473),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b22e),
	.w1(32'hbc3bcc8a),
	.w2(32'hbb95418e),
	.w3(32'hb98a9dc8),
	.w4(32'hbc1862a7),
	.w5(32'hbb602b51),
	.w6(32'hba596808),
	.w7(32'h3b380af9),
	.w8(32'h3aefb98d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17960),
	.w1(32'hbbf2a87e),
	.w2(32'h3b4c9418),
	.w3(32'hb957154f),
	.w4(32'h3b99fc2a),
	.w5(32'h3bb60692),
	.w6(32'hba144e89),
	.w7(32'hba1ab4ae),
	.w8(32'h3b1eb618),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2830da),
	.w1(32'hbc4fca44),
	.w2(32'hbaed77ab),
	.w3(32'h3b9c8e70),
	.w4(32'hbb717f89),
	.w5(32'h3ba39797),
	.w6(32'hbbf037e6),
	.w7(32'h3b82846d),
	.w8(32'h3a8f07cf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf68bfd),
	.w1(32'h3c3631a4),
	.w2(32'h3c72f004),
	.w3(32'h3bf036ac),
	.w4(32'h3c4f0652),
	.w5(32'h3c755774),
	.w6(32'h3c018e50),
	.w7(32'h3c0a7844),
	.w8(32'hbb3afb82),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be198),
	.w1(32'hbbbcc3cc),
	.w2(32'hbb5bb14e),
	.w3(32'hbb1118ee),
	.w4(32'hbb53804a),
	.w5(32'hba9063ae),
	.w6(32'hbb32bf7b),
	.w7(32'h3a06a75d),
	.w8(32'h39688ea6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889e958),
	.w1(32'h3b4ab962),
	.w2(32'h3a4bd750),
	.w3(32'hb9c525df),
	.w4(32'h3a824ba1),
	.w5(32'hb95069d4),
	.w6(32'h3ad32aa2),
	.w7(32'h39edb83c),
	.w8(32'h3aa62746),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb84a),
	.w1(32'h3bdd26cb),
	.w2(32'h3adf198c),
	.w3(32'h3a94d0ca),
	.w4(32'h3b865ba3),
	.w5(32'h39faa253),
	.w6(32'h3b8d3838),
	.w7(32'h3ad5b037),
	.w8(32'hbb81859b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707b73),
	.w1(32'hbb5b4785),
	.w2(32'hbb8103f8),
	.w3(32'hbc3e6e2c),
	.w4(32'hbbc3d744),
	.w5(32'hbc0f9711),
	.w6(32'hbb47c27b),
	.w7(32'hbbd5950a),
	.w8(32'h3c680672),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87871a),
	.w1(32'h3c74d369),
	.w2(32'h3c6e6a9c),
	.w3(32'h3c6c31b9),
	.w4(32'h3c65b5a4),
	.w5(32'h3c6394b1),
	.w6(32'h3c3e6aab),
	.w7(32'h3c421ffa),
	.w8(32'h3b7abf41),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70c3b0),
	.w1(32'hbb9bb577),
	.w2(32'h3bd9a036),
	.w3(32'h3bc890de),
	.w4(32'hba71f9cf),
	.w5(32'h3bb5ce97),
	.w6(32'hbb042333),
	.w7(32'h3b3197b9),
	.w8(32'hbb656609),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3706b1),
	.w1(32'h3b06018f),
	.w2(32'h3b1035da),
	.w3(32'hba881887),
	.w4(32'hbafd6050),
	.w5(32'hbb0eaac3),
	.w6(32'h3afa5388),
	.w7(32'h3916df60),
	.w8(32'h3b744b3b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea3910),
	.w1(32'hbb40d2ae),
	.w2(32'h3a0db401),
	.w3(32'h393a3254),
	.w4(32'hbb1b4692),
	.w5(32'hba7a1c33),
	.w6(32'h3ac93c52),
	.w7(32'h3c0d427a),
	.w8(32'h3afcc26c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac83b46),
	.w1(32'hbb9ce45d),
	.w2(32'hbace79f8),
	.w3(32'hbb071557),
	.w4(32'hba37d102),
	.w5(32'h3ab2f7ab),
	.w6(32'h3998ef60),
	.w7(32'hbb2ce3be),
	.w8(32'hbc86b658),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc172144),
	.w1(32'h39aa2b2a),
	.w2(32'hbb2309ad),
	.w3(32'hbc3a2e10),
	.w4(32'hbb3d9c7c),
	.w5(32'hbb85d12b),
	.w6(32'hbbd2a917),
	.w7(32'hbc100906),
	.w8(32'h3bb03bcb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3233),
	.w1(32'h3c8eb017),
	.w2(32'h3c140a72),
	.w3(32'h3ba2b79c),
	.w4(32'h3c856882),
	.w5(32'h3c0b7aaf),
	.w6(32'h3c48a1d7),
	.w7(32'h3bb8a265),
	.w8(32'hbbd550d7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba471af),
	.w1(32'hb88c1bad),
	.w2(32'hbbb79784),
	.w3(32'hbb82ce65),
	.w4(32'hbac8a484),
	.w5(32'hbc269e9e),
	.w6(32'hba98242c),
	.w7(32'h3b0ff6ec),
	.w8(32'hbb8ff7b1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbebff5),
	.w1(32'hbc4a3def),
	.w2(32'hba3c4afa),
	.w3(32'h3c0ad07c),
	.w4(32'h3bafc155),
	.w5(32'h3c254fcd),
	.w6(32'hbba7e6bd),
	.w7(32'h3bb5c44c),
	.w8(32'h3b4854c0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f68eb),
	.w1(32'h3b4f064a),
	.w2(32'h3bd02355),
	.w3(32'h3b6ff813),
	.w4(32'h3b2b6469),
	.w5(32'h3be5486e),
	.w6(32'h3b86a1a4),
	.w7(32'h3c1461a9),
	.w8(32'hbc072e16),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5930b9),
	.w1(32'h3a5254a6),
	.w2(32'hbb6989db),
	.w3(32'hbbdf1ba5),
	.w4(32'hbb431e62),
	.w5(32'hbc067dd4),
	.w6(32'hbc37c46d),
	.w7(32'hbc12e4ca),
	.w8(32'h39b76692),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a34e7),
	.w1(32'h3af30506),
	.w2(32'h3af26249),
	.w3(32'h3931094d),
	.w4(32'h3a70b7a6),
	.w5(32'h3b0d63c1),
	.w6(32'h3b19a23e),
	.w7(32'h3b668d60),
	.w8(32'h3aa0ce3a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e6ca9),
	.w1(32'h3bce6643),
	.w2(32'h3b0d6de8),
	.w3(32'h3a4ed049),
	.w4(32'h3b3c5eb5),
	.w5(32'h3a62475b),
	.w6(32'h3b6f4e3b),
	.w7(32'h3a82ad18),
	.w8(32'h3a35ada5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71c7eb),
	.w1(32'h3b6144d9),
	.w2(32'h3a81884b),
	.w3(32'h3a2e3b09),
	.w4(32'h3afb019f),
	.w5(32'h39a74d96),
	.w6(32'h3b0533cd),
	.w7(32'h3a33d161),
	.w8(32'h3a9f4f28),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e0d58),
	.w1(32'hbb2902e4),
	.w2(32'hbb4d25bc),
	.w3(32'h3b3005ba),
	.w4(32'h3b318105),
	.w5(32'h3b1616b8),
	.w6(32'h3b0135b7),
	.w7(32'h3b769027),
	.w8(32'hbb3164fd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7be839),
	.w1(32'hbbb46dc8),
	.w2(32'hbb955712),
	.w3(32'hbb3a2024),
	.w4(32'hbb58a227),
	.w5(32'hbb1085fc),
	.w6(32'hbb876672),
	.w7(32'hbb2733ae),
	.w8(32'hbcfb83cb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb94bb),
	.w1(32'hbc3bf215),
	.w2(32'hbc9f923c),
	.w3(32'hbce164d2),
	.w4(32'hbc8ee991),
	.w5(32'hbcaf8151),
	.w6(32'hbca737c9),
	.w7(32'hbcc26e95),
	.w8(32'h3a693b07),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e1a8e),
	.w1(32'h3b30d9bf),
	.w2(32'h39a213f9),
	.w3(32'hb7da2d4d),
	.w4(32'h3abadd1c),
	.w5(32'h3a1b0677),
	.w6(32'h3afc41c8),
	.w7(32'hb88b752a),
	.w8(32'hbb3e2ae3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd513fe),
	.w1(32'hbc1ef728),
	.w2(32'hbbcd0255),
	.w3(32'hbb892ab7),
	.w4(32'hbbc5ae80),
	.w5(32'hbb2d393c),
	.w6(32'hbb9ce8cb),
	.w7(32'hbb21d2c6),
	.w8(32'h3af7e6bc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bfddd),
	.w1(32'h3c08498d),
	.w2(32'h3b203a71),
	.w3(32'h3b1c072b),
	.w4(32'h3ba66d02),
	.w5(32'h3a60d846),
	.w6(32'h3b976bfc),
	.w7(32'h3abb4170),
	.w8(32'h3b09431e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8103f6),
	.w1(32'hbc1e629b),
	.w2(32'hbbf28670),
	.w3(32'h3b041e52),
	.w4(32'hbb0822bc),
	.w5(32'hbabe4716),
	.w6(32'h3ba3bd60),
	.w7(32'hba4061c2),
	.w8(32'hba755bf8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d670),
	.w1(32'hbb779fdf),
	.w2(32'hbbc3da13),
	.w3(32'hba59684d),
	.w4(32'hbb0ec8a0),
	.w5(32'hbb6d7bc0),
	.w6(32'hba6c0d67),
	.w7(32'hbb5e4358),
	.w8(32'h3a296183),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cec6ce),
	.w1(32'h3b6c2d3b),
	.w2(32'h3ad56d69),
	.w3(32'h3a31ec39),
	.w4(32'h3af78a9e),
	.w5(32'h3aa1dcf9),
	.w6(32'h3b061bea),
	.w7(32'h3a978e48),
	.w8(32'h390e1af7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ea2f7),
	.w1(32'h3a482b7a),
	.w2(32'hba986c7a),
	.w3(32'h3afdc2f1),
	.w4(32'h3b4f22b4),
	.w5(32'h3ab10930),
	.w6(32'h3acb4cc8),
	.w7(32'h38bc3bc9),
	.w8(32'hbd18292e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec01d4),
	.w1(32'hbc4c3ba0),
	.w2(32'hbcb15b8f),
	.w3(32'hbd03d397),
	.w4(32'hbca00679),
	.w5(32'hbcc3fa2a),
	.w6(32'hbcc147a8),
	.w7(32'hbce3b739),
	.w8(32'hbc869337),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc760938),
	.w1(32'hbc3620b3),
	.w2(32'hbc746c5e),
	.w3(32'hbc81b2af),
	.w4(32'hbc5d5275),
	.w5(32'hbc7a74d2),
	.w6(32'hbc67c14e),
	.w7(32'hbc7313b2),
	.w8(32'hba612fad),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6a673),
	.w1(32'h3a4f86e4),
	.w2(32'hb7069582),
	.w3(32'hba9f59ac),
	.w4(32'hb98e4ed3),
	.w5(32'h39f52158),
	.w6(32'h3b08b594),
	.w7(32'h3a9cb83e),
	.w8(32'hba8d84ea),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d95a8),
	.w1(32'h3c0b1d0d),
	.w2(32'h3b0a94cd),
	.w3(32'hbbc8ffa5),
	.w4(32'hbb83c132),
	.w5(32'hbbef44c3),
	.w6(32'h3a9bb3b6),
	.w7(32'hbbf72805),
	.w8(32'hba37791b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4778fc),
	.w1(32'hbb41bb05),
	.w2(32'hbadcdd43),
	.w3(32'h3a8d0ce8),
	.w4(32'h3afa39f9),
	.w5(32'h3aff69d7),
	.w6(32'hba2db3e8),
	.w7(32'h3adf3904),
	.w8(32'hbbd04671),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d244),
	.w1(32'hbc4a2938),
	.w2(32'hbb1cac08),
	.w3(32'hbb259194),
	.w4(32'hbb87661c),
	.w5(32'h3a9c044d),
	.w6(32'hbb18e652),
	.w7(32'h3bd0f07f),
	.w8(32'hbc4a01a1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39d4fc),
	.w1(32'hbc41bdbb),
	.w2(32'hbba706cf),
	.w3(32'hbc27c4fb),
	.w4(32'hbc0bbe55),
	.w5(32'hba85924f),
	.w6(32'hbc5af7e4),
	.w7(32'hbc2f7246),
	.w8(32'h3c2491fc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38b0da),
	.w1(32'h3c2f7b7b),
	.w2(32'h3c10af80),
	.w3(32'h3c2fdfd1),
	.w4(32'h3c231ec1),
	.w5(32'h3bfaa23c),
	.w6(32'h3c1d7462),
	.w7(32'h3bed5763),
	.w8(32'hbb7633f6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93915e),
	.w1(32'hbb3396ab),
	.w2(32'hbb645dad),
	.w3(32'hbb48ecc8),
	.w4(32'hba539548),
	.w5(32'hba34e6a3),
	.w6(32'hbb4faf07),
	.w7(32'hbae8c208),
	.w8(32'h3aa5a7c6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b6c5),
	.w1(32'h3c717dbf),
	.w2(32'h3ca16397),
	.w3(32'h3c1e23e7),
	.w4(32'h3c885058),
	.w5(32'h3ca25e89),
	.w6(32'h3c2bd77e),
	.w7(32'h3c361170),
	.w8(32'h3b9bff67),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab00867),
	.w1(32'hbbbda4f4),
	.w2(32'hbb2e8f20),
	.w3(32'h3a9c984e),
	.w4(32'hbbb6a767),
	.w5(32'hbab7821b),
	.w6(32'hba9f164a),
	.w7(32'h3b1c7a5d),
	.w8(32'h3c536024),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c502eea),
	.w1(32'h3b5f3543),
	.w2(32'h39bdc4fc),
	.w3(32'h3b8b8f50),
	.w4(32'h3a584a93),
	.w5(32'hbb92d4d7),
	.w6(32'h3b576e68),
	.w7(32'hbb0fd065),
	.w8(32'h3a90da1c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d66a),
	.w1(32'h3c613d77),
	.w2(32'h3c96cb98),
	.w3(32'h3c13bb24),
	.w4(32'h3c7fb3dd),
	.w5(32'h3c984e5b),
	.w6(32'h3c1fa729),
	.w7(32'h3c2abc58),
	.w8(32'h3a8316d3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037225),
	.w1(32'h3c414999),
	.w2(32'h3c80f13f),
	.w3(32'h3bffa7c4),
	.w4(32'h3c5c14ed),
	.w5(32'h3c825665),
	.w6(32'h3c0a7e34),
	.w7(32'h3c13e258),
	.w8(32'h3c986425),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc062cf),
	.w1(32'h3cc1c979),
	.w2(32'h3c56921f),
	.w3(32'h3c8f08b8),
	.w4(32'h3c94f8b0),
	.w5(32'h3c29f63e),
	.w6(32'h3c8f4045),
	.w7(32'h3c242207),
	.w8(32'h3c5f76b8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29fd99),
	.w1(32'hbbe4aa10),
	.w2(32'h3b38a900),
	.w3(32'h3c72e7ad),
	.w4(32'hbb4bcb88),
	.w5(32'h3bca61ce),
	.w6(32'hbaa3c5a1),
	.w7(32'h3adfc642),
	.w8(32'h3894a2eb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37decd5e),
	.w1(32'h3b0c6b79),
	.w2(32'h39f75191),
	.w3(32'h3909a647),
	.w4(32'h3a9e2052),
	.w5(32'h38a22122),
	.w6(32'h3aa38116),
	.w7(32'h3a1bc9f2),
	.w8(32'h3c034454),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8ec2),
	.w1(32'hbbd13074),
	.w2(32'hbb0f5ff1),
	.w3(32'h3c1e0164),
	.w4(32'h3c09345d),
	.w5(32'h3b892bc8),
	.w6(32'h3b8764ba),
	.w7(32'h3bb7ad0b),
	.w8(32'h3c768aab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c454875),
	.w1(32'h3c0fc1f6),
	.w2(32'h3bec6e21),
	.w3(32'h3c3ccdd7),
	.w4(32'h3c12bdfb),
	.w5(32'h3bc7ffce),
	.w6(32'h3c3867b6),
	.w7(32'h3c0cf637),
	.w8(32'h3c4a2717),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ffea),
	.w1(32'hbc744914),
	.w2(32'hbc3a72ee),
	.w3(32'h3bc73476),
	.w4(32'hbbb0e2a4),
	.w5(32'h3a1da8c6),
	.w6(32'h3b691bbe),
	.w7(32'h3c231866),
	.w8(32'hbc066928),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947f939),
	.w1(32'h3b963511),
	.w2(32'h3bb6eba8),
	.w3(32'hbb1562b4),
	.w4(32'h3b1f6911),
	.w5(32'hb95c27f4),
	.w6(32'hbc137512),
	.w7(32'hbbab2a04),
	.w8(32'hbd050de1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce042c),
	.w1(32'hbc33f1d3),
	.w2(32'hbc9aaac5),
	.w3(32'hbce6c1e9),
	.w4(32'hbc8d7f58),
	.w5(32'hbcac22d1),
	.w6(32'hbca8f18e),
	.w7(32'hbcc83d00),
	.w8(32'hb9ddc7f1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5b5ec),
	.w1(32'hbb6db360),
	.w2(32'hba6fc8ff),
	.w3(32'hb9cd18c6),
	.w4(32'hbacca79f),
	.w5(32'h3a9d176e),
	.w6(32'hba3ba260),
	.w7(32'h3b5d76b8),
	.w8(32'h3b80cf6b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6f1b5),
	.w1(32'h3be9665f),
	.w2(32'hba90a52d),
	.w3(32'hba21fc17),
	.w4(32'h3aed46c6),
	.w5(32'hbacf7d32),
	.w6(32'h3b747196),
	.w7(32'hba6b739c),
	.w8(32'h380d9714),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ad88),
	.w1(32'h3b8a56ad),
	.w2(32'h3a95f9c7),
	.w3(32'h393747b5),
	.w4(32'h3aec9c76),
	.w5(32'h389966cf),
	.w6(32'h3b159c8b),
	.w7(32'h3a497523),
	.w8(32'hbcbf4a2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe16de),
	.w1(32'hbcb0b086),
	.w2(32'hbce6cc0d),
	.w3(32'hbcc8f91c),
	.w4(32'hbcc5082e),
	.w5(32'hbce33cd6),
	.w6(32'hbcc99e6d),
	.w7(32'hbcca6b19),
	.w8(32'h3c567391),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d8257),
	.w1(32'h3c30555d),
	.w2(32'h3b147800),
	.w3(32'h3c0c6d6c),
	.w4(32'h3bac99c6),
	.w5(32'hb9abdbca),
	.w6(32'h3bfcb433),
	.w7(32'h39619e6f),
	.w8(32'h3aaf70d8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f11e2),
	.w1(32'h3bb8add4),
	.w2(32'h3bfa95d2),
	.w3(32'h3b8e3064),
	.w4(32'h3bd54d40),
	.w5(32'h3bfe2fba),
	.w6(32'h3b904df0),
	.w7(32'h3b9b562d),
	.w8(32'h3b55e751),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b312ee5),
	.w1(32'hbb5c0f5a),
	.w2(32'hbae46503),
	.w3(32'h3b98fca8),
	.w4(32'h3c3b8d81),
	.w5(32'h3be9130e),
	.w6(32'h3a8e3f95),
	.w7(32'h3b4fee2e),
	.w8(32'hbbe793e0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8b0bb),
	.w1(32'h3c5eb05d),
	.w2(32'h3b0b453b),
	.w3(32'hbcaf4cbe),
	.w4(32'hbd069904),
	.w5(32'h3b9f8715),
	.w6(32'hbc2200bd),
	.w7(32'hbc4bc316),
	.w8(32'hbb6fec00),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57de22),
	.w1(32'hbb9e186c),
	.w2(32'hbb61eaf8),
	.w3(32'h3b360f3f),
	.w4(32'h3a5a4ea4),
	.w5(32'hba3e822a),
	.w6(32'hbb96e9c0),
	.w7(32'hbb4f3954),
	.w8(32'h3a8d8f06),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba835fba),
	.w1(32'hbb5ef6fc),
	.w2(32'hbaa497e1),
	.w3(32'h3bbd3502),
	.w4(32'h3b4c4f6f),
	.w5(32'h3b0c0c3d),
	.w6(32'h3aded689),
	.w7(32'hba5a1b8c),
	.w8(32'hbcad32e5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c6377),
	.w1(32'hbc04b9e6),
	.w2(32'hbb5b63af),
	.w3(32'hbc263a44),
	.w4(32'hbb883986),
	.w5(32'hbbdb1c5d),
	.w6(32'hbc4bcb81),
	.w7(32'hbc5a94ec),
	.w8(32'h3c349729),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b732506),
	.w1(32'hbbc956b0),
	.w2(32'hbb9a087b),
	.w3(32'hbbda9856),
	.w4(32'hbc990a74),
	.w5(32'h3c1ad51a),
	.w6(32'h3cbccedd),
	.w7(32'h3c697814),
	.w8(32'hbbcd24b4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48d33d),
	.w1(32'hbbb58c44),
	.w2(32'hbc53895b),
	.w3(32'hbad4091a),
	.w4(32'h3b5935ee),
	.w5(32'hbbfaac44),
	.w6(32'h39a8a8d3),
	.w7(32'hbba76369),
	.w8(32'h3c1af6ca),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e07b),
	.w1(32'h3b6f76b2),
	.w2(32'h3bfb7eb8),
	.w3(32'hbb9fe656),
	.w4(32'hbb0cf678),
	.w5(32'h3a8abb46),
	.w6(32'h3b9da83b),
	.w7(32'h3c58e90c),
	.w8(32'hbb4b194f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38bbd3),
	.w1(32'hbb9c905f),
	.w2(32'hbb30f14e),
	.w3(32'h3a485412),
	.w4(32'h3a74e6d8),
	.w5(32'hbb3b40a3),
	.w6(32'h3ab347f1),
	.w7(32'hbb649ef4),
	.w8(32'hbb58ea30),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1acca9),
	.w1(32'hbb460cb6),
	.w2(32'hba8bf80c),
	.w3(32'h3aba44b1),
	.w4(32'h39b5e303),
	.w5(32'h393bac96),
	.w6(32'hbac56abd),
	.w7(32'hbb314590),
	.w8(32'hbbcfbf14),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d253),
	.w1(32'hbbcccfb9),
	.w2(32'hbb621186),
	.w3(32'h3b51ee40),
	.w4(32'h3b037994),
	.w5(32'hba64c9cd),
	.w6(32'hbb8c23e9),
	.w7(32'hbbc62f38),
	.w8(32'hbbafd1bd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9deb0f),
	.w1(32'h3c2943d6),
	.w2(32'h3b922331),
	.w3(32'hbc65a261),
	.w4(32'hbcfb52e1),
	.w5(32'hbcaf6f21),
	.w6(32'h3b654b8a),
	.w7(32'hbbf6d6f7),
	.w8(32'h3b9c20cf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac63ba2),
	.w1(32'h3bc93872),
	.w2(32'h392fe3d2),
	.w3(32'hbbcf5040),
	.w4(32'hbb2e6b66),
	.w5(32'hba0d4680),
	.w6(32'h3c274d98),
	.w7(32'h3c164947),
	.w8(32'h3b9f407d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb56bf9f6),
	.w1(32'h3c48bf8f),
	.w2(32'hbbeee9be),
	.w3(32'hbc461447),
	.w4(32'hbc53f045),
	.w5(32'h3b21b3ae),
	.w6(32'hbcc62c4a),
	.w7(32'hbbaf6f32),
	.w8(32'hbc539f23),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b9443),
	.w1(32'hbc7097a4),
	.w2(32'hbcb4ee07),
	.w3(32'hbc195c30),
	.w4(32'hbc8eb609),
	.w5(32'hbba8de94),
	.w6(32'hbb7aef53),
	.w7(32'hbc4202d4),
	.w8(32'hb9f0798d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bb93),
	.w1(32'h3c9983f7),
	.w2(32'h3c8cac3b),
	.w3(32'h3b3ff51f),
	.w4(32'h3c038f1d),
	.w5(32'hbb556969),
	.w6(32'hbbec7784),
	.w7(32'h3bb190ea),
	.w8(32'h3c303f85),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9d92),
	.w1(32'h3d17ddb9),
	.w2(32'hbc04b998),
	.w3(32'hbcf194a5),
	.w4(32'hbc1acff0),
	.w5(32'hbaa08c75),
	.w6(32'h3c6a90d5),
	.w7(32'h3b7a3fde),
	.w8(32'h3bf8de5a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108ce8),
	.w1(32'h3aafb2be),
	.w2(32'h3b9aed56),
	.w3(32'h3c21c6f7),
	.w4(32'h3bf2b7a1),
	.w5(32'h3c14dd6c),
	.w6(32'h3b8b757a),
	.w7(32'h3bf50931),
	.w8(32'hbbfffc20),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4535d6),
	.w1(32'h39aac405),
	.w2(32'hbb1c7150),
	.w3(32'hbb6ad80f),
	.w4(32'hbbb24616),
	.w5(32'hb861fc9e),
	.w6(32'h39e1fd9e),
	.w7(32'h376c49dc),
	.w8(32'hbb017c85),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16d573),
	.w1(32'h3c3a3178),
	.w2(32'hbbedff2c),
	.w3(32'hbc7f390f),
	.w4(32'hbccb7899),
	.w5(32'hbbab1a01),
	.w6(32'hbad0acdd),
	.w7(32'h3ac7af04),
	.w8(32'hbbe40f30),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb15dff),
	.w1(32'hbb986069),
	.w2(32'hbc312559),
	.w3(32'hbc49493e),
	.w4(32'hbc3a5299),
	.w5(32'hbcaff0ec),
	.w6(32'hbb27afe7),
	.w7(32'hbbf0bc79),
	.w8(32'hbb158620),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956ebf9),
	.w1(32'hbbc0e1fd),
	.w2(32'hbb7d049c),
	.w3(32'h3c5d4567),
	.w4(32'h3c06e862),
	.w5(32'h3bdb705d),
	.w6(32'hbb801ef3),
	.w7(32'hbb9e2f44),
	.w8(32'h3bb3e265),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2dd2),
	.w1(32'h3d1c239b),
	.w2(32'h3c8febcb),
	.w3(32'hbba6efb1),
	.w4(32'hbc9c5402),
	.w5(32'h3caa2d75),
	.w6(32'h3ce681c6),
	.w7(32'hbc33980e),
	.w8(32'hb9f0b9fc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule