module layer_10_featuremap_323(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8afb67),
	.w1(32'hbbdce1da),
	.w2(32'hba9b4e54),
	.w3(32'hb9e833ab),
	.w4(32'hbb2f8477),
	.w5(32'hbbad3ccb),
	.w6(32'hbba7da19),
	.w7(32'hbb9c7347),
	.w8(32'hbb09a03b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf733f3),
	.w1(32'hbbabff8c),
	.w2(32'h3bbe96a3),
	.w3(32'hbbad80c9),
	.w4(32'hbaa2b47b),
	.w5(32'hbc5a19ac),
	.w6(32'hbbab5cb4),
	.w7(32'hbb572c77),
	.w8(32'hb99e4b51),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc134e5),
	.w1(32'h3ba04397),
	.w2(32'h3ac48a37),
	.w3(32'hbabfc31b),
	.w4(32'hbad72a84),
	.w5(32'hbab9930b),
	.w6(32'h3c894300),
	.w7(32'h3c487505),
	.w8(32'hbbbdf55f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6989b5),
	.w1(32'hbab3a8fe),
	.w2(32'h3ac09177),
	.w3(32'hbb948e6d),
	.w4(32'hbbfb2e55),
	.w5(32'hbbb8a8dd),
	.w6(32'hba6aa6aa),
	.w7(32'hb9dde680),
	.w8(32'hbc2445c6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5861),
	.w1(32'hb894b563),
	.w2(32'h3b84f6c2),
	.w3(32'hba959e79),
	.w4(32'h3984fe32),
	.w5(32'h3b5b0dc1),
	.w6(32'h3a8475a2),
	.w7(32'h3a3edee0),
	.w8(32'hb9fffab5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39102d78),
	.w1(32'h3b8aab12),
	.w2(32'h3b0a1031),
	.w3(32'hbb15c8c3),
	.w4(32'hbad5335f),
	.w5(32'hbb0e264f),
	.w6(32'h3a872e43),
	.w7(32'h3af89c53),
	.w8(32'hbac95c12),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3ff6),
	.w1(32'h3a2ef675),
	.w2(32'h3b458d18),
	.w3(32'hbb08e38a),
	.w4(32'h3b00839c),
	.w5(32'h3c6cb91a),
	.w6(32'h39c5589d),
	.w7(32'h3a17801d),
	.w8(32'h3c2eb887),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c935b),
	.w1(32'h3b84c6f4),
	.w2(32'h3c5938e8),
	.w3(32'h3cb4c1ff),
	.w4(32'h3bb2f899),
	.w5(32'hb9b68b6f),
	.w6(32'h3bde5d85),
	.w7(32'h3c22c223),
	.w8(32'h3ae31429),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d348),
	.w1(32'h3b9889cb),
	.w2(32'h3b77a9fa),
	.w3(32'h3989e09e),
	.w4(32'h3b0c4904),
	.w5(32'h3ac98fb3),
	.w6(32'hb9ca1583),
	.w7(32'hba4dde2a),
	.w8(32'h382809b0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2be068),
	.w1(32'hb935a57b),
	.w2(32'h3a3539d7),
	.w3(32'hbaf065c0),
	.w4(32'hbbac9cd0),
	.w5(32'h3c030029),
	.w6(32'h3c011062),
	.w7(32'h3ba599e8),
	.w8(32'h3c5639c0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a4773),
	.w1(32'h3bdcde3f),
	.w2(32'h3bf2e139),
	.w3(32'hbb203365),
	.w4(32'hbba15e72),
	.w5(32'h3bed38f1),
	.w6(32'h3b23a777),
	.w7(32'h3b1385d6),
	.w8(32'h3c324836),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891060),
	.w1(32'h3bfd2e7c),
	.w2(32'h3bcb03bd),
	.w3(32'h3b68868d),
	.w4(32'hbc07394a),
	.w5(32'hbc217291),
	.w6(32'hbc40ef61),
	.w7(32'hbbfae862),
	.w8(32'hbc07acce),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc455),
	.w1(32'h3b38c95f),
	.w2(32'h3b45ce51),
	.w3(32'h3be9f148),
	.w4(32'h3b5c795b),
	.w5(32'hbc16d08b),
	.w6(32'h3c3a997a),
	.w7(32'h3ba6db07),
	.w8(32'hbb952091),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc814ee3),
	.w1(32'hbc0a98cb),
	.w2(32'h3b89034a),
	.w3(32'hbac052d0),
	.w4(32'hba7de248),
	.w5(32'h3c09006b),
	.w6(32'h3aad5e95),
	.w7(32'h3b2febc8),
	.w8(32'h3b5b8edd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de3682),
	.w1(32'h3bddb7a7),
	.w2(32'h3ab71b81),
	.w3(32'hbaa65599),
	.w4(32'h3a204683),
	.w5(32'hba70bfec),
	.w6(32'h3b9c6fe7),
	.w7(32'h3b753ede),
	.w8(32'h3b8f074a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406506),
	.w1(32'hbc3ea31a),
	.w2(32'h3ab1e9be),
	.w3(32'hbaa6f018),
	.w4(32'hbbc1f145),
	.w5(32'h372e4f6c),
	.w6(32'h3aec41b1),
	.w7(32'h3b4a408b),
	.w8(32'h3bf63bf9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05a08c),
	.w1(32'h3c0a3b31),
	.w2(32'h3c1ec9f8),
	.w3(32'h3ba2a65b),
	.w4(32'h3b0d5dd8),
	.w5(32'hbb950477),
	.w6(32'h3c0f8a07),
	.w7(32'h3b7b3a5a),
	.w8(32'hbbab806c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71ae79),
	.w1(32'h3bbf3338),
	.w2(32'h3b32c552),
	.w3(32'h3c803279),
	.w4(32'h3bc5f69d),
	.w5(32'hbbc732b0),
	.w6(32'h3c3867ab),
	.w7(32'h3c5a8a53),
	.w8(32'h3b168ea8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dff73),
	.w1(32'h3add9643),
	.w2(32'hba4a5088),
	.w3(32'h3c8d495c),
	.w4(32'h3c0d5739),
	.w5(32'h3c6c3887),
	.w6(32'h3c141174),
	.w7(32'h3bf089ad),
	.w8(32'h3b4c76ea),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbff5f0),
	.w1(32'h3c20822f),
	.w2(32'hba9e101a),
	.w3(32'h3c430259),
	.w4(32'hbae9b29a),
	.w5(32'hbb6790e3),
	.w6(32'hbb1f0660),
	.w7(32'hbba7098f),
	.w8(32'hbbd93c39),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140bef),
	.w1(32'h3914440f),
	.w2(32'h3b576068),
	.w3(32'h3b98539f),
	.w4(32'hbbc1a1c9),
	.w5(32'h39a8210c),
	.w6(32'h3af45ba8),
	.w7(32'hbba81d92),
	.w8(32'hbba405cd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fc57),
	.w1(32'hbbca9ac3),
	.w2(32'h3ab16c76),
	.w3(32'hbbe7ce73),
	.w4(32'h38209fd1),
	.w5(32'h3c4ffbdc),
	.w6(32'hbbf12d33),
	.w7(32'hba7097f1),
	.w8(32'h3bc70943),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd5ba),
	.w1(32'h3c3c248d),
	.w2(32'h3ad5134a),
	.w3(32'h3c653277),
	.w4(32'hbb7c68b6),
	.w5(32'h3bc26fad),
	.w6(32'h3cbd1c99),
	.w7(32'hbb98eb9e),
	.w8(32'h3c41c65b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de38f),
	.w1(32'h3b37c1eb),
	.w2(32'h3b87be2c),
	.w3(32'hbbbbcfb5),
	.w4(32'hbb91e8ed),
	.w5(32'h3c8e2a21),
	.w6(32'hba03f325),
	.w7(32'h3c7f7e36),
	.w8(32'h3d3ccecc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbebbba),
	.w1(32'hbbccc50e),
	.w2(32'h3c159fdb),
	.w3(32'h3c314996),
	.w4(32'h3bf00a4b),
	.w5(32'h3bff7761),
	.w6(32'h3d1c048d),
	.w7(32'h3cb1795c),
	.w8(32'h3b297a7e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f1ab),
	.w1(32'hb94dbdf4),
	.w2(32'h3bad796b),
	.w3(32'h3b7dd725),
	.w4(32'h3aab79c0),
	.w5(32'h3ab48393),
	.w6(32'hbb84cfb0),
	.w7(32'hb8c1ae9c),
	.w8(32'hbae7a251),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20c8c3),
	.w1(32'h3c10db93),
	.w2(32'hbb32840c),
	.w3(32'h3b63254e),
	.w4(32'h3a3ecdb1),
	.w5(32'h3b666b78),
	.w6(32'h3b9f7101),
	.w7(32'h3ab6d91e),
	.w8(32'h3a3774bc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b896e39),
	.w1(32'h3b54aa4e),
	.w2(32'hbab60e85),
	.w3(32'hb9b3ee18),
	.w4(32'hbbd11f45),
	.w5(32'hb872c293),
	.w6(32'h3a1425a8),
	.w7(32'hbc0d6fdd),
	.w8(32'h3b91f883),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf207ce),
	.w1(32'hbca4bd53),
	.w2(32'hbb9b58e6),
	.w3(32'hbc814d08),
	.w4(32'hbaa35659),
	.w5(32'hbbcf7f97),
	.w6(32'hbc81bc4e),
	.w7(32'hbb932781),
	.w8(32'hbc273123),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdeb4d),
	.w1(32'hbc348bee),
	.w2(32'hbb62e411),
	.w3(32'hba251454),
	.w4(32'hbba40f23),
	.w5(32'hbb7b4a2d),
	.w6(32'h3a02211e),
	.w7(32'hbbf14bfd),
	.w8(32'hbb8ca902),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23148d),
	.w1(32'h3af88f68),
	.w2(32'hbc308222),
	.w3(32'h3c1afa36),
	.w4(32'h3abd8c84),
	.w5(32'hbc0b9428),
	.w6(32'hb6e887ec),
	.w7(32'h3a3d520f),
	.w8(32'hbbca8cd5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad1b88),
	.w1(32'hbbd500c9),
	.w2(32'hbb1e33b2),
	.w3(32'hbc360ac1),
	.w4(32'hbba01c9a),
	.w5(32'h3bfcb50c),
	.w6(32'h3b4a2c2c),
	.w7(32'h3c181afc),
	.w8(32'h3cfda1c1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf57182),
	.w1(32'hbc6500d1),
	.w2(32'hbbf17040),
	.w3(32'h3c755b8d),
	.w4(32'h3bec0ec6),
	.w5(32'hbaf8b3cf),
	.w6(32'h3bc6e248),
	.w7(32'hbbbd9a42),
	.w8(32'h3c10fe62),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118974),
	.w1(32'hbc38320b),
	.w2(32'hb976a2c3),
	.w3(32'hbc005ef4),
	.w4(32'hbb4b2480),
	.w5(32'h3bbe6c4c),
	.w6(32'hbc58598c),
	.w7(32'h3b52b515),
	.w8(32'h3bda5560),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d304a),
	.w1(32'hbc52907a),
	.w2(32'hbb8d3dbe),
	.w3(32'hbc1f6884),
	.w4(32'hbb3cecba),
	.w5(32'hbbe29954),
	.w6(32'hbb73b8ff),
	.w7(32'h3c27895d),
	.w8(32'h3b67d7fe),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22427d),
	.w1(32'h3c4ac3dc),
	.w2(32'h3ad7e173),
	.w3(32'h3c093d80),
	.w4(32'h3bad59c7),
	.w5(32'hbba12ee9),
	.w6(32'h3cb21eb7),
	.w7(32'h3a7ae3c1),
	.w8(32'h3bedde66),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3933c),
	.w1(32'h3bde4569),
	.w2(32'hbaba83b9),
	.w3(32'hbbbec2eb),
	.w4(32'h3c8d9966),
	.w5(32'hbbb3f230),
	.w6(32'hbb92a842),
	.w7(32'h3b9de540),
	.w8(32'hbba122be),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8ee5e),
	.w1(32'hbb90b972),
	.w2(32'h3bea1b79),
	.w3(32'hbc9c0274),
	.w4(32'hbc30279a),
	.w5(32'hbb71cc92),
	.w6(32'hbc7b1282),
	.w7(32'hbba8e418),
	.w8(32'hbb33846a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf879),
	.w1(32'hbbd6e302),
	.w2(32'h3bfeff0e),
	.w3(32'hbc84be23),
	.w4(32'hbc1602cc),
	.w5(32'h3c2d4b43),
	.w6(32'hbc8b32b6),
	.w7(32'hbc24fabc),
	.w8(32'hbbb081c2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3e1e0),
	.w1(32'hb939f399),
	.w2(32'h3b44cab6),
	.w3(32'hbbafd385),
	.w4(32'hbaad595a),
	.w5(32'h3c87b074),
	.w6(32'hbbe5b998),
	.w7(32'h3b8bffdf),
	.w8(32'h3c9f6155),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15157b),
	.w1(32'h3b9cd80a),
	.w2(32'h3cc3b10d),
	.w3(32'hb9162362),
	.w4(32'h3c0580ae),
	.w5(32'hbac35f06),
	.w6(32'hbc5bf35b),
	.w7(32'h3cb8086e),
	.w8(32'hbb9524a8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046a95),
	.w1(32'hb80a9c8a),
	.w2(32'h3be30764),
	.w3(32'hbb4f53b4),
	.w4(32'h3b3fd1c5),
	.w5(32'h3a877a9a),
	.w6(32'hbba637ea),
	.w7(32'h3b959ce6),
	.w8(32'hbb1a902a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3652d),
	.w1(32'hbb3042a6),
	.w2(32'hbbbed919),
	.w3(32'hbb9b3666),
	.w4(32'hbab1b737),
	.w5(32'hbb820d79),
	.w6(32'hbb902bee),
	.w7(32'h3a27831c),
	.w8(32'h3b6f7151),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94d72b),
	.w1(32'h3b4f33dc),
	.w2(32'h3b9badd2),
	.w3(32'h3c433227),
	.w4(32'h3b5932b0),
	.w5(32'hbb2fc753),
	.w6(32'h3c281ad3),
	.w7(32'h3c326188),
	.w8(32'h3a9e47b9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001e55),
	.w1(32'hbb858864),
	.w2(32'h3aa4658b),
	.w3(32'hbb733b33),
	.w4(32'hbaf4197e),
	.w5(32'h3c06d5fa),
	.w6(32'hbbb0691e),
	.w7(32'h3b9bfcb4),
	.w8(32'h3bca3a1c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947afcb),
	.w1(32'hbbfca475),
	.w2(32'hbb820a53),
	.w3(32'h3bb29bec),
	.w4(32'h3a6e740b),
	.w5(32'h3a5ef9f0),
	.w6(32'hbb1121f4),
	.w7(32'h3ab55092),
	.w8(32'h3bbb8d98),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5719d6),
	.w1(32'hb772d9bc),
	.w2(32'hba82988e),
	.w3(32'hba921551),
	.w4(32'hbad60da8),
	.w5(32'h3b6a40fa),
	.w6(32'h3b7d57ae),
	.w7(32'h3b13b011),
	.w8(32'h3b555d65),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb54282),
	.w1(32'h3b298a0d),
	.w2(32'h3b9d3309),
	.w3(32'h3c8c8ecc),
	.w4(32'h3c8fdea0),
	.w5(32'hb894e27c),
	.w6(32'h3c7ad6d3),
	.w7(32'h3c2f1feb),
	.w8(32'h3a44bf42),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07b170),
	.w1(32'h3ad08fe5),
	.w2(32'hbaf65622),
	.w3(32'hb9fca1df),
	.w4(32'hb9d41584),
	.w5(32'hbb8932fa),
	.w6(32'hbb8092dd),
	.w7(32'h3b0f7e60),
	.w8(32'hbc243212),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045ff7),
	.w1(32'hbc0625ee),
	.w2(32'hbae30d62),
	.w3(32'hbbc997fe),
	.w4(32'h3a69ba11),
	.w5(32'hbbf7af87),
	.w6(32'hbc117aae),
	.w7(32'hba4c5164),
	.w8(32'hbc66ee15),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3171f6),
	.w1(32'h3c8b68a8),
	.w2(32'hbbc3fff6),
	.w3(32'h3cb8bcd4),
	.w4(32'hba9b8bd2),
	.w5(32'hbb2f500f),
	.w6(32'h3d12d2c5),
	.w7(32'hbc0b154c),
	.w8(32'hbb247705),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb626607),
	.w1(32'h3925fa38),
	.w2(32'hbb31a175),
	.w3(32'h3b3476b5),
	.w4(32'h384f10e8),
	.w5(32'h3c687eb1),
	.w6(32'h3a809b93),
	.w7(32'hb8c40cbd),
	.w8(32'h3c175329),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5c72e),
	.w1(32'hba7c6695),
	.w2(32'h3a9ea714),
	.w3(32'h3b45602b),
	.w4(32'hbc4ac9f9),
	.w5(32'h3b33f46a),
	.w6(32'hbafa58b2),
	.w7(32'hbc26db04),
	.w8(32'h3bc72029),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ac78),
	.w1(32'hbbd474d2),
	.w2(32'h3babde28),
	.w3(32'h3a2019f6),
	.w4(32'h3b8928d1),
	.w5(32'h3c8c4ed3),
	.w6(32'h3c5ddd99),
	.w7(32'h3bef2776),
	.w8(32'h3c146f4b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c029b68),
	.w1(32'h3c5507dc),
	.w2(32'h3baaacdc),
	.w3(32'h3a2c75a8),
	.w4(32'hbb613b75),
	.w5(32'hbb9be3ef),
	.w6(32'hbbe630fd),
	.w7(32'hbba85d1c),
	.w8(32'hbc08844e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32c009),
	.w1(32'hbcb2f0c5),
	.w2(32'h3b2e556b),
	.w3(32'hbc5074f0),
	.w4(32'hbc1d994d),
	.w5(32'h3c7e1c58),
	.w6(32'hbc864b9e),
	.w7(32'h3aaf9cf3),
	.w8(32'h3cd21ea1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38124c),
	.w1(32'hbb7fed34),
	.w2(32'h3c8c1f3b),
	.w3(32'h3b950920),
	.w4(32'h3c8903c4),
	.w5(32'hbb0f4b93),
	.w6(32'hbaa7f5dc),
	.w7(32'h3ce2a803),
	.w8(32'hbb681c98),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50012c),
	.w1(32'h3c84265a),
	.w2(32'h3c0e5dd5),
	.w3(32'h3be739df),
	.w4(32'hbadd9270),
	.w5(32'hbb37784f),
	.w6(32'h3c3b3350),
	.w7(32'hbb150bef),
	.w8(32'hbbfb0a75),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0ee7f),
	.w1(32'hbb483867),
	.w2(32'h3a4a3061),
	.w3(32'hbb861592),
	.w4(32'hbacaf255),
	.w5(32'h399c52d9),
	.w6(32'hbc1160ee),
	.w7(32'hbb63628f),
	.w8(32'hbc2d1bb7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5c373),
	.w1(32'hbc366736),
	.w2(32'hbadf249d),
	.w3(32'hbb5e0485),
	.w4(32'h3bafc365),
	.w5(32'hbb756040),
	.w6(32'hbc4f0e52),
	.w7(32'hbad8782c),
	.w8(32'hbba055c5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ce9f4),
	.w1(32'hbb23bda5),
	.w2(32'hbb938b9d),
	.w3(32'h3b1ddad0),
	.w4(32'h3943edb2),
	.w5(32'hb963b091),
	.w6(32'h399cddab),
	.w7(32'hbb191d13),
	.w8(32'hbb89e0a9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53d14),
	.w1(32'hbb219613),
	.w2(32'hbad7a7c4),
	.w3(32'h3c141d1b),
	.w4(32'hbb4cf552),
	.w5(32'hbbce86f9),
	.w6(32'h3b0d5959),
	.w7(32'hbadcfe62),
	.w8(32'hbc2b9124),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f58e),
	.w1(32'hba20a50b),
	.w2(32'hbb42c422),
	.w3(32'hbbf7a2dd),
	.w4(32'hbc1b5409),
	.w5(32'h3c52b8aa),
	.w6(32'hbbf3ce16),
	.w7(32'hbaf301ca),
	.w8(32'h3c4d2b03),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcce2f7),
	.w1(32'hbc4ed04c),
	.w2(32'h3be928e1),
	.w3(32'hbc0a9de4),
	.w4(32'h3b5cae06),
	.w5(32'hbbfae769),
	.w6(32'hbb939e07),
	.w7(32'h3b624b43),
	.w8(32'hbc8595eb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75164d),
	.w1(32'hbbebdc9e),
	.w2(32'hbc6e192e),
	.w3(32'hbb934a20),
	.w4(32'hbb86c6be),
	.w5(32'h3b1cfad5),
	.w6(32'hbb82a31c),
	.w7(32'hbbe213ec),
	.w8(32'hbbd9e61b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97fd8c),
	.w1(32'h3c159abf),
	.w2(32'h3992718e),
	.w3(32'hbb4b7f5a),
	.w4(32'hbb88bb44),
	.w5(32'h3ad269cd),
	.w6(32'hbc8b5b6b),
	.w7(32'hbc2b7bec),
	.w8(32'h3a048beb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae8ba),
	.w1(32'hbafbc127),
	.w2(32'hbb9c2852),
	.w3(32'h3bb4fe61),
	.w4(32'hbbd1485e),
	.w5(32'hbbef555e),
	.w6(32'h3c350df4),
	.w7(32'h3b0124ea),
	.w8(32'hbc498c62),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab27179),
	.w1(32'h3b7e1ddc),
	.w2(32'h3aed257e),
	.w3(32'h3b2ec88b),
	.w4(32'h3baccbd1),
	.w5(32'h3cb8384f),
	.w6(32'h3c257eff),
	.w7(32'h393ec539),
	.w8(32'h3ce39846),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cf1ca),
	.w1(32'h3ce1a03b),
	.w2(32'hbb154258),
	.w3(32'h3cf83e4a),
	.w4(32'hb99024b4),
	.w5(32'hbb3ea807),
	.w6(32'h3c966b56),
	.w7(32'hbc3a51e2),
	.w8(32'hbb18e43e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9cd9),
	.w1(32'hbb960544),
	.w2(32'h3b95a21c),
	.w3(32'hbc9204b0),
	.w4(32'hbb9c5fef),
	.w5(32'h3bbc5078),
	.w6(32'hbc990002),
	.w7(32'hbad7ecf6),
	.w8(32'h3b640846),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3065c),
	.w1(32'h3b06c990),
	.w2(32'hba672eb7),
	.w3(32'h3b5d4e8c),
	.w4(32'hbac401e9),
	.w5(32'hbb0770e8),
	.w6(32'hbb3735f3),
	.w7(32'hbb234eef),
	.w8(32'hbc23640d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3d1e),
	.w1(32'hb99c1ce3),
	.w2(32'h3ad72253),
	.w3(32'hba603eea),
	.w4(32'hbbbfc42f),
	.w5(32'hbb92ea83),
	.w6(32'h3b6366d9),
	.w7(32'hba8f6714),
	.w8(32'h3b18918a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f030ef),
	.w1(32'hbb3ea15a),
	.w2(32'h3984137e),
	.w3(32'hbb4abf24),
	.w4(32'hb8282974),
	.w5(32'h3a200234),
	.w6(32'h3b8a57f4),
	.w7(32'h3b2e4ff4),
	.w8(32'h3a1cd9db),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade15d5),
	.w1(32'hbb80d8e7),
	.w2(32'hba9f084d),
	.w3(32'hbbc544df),
	.w4(32'hba43482c),
	.w5(32'hbb7a7aed),
	.w6(32'hbc1869de),
	.w7(32'h396df9f6),
	.w8(32'h3b2cbe7a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7863d4),
	.w1(32'hb9f4d7fc),
	.w2(32'h3aa67549),
	.w3(32'hba254d1d),
	.w4(32'hbac757e2),
	.w5(32'hbbec5b22),
	.w6(32'hba114a71),
	.w7(32'h3a3cfcdb),
	.w8(32'hbbd8ea1a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab3e2e),
	.w1(32'h3c00c747),
	.w2(32'h3b358eab),
	.w3(32'h3c128e4f),
	.w4(32'h3bd437a5),
	.w5(32'h3c0a8a50),
	.w6(32'h3c3bac60),
	.w7(32'h3c2c78fa),
	.w8(32'h38870dd5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121898),
	.w1(32'h3c81e790),
	.w2(32'h3ca12988),
	.w3(32'h3c14dbb5),
	.w4(32'h3c1f38bf),
	.w5(32'hbba003e9),
	.w6(32'hbc3eec42),
	.w7(32'h3ba4a1f7),
	.w8(32'h36d8c92b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0f9c8),
	.w1(32'h3a3b5f9a),
	.w2(32'h3b72d254),
	.w3(32'h3c0817b1),
	.w4(32'h3b3f06e6),
	.w5(32'h3c1e08ca),
	.w6(32'h3bcd5efb),
	.w7(32'h3bf12f3b),
	.w8(32'h3b109879),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74279d),
	.w1(32'hbada27e5),
	.w2(32'hbb7467d2),
	.w3(32'h3b771308),
	.w4(32'hba7780ca),
	.w5(32'h3b11992d),
	.w6(32'h3b3b93df),
	.w7(32'h3b5d8e55),
	.w8(32'h3b10eb4f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b3ff),
	.w1(32'h3bcd15b8),
	.w2(32'h3b30833c),
	.w3(32'h39fd7dc8),
	.w4(32'h3b13de50),
	.w5(32'h3c2eddd0),
	.w6(32'h3a94abbe),
	.w7(32'h3b368225),
	.w8(32'hbb39e735),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9890c6),
	.w1(32'h3a869afe),
	.w2(32'h3b7a861d),
	.w3(32'h3aea58f6),
	.w4(32'hbb31f725),
	.w5(32'hb98d8b63),
	.w6(32'h3aaf3376),
	.w7(32'h3a0caff2),
	.w8(32'hbb358c1e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76ce8a),
	.w1(32'h3bc41280),
	.w2(32'h3a01f19c),
	.w3(32'h3b67252b),
	.w4(32'h3bb85a30),
	.w5(32'hbbe009d8),
	.w6(32'h3bfbca71),
	.w7(32'h3c0ef171),
	.w8(32'h3bad5dab),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3799a2c1),
	.w1(32'h3bb484d6),
	.w2(32'h3b6dff53),
	.w3(32'h3bec2c0d),
	.w4(32'h3c0caec8),
	.w5(32'hba30001f),
	.w6(32'h3d190984),
	.w7(32'h3bc5bef0),
	.w8(32'hbb30fbb0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd52bd),
	.w1(32'hba753642),
	.w2(32'hbc055741),
	.w3(32'h39c1dcfc),
	.w4(32'hbbe4d90d),
	.w5(32'hbc1df6af),
	.w6(32'h3bacc234),
	.w7(32'hba51c590),
	.w8(32'hbb959a73),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0710dd),
	.w1(32'hb86b407c),
	.w2(32'hbb0fd74b),
	.w3(32'h3a14c393),
	.w4(32'h3bed12a3),
	.w5(32'h3b33b0e0),
	.w6(32'h3cb71f98),
	.w7(32'h3b6de563),
	.w8(32'h3b16580c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b0af),
	.w1(32'h396edfe2),
	.w2(32'hbb8b1ffd),
	.w3(32'h3b88d9c5),
	.w4(32'hbad8d512),
	.w5(32'hbb6bc684),
	.w6(32'h3b35236a),
	.w7(32'hbb47fa82),
	.w8(32'hbbc78b2c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08b593),
	.w1(32'h3c83e32b),
	.w2(32'hbb6a1c4b),
	.w3(32'h3ba4d117),
	.w4(32'h3bca0983),
	.w5(32'hbb925d9c),
	.w6(32'h3c52ae92),
	.w7(32'h3c11a8b2),
	.w8(32'h368100a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8eb3d),
	.w1(32'hbbd98ffe),
	.w2(32'hbc5d5de0),
	.w3(32'hbc0d7346),
	.w4(32'hbb86c990),
	.w5(32'hb9d846d4),
	.w6(32'hbc08961b),
	.w7(32'hbc584b0d),
	.w8(32'hba9d3f2a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966995b),
	.w1(32'h3b8fa19e),
	.w2(32'h3bb70c63),
	.w3(32'h3a69646a),
	.w4(32'h3b927cba),
	.w5(32'hb9fa92f9),
	.w6(32'h3ba84b03),
	.w7(32'h3b8cce92),
	.w8(32'hbbd948a2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a59d),
	.w1(32'hbb71290f),
	.w2(32'h3bfa9380),
	.w3(32'h3b740fa6),
	.w4(32'h3c24462b),
	.w5(32'h3ab05c6b),
	.w6(32'h3c86f02a),
	.w7(32'h3c1bb33d),
	.w8(32'h3b9c3d37),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9242c8),
	.w1(32'hba259724),
	.w2(32'h3ae8c7fa),
	.w3(32'hbc1a2671),
	.w4(32'hbc2206b5),
	.w5(32'hbb974230),
	.w6(32'hbb9cee1e),
	.w7(32'hbbc150d3),
	.w8(32'hbc5830bf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f06a4),
	.w1(32'hbbfbcec8),
	.w2(32'h3a7c8e37),
	.w3(32'hbca19dbb),
	.w4(32'h3a28f6f9),
	.w5(32'hbc57a6d0),
	.w6(32'hba69d36c),
	.w7(32'h3ac34563),
	.w8(32'hbb5e7349),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5862af),
	.w1(32'hbbe26a6a),
	.w2(32'h3aa8db43),
	.w3(32'hbc3ed74b),
	.w4(32'hbb0a4b5f),
	.w5(32'h3af7b8bf),
	.w6(32'hbb9954a6),
	.w7(32'hba425dd1),
	.w8(32'h3b258dc0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cd07),
	.w1(32'h3ca47bb5),
	.w2(32'hbb54c477),
	.w3(32'h3ca3eb19),
	.w4(32'hbc2398ab),
	.w5(32'hbabdae23),
	.w6(32'h3cc30849),
	.w7(32'hbc282a73),
	.w8(32'h3abf00b1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869f60),
	.w1(32'hbc38b83e),
	.w2(32'hbbc2fa93),
	.w3(32'hbba03827),
	.w4(32'hbc15a92d),
	.w5(32'hbbfcf161),
	.w6(32'hbbe46222),
	.w7(32'hbb64ab16),
	.w8(32'h3b502db9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3baa0),
	.w1(32'hbb06c242),
	.w2(32'h380227e1),
	.w3(32'hbb261016),
	.w4(32'hbbc0da33),
	.w5(32'h3ba6adb0),
	.w6(32'h3bd8788a),
	.w7(32'h3bc2333b),
	.w8(32'hbae6164a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09fe6e),
	.w1(32'h3b233164),
	.w2(32'h3b66aaca),
	.w3(32'h39efb955),
	.w4(32'h38df39f7),
	.w5(32'hbaec9487),
	.w6(32'h3a8ff5d0),
	.w7(32'h3c07c88d),
	.w8(32'hbc85a1f2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc491e03),
	.w1(32'h39948e2c),
	.w2(32'h3c14f89a),
	.w3(32'hbbe72786),
	.w4(32'h3b3fe0e9),
	.w5(32'h3b69f207),
	.w6(32'hbb436efc),
	.w7(32'h3c06def4),
	.w8(32'h3c192a1d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb95d80),
	.w1(32'h3c00d721),
	.w2(32'h3c10e6a2),
	.w3(32'h3aca0ab3),
	.w4(32'h3a9716b1),
	.w5(32'hba68dcac),
	.w6(32'h3b818847),
	.w7(32'h3bb41bb3),
	.w8(32'hbb158e6b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fa7ea),
	.w1(32'h3be2bdc4),
	.w2(32'h3bc4bb82),
	.w3(32'h3bfa62bf),
	.w4(32'h3c31bd10),
	.w5(32'h39e7a63b),
	.w6(32'hb9742a2c),
	.w7(32'h3c03587a),
	.w8(32'hb95eb9d2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4c4b6),
	.w1(32'hbba59389),
	.w2(32'h3b9ad944),
	.w3(32'hbba313c5),
	.w4(32'hbb8961f4),
	.w5(32'hb9b9d420),
	.w6(32'h3bb1b100),
	.w7(32'hbbc12295),
	.w8(32'h393cdd11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8c5d),
	.w1(32'hbaa72b1e),
	.w2(32'h3b7dcd7c),
	.w3(32'hbb8b20b7),
	.w4(32'hbbcd4556),
	.w5(32'h3c332c6e),
	.w6(32'hbc1762cb),
	.w7(32'hbba8782f),
	.w8(32'h3c741d06),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73ff22),
	.w1(32'h3b77f53a),
	.w2(32'hbab6bcdb),
	.w3(32'hbb3e4542),
	.w4(32'hbb125071),
	.w5(32'h3b20e4df),
	.w6(32'h3a3d60e7),
	.w7(32'hb9a9bc29),
	.w8(32'h3be198be),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b174d7a),
	.w1(32'hbbbd746a),
	.w2(32'hbc2a380a),
	.w3(32'hba42662b),
	.w4(32'hbb91f992),
	.w5(32'hbaefb245),
	.w6(32'hbb1810d1),
	.w7(32'hbb87dc7a),
	.w8(32'hbbacc33b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c072f),
	.w1(32'h3caf1017),
	.w2(32'h3c63f531),
	.w3(32'h3c5b754f),
	.w4(32'h3caec47b),
	.w5(32'h3b7e8786),
	.w6(32'h3bb92472),
	.w7(32'h3c031b77),
	.w8(32'h3bfcf776),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fc4e2),
	.w1(32'h3b642122),
	.w2(32'h3a98156b),
	.w3(32'hbbe0bd3d),
	.w4(32'h3ab9f45a),
	.w5(32'h3c260bb0),
	.w6(32'hb8e5525d),
	.w7(32'hbbe841ae),
	.w8(32'h3be69de6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc17bc6),
	.w1(32'hbc2d201e),
	.w2(32'hbc427b4b),
	.w3(32'hbb94ac93),
	.w4(32'hbc279c64),
	.w5(32'h3aadd287),
	.w6(32'hbbcf3f41),
	.w7(32'hbc268f40),
	.w8(32'h39f68857),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24fff9),
	.w1(32'h3affdafe),
	.w2(32'hba39b7ad),
	.w3(32'h3b127ca6),
	.w4(32'h3a37a847),
	.w5(32'h3ae5a3e6),
	.w6(32'h3b9d99bf),
	.w7(32'h3a7e3ada),
	.w8(32'h3b413583),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00445c),
	.w1(32'h3a94b1f9),
	.w2(32'h3c0beca9),
	.w3(32'h3bdc609d),
	.w4(32'h3c3529f5),
	.w5(32'hbb44d10a),
	.w6(32'h3c10d29c),
	.w7(32'h3c31f69b),
	.w8(32'hb9da30d7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b5de6),
	.w1(32'hba7e024b),
	.w2(32'h3adef2e4),
	.w3(32'hbb597496),
	.w4(32'hba1b2275),
	.w5(32'h3b0d294e),
	.w6(32'h383d7d76),
	.w7(32'h3650e790),
	.w8(32'h3b5f9dc7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1929d),
	.w1(32'hbaea12fa),
	.w2(32'h3be8dd3d),
	.w3(32'hbbb305b1),
	.w4(32'hbbc62626),
	.w5(32'h3b60b6d9),
	.w6(32'hbbe77e30),
	.w7(32'hbb9892ce),
	.w8(32'h3abe8a34),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc689f7),
	.w1(32'h3c617398),
	.w2(32'h3ce0ef12),
	.w3(32'hbb276bda),
	.w4(32'h3c1b1621),
	.w5(32'h3a8ce98e),
	.w6(32'h3bee7276),
	.w7(32'h3cd90656),
	.w8(32'h3bc12f40),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e70f0),
	.w1(32'h3aaa55ae),
	.w2(32'hba4b7b17),
	.w3(32'h3b6152c2),
	.w4(32'hb99ee0bc),
	.w5(32'h3bec29a8),
	.w6(32'h3a737cc9),
	.w7(32'hbad4de86),
	.w8(32'h3c456e26),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989a499),
	.w1(32'h3baa5c2a),
	.w2(32'h3bee2b3f),
	.w3(32'h3cbef84e),
	.w4(32'h3c3c5dd0),
	.w5(32'h39edd0e2),
	.w6(32'h3d068d65),
	.w7(32'h3ca6211f),
	.w8(32'hbb072de6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac55b65),
	.w1(32'hbbe641ee),
	.w2(32'h3bd863a9),
	.w3(32'h3bcc2cce),
	.w4(32'h3c0b6cf7),
	.w5(32'h3ace75b6),
	.w6(32'hba5b7e3e),
	.w7(32'h3c25e8ad),
	.w8(32'h3ae6a7a6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122754),
	.w1(32'h3c988a12),
	.w2(32'h3cb0ecf6),
	.w3(32'hbb0c21ae),
	.w4(32'h39f69ebe),
	.w5(32'h3a604b04),
	.w6(32'h3b81237f),
	.w7(32'h3c5970cb),
	.w8(32'h3b1c4f2f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa33145),
	.w1(32'h3bcfcac1),
	.w2(32'h3be730d5),
	.w3(32'h3bb27c35),
	.w4(32'h3b57b25b),
	.w5(32'hbb9076fc),
	.w6(32'h3c378ecf),
	.w7(32'h3c04410f),
	.w8(32'h3b84533f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c7a3),
	.w1(32'h3be65aed),
	.w2(32'h3b0c44ea),
	.w3(32'hbbf444b8),
	.w4(32'h3b498646),
	.w5(32'h39ae1d61),
	.w6(32'hbc02e8ab),
	.w7(32'hbb7303a2),
	.w8(32'hb9ae5663),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf613),
	.w1(32'hbb13999e),
	.w2(32'hbb8d7cec),
	.w3(32'h399a9b6f),
	.w4(32'hbb340992),
	.w5(32'h3a9354c8),
	.w6(32'hbb14b3a9),
	.w7(32'hbb867d05),
	.w8(32'hbb14d398),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe1d23),
	.w1(32'hbc30a21c),
	.w2(32'hbba2995d),
	.w3(32'hbb8f3579),
	.w4(32'hbbac4e66),
	.w5(32'hbb7f5c75),
	.w6(32'hbc26baac),
	.w7(32'hbbc79ab4),
	.w8(32'h38eadccb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a41d0),
	.w1(32'h3bbfb659),
	.w2(32'h3bfcb43f),
	.w3(32'hbbb01581),
	.w4(32'h3bb07801),
	.w5(32'h3c0760a3),
	.w6(32'hbb5b548c),
	.w7(32'h3b1d5f17),
	.w8(32'h3be3f020),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c360e5c),
	.w1(32'h3b7f5290),
	.w2(32'h3b0650ae),
	.w3(32'h3bc9a1ec),
	.w4(32'h3be274d1),
	.w5(32'hbbdd11b9),
	.w6(32'h3b85b540),
	.w7(32'h3b34bd47),
	.w8(32'hbb57e345),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c30e0),
	.w1(32'h3b5d43e8),
	.w2(32'h3bf6c110),
	.w3(32'hbc3fe5c4),
	.w4(32'hbbeb0b6c),
	.w5(32'h3b70a042),
	.w6(32'hbbe6c4f0),
	.w7(32'hbb2c2742),
	.w8(32'h3b762e24),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8f37b),
	.w1(32'hbbc74ed3),
	.w2(32'hbb87ea5c),
	.w3(32'h3afbdc17),
	.w4(32'hba0fd041),
	.w5(32'h3b818b71),
	.w6(32'hbb6bd36b),
	.w7(32'h38029aa3),
	.w8(32'hbb1b046d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658dc4),
	.w1(32'h3ac2a0bf),
	.w2(32'h3ac32d4f),
	.w3(32'h396c7a3e),
	.w4(32'hba43d030),
	.w5(32'hbb0a5edf),
	.w6(32'hbb7a8a65),
	.w7(32'hbb97b53f),
	.w8(32'hbbc1f5a4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280417),
	.w1(32'hbb25b4f2),
	.w2(32'h3b783bdf),
	.w3(32'h3b945e5f),
	.w4(32'h3be415f3),
	.w5(32'hbae09701),
	.w6(32'hbb3cf388),
	.w7(32'h3c26f26d),
	.w8(32'hbba0325e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba091293),
	.w1(32'h3af6d1f1),
	.w2(32'h3ab5c922),
	.w3(32'hbb4e5ad8),
	.w4(32'hbb632a26),
	.w5(32'h3a569feb),
	.w6(32'hbb90ecbd),
	.w7(32'hbb68ff68),
	.w8(32'hba1a3861),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035257),
	.w1(32'hbc338e9b),
	.w2(32'h370df2d8),
	.w3(32'h3b0fcd52),
	.w4(32'h3c20a2de),
	.w5(32'hbb0b945a),
	.w6(32'h3c25c6f0),
	.w7(32'h3c33c6fc),
	.w8(32'h3b5fc31e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd596d),
	.w1(32'hbb44c369),
	.w2(32'hbb8d4ea1),
	.w3(32'h3bde4fb6),
	.w4(32'h3b6a0850),
	.w5(32'hba7bcd32),
	.w6(32'h3c07ee97),
	.w7(32'h3b709268),
	.w8(32'hbafa1484),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85058),
	.w1(32'hba7f34c4),
	.w2(32'hb90508ad),
	.w3(32'h3aa3ddc1),
	.w4(32'h39644e32),
	.w5(32'h3b4c4ac6),
	.w6(32'h37c89f7e),
	.w7(32'hb984c2cf),
	.w8(32'h3b3b7f9f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5500b),
	.w1(32'hbb9d6c06),
	.w2(32'hbbe5a480),
	.w3(32'h3ad75541),
	.w4(32'hbaf3e72b),
	.w5(32'h3b167ddd),
	.w6(32'hbb190852),
	.w7(32'hbc0d321a),
	.w8(32'h3972e28d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c57811),
	.w1(32'hbaf09bde),
	.w2(32'h39b746eb),
	.w3(32'hba43d8bb),
	.w4(32'h3a2c9d9e),
	.w5(32'hbc073795),
	.w6(32'hbbb9d127),
	.w7(32'hbb06e0f7),
	.w8(32'hbbd07ce2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806305c),
	.w1(32'h3c2125a5),
	.w2(32'hbba60a6d),
	.w3(32'h3c2f0b0a),
	.w4(32'h3b3b03a2),
	.w5(32'hbb8d04a0),
	.w6(32'h3b40209b),
	.w7(32'h3b42766e),
	.w8(32'hba84f988),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc480),
	.w1(32'hbb46b4b4),
	.w2(32'hbb49715f),
	.w3(32'hbb6a7b62),
	.w4(32'hbbd032b0),
	.w5(32'hbabbf752),
	.w6(32'h3a4f6f01),
	.w7(32'hbad61fd6),
	.w8(32'hba2cfce7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59a8c5),
	.w1(32'h3c15d017),
	.w2(32'h3c077a8c),
	.w3(32'h3c845eca),
	.w4(32'h3c34aa37),
	.w5(32'hbb61742b),
	.w6(32'h3ca3adb9),
	.w7(32'h3c80c754),
	.w8(32'h3b11b9ae),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac30ac1),
	.w1(32'h3a2dbd98),
	.w2(32'hbb0e8300),
	.w3(32'hbb3fd8ae),
	.w4(32'hba6dac0d),
	.w5(32'hbaef8a35),
	.w6(32'hba9a8d4a),
	.w7(32'hbb067d79),
	.w8(32'h3719413f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47718d),
	.w1(32'h3aa4d8a9),
	.w2(32'h3b3c1dcb),
	.w3(32'h395f5168),
	.w4(32'hbac2a55e),
	.w5(32'hbb5f7a69),
	.w6(32'h3bd3bafe),
	.w7(32'h3ba70c87),
	.w8(32'h3a4dc111),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f3dbb),
	.w1(32'h3ba405c0),
	.w2(32'hba1de563),
	.w3(32'h3b850d61),
	.w4(32'h3a37148f),
	.w5(32'hbb3b4da7),
	.w6(32'h3bb679b9),
	.w7(32'h3a466599),
	.w8(32'hbb50e43a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87dc90),
	.w1(32'hbb2fd83d),
	.w2(32'hbb003246),
	.w3(32'hbb6225fc),
	.w4(32'hbb1c107c),
	.w5(32'hb93adfb8),
	.w6(32'hbb900e9f),
	.w7(32'hbb30e279),
	.w8(32'h3c09f002),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d181),
	.w1(32'hbad74516),
	.w2(32'h3b033157),
	.w3(32'h3c19064b),
	.w4(32'h3a704fe4),
	.w5(32'hbbb7db3f),
	.w6(32'h3c4c7dfb),
	.w7(32'h3a7a1a9f),
	.w8(32'hbb9f2e34),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c174),
	.w1(32'hbbf2c8c8),
	.w2(32'hbb57affd),
	.w3(32'hbbbb321e),
	.w4(32'hb88ad1b6),
	.w5(32'hbbd9eda0),
	.w6(32'hbc27edeb),
	.w7(32'hbacca923),
	.w8(32'hbbd0048c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc82e22),
	.w1(32'hbb3a7c13),
	.w2(32'h3c147ec2),
	.w3(32'hbc0aa549),
	.w4(32'hbb0720af),
	.w5(32'h3b7edaef),
	.w6(32'hbc06f88a),
	.w7(32'h3be1fec2),
	.w8(32'h3bee9db2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cd7da),
	.w1(32'h3b2f9cb9),
	.w2(32'h3aa10144),
	.w3(32'h3a6817e2),
	.w4(32'hba243ae1),
	.w5(32'hbb3fcb0d),
	.w6(32'h3b494d47),
	.w7(32'hb970ba30),
	.w8(32'hbb048364),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432586),
	.w1(32'hbb67b9b6),
	.w2(32'hbc17c1a1),
	.w3(32'hbc0c4049),
	.w4(32'hbc10dc76),
	.w5(32'h39ae520e),
	.w6(32'hbc12b89c),
	.w7(32'hbc550245),
	.w8(32'h39a5efaa),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32a175),
	.w1(32'h3b86392c),
	.w2(32'h3b12ca94),
	.w3(32'h3b8458eb),
	.w4(32'h3b230f3e),
	.w5(32'hbae133d5),
	.w6(32'h3bfe49d0),
	.w7(32'h3adb18ba),
	.w8(32'hbb7d4bb1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb197b65),
	.w1(32'hbb700f2a),
	.w2(32'hba86f8f1),
	.w3(32'hbb5d8285),
	.w4(32'h3b07fae6),
	.w5(32'h3aa541f6),
	.w6(32'hbbe916bf),
	.w7(32'hbb03cffd),
	.w8(32'hbb4c1a72),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964b5a8),
	.w1(32'h3bc2bd00),
	.w2(32'h3c37c4e8),
	.w3(32'hbb95cc4d),
	.w4(32'hbaa229d1),
	.w5(32'h3c39db14),
	.w6(32'hbbf41f18),
	.w7(32'hb9b3885c),
	.w8(32'h3bd8fc05),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba377be),
	.w1(32'h3bb850a8),
	.w2(32'h3c69a3a2),
	.w3(32'h3cd4033d),
	.w4(32'h3cf11ebd),
	.w5(32'h3b82b909),
	.w6(32'h3cadb6f4),
	.w7(32'h3d0ffa24),
	.w8(32'h3bb83ca3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb151),
	.w1(32'h3b9cdeb5),
	.w2(32'hba17eff9),
	.w3(32'hbb0e9c8f),
	.w4(32'hbad7b978),
	.w5(32'h3be51436),
	.w6(32'hba019b96),
	.w7(32'hbb38fc75),
	.w8(32'h3c1c4f84),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4acf8),
	.w1(32'h3bdc2b7e),
	.w2(32'h3b73369b),
	.w3(32'h3c23d7b7),
	.w4(32'h3b77d228),
	.w5(32'h3c9278fe),
	.w6(32'h3ca15aa9),
	.w7(32'h3c286a50),
	.w8(32'h3cd03de8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af07776),
	.w1(32'h3a99dde4),
	.w2(32'hbadd9df8),
	.w3(32'h3c4e766a),
	.w4(32'hbac2cb89),
	.w5(32'hbaa89e2e),
	.w6(32'h3c9778ae),
	.w7(32'h3b35d99c),
	.w8(32'h3ab8bbcc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c8aaf),
	.w1(32'hbb927cf2),
	.w2(32'hbb690367),
	.w3(32'hbb832434),
	.w4(32'h3b1a0f82),
	.w5(32'hbb17d9a4),
	.w6(32'hbaef84bf),
	.w7(32'h3badec2b),
	.w8(32'h3be93abe),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0591f),
	.w1(32'h3c8f4cfc),
	.w2(32'h3c7b449f),
	.w3(32'hbb187a41),
	.w4(32'hbbd2c839),
	.w5(32'h38616db8),
	.w6(32'h3b23ba1c),
	.w7(32'h3a261b95),
	.w8(32'hb9af0162),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5acaa3),
	.w1(32'h3a8e78e4),
	.w2(32'h3b4a610d),
	.w3(32'hbb9da762),
	.w4(32'hbb69ccfa),
	.w5(32'hbaf87034),
	.w6(32'hbb45816d),
	.w7(32'hbb0df0f2),
	.w8(32'hbb80b8d2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89dd34),
	.w1(32'hbb1a2444),
	.w2(32'h3bab360f),
	.w3(32'hba403319),
	.w4(32'h3be9e520),
	.w5(32'hbb41cfdd),
	.w6(32'hbbc366f7),
	.w7(32'h3b1d03c6),
	.w8(32'hbb7158dc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5db16),
	.w1(32'h3ac54b0a),
	.w2(32'h3b7f190e),
	.w3(32'hbaeb0c3b),
	.w4(32'hba0ddf17),
	.w5(32'hbc149e5d),
	.w6(32'h3a776bcd),
	.w7(32'h3a6bfcda),
	.w8(32'hbbf9b3f0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa98db),
	.w1(32'hbc172187),
	.w2(32'h3aa5fab7),
	.w3(32'hbb16cd37),
	.w4(32'h3c26c8e2),
	.w5(32'hb7d757ad),
	.w6(32'hbc33a37b),
	.w7(32'h3c43e838),
	.w8(32'h3ae62f0b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f05bec),
	.w1(32'hbba66e45),
	.w2(32'hba97065e),
	.w3(32'hbb80c7f4),
	.w4(32'hbabf9182),
	.w5(32'hbc2ac989),
	.w6(32'hbb75a478),
	.w7(32'h3b28eb96),
	.w8(32'hba1bb795),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aceb0),
	.w1(32'h3c2cfecb),
	.w2(32'h3bc5b8a7),
	.w3(32'hbba575b9),
	.w4(32'hbb57678d),
	.w5(32'h3bc15d8c),
	.w6(32'h3be07870),
	.w7(32'h3bae3682),
	.w8(32'hba1d6e42),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139274),
	.w1(32'hbc29bad3),
	.w2(32'hbb9f038d),
	.w3(32'h3c10bc64),
	.w4(32'h3bb0dbc5),
	.w5(32'h3ab2329b),
	.w6(32'h3ba23b38),
	.w7(32'hbb25cf65),
	.w8(32'hbb806b99),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e43ea),
	.w1(32'h3c088377),
	.w2(32'h3c6dcd38),
	.w3(32'hbb16043d),
	.w4(32'h3bc255c0),
	.w5(32'hbb94faaa),
	.w6(32'h3bb9745d),
	.w7(32'h3c7fcdf3),
	.w8(32'hbb3bf277),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5dd11),
	.w1(32'hbb9dc822),
	.w2(32'hbbafc003),
	.w3(32'hbc1ee882),
	.w4(32'hbba43496),
	.w5(32'h3b8dbabf),
	.w6(32'hbc222878),
	.w7(32'hbc1f74fc),
	.w8(32'h3ca27979),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d19eefa),
	.w1(32'h3cd60aa6),
	.w2(32'h3c8201cc),
	.w3(32'h3bcc6c4f),
	.w4(32'h3b16f6e2),
	.w5(32'h3c08ff57),
	.w6(32'h3c82d74b),
	.w7(32'h3bd94e0a),
	.w8(32'h3c3a3fe3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eccae),
	.w1(32'hba76dc2b),
	.w2(32'h3b8a2c7f),
	.w3(32'h3bb7a7ab),
	.w4(32'hba261bb2),
	.w5(32'h393288a1),
	.w6(32'h3bad40c6),
	.w7(32'h3a4d6a8b),
	.w8(32'h3c2daf74),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53110),
	.w1(32'h3c529f72),
	.w2(32'hbac7b72a),
	.w3(32'hbbb1adbd),
	.w4(32'h3898f1f5),
	.w5(32'hbc1fb7c8),
	.w6(32'h3b7e97aa),
	.w7(32'h3ae48f8f),
	.w8(32'hbbd7df06),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a957),
	.w1(32'hbb4b2915),
	.w2(32'hba70aacc),
	.w3(32'hbbaa05c5),
	.w4(32'hba34bf4e),
	.w5(32'h39ec5b50),
	.w6(32'hbbedde26),
	.w7(32'hbb863b66),
	.w8(32'hbbb5f220),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5b13a),
	.w1(32'hbb8c8838),
	.w2(32'hbb967e8a),
	.w3(32'h3b321e34),
	.w4(32'h3b2739d1),
	.w5(32'hbb143faf),
	.w6(32'hbb7f58dc),
	.w7(32'hbb14c8cd),
	.w8(32'hba3652ba),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0d190),
	.w1(32'hbbdc8ff7),
	.w2(32'hbc019898),
	.w3(32'hbb0652e4),
	.w4(32'hbc53d6ab),
	.w5(32'h3b526f69),
	.w6(32'h3b05b3b1),
	.w7(32'hbc0ab5aa),
	.w8(32'h3b683f6a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a3f9),
	.w1(32'hbb5a5fbb),
	.w2(32'h3b76b4ce),
	.w3(32'h3b110980),
	.w4(32'hbb0b771f),
	.w5(32'hbc0129ce),
	.w6(32'h3bf069c2),
	.w7(32'h3b8c3ca5),
	.w8(32'hbb3d9fd5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4e565),
	.w1(32'hbb862fa1),
	.w2(32'hbae2f31e),
	.w3(32'hbb912b54),
	.w4(32'hbabe2225),
	.w5(32'hbaeff92f),
	.w6(32'hbbf0dbd6),
	.w7(32'hbb92eb36),
	.w8(32'hbb8e4cd3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20b306),
	.w1(32'h3af7289f),
	.w2(32'h3c7ebfd2),
	.w3(32'hb9638dae),
	.w4(32'h3bd799b9),
	.w5(32'hbb7a1fef),
	.w6(32'hbc38c3f8),
	.w7(32'h3b5943a3),
	.w8(32'hbba46c71),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb033fab),
	.w1(32'hbaa0adb7),
	.w2(32'h3c295535),
	.w3(32'hb9d95180),
	.w4(32'h3ac30c20),
	.w5(32'hbb6fb4c4),
	.w6(32'hbc13cbd6),
	.w7(32'hba56288d),
	.w8(32'hbbf701a3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba339ac6),
	.w1(32'hbc5732f8),
	.w2(32'hbc11681d),
	.w3(32'hbb42b099),
	.w4(32'hbbf8ae14),
	.w5(32'h3b7c5149),
	.w6(32'hbbb9661c),
	.w7(32'hbc27703a),
	.w8(32'h3b10bb59),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fed04),
	.w1(32'h3bc1cce7),
	.w2(32'h3b8a4d47),
	.w3(32'h3a8e98c1),
	.w4(32'h3badba8d),
	.w5(32'h3b5870a3),
	.w6(32'h3b910c4d),
	.w7(32'h3b963e8a),
	.w8(32'h3b18ec5d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b518bae),
	.w1(32'hbbcb33f1),
	.w2(32'hbb7e8cca),
	.w3(32'h3ade4892),
	.w4(32'h392d003f),
	.w5(32'h3a04854b),
	.w6(32'h3adc1089),
	.w7(32'h3a2e17d5),
	.w8(32'h3c1e8777),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b77f),
	.w1(32'h3c05e376),
	.w2(32'h3ba29868),
	.w3(32'h3bd74270),
	.w4(32'h3b998794),
	.w5(32'hbbc3b8f5),
	.w6(32'h3c5534f2),
	.w7(32'h3be6b2ab),
	.w8(32'hbc0796b2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7274a5),
	.w1(32'hbbc3c6b3),
	.w2(32'hbb87183c),
	.w3(32'hbbd00981),
	.w4(32'hbaa32527),
	.w5(32'h3b4e9687),
	.w6(32'hbc035bbb),
	.w7(32'hbb75bf61),
	.w8(32'h3bf40d88),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0005f2),
	.w1(32'h3c04d6bf),
	.w2(32'h3b6cd73e),
	.w3(32'h3bd66a30),
	.w4(32'h3adf1fb7),
	.w5(32'h3b326267),
	.w6(32'h3c4bbbb9),
	.w7(32'h3b7d6ed9),
	.w8(32'hbb04e813),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2620),
	.w1(32'h3c4bd0fd),
	.w2(32'h3cab9843),
	.w3(32'h3bdbc05b),
	.w4(32'h3c3b887e),
	.w5(32'hbbda1b89),
	.w6(32'h3b4b55ac),
	.w7(32'h3cdb6bce),
	.w8(32'hbb8ec238),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa57af6),
	.w1(32'h3ac29860),
	.w2(32'h3b238b6c),
	.w3(32'h3a7afde3),
	.w4(32'h3bbb26cf),
	.w5(32'hbbba995d),
	.w6(32'hbb6d0878),
	.w7(32'h3b6bdd0c),
	.w8(32'hbc36a142),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26253),
	.w1(32'hbb3837f4),
	.w2(32'h3c64e23f),
	.w3(32'hbbdb57c6),
	.w4(32'h3a15c600),
	.w5(32'h3b7d6b6c),
	.w6(32'hbc0da365),
	.w7(32'h3bd17f3e),
	.w8(32'h3c4002c7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9b8c),
	.w1(32'h3c76d10c),
	.w2(32'h3ab625d2),
	.w3(32'h3c3dc4c1),
	.w4(32'h3a98c7d8),
	.w5(32'h3a297bdf),
	.w6(32'h3c46345f),
	.w7(32'h3958c1fa),
	.w8(32'h3a190040),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdced0c),
	.w1(32'h3b516b97),
	.w2(32'h3b6d231b),
	.w3(32'hba24fbc2),
	.w4(32'h3bb0b7fa),
	.w5(32'hbbe2e76c),
	.w6(32'hbb37ebd9),
	.w7(32'h3b893531),
	.w8(32'hbba38c10),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35ab99),
	.w1(32'h39d1146d),
	.w2(32'hbb0e9252),
	.w3(32'hba975c63),
	.w4(32'h3af8c7c6),
	.w5(32'hba815ddd),
	.w6(32'hbb057e71),
	.w7(32'hbb05a5d6),
	.w8(32'h3b925317),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb6919),
	.w1(32'h3c12b044),
	.w2(32'h3bc004e5),
	.w3(32'hbb46f8c5),
	.w4(32'h39a5e30b),
	.w5(32'h3b6e0dc0),
	.w6(32'h3a6dec98),
	.w7(32'h3b4e8da1),
	.w8(32'h3c265872),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ef46),
	.w1(32'hb9f90d3e),
	.w2(32'hbb6f14a0),
	.w3(32'hbadc57e1),
	.w4(32'hbb6d7696),
	.w5(32'hbb4eb0be),
	.w6(32'hb99f0518),
	.w7(32'hba3d803e),
	.w8(32'h3a3f9c8b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b6b1c),
	.w1(32'h3bd696d5),
	.w2(32'h3b2fead7),
	.w3(32'h3c02e3e6),
	.w4(32'h3a81921a),
	.w5(32'hbbe2d7ad),
	.w6(32'h3c31d550),
	.w7(32'h3b4cf7fa),
	.w8(32'hbb61dad3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34c899),
	.w1(32'hbba2e600),
	.w2(32'hbc26fd96),
	.w3(32'h3bf1fb44),
	.w4(32'h3a802eb8),
	.w5(32'hbba1ee16),
	.w6(32'h3bd1b0fe),
	.w7(32'hbbb28c5e),
	.w8(32'hbb72cfd6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb576c0c),
	.w1(32'hbbcab811),
	.w2(32'hbaa97082),
	.w3(32'hbbbb715e),
	.w4(32'hbc23e313),
	.w5(32'h3a8a27a0),
	.w6(32'hbb582516),
	.w7(32'hbbb9e9e5),
	.w8(32'hbb0017eb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafda4f),
	.w1(32'h3b13be04),
	.w2(32'h3b4aa74a),
	.w3(32'hbb1be931),
	.w4(32'h3afbc96d),
	.w5(32'hbba4ddd4),
	.w6(32'hbb5e5249),
	.w7(32'h3b2d5239),
	.w8(32'hba0f1f3e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9401d9),
	.w1(32'h3c6dc83b),
	.w2(32'h3c549e2a),
	.w3(32'hbb595a36),
	.w4(32'hba2cb63b),
	.w5(32'hbb3024d3),
	.w6(32'hbb0d5376),
	.w7(32'h39de64b4),
	.w8(32'h3b1ee1fd),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3a248),
	.w1(32'h3b1c36bb),
	.w2(32'hbb65fb0e),
	.w3(32'hb9e5c085),
	.w4(32'hbb75dfdc),
	.w5(32'hbbf0efa8),
	.w6(32'h38acf558),
	.w7(32'hbb47c04c),
	.w8(32'hbb8d639b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7fdcd),
	.w1(32'hbc0ab9a8),
	.w2(32'hbbf15fb2),
	.w3(32'hbc7bc0f1),
	.w4(32'hbc1febbf),
	.w5(32'hbb38ab67),
	.w6(32'hbc8a69a7),
	.w7(32'hbc0bc242),
	.w8(32'hbb956296),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae17981),
	.w1(32'h3b9563aa),
	.w2(32'h3c0dfc4f),
	.w3(32'hbabdf4ae),
	.w4(32'hbb1bd61b),
	.w5(32'hba1be3a7),
	.w6(32'hbb9c24a7),
	.w7(32'hbb85dd0e),
	.w8(32'h3aaef153),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398a54),
	.w1(32'h3b3e9115),
	.w2(32'hbaa37e6b),
	.w3(32'hba1f6821),
	.w4(32'hbb778294),
	.w5(32'hbc101dad),
	.w6(32'h39a2f235),
	.w7(32'hbb0a4bc1),
	.w8(32'hbb70fc04),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3035a5),
	.w1(32'hba38e64d),
	.w2(32'h3bdcde55),
	.w3(32'hbb768815),
	.w4(32'h3bf5f8c1),
	.w5(32'h3a38e47c),
	.w6(32'hbb95f6cf),
	.w7(32'h3bffb4c5),
	.w8(32'hbad7115d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a4dd),
	.w1(32'hbc127e30),
	.w2(32'h3b14eb2c),
	.w3(32'hbbfc3b14),
	.w4(32'hbb52ac2a),
	.w5(32'hba3122dc),
	.w6(32'hbc4ded02),
	.w7(32'h3bb7b3fe),
	.w8(32'h3aa9a16c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a922ce4),
	.w1(32'hbb486fd6),
	.w2(32'h3be103f3),
	.w3(32'h3bace70d),
	.w4(32'h3bbe4da0),
	.w5(32'h3b898ddb),
	.w6(32'h3add752f),
	.w7(32'h3b27f789),
	.w8(32'h3c2979cf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed2c8),
	.w1(32'h3be0dd10),
	.w2(32'h3bf3488e),
	.w3(32'h3b0a265e),
	.w4(32'h3c038a45),
	.w5(32'h3a974a65),
	.w6(32'h3b08ed8d),
	.w7(32'h3bb17433),
	.w8(32'h3b062788),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19b21),
	.w1(32'h3a68db06),
	.w2(32'hbb74ef40),
	.w3(32'h3a82db5e),
	.w4(32'hbb8ad569),
	.w5(32'hbb905804),
	.w6(32'hbab616d6),
	.w7(32'hbb723e6b),
	.w8(32'h3a8ed654),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31c7e),
	.w1(32'hbb502309),
	.w2(32'hbbb5dc47),
	.w3(32'h3af0478b),
	.w4(32'h3ba11270),
	.w5(32'hbbbdc0f3),
	.w6(32'h3b22d5bf),
	.w7(32'h3b57ecc2),
	.w8(32'hbb2c9b2a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f1f44),
	.w1(32'hbb575235),
	.w2(32'hbc018310),
	.w3(32'hbba8973d),
	.w4(32'hbbd07331),
	.w5(32'h3a883b59),
	.w6(32'hbb9cc41b),
	.w7(32'hbbcadf82),
	.w8(32'h3a3604ef),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394539d3),
	.w1(32'hbae75377),
	.w2(32'hbaee583d),
	.w3(32'h3bbc1622),
	.w4(32'hbaaa0d08),
	.w5(32'hbb049590),
	.w6(32'h3afc1c61),
	.w7(32'hbac458f9),
	.w8(32'h39b9b32a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b817),
	.w1(32'hbb93e7c2),
	.w2(32'hbaf5ecfc),
	.w3(32'hbbb43aca),
	.w4(32'hbb6daffa),
	.w5(32'h3bf1ed82),
	.w6(32'hbc13f061),
	.w7(32'hbab9ad33),
	.w8(32'h3c2758ce),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8590c9),
	.w1(32'h3bbd8034),
	.w2(32'h3bf7078b),
	.w3(32'h3b8effa1),
	.w4(32'hbba1fb6a),
	.w5(32'h3b2c6bbe),
	.w6(32'h3be1f92c),
	.w7(32'h39d6ea84),
	.w8(32'h3badf53f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d6dd9),
	.w1(32'hbaf12168),
	.w2(32'h3a20cfe9),
	.w3(32'h397a582e),
	.w4(32'h3b59b398),
	.w5(32'h3bb12fed),
	.w6(32'hbb148d4e),
	.w7(32'h3b002a33),
	.w8(32'h3bc3c58e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeac35),
	.w1(32'h3b748b7f),
	.w2(32'h3b86b979),
	.w3(32'h3a454106),
	.w4(32'h3ab0e77f),
	.w5(32'h39bbb174),
	.w6(32'h3b8856a9),
	.w7(32'h3b932760),
	.w8(32'h3b52db03),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f2200),
	.w1(32'h3b5b6495),
	.w2(32'hb9a3a3c3),
	.w3(32'hbad62745),
	.w4(32'hbb3064dd),
	.w5(32'h3b6e50a5),
	.w6(32'h3b84c41f),
	.w7(32'hba2c5dd3),
	.w8(32'h3bbc88f6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35cc9e),
	.w1(32'h3ac3dd67),
	.w2(32'h3a240081),
	.w3(32'h3c2a4025),
	.w4(32'h3b938294),
	.w5(32'hbb81c314),
	.w6(32'h3b41c8e1),
	.w7(32'h3b876da3),
	.w8(32'h3a1117f7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a739),
	.w1(32'hbafd7ec0),
	.w2(32'hb9b679de),
	.w3(32'hbb881154),
	.w4(32'hbafab12e),
	.w5(32'hbb554d01),
	.w6(32'hbbb0c801),
	.w7(32'hbb5ea89f),
	.w8(32'hbbba6f54),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139d22),
	.w1(32'hbc554aea),
	.w2(32'hbc22c061),
	.w3(32'hbc2acfb9),
	.w4(32'hbc33acc5),
	.w5(32'h3929054e),
	.w6(32'hbc5fc467),
	.w7(32'hbc264015),
	.w8(32'hbb1c03ad),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21c020),
	.w1(32'hbc18eb72),
	.w2(32'hbbc56f5c),
	.w3(32'hbbd6a12e),
	.w4(32'h3ab7f3c3),
	.w5(32'h3bbb1c5e),
	.w6(32'hbc39c5b0),
	.w7(32'hbafb202d),
	.w8(32'h3b99910e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a041134),
	.w1(32'hb90ef6a4),
	.w2(32'hbb8d5daa),
	.w3(32'h3be6d730),
	.w4(32'h390573e7),
	.w5(32'h3ad1207f),
	.w6(32'h3c2f5955),
	.w7(32'h3b87069a),
	.w8(32'h3ac2d87a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e53d3),
	.w1(32'hbab05626),
	.w2(32'h3a2fcc21),
	.w3(32'hbad6b538),
	.w4(32'h3a63d7f6),
	.w5(32'h3c2738fd),
	.w6(32'hbb9fe37a),
	.w7(32'h39355d46),
	.w8(32'h3c838f5c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c214d),
	.w1(32'h3c38e0c1),
	.w2(32'h3b9e8165),
	.w3(32'h3c099b54),
	.w4(32'h3c0034ea),
	.w5(32'hbbcd7fd5),
	.w6(32'h3c49d9af),
	.w7(32'h3c0a73bb),
	.w8(32'hbbd687a9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08b6d6),
	.w1(32'hb937babe),
	.w2(32'h3aad8177),
	.w3(32'h3bfcbf30),
	.w4(32'h3bd400ef),
	.w5(32'hbb82ccb0),
	.w6(32'hb9c62d8b),
	.w7(32'h3ba4dc2d),
	.w8(32'hbb62dde4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ddfb0),
	.w1(32'h3ba70439),
	.w2(32'h3babd987),
	.w3(32'h3b398bec),
	.w4(32'h3adf8d49),
	.w5(32'hbb8fe0f4),
	.w6(32'h3bec2aba),
	.w7(32'h3b782ed0),
	.w8(32'hbb7cbe3f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3d56e),
	.w1(32'hbb8dd2d5),
	.w2(32'h3b003135),
	.w3(32'hbbb96b22),
	.w4(32'hbb1bfa63),
	.w5(32'h3abc647d),
	.w6(32'hbbf15bfc),
	.w7(32'hb99e0b52),
	.w8(32'h3aae90ad),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1da539),
	.w1(32'h3b3851d7),
	.w2(32'hbb2d1d5e),
	.w3(32'h3c56db44),
	.w4(32'h3b04d1fb),
	.w5(32'hbb42959a),
	.w6(32'h3c038cc8),
	.w7(32'h3a95a573),
	.w8(32'hbbd7abd5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bcee8),
	.w1(32'hbaeea0eb),
	.w2(32'h3b6fe598),
	.w3(32'h3b4a9fc0),
	.w4(32'h3bbf0cea),
	.w5(32'hbadcbfa0),
	.w6(32'h3a771806),
	.w7(32'h3c8508ab),
	.w8(32'hbbdba8f7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc298195),
	.w1(32'hbc05a758),
	.w2(32'h3ae85d5d),
	.w3(32'h3ba0c621),
	.w4(32'h3baf4967),
	.w5(32'hbb593acc),
	.w6(32'hb8a68c62),
	.w7(32'h3b3ffb73),
	.w8(32'hbbba6aa3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f165),
	.w1(32'hbbd8e1be),
	.w2(32'hbb60d154),
	.w3(32'hbbe8d3ed),
	.w4(32'hbc448b60),
	.w5(32'h3b002305),
	.w6(32'hbc23c910),
	.w7(32'hbc364d15),
	.w8(32'h3abe863b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cc1d3),
	.w1(32'hbb543b8c),
	.w2(32'hbb6deaf8),
	.w3(32'hbb50f307),
	.w4(32'hbacc1451),
	.w5(32'hbaf51950),
	.w6(32'hbb897998),
	.w7(32'hbb785e1d),
	.w8(32'h3afed94f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39941275),
	.w1(32'hbb3bf6f9),
	.w2(32'h3b82e1d6),
	.w3(32'h3bcfd2c4),
	.w4(32'h3c077186),
	.w5(32'h3c0a8174),
	.w6(32'hbadde6c3),
	.w7(32'h3b5d718d),
	.w8(32'h3c285aba),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9df00d),
	.w1(32'h3b281040),
	.w2(32'hbb32d36b),
	.w3(32'h3bd0f308),
	.w4(32'h39d11692),
	.w5(32'hbc264bcf),
	.w6(32'h3c2975dd),
	.w7(32'h3bad5d79),
	.w8(32'hbc2833ce),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacc564),
	.w1(32'h3b828276),
	.w2(32'h3bc24759),
	.w3(32'hbb72ecf8),
	.w4(32'h3a186e7e),
	.w5(32'h3ba99bcc),
	.w6(32'h3b9b1753),
	.w7(32'h3bc002d9),
	.w8(32'h3ba6cd2d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822ff8),
	.w1(32'h3b46c705),
	.w2(32'h3b1b6a17),
	.w3(32'h39e526a2),
	.w4(32'hba4f8ef1),
	.w5(32'h3ba9601a),
	.w6(32'h3ac71d73),
	.w7(32'hba598934),
	.w8(32'h3a85ce14),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9af51a),
	.w1(32'hba5ba326),
	.w2(32'hb8db584c),
	.w3(32'h3bd629ff),
	.w4(32'h3bc45ae5),
	.w5(32'h3a66d7eb),
	.w6(32'h3be21d54),
	.w7(32'h3b899f65),
	.w8(32'h3be88c12),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b5474),
	.w1(32'hb9cbfced),
	.w2(32'h3b155d37),
	.w3(32'hbb0c3574),
	.w4(32'hba4171ec),
	.w5(32'h3b4aa664),
	.w6(32'h3b4223a0),
	.w7(32'h3ac9d0d2),
	.w8(32'h3ba9bbb1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ea462),
	.w1(32'hbb0ee5aa),
	.w2(32'hba5eb10b),
	.w3(32'h3b2136e1),
	.w4(32'h39d931d3),
	.w5(32'hba5eba80),
	.w6(32'hbab0b48e),
	.w7(32'hbb82ebec),
	.w8(32'hba17fda5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3da1d8),
	.w1(32'h3b8b687d),
	.w2(32'h3b1c5bea),
	.w3(32'h3c152036),
	.w4(32'h3c346102),
	.w5(32'hbbb3d818),
	.w6(32'h3c0f2239),
	.w7(32'h3c1915e6),
	.w8(32'h3a4532e7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa6b4),
	.w1(32'hbb67680d),
	.w2(32'hbc02d1bf),
	.w3(32'h392d41f0),
	.w4(32'hbb1d8342),
	.w5(32'hbbc8746b),
	.w6(32'h389c7a6d),
	.w7(32'hbabfaa9b),
	.w8(32'hbb835446),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ec23),
	.w1(32'hbb828b00),
	.w2(32'hba4cf576),
	.w3(32'hbba0bf67),
	.w4(32'hbb8028a4),
	.w5(32'h3b16427f),
	.w6(32'hbbecd66d),
	.w7(32'hbb868332),
	.w8(32'h3af8cae1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7e5e5),
	.w1(32'h3ba36358),
	.w2(32'h3acd5c4c),
	.w3(32'h3bb4a59f),
	.w4(32'h39a6da53),
	.w5(32'hbb9a7b7e),
	.w6(32'h3bd37834),
	.w7(32'h3a32f667),
	.w8(32'hbb75161c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2962bd),
	.w1(32'h39a4b2e0),
	.w2(32'h3abfcbfa),
	.w3(32'hba727dd6),
	.w4(32'h3b82d9c4),
	.w5(32'hba55eef9),
	.w6(32'h3ab30f3e),
	.w7(32'h3b0320b0),
	.w8(32'hba4dfd57),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54093e),
	.w1(32'hbaafa931),
	.w2(32'hb9f83c18),
	.w3(32'hb99baad0),
	.w4(32'h398c6452),
	.w5(32'h3b1781a0),
	.w6(32'h3af74762),
	.w7(32'h3b423433),
	.w8(32'h3b0e1b05),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7b1b8),
	.w1(32'h3b122467),
	.w2(32'hbb864e45),
	.w3(32'h3ad10c42),
	.w4(32'hbb9711cd),
	.w5(32'h395c6ed1),
	.w6(32'h3a8b4182),
	.w7(32'hbbad6f42),
	.w8(32'h3b3dd863),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02196c),
	.w1(32'h3b6c20a9),
	.w2(32'h3b0894f0),
	.w3(32'h3b022127),
	.w4(32'hb9b9e0bd),
	.w5(32'h3aad0da8),
	.w6(32'h3bb6f280),
	.w7(32'h3b4f46cb),
	.w8(32'h3a6e89a7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8324d8),
	.w1(32'hba763543),
	.w2(32'hbb4067f3),
	.w3(32'hba10645a),
	.w4(32'h3b4a1400),
	.w5(32'hbafaf230),
	.w6(32'h3ab61c64),
	.w7(32'hba8c7bca),
	.w8(32'hbb04a4e9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7046b),
	.w1(32'hbb1bbdaf),
	.w2(32'hbaaeb136),
	.w3(32'h3b8b09a1),
	.w4(32'hb97eece7),
	.w5(32'h3c08fc49),
	.w6(32'h3c2add74),
	.w7(32'h3b8c6713),
	.w8(32'h3c2ad8e0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62ebb5),
	.w1(32'h3bbcbc77),
	.w2(32'h3bd49737),
	.w3(32'h3bf788dc),
	.w4(32'h3bca1ef8),
	.w5(32'h3ab5a240),
	.w6(32'h3b9b59a1),
	.w7(32'h3b932dc7),
	.w8(32'h3af4f7bc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a1937),
	.w1(32'hbb335cd6),
	.w2(32'hbb6ce725),
	.w3(32'h3b251334),
	.w4(32'hbb661abc),
	.w5(32'hbb806911),
	.w6(32'h3ba0bc20),
	.w7(32'hba870494),
	.w8(32'h3ab41fd4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b537cd1),
	.w1(32'h3ba390da),
	.w2(32'h3bc7effa),
	.w3(32'hbb68617a),
	.w4(32'hbb88f395),
	.w5(32'h3983bcbd),
	.w6(32'hba7f03fe),
	.w7(32'hbaf1110e),
	.w8(32'hb9aacd05),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbba5b),
	.w1(32'h3a54b332),
	.w2(32'h39b16128),
	.w3(32'h3b586455),
	.w4(32'h3b1e967c),
	.w5(32'hba601697),
	.w6(32'h3ae287db),
	.w7(32'h39fbbac0),
	.w8(32'hbaacb9e7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e45e8),
	.w1(32'h3addc4f8),
	.w2(32'hba78250b),
	.w3(32'h3a1db45a),
	.w4(32'hba330bf7),
	.w5(32'h39be076c),
	.w6(32'hbafd7b67),
	.w7(32'hbb0f2675),
	.w8(32'hbb614178),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a477a),
	.w1(32'hba88e9f0),
	.w2(32'h3b05f489),
	.w3(32'h39aa9d7d),
	.w4(32'h3925d808),
	.w5(32'h3b82ad0d),
	.w6(32'hbb5c819e),
	.w7(32'hb987f83d),
	.w8(32'h3adadb15),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b46d),
	.w1(32'hb968c0cb),
	.w2(32'h3918ab68),
	.w3(32'h3b52befb),
	.w4(32'hb91dd977),
	.w5(32'hbbd4a554),
	.w6(32'h3a94a329),
	.w7(32'hb9cf01c4),
	.w8(32'hbb526457),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32207),
	.w1(32'hbb20a827),
	.w2(32'hbbb4cdea),
	.w3(32'hbb9134d2),
	.w4(32'hbbe64f9e),
	.w5(32'hbb89b79f),
	.w6(32'hbb8584f2),
	.w7(32'hbc1560ff),
	.w8(32'hbb2b3baa),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00817f),
	.w1(32'h3b35ef1d),
	.w2(32'hba68150a),
	.w3(32'h39dab2dc),
	.w4(32'h38d2bcd9),
	.w5(32'h3ac20665),
	.w6(32'h3a3446d4),
	.w7(32'h3acff5d3),
	.w8(32'h3b1e3c0d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3601c),
	.w1(32'h3bec9579),
	.w2(32'h3c414201),
	.w3(32'h3ba704f3),
	.w4(32'h3c24033c),
	.w5(32'h3c0ce6ee),
	.w6(32'h3b8ea866),
	.w7(32'h3c261a87),
	.w8(32'h3a7f7cd9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61c6cb),
	.w1(32'h3b2805e8),
	.w2(32'h3bd45168),
	.w3(32'h3c12a577),
	.w4(32'h3bf5c577),
	.w5(32'h3acd8831),
	.w6(32'h3b9c3f33),
	.w7(32'h3b05659e),
	.w8(32'h3b2aba9c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71fd9),
	.w1(32'h3c025af9),
	.w2(32'h3c32e5e0),
	.w3(32'hba10865d),
	.w4(32'h3a2b4a51),
	.w5(32'h3c1db6bc),
	.w6(32'h3acf705d),
	.w7(32'h3ba599ca),
	.w8(32'h3c1f9271),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b35ed),
	.w1(32'h3b113a64),
	.w2(32'h3b6817fa),
	.w3(32'h3bc53734),
	.w4(32'h3c2ad0b8),
	.w5(32'hbb12a168),
	.w6(32'h3c156cfc),
	.w7(32'h3bcbb27d),
	.w8(32'hbb7149b1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dfdc6),
	.w1(32'h3a9a68f1),
	.w2(32'h3aa66ed0),
	.w3(32'h3bed08d0),
	.w4(32'hbbc1901f),
	.w5(32'hbb37e18b),
	.w6(32'h3c5cb899),
	.w7(32'h3b8bd44d),
	.w8(32'hbb0b9ae6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fdeea),
	.w1(32'h3b1f89bf),
	.w2(32'h3b711897),
	.w3(32'hba9c3a4e),
	.w4(32'hbb26674b),
	.w5(32'hbb18f196),
	.w6(32'h3b660d97),
	.w7(32'h3b259956),
	.w8(32'hba85deac),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f483f),
	.w1(32'h3abb1b2d),
	.w2(32'hbacfcabe),
	.w3(32'h3b1f8548),
	.w4(32'hbaeae31d),
	.w5(32'h3c5c2d7c),
	.w6(32'hb92a6344),
	.w7(32'hbb701f3e),
	.w8(32'h3c81843e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule