module layer_8_featuremap_222(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2796fe),
	.w1(32'hbc08fc02),
	.w2(32'hbc3538df),
	.w3(32'h3c693636),
	.w4(32'hbb2de03d),
	.w5(32'hbc0ef3b4),
	.w6(32'h3a6e6209),
	.w7(32'hbb0d21f5),
	.w8(32'hbba034dd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28c1a6),
	.w1(32'h3b6ec060),
	.w2(32'h3ac257cf),
	.w3(32'hbc71dfd9),
	.w4(32'h39e786b3),
	.w5(32'hbb14fae1),
	.w6(32'h3b6fb0f8),
	.w7(32'h3abbde74),
	.w8(32'hbaa1b26a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800413),
	.w1(32'h3b40ac1f),
	.w2(32'hbb077722),
	.w3(32'hbbccaeab),
	.w4(32'hbb2116cd),
	.w5(32'h3ab0ac5f),
	.w6(32'hba178f70),
	.w7(32'h3a98be6f),
	.w8(32'h3b81de12),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ac1a8),
	.w1(32'hba9d379c),
	.w2(32'hbb6af32e),
	.w3(32'h3ba2258d),
	.w4(32'h3b5e442f),
	.w5(32'hbb304a61),
	.w6(32'hbbe1f886),
	.w7(32'hbc103e50),
	.w8(32'hbbdc98ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109db4),
	.w1(32'h38980e42),
	.w2(32'hbaaa5db8),
	.w3(32'hbbbebc91),
	.w4(32'h3a885562),
	.w5(32'hbb4d9f1a),
	.w6(32'h3a12c0da),
	.w7(32'h39bb0e2a),
	.w8(32'hbb1e2640),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9046ac),
	.w1(32'hbb934344),
	.w2(32'hbbe617ae),
	.w3(32'hbc0c9406),
	.w4(32'hbbeaa065),
	.w5(32'hbc3b4fcc),
	.w6(32'hbb3b7337),
	.w7(32'hbc23a18b),
	.w8(32'hbbf8b2fe),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f101),
	.w1(32'hbb441565),
	.w2(32'hbaf143bf),
	.w3(32'h3a77e12c),
	.w4(32'h3a693e59),
	.w5(32'h3ab969ef),
	.w6(32'hbb4cc425),
	.w7(32'hbb331347),
	.w8(32'hba2a7b0c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0709a0),
	.w1(32'h3b5b32ac),
	.w2(32'hbaf980c0),
	.w3(32'h3af09928),
	.w4(32'h3acb856b),
	.w5(32'h3aba25f6),
	.w6(32'h3ba29668),
	.w7(32'h3a90fa77),
	.w8(32'h3ae1cabc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a236e),
	.w1(32'h3b31d889),
	.w2(32'hba278101),
	.w3(32'h3c0d2da5),
	.w4(32'h3b7d2f14),
	.w5(32'hbb0de32a),
	.w6(32'h3b55c219),
	.w7(32'h3ab6c4af),
	.w8(32'h3abe20a2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117eab),
	.w1(32'hbc1cb962),
	.w2(32'hbbe4237b),
	.w3(32'hbc133d42),
	.w4(32'h3b950d63),
	.w5(32'h3ae0278a),
	.w6(32'hbb133e90),
	.w7(32'hb99e0a1a),
	.w8(32'h3aac0c04),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5678ee),
	.w1(32'h3c21df0c),
	.w2(32'h3bf0e37b),
	.w3(32'h3bc11824),
	.w4(32'h3c05737e),
	.w5(32'h3c0cef9d),
	.w6(32'h3bdbab10),
	.w7(32'h3b99dec7),
	.w8(32'h3b453570),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c378245),
	.w1(32'hbaecb6b1),
	.w2(32'hbaa120c2),
	.w3(32'h3c4cb15a),
	.w4(32'hbbc0d06c),
	.w5(32'hbb1c55ed),
	.w6(32'hbaa18384),
	.w7(32'hbb15f6ba),
	.w8(32'hbb7a9b44),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081ae4),
	.w1(32'hbb9cdd82),
	.w2(32'hbba72480),
	.w3(32'h3a8784e5),
	.w4(32'h3a739295),
	.w5(32'hbacef82f),
	.w6(32'h3b9c7744),
	.w7(32'hbb3752eb),
	.w8(32'hbbaef08f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0e969),
	.w1(32'hbafe903a),
	.w2(32'hbbd51a90),
	.w3(32'h3ac4ea62),
	.w4(32'hbba470af),
	.w5(32'hbadb06b8),
	.w6(32'h37c7b7e1),
	.w7(32'hba81c1fd),
	.w8(32'hbb997e3a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d1e1),
	.w1(32'hb98564c4),
	.w2(32'hbabd8a3f),
	.w3(32'h39569011),
	.w4(32'h3abaf194),
	.w5(32'h3a113754),
	.w6(32'h3a72aaa2),
	.w7(32'h382e1cc1),
	.w8(32'h3aeec263),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ea79),
	.w1(32'hbc53ac0f),
	.w2(32'hbb7dc5ce),
	.w3(32'hba191d01),
	.w4(32'hbb688b2b),
	.w5(32'hbb9a5ec5),
	.w6(32'hbc2eeab6),
	.w7(32'hbb3bbbe5),
	.w8(32'hbbe7559a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc612d92),
	.w1(32'h3ac67805),
	.w2(32'hbafcedfe),
	.w3(32'hbc4ba5f8),
	.w4(32'h3b9e6ac2),
	.w5(32'h3b5ed3bc),
	.w6(32'h3ac44360),
	.w7(32'hbb81adea),
	.w8(32'hbbaf156c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98fb12),
	.w1(32'hbb3fcb4b),
	.w2(32'hbb8eddda),
	.w3(32'hbb9ee72c),
	.w4(32'hbaec9c17),
	.w5(32'hbb9e040d),
	.w6(32'hbb2e91ae),
	.w7(32'hbbc06d9b),
	.w8(32'hbb9a94d7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfdfbb),
	.w1(32'hbbc476e7),
	.w2(32'hbbc906d7),
	.w3(32'hbbaa0470),
	.w4(32'hbc0a15c9),
	.w5(32'hbc320ce9),
	.w6(32'hbaf2bb32),
	.w7(32'hbb3161ac),
	.w8(32'hbbe67c94),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1004),
	.w1(32'hb97a97b6),
	.w2(32'h39854fa1),
	.w3(32'hbb384c4e),
	.w4(32'h3a928e97),
	.w5(32'h3b2d67c0),
	.w6(32'h3a062a13),
	.w7(32'h388189ab),
	.w8(32'h3b1a7b7f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a81c6),
	.w1(32'h3a93521d),
	.w2(32'hbbc42d6f),
	.w3(32'h3b4376b9),
	.w4(32'h3b0e1a5f),
	.w5(32'hba1c8347),
	.w6(32'h3b801de8),
	.w7(32'h3bf8d975),
	.w8(32'hb99563fe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b537da0),
	.w1(32'hbc16523e),
	.w2(32'hbc42dd7c),
	.w3(32'h3b0029dd),
	.w4(32'hbc01dd34),
	.w5(32'hbbe09168),
	.w6(32'hbbf4cdaf),
	.w7(32'hbc18a27e),
	.w8(32'hbaccd433),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2479f0),
	.w1(32'hbb7c65ed),
	.w2(32'hbc5819f0),
	.w3(32'hbc03647c),
	.w4(32'hbab7d754),
	.w5(32'hbb531cca),
	.w6(32'hba850d6e),
	.w7(32'hbb846415),
	.w8(32'h3bf515aa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb672b09),
	.w1(32'hbbf3402f),
	.w2(32'hbc05e0f8),
	.w3(32'h3a779eb4),
	.w4(32'hbc01f55f),
	.w5(32'hba7e8694),
	.w6(32'hbc310ca6),
	.w7(32'hbc2e1d86),
	.w8(32'hbba24c4a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6664f),
	.w1(32'hbc05f3b6),
	.w2(32'hbbf347ee),
	.w3(32'hbbb7df6e),
	.w4(32'h398fdc7b),
	.w5(32'h3b4a66e4),
	.w6(32'hbc24aa8b),
	.w7(32'hbc0c9b54),
	.w8(32'hbbd7f44c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6f02),
	.w1(32'h3bc534d1),
	.w2(32'h3b6e5f70),
	.w3(32'h3b3a9af5),
	.w4(32'h3b14b9cd),
	.w5(32'h3c05f5f0),
	.w6(32'h3bd001ae),
	.w7(32'h3c19b393),
	.w8(32'h3b511f68),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba80e44),
	.w1(32'h3afdd896),
	.w2(32'h3b53bd90),
	.w3(32'h3bb38790),
	.w4(32'h36fa8889),
	.w5(32'h3a92d652),
	.w6(32'hbbf426bd),
	.w7(32'hbb70e6ad),
	.w8(32'hbbb651af),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e37a4),
	.w1(32'hba424414),
	.w2(32'hbbbcfc31),
	.w3(32'h3997cccb),
	.w4(32'h3a21ada3),
	.w5(32'hbab1a610),
	.w6(32'hbaaad5db),
	.w7(32'hbbbb8344),
	.w8(32'hbb8897e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695a51),
	.w1(32'h3bd97c40),
	.w2(32'h3b845904),
	.w3(32'hbb4d413e),
	.w4(32'h3bc3bacf),
	.w5(32'h3be170eb),
	.w6(32'h3c26c2d9),
	.w7(32'h3b68313a),
	.w8(32'h3ba1a3eb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33f9a9),
	.w1(32'hbb28469f),
	.w2(32'hbb13b5a6),
	.w3(32'h3cbc7497),
	.w4(32'hbb35a9de),
	.w5(32'hbafc3627),
	.w6(32'hbaac09bb),
	.w7(32'hba8dcc0c),
	.w8(32'hbba2d720),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08e09),
	.w1(32'hbb448247),
	.w2(32'h3ac2e14f),
	.w3(32'hbbc9721b),
	.w4(32'hbae7aed9),
	.w5(32'h3bbe0a41),
	.w6(32'h3ba33c16),
	.w7(32'h3ae5bd47),
	.w8(32'h3b265c24),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54aaa7),
	.w1(32'h3b9d7bca),
	.w2(32'h3b2a0ef9),
	.w3(32'h3c9cae2b),
	.w4(32'h3b8dd5c5),
	.w5(32'hbb058d3d),
	.w6(32'h3c376166),
	.w7(32'h3bd54f7c),
	.w8(32'h3c13ee43),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a923fe5),
	.w1(32'h3ab8b090),
	.w2(32'hbb9a0171),
	.w3(32'h39f3fc78),
	.w4(32'hbbd4828a),
	.w5(32'h3ab9f2ac),
	.w6(32'hbb336502),
	.w7(32'h3ab88de5),
	.w8(32'h3a75cd8b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1764f3),
	.w1(32'hbb222020),
	.w2(32'hbb72b0d6),
	.w3(32'h39d37b05),
	.w4(32'hbaa37711),
	.w5(32'hbaeae4c7),
	.w6(32'h3992c905),
	.w7(32'h3b35db3e),
	.w8(32'hbada4de1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc7de),
	.w1(32'hbba5384a),
	.w2(32'hbb408bc8),
	.w3(32'hbbc38386),
	.w4(32'hba0b7098),
	.w5(32'h393600d8),
	.w6(32'h3a068c6e),
	.w7(32'hbb22f145),
	.w8(32'h3b37ff5a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1403d6),
	.w1(32'hbb8674a9),
	.w2(32'h3a80e1bf),
	.w3(32'h3bafc967),
	.w4(32'hbb4c55d1),
	.w5(32'h3a61bda2),
	.w6(32'hbab712ef),
	.w7(32'hbb744c60),
	.w8(32'hbaa5e740),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba403840),
	.w1(32'h3a4b7156),
	.w2(32'h3a5da885),
	.w3(32'h3b8631d9),
	.w4(32'h3aefb9d3),
	.w5(32'h3ae5b65c),
	.w6(32'h3ab27a5e),
	.w7(32'hbafe3445),
	.w8(32'h38a8be3e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecf071),
	.w1(32'h3b9dcc49),
	.w2(32'h3adcce21),
	.w3(32'h3b4281a0),
	.w4(32'h3bc2d283),
	.w5(32'h3b1d5190),
	.w6(32'h3baad617),
	.w7(32'h3b9f665a),
	.w8(32'h3b88af58),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d43974),
	.w1(32'hbb95cd95),
	.w2(32'h3beb806c),
	.w3(32'hbab0bdd4),
	.w4(32'hbafdec2e),
	.w5(32'h3bf8bf4d),
	.w6(32'hba2bc76a),
	.w7(32'h3a4531d5),
	.w8(32'h3a99f4bd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79c40b),
	.w1(32'hbb986d21),
	.w2(32'hbbeae021),
	.w3(32'h3c1e1fc6),
	.w4(32'hba084db1),
	.w5(32'hba5ddd5a),
	.w6(32'hbbda7e6e),
	.w7(32'hbb1d463d),
	.w8(32'hbbac18c1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bb94e),
	.w1(32'h3be916b9),
	.w2(32'h3ba3439d),
	.w3(32'hba9fb277),
	.w4(32'h3b9764fe),
	.w5(32'h3ac65f6c),
	.w6(32'h3c09fd5b),
	.w7(32'h3c0030d1),
	.w8(32'h3be6b39f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f946),
	.w1(32'h3ab10b0b),
	.w2(32'h3b8adf56),
	.w3(32'h3a5d3247),
	.w4(32'hbae6d439),
	.w5(32'hbb72d49a),
	.w6(32'h3b252dfc),
	.w7(32'h3b8a6f91),
	.w8(32'h3c10d9ac),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc962d0),
	.w1(32'hbac48d37),
	.w2(32'hbb886cb5),
	.w3(32'hbb6f6aa3),
	.w4(32'hbb9658dd),
	.w5(32'h3ac1c91c),
	.w6(32'hbb33a13f),
	.w7(32'hbc05ad70),
	.w8(32'hbc0a7c09),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d04982),
	.w1(32'hbbabde23),
	.w2(32'hb7109eb3),
	.w3(32'h3bb242a3),
	.w4(32'hbb9471d9),
	.w5(32'hbb2c3126),
	.w6(32'hbb7f5cd2),
	.w7(32'hba3097a5),
	.w8(32'hbbed458d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e79eb),
	.w1(32'hbb882d44),
	.w2(32'hbbd3477b),
	.w3(32'hbba6543e),
	.w4(32'hbb896328),
	.w5(32'hbb0b4d82),
	.w6(32'hbad2b84f),
	.w7(32'hbb81e367),
	.w8(32'hbb013d5e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e80dd),
	.w1(32'hba3d1c7c),
	.w2(32'hba4dd51d),
	.w3(32'hbace5079),
	.w4(32'hbb127778),
	.w5(32'hbb5318e4),
	.w6(32'h38cd13ab),
	.w7(32'hba8c275d),
	.w8(32'hb82f2ab4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf72a0c),
	.w1(32'hbbcf6857),
	.w2(32'hbbb56ff4),
	.w3(32'hbb7cdce8),
	.w4(32'hbbc3733b),
	.w5(32'hbafaee3b),
	.w6(32'hbb8c5265),
	.w7(32'hbb27831a),
	.w8(32'hbb8edc09),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b07f),
	.w1(32'h3aba4c4a),
	.w2(32'hbb8b6266),
	.w3(32'h3b36c0e4),
	.w4(32'h39a20d22),
	.w5(32'hb92b476b),
	.w6(32'hbba044f3),
	.w7(32'hbb9f6cff),
	.w8(32'h3892a9e9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bd7ff),
	.w1(32'hbb90b6b7),
	.w2(32'hbc23e1be),
	.w3(32'hbbe63db5),
	.w4(32'hbb28e906),
	.w5(32'hbbbc62d7),
	.w6(32'hbb94f594),
	.w7(32'hbbf3ed3a),
	.w8(32'hbb4a5105),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ea41),
	.w1(32'h39a25f18),
	.w2(32'hbb88d677),
	.w3(32'hbbe12b92),
	.w4(32'hbbe618a4),
	.w5(32'hbbaef937),
	.w6(32'hbacbd22b),
	.w7(32'hbb992524),
	.w8(32'hbb81035b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bd89),
	.w1(32'h3a7d948e),
	.w2(32'hbaa6d9b1),
	.w3(32'hba9d639e),
	.w4(32'h3920e9ac),
	.w5(32'hba84c6bf),
	.w6(32'h3aaf10e5),
	.w7(32'h39b70c12),
	.w8(32'h39fe4b7f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59db03),
	.w1(32'hbaf1b455),
	.w2(32'hbb9c39f7),
	.w3(32'hba89ce40),
	.w4(32'hbb6b9841),
	.w5(32'hbc09fe0a),
	.w6(32'hb9ea72d0),
	.w7(32'hbb026bb6),
	.w8(32'hbb63ea23),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b11ec),
	.w1(32'hb92ca9fc),
	.w2(32'hbbad321f),
	.w3(32'hbb98b849),
	.w4(32'hbb1f335b),
	.w5(32'hbbeaf7e3),
	.w6(32'h3abf0860),
	.w7(32'hbae72d53),
	.w8(32'hbbae63e4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d5f05),
	.w1(32'h3b33cc1e),
	.w2(32'h3b14067a),
	.w3(32'hbc47845c),
	.w4(32'h3bbb6b8e),
	.w5(32'h3c0185d0),
	.w6(32'h3ab08421),
	.w7(32'hba2c6ff0),
	.w8(32'hbb80c7a9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8fff),
	.w1(32'hbb8f15b6),
	.w2(32'hbb78989b),
	.w3(32'hbb836d65),
	.w4(32'hbb920ae8),
	.w5(32'hbb31d242),
	.w6(32'hbbd86eb3),
	.w7(32'hbb80e6ed),
	.w8(32'h39dea931),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b409075),
	.w1(32'hbba11cc4),
	.w2(32'hbbc608d2),
	.w3(32'h3ad37245),
	.w4(32'hbaa5b4db),
	.w5(32'hbb76988b),
	.w6(32'h3aa9b66b),
	.w7(32'h3abb0179),
	.w8(32'hb91477dd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb822380),
	.w1(32'hbb4ea2d4),
	.w2(32'h3b0e1600),
	.w3(32'hbb9902b4),
	.w4(32'h3b884fa0),
	.w5(32'h3ca5850b),
	.w6(32'hbba31aba),
	.w7(32'hbbb10de0),
	.w8(32'h3b861680),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c5a61),
	.w1(32'hbaa4c76e),
	.w2(32'hbb0a8c22),
	.w3(32'h3cd10b42),
	.w4(32'hba14333c),
	.w5(32'h3b2690b7),
	.w6(32'hba8c0077),
	.w7(32'hbbad65de),
	.w8(32'hbb408513),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa042),
	.w1(32'hbb1ae79f),
	.w2(32'hbb146ad5),
	.w3(32'h3c3afbf3),
	.w4(32'hbb361dea),
	.w5(32'hba8779a8),
	.w6(32'hbb617fd7),
	.w7(32'hbb486955),
	.w8(32'hbb266b74),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf595),
	.w1(32'hbbfe7aeb),
	.w2(32'hbc18b04a),
	.w3(32'hb9050c2e),
	.w4(32'hbb6cf5c0),
	.w5(32'hbb4e2c0c),
	.w6(32'hbc2ee0bd),
	.w7(32'hbb9ca3b6),
	.w8(32'hbc14a0ae),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98930f),
	.w1(32'hbbb619a7),
	.w2(32'hbb3b4ade),
	.w3(32'hbb809a86),
	.w4(32'hbba15f47),
	.w5(32'h3bc885e2),
	.w6(32'hbbb1dae3),
	.w7(32'hbbae6761),
	.w8(32'hb9fc0574),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac8760),
	.w1(32'h399025be),
	.w2(32'hbb50b699),
	.w3(32'h3b5ecc61),
	.w4(32'hbabe6791),
	.w5(32'hbc2b75ab),
	.w6(32'hbb13f209),
	.w7(32'hbb334a79),
	.w8(32'hbaf10a14),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc345cce),
	.w1(32'h3c16c7e2),
	.w2(32'h3b91fba5),
	.w3(32'hbc9145ed),
	.w4(32'h3c1155cd),
	.w5(32'h3b57e3be),
	.w6(32'h3c1002e9),
	.w7(32'h3b88c7a2),
	.w8(32'h3c0fd248),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fbedf),
	.w1(32'h3b9f4bbe),
	.w2(32'h3b8e6aca),
	.w3(32'h3b5fc656),
	.w4(32'h3b311643),
	.w5(32'h3ac18f85),
	.w6(32'h3bc19523),
	.w7(32'h3baded7f),
	.w8(32'h3b66c907),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4841ec),
	.w1(32'h3bb2d858),
	.w2(32'h3b423b54),
	.w3(32'hb77f7a52),
	.w4(32'h3b632bd0),
	.w5(32'h3af9de07),
	.w6(32'h3bdd2353),
	.w7(32'h3b9c209a),
	.w8(32'h3b63580b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3c2ea),
	.w1(32'hbb293496),
	.w2(32'hb9673d7d),
	.w3(32'h3b47f91b),
	.w4(32'hbb4d9900),
	.w5(32'hbb538266),
	.w6(32'hb4c04256),
	.w7(32'hbb8598d4),
	.w8(32'hba262bcc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe63ce),
	.w1(32'h3b6a0be5),
	.w2(32'hbb0fd3e5),
	.w3(32'hbabcdfba),
	.w4(32'h3aa25751),
	.w5(32'hbbfe3deb),
	.w6(32'hbb778614),
	.w7(32'hbb80ae81),
	.w8(32'hbbb14060),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f8053),
	.w1(32'h3acb1a70),
	.w2(32'hbae6be8b),
	.w3(32'hbc727829),
	.w4(32'h3b4d5888),
	.w5(32'h3b80cb2a),
	.w6(32'h3b8d26e2),
	.w7(32'hba5c5b43),
	.w8(32'h3a40dad8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920ecbf),
	.w1(32'h3abf0cbf),
	.w2(32'hbc27cd03),
	.w3(32'hbb844a27),
	.w4(32'hba25ca9c),
	.w5(32'h3a3b84df),
	.w6(32'h3988f6bb),
	.w7(32'hbae62c5c),
	.w8(32'hba94e8a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8a654),
	.w1(32'hbaca502a),
	.w2(32'hbbc6cc13),
	.w3(32'hbb8ee976),
	.w4(32'h3b5dad8b),
	.w5(32'h3b209634),
	.w6(32'hbbb3b565),
	.w7(32'hbc2e6b0e),
	.w8(32'h3ba210c5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649848),
	.w1(32'hbb9f3831),
	.w2(32'hbb98a41c),
	.w3(32'h3c2d3a74),
	.w4(32'hbb1365de),
	.w5(32'hbbc37799),
	.w6(32'hbbd35910),
	.w7(32'hbb08955a),
	.w8(32'h3a4770ee),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc829),
	.w1(32'hbb22233e),
	.w2(32'hba6a26c3),
	.w3(32'hbc4ffee9),
	.w4(32'hbbacbf1e),
	.w5(32'hbad42d73),
	.w6(32'hbba47f12),
	.w7(32'hbac79b73),
	.w8(32'h3a8ad444),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab871e8),
	.w1(32'hbb9836e6),
	.w2(32'hbb033cfd),
	.w3(32'h3b40a1e0),
	.w4(32'hbb82e423),
	.w5(32'hbba797b2),
	.w6(32'h3b9047dd),
	.w7(32'h3ae776c1),
	.w8(32'hbb0daafd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2767),
	.w1(32'hbc107852),
	.w2(32'hbbdaf3f2),
	.w3(32'hba735d7a),
	.w4(32'hbb5d2352),
	.w5(32'hba802229),
	.w6(32'hbb918a47),
	.w7(32'hbbb89c6d),
	.w8(32'hbb50358e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea4029),
	.w1(32'hbbdc7fe6),
	.w2(32'hbc2bc785),
	.w3(32'h3b3094dd),
	.w4(32'hbbd7aa50),
	.w5(32'hbbfa0517),
	.w6(32'hbc17b3bf),
	.w7(32'hbc0d1632),
	.w8(32'hbb64b60a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f1f8),
	.w1(32'hb90109a9),
	.w2(32'hbb0db5c0),
	.w3(32'hbb84431c),
	.w4(32'hbb5eb942),
	.w5(32'h3aad8947),
	.w6(32'h3b154a35),
	.w7(32'hbabf8d02),
	.w8(32'h3bc37ad5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcd7f7),
	.w1(32'hbbfb9d9b),
	.w2(32'hbbc30bb2),
	.w3(32'hbb564fd3),
	.w4(32'hbb832da5),
	.w5(32'h3addb2cc),
	.w6(32'hbbca2d00),
	.w7(32'hbc0dc826),
	.w8(32'hbb858566),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b640dcd),
	.w1(32'hbbc7fa25),
	.w2(32'hbbbbe578),
	.w3(32'h3c034145),
	.w4(32'hbba715ec),
	.w5(32'h3ac20aa0),
	.w6(32'hbbaa375b),
	.w7(32'hbbfa1a69),
	.w8(32'hbab82a2e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73ba81),
	.w1(32'hbc556328),
	.w2(32'hbc1a5444),
	.w3(32'h3c44a7b4),
	.w4(32'hbc68b730),
	.w5(32'hbbbd08bf),
	.w6(32'hbc1a0e21),
	.w7(32'hbc036a26),
	.w8(32'hbb6854c1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2f0e4),
	.w1(32'h3a38757e),
	.w2(32'hbb69e57e),
	.w3(32'h39945a3d),
	.w4(32'h3a4da51d),
	.w5(32'hbb5891a1),
	.w6(32'hbaae51bc),
	.w7(32'hb8c5c7a5),
	.w8(32'h3a05062a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cf2e),
	.w1(32'h3be0fe5f),
	.w2(32'h3ad3e9b4),
	.w3(32'hb9a22826),
	.w4(32'hbad32f77),
	.w5(32'hba75a74a),
	.w6(32'hba1db7e3),
	.w7(32'hbb5163ae),
	.w8(32'hbb7a8914),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1fef),
	.w1(32'hbaa04875),
	.w2(32'hbb54cd5b),
	.w3(32'h3b5afbba),
	.w4(32'hbb8ef098),
	.w5(32'hbb817133),
	.w6(32'hbbb4f527),
	.w7(32'hbb6bf4f8),
	.w8(32'hbbb292fb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bc8ce),
	.w1(32'h3a8a0a94),
	.w2(32'hbac7ca1f),
	.w3(32'hbbdff482),
	.w4(32'h3b3678e5),
	.w5(32'h3a004a99),
	.w6(32'h3c1efec0),
	.w7(32'h3b1f8906),
	.w8(32'h3b493108),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b1dba),
	.w1(32'hbba9d6ee),
	.w2(32'hbafc767d),
	.w3(32'hbbee395e),
	.w4(32'h3abd8c58),
	.w5(32'hbba700da),
	.w6(32'hbc1a4168),
	.w7(32'hbba840c1),
	.w8(32'hbb4aa7aa),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b590a),
	.w1(32'hbb8212df),
	.w2(32'hba079786),
	.w3(32'hbb5cf580),
	.w4(32'h3a460942),
	.w5(32'h3b8e21bf),
	.w6(32'hbb6ceac6),
	.w7(32'hba401d33),
	.w8(32'hbb2cd83a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e93c),
	.w1(32'hb9380449),
	.w2(32'hbc191a57),
	.w3(32'h3ba58783),
	.w4(32'hbbd6d134),
	.w5(32'hbc324ddc),
	.w6(32'h3a851c31),
	.w7(32'hbbcc147e),
	.w8(32'hbba0b343),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c7c45),
	.w1(32'h393db708),
	.w2(32'h3b85ca27),
	.w3(32'hbc56ad02),
	.w4(32'h3b85ea42),
	.w5(32'h3b4e1637),
	.w6(32'h3abe2ffd),
	.w7(32'h3b67e797),
	.w8(32'h3ba4fccf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a561b),
	.w1(32'h3b4c911d),
	.w2(32'h3944f899),
	.w3(32'h3bbea21e),
	.w4(32'h3b6e43e3),
	.w5(32'hb9b01fa8),
	.w6(32'hb896de91),
	.w7(32'hba61408f),
	.w8(32'hbb4c23ab),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0df1c),
	.w1(32'hbb2ebb4b),
	.w2(32'h39e7ea0b),
	.w3(32'hbb98cc9a),
	.w4(32'h3a0f31d7),
	.w5(32'h3bcad1da),
	.w6(32'h3a356a06),
	.w7(32'hba331779),
	.w8(32'hb8f765a0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a602c),
	.w1(32'h3aa6e736),
	.w2(32'hba70fa97),
	.w3(32'h3c8130d4),
	.w4(32'hbbde60c8),
	.w5(32'h3b2a4fe9),
	.w6(32'hbb8cc796),
	.w7(32'hba8d1499),
	.w8(32'hbb35f948),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be64452),
	.w1(32'h3a10b46c),
	.w2(32'h3a3e3fdc),
	.w3(32'h3bf6f396),
	.w4(32'hbb9b2c3c),
	.w5(32'hbb436f88),
	.w6(32'h39f3ae2e),
	.w7(32'h3af141fe),
	.w8(32'hbae6a874),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c05da),
	.w1(32'hb80bca84),
	.w2(32'hbc059294),
	.w3(32'hbb411e3d),
	.w4(32'h39b7d403),
	.w5(32'h3ab304fc),
	.w6(32'hbbc703bf),
	.w7(32'hbbed1902),
	.w8(32'hbbee230b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587781),
	.w1(32'h3ac4399e),
	.w2(32'h3ad62f29),
	.w3(32'hbaecfcf8),
	.w4(32'h3a252ac2),
	.w5(32'h39a46f90),
	.w6(32'h3a8b3ae6),
	.w7(32'h3ae33fb2),
	.w8(32'h39facb89),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c7a26),
	.w1(32'hbacb5274),
	.w2(32'hba2560be),
	.w3(32'h3a8335a0),
	.w4(32'hbb11f9a2),
	.w5(32'hbad210ae),
	.w6(32'hbac4eaae),
	.w7(32'hba31d980),
	.w8(32'hbb1b63a3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d229),
	.w1(32'hbc4830e7),
	.w2(32'hbc87d4fc),
	.w3(32'hba7a8f18),
	.w4(32'hbbe33ac6),
	.w5(32'hbc11773c),
	.w6(32'hbbbc0180),
	.w7(32'hbc4b362f),
	.w8(32'hbc2c772c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128ef5),
	.w1(32'h3b22dcdb),
	.w2(32'h3ba04fb1),
	.w3(32'h3b8d9233),
	.w4(32'h3bd8ab12),
	.w5(32'h3c35a0d0),
	.w6(32'h3ab7a12a),
	.w7(32'h3a92cd7a),
	.w8(32'h3bb20065),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c604456),
	.w1(32'hbb6aca0b),
	.w2(32'hbab4898a),
	.w3(32'h3c9ddb2a),
	.w4(32'hbb673bbc),
	.w5(32'h3bc068d8),
	.w6(32'hbb60ef38),
	.w7(32'h3ae8ec10),
	.w8(32'h3b63bafd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30d4f3),
	.w1(32'hb5b0f519),
	.w2(32'hbaccafe7),
	.w3(32'h3c2483cc),
	.w4(32'h3b9ad2db),
	.w5(32'h39404b45),
	.w6(32'hbc12f5ff),
	.w7(32'hba03b386),
	.w8(32'h3be9f8ba),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b620b9d),
	.w1(32'hbbb40983),
	.w2(32'h3aab94d1),
	.w3(32'hba2434a9),
	.w4(32'hbba23743),
	.w5(32'hb9ed4676),
	.w6(32'h39a40f8b),
	.w7(32'hbb02cb1f),
	.w8(32'hbb1c2ee9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6776f),
	.w1(32'hbbb3dd07),
	.w2(32'hbc431d5f),
	.w3(32'hba505ce0),
	.w4(32'hbbd699dc),
	.w5(32'hba1fe8b1),
	.w6(32'hbaf18efb),
	.w7(32'hbc34cdb0),
	.w8(32'hbb713828),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990e602),
	.w1(32'h395d8490),
	.w2(32'hba8313af),
	.w3(32'hbad2b0bb),
	.w4(32'h3b92d27b),
	.w5(32'hbb2ad2e2),
	.w6(32'hbb7b8ddb),
	.w7(32'hbbc5afbc),
	.w8(32'h3ae79267),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20628b),
	.w1(32'h3aaebf23),
	.w2(32'h3a651812),
	.w3(32'hb70760a4),
	.w4(32'hbaf1b341),
	.w5(32'hbbaef63e),
	.w6(32'hbaf205e1),
	.w7(32'h3a072256),
	.w8(32'hb987fbf7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25399),
	.w1(32'hbbd60952),
	.w2(32'hbbfd11ad),
	.w3(32'hbc00b2f8),
	.w4(32'hba3db14d),
	.w5(32'hbb44212e),
	.w6(32'hbb76e7b2),
	.w7(32'hbbb3ce03),
	.w8(32'hbb6b1762),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb224d71),
	.w1(32'h3a437ebe),
	.w2(32'h3c87fb8d),
	.w3(32'hbb7a3d73),
	.w4(32'hb98c4d5e),
	.w5(32'h3c2a844d),
	.w6(32'h3b254166),
	.w7(32'h3bd436d7),
	.w8(32'h3c8d5721),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d098c54),
	.w1(32'hbab3c9c5),
	.w2(32'hba927b90),
	.w3(32'h3ba4b5ac),
	.w4(32'h388fb55b),
	.w5(32'h3afe44b7),
	.w6(32'h3ab6fca4),
	.w7(32'hb920bebc),
	.w8(32'h3a144d06),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3775c350),
	.w1(32'h3a30fb42),
	.w2(32'hba4927a6),
	.w3(32'hbb94d7a0),
	.w4(32'h3a9de928),
	.w5(32'h395560f4),
	.w6(32'h3b2c95f5),
	.w7(32'h3a921146),
	.w8(32'h3a959524),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb83c),
	.w1(32'hbc50dd3f),
	.w2(32'hbbe0c778),
	.w3(32'hbb05f268),
	.w4(32'hb9a85830),
	.w5(32'h3b641f5e),
	.w6(32'hbbfb1222),
	.w7(32'hbc0762b9),
	.w8(32'hbb481ca9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54c99),
	.w1(32'hbb6599ff),
	.w2(32'hbb2894f3),
	.w3(32'h3c0f790e),
	.w4(32'hbbca2fe3),
	.w5(32'h39a9f494),
	.w6(32'hbba204a8),
	.w7(32'hbc18e29d),
	.w8(32'hbc297dc3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec6828),
	.w1(32'h3b0750df),
	.w2(32'h3b839223),
	.w3(32'h3a2faaa2),
	.w4(32'h3bacfe50),
	.w5(32'h3b3ffeb9),
	.w6(32'h3b13a624),
	.w7(32'h3a13f9ff),
	.w8(32'h3b18630e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfba15),
	.w1(32'h3b3fe5db),
	.w2(32'h3b4df68f),
	.w3(32'hb8b7ae96),
	.w4(32'h3b098cbf),
	.w5(32'h3ab160a7),
	.w6(32'h3b222775),
	.w7(32'h3b20cafb),
	.w8(32'h3abafe11),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92d12f),
	.w1(32'hbae26fad),
	.w2(32'hbbea8fa3),
	.w3(32'h3a2334d2),
	.w4(32'hbb25d062),
	.w5(32'hbb0c6333),
	.w6(32'hbb29f225),
	.w7(32'hba11762b),
	.w8(32'hbb0f639b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad49ee6),
	.w1(32'hba22b414),
	.w2(32'hb9c6d702),
	.w3(32'hbacbe4f6),
	.w4(32'hba99a5c1),
	.w5(32'hb93319ba),
	.w6(32'h3a931154),
	.w7(32'h367ba237),
	.w8(32'h3a84293f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e3aaa),
	.w1(32'hbb618b09),
	.w2(32'hbc362d1c),
	.w3(32'h3b0c029c),
	.w4(32'hbadbc614),
	.w5(32'hbba8a1ca),
	.w6(32'hbb9c06c7),
	.w7(32'hbb494ec6),
	.w8(32'hbb6220aa),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02a409),
	.w1(32'h3b50383d),
	.w2(32'hbaaab8be),
	.w3(32'hba86f3ed),
	.w4(32'h3b19e072),
	.w5(32'h3a0a7800),
	.w6(32'h3b189843),
	.w7(32'hbbda33b7),
	.w8(32'hbba4daa5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84785d),
	.w1(32'hbaa1568e),
	.w2(32'hb97e6544),
	.w3(32'hbb809a0a),
	.w4(32'hbb5da7a1),
	.w5(32'hbb46836b),
	.w6(32'h3b60eb6a),
	.w7(32'h3a474c09),
	.w8(32'hba8c4584),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cbad9),
	.w1(32'h3b582bdd),
	.w2(32'h3a7f77c0),
	.w3(32'h3ae26d4c),
	.w4(32'h3ab8eca1),
	.w5(32'h381bade0),
	.w6(32'h3b6f8aa4),
	.w7(32'h3ad7e890),
	.w8(32'h38e14cfb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36fd61),
	.w1(32'h3a4ef94a),
	.w2(32'hb95e2baf),
	.w3(32'hb9af1541),
	.w4(32'h3baa38d9),
	.w5(32'hbb381a91),
	.w6(32'h3bb6deb7),
	.w7(32'h3b4d69b3),
	.w8(32'h3b5b7199),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23c5a8),
	.w1(32'hbb4eac94),
	.w2(32'hbb7bee59),
	.w3(32'hbc69a720),
	.w4(32'hbb5f4b3c),
	.w5(32'hbb7935d9),
	.w6(32'hbb577705),
	.w7(32'hbb647d6e),
	.w8(32'h38f1ef5e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897f2c),
	.w1(32'h3ab4a3d0),
	.w2(32'h3b18885e),
	.w3(32'hbbbf01bb),
	.w4(32'hbb0e8fcc),
	.w5(32'h3a2b987f),
	.w6(32'hbba4e355),
	.w7(32'hbbeaadf5),
	.w8(32'hbb5f2e4f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa86110),
	.w1(32'hba8b1348),
	.w2(32'hba9d8a71),
	.w3(32'h3b6f1ba2),
	.w4(32'hbb1ba98d),
	.w5(32'hbaef8fdf),
	.w6(32'hb9b63c21),
	.w7(32'hb990324d),
	.w8(32'h3a3bfab3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79797),
	.w1(32'hbc134071),
	.w2(32'hbc0ff9fb),
	.w3(32'h39da6c96),
	.w4(32'hbc2c2da8),
	.w5(32'hbc1da8b0),
	.w6(32'hba378ba9),
	.w7(32'hbba51759),
	.w8(32'hb9b8cf4e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c4c4),
	.w1(32'hbb011bc2),
	.w2(32'h3b59926f),
	.w3(32'hbbe71062),
	.w4(32'hb95d27fe),
	.w5(32'h385748ba),
	.w6(32'h3b9b94df),
	.w7(32'hb96afa69),
	.w8(32'hba5d7b39),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d112),
	.w1(32'h3b2391fc),
	.w2(32'h3b094887),
	.w3(32'h38f6f7d1),
	.w4(32'h3b385e47),
	.w5(32'h3a90980b),
	.w6(32'h3b2d9f22),
	.w7(32'h3b140251),
	.w8(32'h3b07e07d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ba06b),
	.w1(32'hbb777c5c),
	.w2(32'hbbd50374),
	.w3(32'h3a009bcc),
	.w4(32'hbb1288ad),
	.w5(32'hbc0933c8),
	.w6(32'hbb6d42ed),
	.w7(32'hbb508550),
	.w8(32'hba337b06),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034fa1),
	.w1(32'hbbd98c59),
	.w2(32'hbba2a017),
	.w3(32'hbbc7d71a),
	.w4(32'hbb206400),
	.w5(32'hbaf1789e),
	.w6(32'hbc35d2df),
	.w7(32'hbc29e7a9),
	.w8(32'hbb3aac98),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a36b2),
	.w1(32'hbc09fb9c),
	.w2(32'hbb7a6ee0),
	.w3(32'hbbd1fce5),
	.w4(32'hb992f4f0),
	.w5(32'hbc233d47),
	.w6(32'hbc20e549),
	.w7(32'hbb775b97),
	.w8(32'hbbac0bb3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa162),
	.w1(32'hb5adb0b4),
	.w2(32'h3adb0414),
	.w3(32'hb536ce4d),
	.w4(32'hb937733e),
	.w5(32'h3a8ec0e3),
	.w6(32'hb9866dfa),
	.w7(32'h3a87d16b),
	.w8(32'hb847a02f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977fb23),
	.w1(32'hbbc6297d),
	.w2(32'hbb4b90d5),
	.w3(32'hb8f7e7b1),
	.w4(32'hbbbce358),
	.w5(32'hbb397020),
	.w6(32'hbbb4385f),
	.w7(32'hbb2d0385),
	.w8(32'h3a1bda19),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule