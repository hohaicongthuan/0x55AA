module layer_10_featuremap_82(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9602e7d),
	.w1(32'hbaccf0fe),
	.w2(32'hb86c6508),
	.w3(32'hb8a90f99),
	.w4(32'h3a694f39),
	.w5(32'hbb1729b8),
	.w6(32'hba8d2f41),
	.w7(32'h3a9d50ca),
	.w8(32'hbaf01d42),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc40bb),
	.w1(32'h3a966ff5),
	.w2(32'h3addfdea),
	.w3(32'h38349a77),
	.w4(32'hbaa97150),
	.w5(32'h3b5acf09),
	.w6(32'hbb1ddfb1),
	.w7(32'h3adac5ac),
	.w8(32'hbac7710b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223215),
	.w1(32'h3a937330),
	.w2(32'h3b4a7544),
	.w3(32'hb9ccaa63),
	.w4(32'h3ba6d432),
	.w5(32'hbb37a701),
	.w6(32'h3b040a21),
	.w7(32'hbaff66cf),
	.w8(32'h3a7b8bfa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a00a9),
	.w1(32'h3bea0115),
	.w2(32'h3934324e),
	.w3(32'h3b6b1b4f),
	.w4(32'h3b2adff3),
	.w5(32'h39d2da0a),
	.w6(32'h39add518),
	.w7(32'h3b3cedff),
	.w8(32'hba37b279),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab109eb),
	.w1(32'h3a9ab113),
	.w2(32'h3ae9061a),
	.w3(32'hbaf6af00),
	.w4(32'h3a79e2a6),
	.w5(32'hb93923b2),
	.w6(32'h3b7ef634),
	.w7(32'hba1a48b2),
	.w8(32'hbb2f6056),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bffef),
	.w1(32'hbad8846b),
	.w2(32'h3a8dad71),
	.w3(32'h3a47a3e6),
	.w4(32'h3a60b6f9),
	.w5(32'hba669116),
	.w6(32'h3a673d72),
	.w7(32'hba9b3b56),
	.w8(32'hbaa24a80),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d94a),
	.w1(32'hbbcce91d),
	.w2(32'hbb0c8b4d),
	.w3(32'hbaf4587b),
	.w4(32'hba48bb7b),
	.w5(32'h3c704fac),
	.w6(32'hbb812885),
	.w7(32'hbb23ac45),
	.w8(32'h3c79ac5c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59acc2),
	.w1(32'h38c322c7),
	.w2(32'hb8df3acd),
	.w3(32'h3a12fc41),
	.w4(32'hbaa74d7c),
	.w5(32'h3b485753),
	.w6(32'h3b993aa2),
	.w7(32'hb98c0119),
	.w8(32'h3bc08d56),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1470),
	.w1(32'h3c5669ef),
	.w2(32'h3b511640),
	.w3(32'hbb18af26),
	.w4(32'hbbb78f2e),
	.w5(32'hb9c70544),
	.w6(32'h39fb6a55),
	.w7(32'hbad95966),
	.w8(32'h37af0eb9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101a27),
	.w1(32'h389ba79e),
	.w2(32'h3b73dd09),
	.w3(32'hbafd105a),
	.w4(32'h3b4aecea),
	.w5(32'hb7724761),
	.w6(32'h39980d22),
	.w7(32'hbc107af7),
	.w8(32'hbb253096),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c272c),
	.w1(32'hbae6a995),
	.w2(32'h3b265b0e),
	.w3(32'h3a536e32),
	.w4(32'h3b70115c),
	.w5(32'hbb71c4db),
	.w6(32'hba67a86d),
	.w7(32'hbb835f8f),
	.w8(32'hba7bbc0a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c16af),
	.w1(32'hba945945),
	.w2(32'hba4053ea),
	.w3(32'h3a870445),
	.w4(32'h3b4548f7),
	.w5(32'hb9039b62),
	.w6(32'hbaae28af),
	.w7(32'hb85f9f67),
	.w8(32'hba7ec3fa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc30c),
	.w1(32'h3a0fcd06),
	.w2(32'hbb94b7f0),
	.w3(32'hbab704d5),
	.w4(32'h39b43581),
	.w5(32'hbaa3ae27),
	.w6(32'hbb64e208),
	.w7(32'hbaa51e9c),
	.w8(32'h3b02b0c2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced0579),
	.w1(32'hbb078924),
	.w2(32'hbb21017e),
	.w3(32'h3ae74b5d),
	.w4(32'h3ad0624a),
	.w5(32'hb9e586c8),
	.w6(32'hbba19fb1),
	.w7(32'h3b39c3a0),
	.w8(32'h37b1b202),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb191a3),
	.w1(32'h3b2830fd),
	.w2(32'hbacf4ec9),
	.w3(32'h398e2735),
	.w4(32'h3a8d18e3),
	.w5(32'h3a78de5d),
	.w6(32'h39d29c9f),
	.w7(32'h3b985cb6),
	.w8(32'h3a78484f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3619f3),
	.w1(32'hb99eaaa8),
	.w2(32'h3b119f57),
	.w3(32'h3c6871e9),
	.w4(32'hba898e14),
	.w5(32'hbac61154),
	.w6(32'hba136b73),
	.w7(32'h3a0b230d),
	.w8(32'h3c46276a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a97f),
	.w1(32'h3c15010c),
	.w2(32'h3b357327),
	.w3(32'hbb1b114d),
	.w4(32'h383653d6),
	.w5(32'hbbe3e85a),
	.w6(32'hb9be1f26),
	.w7(32'hbb4426f6),
	.w8(32'hbb1cac1b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf20925),
	.w1(32'hbbeaff30),
	.w2(32'h3a9df150),
	.w3(32'hb94e6995),
	.w4(32'h3b3194ae),
	.w5(32'h39a05d0e),
	.w6(32'h3b9cd30d),
	.w7(32'hbbf30d0d),
	.w8(32'hba81863e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0903d4),
	.w1(32'hbb51aca5),
	.w2(32'hba5312a7),
	.w3(32'h3ba64037),
	.w4(32'hbb301017),
	.w5(32'h3b636cd3),
	.w6(32'hba9b48b6),
	.w7(32'hbb549c70),
	.w8(32'h3993b868),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41d0ac),
	.w1(32'hbb780cf3),
	.w2(32'hbaf89a72),
	.w3(32'h3a04c7b6),
	.w4(32'h3bb62500),
	.w5(32'hb99a2c0c),
	.w6(32'hba9f25c7),
	.w7(32'hba91ba53),
	.w8(32'hbb1d3201),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11398),
	.w1(32'h3ad75732),
	.w2(32'h3a7a1d5a),
	.w3(32'hb9411abe),
	.w4(32'h3b567b22),
	.w5(32'h3b40ac0f),
	.w6(32'h3bf4e9c8),
	.w7(32'h3b89ad89),
	.w8(32'hba6a9e4c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa57d44),
	.w1(32'hbad0aa71),
	.w2(32'hbb847594),
	.w3(32'h37931868),
	.w4(32'h3a56eca8),
	.w5(32'h3a5fe4b0),
	.w6(32'hb9b96402),
	.w7(32'hb8b165d6),
	.w8(32'h3795d118),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abef0d7),
	.w1(32'h39aae01b),
	.w2(32'hbc2c79f9),
	.w3(32'h39f0fe92),
	.w4(32'h3a9c92cc),
	.w5(32'hbc6ab1f3),
	.w6(32'hbace5634),
	.w7(32'h3b7da931),
	.w8(32'h3961359d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4a748),
	.w1(32'h3a6689df),
	.w2(32'hb90cfdb7),
	.w3(32'h3aa49512),
	.w4(32'hba0fd96f),
	.w5(32'h3b3756a8),
	.w6(32'h3b0a3f11),
	.w7(32'hb9258fa2),
	.w8(32'hb9ade3cb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968418),
	.w1(32'h3b472e33),
	.w2(32'h3bd7dbe9),
	.w3(32'h3af7039f),
	.w4(32'h3ac76f4d),
	.w5(32'h3b4a1720),
	.w6(32'hba660741),
	.w7(32'hbad32391),
	.w8(32'hbb249639),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e84b9),
	.w1(32'hbacca146),
	.w2(32'hbb38e7ba),
	.w3(32'h3b196bad),
	.w4(32'hbc43d4b2),
	.w5(32'hba643137),
	.w6(32'hbb75ce95),
	.w7(32'hbaf2b91b),
	.w8(32'h390bae7c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175222),
	.w1(32'h39f6e00c),
	.w2(32'hbb9abe30),
	.w3(32'hba1ff6da),
	.w4(32'h3af12787),
	.w5(32'hba691fa1),
	.w6(32'hb92194cd),
	.w7(32'hba65d2ae),
	.w8(32'hbb6b8ffe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aee5c),
	.w1(32'h3b4828be),
	.w2(32'h3c89b03e),
	.w3(32'hbb40de27),
	.w4(32'hbc614dd3),
	.w5(32'h3c9bea73),
	.w6(32'hba6bb64d),
	.w7(32'h3badc514),
	.w8(32'hbb8dc503),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62673b),
	.w1(32'h3bb0453f),
	.w2(32'hbbc7e0f8),
	.w3(32'hbb6d8fda),
	.w4(32'h398d0c33),
	.w5(32'h3b8cbb97),
	.w6(32'hbb2c1f6b),
	.w7(32'hbb0ce0e4),
	.w8(32'hbbc2a3de),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80791c),
	.w1(32'hbb53cb93),
	.w2(32'h3bdb1525),
	.w3(32'hbb85edc0),
	.w4(32'hbb846beb),
	.w5(32'h3bc612e2),
	.w6(32'h3c41c3b1),
	.w7(32'h39e797b8),
	.w8(32'hbb92bebf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c05b),
	.w1(32'h3b987613),
	.w2(32'hbc10c69f),
	.w3(32'hba22eb92),
	.w4(32'hbb2e577f),
	.w5(32'hbb265b9b),
	.w6(32'hbb4291ee),
	.w7(32'hbb9e4edd),
	.w8(32'hbc4af91e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3acbbd),
	.w1(32'hba636ade),
	.w2(32'hbb5df5f7),
	.w3(32'hbb43311b),
	.w4(32'h3b224cde),
	.w5(32'h3bd039f8),
	.w6(32'hbb8ea8d3),
	.w7(32'hbb922f2b),
	.w8(32'h3c68ff9e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1775ee),
	.w1(32'hbc0b9bf6),
	.w2(32'hbbb513ac),
	.w3(32'hbbfc4faf),
	.w4(32'h3b23157d),
	.w5(32'h3bf2585c),
	.w6(32'h3b0e083e),
	.w7(32'h3bf44c94),
	.w8(32'hbae4892e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0b55),
	.w1(32'h3d386401),
	.w2(32'hbbf567b8),
	.w3(32'hbad141c0),
	.w4(32'h3b06052f),
	.w5(32'h3a826601),
	.w6(32'h38a29a8f),
	.w7(32'h3b95627a),
	.w8(32'h398d33d9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d49b8),
	.w1(32'hbbdd789f),
	.w2(32'hbb59d669),
	.w3(32'h3a8fa7a7),
	.w4(32'h3aa15115),
	.w5(32'h3a7469ff),
	.w6(32'hbb50be3c),
	.w7(32'h3c5b0f7b),
	.w8(32'h3b7a3054),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2563fc),
	.w1(32'h3c2cc570),
	.w2(32'hbc6da9a1),
	.w3(32'h3c235d8a),
	.w4(32'hbb78f8b5),
	.w5(32'hbb8a0335),
	.w6(32'hbb5c3385),
	.w7(32'h39ddf432),
	.w8(32'h3bf3373b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8c59),
	.w1(32'hba481d38),
	.w2(32'h3b7be7e7),
	.w3(32'h3b974e9b),
	.w4(32'h3b75a76f),
	.w5(32'hbbc16fd6),
	.w6(32'h3afd4ec8),
	.w7(32'hbbe35d1f),
	.w8(32'h3a94956b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389de262),
	.w1(32'h3864ade0),
	.w2(32'h3c5ddd02),
	.w3(32'h3bf7968e),
	.w4(32'h3b2b2704),
	.w5(32'h3850cb5d),
	.w6(32'hbbc9254e),
	.w7(32'h3ac68596),
	.w8(32'h397a4d00),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a831857),
	.w1(32'h3c0d727f),
	.w2(32'h3b05a038),
	.w3(32'hbb50f58c),
	.w4(32'h3aed0281),
	.w5(32'hbb193eb3),
	.w6(32'hbc0136f1),
	.w7(32'hbc255a93),
	.w8(32'h3b5fe52e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7f0cd),
	.w1(32'h3abc0f22),
	.w2(32'hbae913df),
	.w3(32'hba4f53a9),
	.w4(32'h394d1ab5),
	.w5(32'hba6359ac),
	.w6(32'hbb604a0d),
	.w7(32'h3a377eb5),
	.w8(32'h3b1e41c0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h32bd686d),
	.w1(32'hbb6a0670),
	.w2(32'hbc1b9a7f),
	.w3(32'h3c01b91b),
	.w4(32'h3aaa45e5),
	.w5(32'hbba475cf),
	.w6(32'h3892ab28),
	.w7(32'hbb957f4b),
	.w8(32'hba70679c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a698b5b),
	.w1(32'hb8d0ec11),
	.w2(32'hbbd71963),
	.w3(32'hb811f81c),
	.w4(32'hbb14a422),
	.w5(32'h3af02546),
	.w6(32'hbbbc18ae),
	.w7(32'hbbdb5ebb),
	.w8(32'h3c3e14cd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd2ec0),
	.w1(32'hb9c0b79e),
	.w2(32'hbc1070bd),
	.w3(32'h3cabb0ac),
	.w4(32'hbb2b7264),
	.w5(32'hbbd2babc),
	.w6(32'h3bc261cc),
	.w7(32'hbbad3df6),
	.w8(32'h3bb87afd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7334f2),
	.w1(32'hbb8a8751),
	.w2(32'h3b0e0052),
	.w3(32'hbab32bb6),
	.w4(32'hbc807688),
	.w5(32'h3a2f4bda),
	.w6(32'hbb351687),
	.w7(32'hbb5fae02),
	.w8(32'hbb9cf1b7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcc819),
	.w1(32'hbc5fba49),
	.w2(32'h3baef033),
	.w3(32'hb9725d81),
	.w4(32'hbb7a7ddf),
	.w5(32'h3c2f1a06),
	.w6(32'hbaa8b190),
	.w7(32'hbad88ab8),
	.w8(32'hb80a6295),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83241b),
	.w1(32'hbab73133),
	.w2(32'hbc344bb0),
	.w3(32'h3b2542f1),
	.w4(32'hbc1612f3),
	.w5(32'h3cb4d0d9),
	.w6(32'hbbec82b8),
	.w7(32'hbb98ae62),
	.w8(32'h3bb766ec),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d569073),
	.w1(32'hbae04bbe),
	.w2(32'h3af1467b),
	.w3(32'h3c1f43e3),
	.w4(32'hbb1047a6),
	.w5(32'hba85ef2c),
	.w6(32'hba8e843c),
	.w7(32'h3aeb508c),
	.w8(32'hbbb7af08),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ba2f7),
	.w1(32'h39183be5),
	.w2(32'hbba5debd),
	.w3(32'hb90621b8),
	.w4(32'hbb488f54),
	.w5(32'hbbf87252),
	.w6(32'hbbd041a9),
	.w7(32'h39a67347),
	.w8(32'h3b49eb41),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b424bba),
	.w1(32'h3b7d62e9),
	.w2(32'hbb5413dd),
	.w3(32'h39a0057c),
	.w4(32'hbb9f6088),
	.w5(32'h3bef1896),
	.w6(32'hbb7457a8),
	.w7(32'hbb6968b0),
	.w8(32'hbbc78dc4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba454ab),
	.w1(32'hba9b4aa6),
	.w2(32'h3a2cbc9a),
	.w3(32'hbbc4578c),
	.w4(32'h3bffa4c1),
	.w5(32'h3b6b3f8f),
	.w6(32'hbbd63584),
	.w7(32'hbaa57269),
	.w8(32'h3a520352),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836cd19),
	.w1(32'hbb210fd4),
	.w2(32'h3b04eb41),
	.w3(32'h3bb4c57f),
	.w4(32'hbaee44f0),
	.w5(32'h38a0a956),
	.w6(32'hb9f38129),
	.w7(32'h38c35e84),
	.w8(32'hbb9acf75),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22fc3),
	.w1(32'h3906d562),
	.w2(32'hbc11ae3c),
	.w3(32'hbab37c7c),
	.w4(32'h3c37acd2),
	.w5(32'hb91ee6f3),
	.w6(32'hbbefb288),
	.w7(32'h3c366ac5),
	.w8(32'h38c13264),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf1bd6),
	.w1(32'hbb0bff94),
	.w2(32'h3816c85c),
	.w3(32'hbc31059a),
	.w4(32'hbb8f9bfc),
	.w5(32'h3b5b23c4),
	.w6(32'h3a5e10fc),
	.w7(32'h3bb4f0b8),
	.w8(32'h3c6151ec),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2d2f),
	.w1(32'h3d05fbde),
	.w2(32'hbb1bd8ae),
	.w3(32'hbb6e016a),
	.w4(32'hbb9665ab),
	.w5(32'h3c09d35b),
	.w6(32'hbc03f72f),
	.w7(32'h3ae30532),
	.w8(32'hbc7317f6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e162),
	.w1(32'h3b2e79c3),
	.w2(32'hbc280f4e),
	.w3(32'hbc58e474),
	.w4(32'hba21dad6),
	.w5(32'h3a32a803),
	.w6(32'h3bf8f587),
	.w7(32'h3bd3d5cd),
	.w8(32'hbb73c09a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82afb0),
	.w1(32'h3ad04f08),
	.w2(32'hbac2d59e),
	.w3(32'hbb4bba43),
	.w4(32'h3b12794f),
	.w5(32'hbb88ff0e),
	.w6(32'h3ae10f9b),
	.w7(32'h3bd2c989),
	.w8(32'hbbdf2b01),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07fea2),
	.w1(32'hbb68d990),
	.w2(32'h3ccb3a49),
	.w3(32'hbb59f89e),
	.w4(32'h39b7b374),
	.w5(32'h3a47f1d7),
	.w6(32'h3c4235b4),
	.w7(32'hbb5b8214),
	.w8(32'hba799388),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab993dd),
	.w1(32'hbacd018b),
	.w2(32'hba0730c5),
	.w3(32'h3bb256f0),
	.w4(32'h3c398762),
	.w5(32'hbb87192c),
	.w6(32'hbb36fa05),
	.w7(32'h3bf5980d),
	.w8(32'hbb97153c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1045e),
	.w1(32'h3aa5eab5),
	.w2(32'hbba15991),
	.w3(32'h3c2f8c6d),
	.w4(32'h3bcb659d),
	.w5(32'hbb8c407d),
	.w6(32'h3ba509ad),
	.w7(32'h398ed256),
	.w8(32'h3b0d3fbf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45b472),
	.w1(32'hbb956f0d),
	.w2(32'h3b7d7961),
	.w3(32'hba9020bd),
	.w4(32'hba9c439c),
	.w5(32'h3b9eb153),
	.w6(32'h3abc4e13),
	.w7(32'hbc2db008),
	.w8(32'hbb637ce2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b4217),
	.w1(32'h3ab06504),
	.w2(32'hba943c49),
	.w3(32'h3ac2e19b),
	.w4(32'hbbca3c39),
	.w5(32'hba96d8b5),
	.w6(32'h3c99e503),
	.w7(32'h3960b592),
	.w8(32'hbc5b8f71),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9da8),
	.w1(32'hbb1d36fc),
	.w2(32'hb9c4a413),
	.w3(32'h3bb0281e),
	.w4(32'hbb737d41),
	.w5(32'h3cf3c784),
	.w6(32'hbbc2497f),
	.w7(32'hbb5286ae),
	.w8(32'h3b021323),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6480b),
	.w1(32'h3a50c84a),
	.w2(32'hbb800378),
	.w3(32'h3bfbb4ed),
	.w4(32'hbba93e90),
	.w5(32'hbb7e542b),
	.w6(32'hbb2aa188),
	.w7(32'hbbbc7e95),
	.w8(32'h3b42bea7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa67e),
	.w1(32'h3c69aeaf),
	.w2(32'h3b59dd24),
	.w3(32'h3bef433f),
	.w4(32'hbc298298),
	.w5(32'h3c113ae8),
	.w6(32'hbb6bf8b3),
	.w7(32'h3a8766c6),
	.w8(32'hbc0f9279),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b6c7),
	.w1(32'h3be29d1a),
	.w2(32'hb9b453cd),
	.w3(32'hba348052),
	.w4(32'hbbc98db5),
	.w5(32'h39abc9c4),
	.w6(32'hbb33c47d),
	.w7(32'h3cb5ab11),
	.w8(32'h3af5636b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c6a95),
	.w1(32'h3b01f68f),
	.w2(32'hbad23ef7),
	.w3(32'h3ab5c9cd),
	.w4(32'hba91f7c4),
	.w5(32'h364cacd2),
	.w6(32'h3bbbe50b),
	.w7(32'hbc4f08a5),
	.w8(32'hbbc63044),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf54052),
	.w1(32'h3b608ef4),
	.w2(32'hbbc353dc),
	.w3(32'h3d1bf575),
	.w4(32'hbc02385d),
	.w5(32'h3bde80a2),
	.w6(32'hb6c397aa),
	.w7(32'h390eda29),
	.w8(32'h3b86bd4f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75aebf),
	.w1(32'h3b9f438d),
	.w2(32'hbb3b04c3),
	.w3(32'h3b3d0fc2),
	.w4(32'hbc0362f7),
	.w5(32'hbb7b5433),
	.w6(32'h3be77287),
	.w7(32'hbacc16d8),
	.w8(32'h3b4c9d7a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cda85),
	.w1(32'h3c485deb),
	.w2(32'h384ac8a6),
	.w3(32'hbb5be10f),
	.w4(32'hb8045606),
	.w5(32'h3b299a8e),
	.w6(32'hbb0ba526),
	.w7(32'h3a563911),
	.w8(32'hbbbbd4d1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba453277),
	.w1(32'hbba7344c),
	.w2(32'h3b8d9383),
	.w3(32'hbb5d54a2),
	.w4(32'hbc08de07),
	.w5(32'h3aaa29a0),
	.w6(32'h3ac688b8),
	.w7(32'hbb2301d1),
	.w8(32'h3bd9f273),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91668f),
	.w1(32'h3ab8f7e0),
	.w2(32'hbb7dfc18),
	.w3(32'hbc110311),
	.w4(32'hbb6f87f4),
	.w5(32'hbbbd9278),
	.w6(32'h3bb52dfd),
	.w7(32'hbbf0d31c),
	.w8(32'hbabf3f0e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c224),
	.w1(32'h398ef52f),
	.w2(32'h3b9a96d3),
	.w3(32'hba88d5e4),
	.w4(32'hbc02bef9),
	.w5(32'h3a0c08dd),
	.w6(32'hbb1a9554),
	.w7(32'hbba4c994),
	.w8(32'hbc07917c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36cece),
	.w1(32'hbb03362f),
	.w2(32'h3a9ae0c5),
	.w3(32'h3b8a0520),
	.w4(32'h3b2f7c30),
	.w5(32'h3a930bd6),
	.w6(32'hbaf74922),
	.w7(32'hbc088943),
	.w8(32'h3b9d6099),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae96934),
	.w1(32'hb5494981),
	.w2(32'hbb093838),
	.w3(32'h3a7c3478),
	.w4(32'h3bc14874),
	.w5(32'hbb29ca73),
	.w6(32'h3a53524e),
	.w7(32'h3bc6f732),
	.w8(32'hbb805c8c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5538),
	.w1(32'hbb85cc5c),
	.w2(32'h3a103dc5),
	.w3(32'h3c1d4fce),
	.w4(32'h3b47da99),
	.w5(32'hb940af17),
	.w6(32'h3c4c1b91),
	.w7(32'h3c20704d),
	.w8(32'h3bf3fbd2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388869aa),
	.w1(32'h3bb7fe28),
	.w2(32'h3b386228),
	.w3(32'h3a9ad4a5),
	.w4(32'hbbcf96c8),
	.w5(32'hbb103b16),
	.w6(32'hbb4ffc46),
	.w7(32'hbc47ea9c),
	.w8(32'hba74e6c2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72356c),
	.w1(32'hbc541332),
	.w2(32'hbbb5c209),
	.w3(32'hbb5b2ce2),
	.w4(32'h3a7ba6e1),
	.w5(32'hbb21e05b),
	.w6(32'hbb9a40ef),
	.w7(32'hbb937aee),
	.w8(32'h3bdf881d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3a677),
	.w1(32'hba7a96b8),
	.w2(32'hbb73b284),
	.w3(32'h3b637d29),
	.w4(32'h3b51b6e4),
	.w5(32'hbbbfadf7),
	.w6(32'hbadc032e),
	.w7(32'hbb2e05c3),
	.w8(32'hbbd2710e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca8fcc),
	.w1(32'hbae8f785),
	.w2(32'h3b50b001),
	.w3(32'hb93ad137),
	.w4(32'hb90ba12c),
	.w5(32'hbb57d6b3),
	.w6(32'hbc2fb981),
	.w7(32'hba5c827b),
	.w8(32'h3ae4b9e4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c3564),
	.w1(32'h3ac16a88),
	.w2(32'hbbf94164),
	.w3(32'h3b6ae8fe),
	.w4(32'h3b2ff1fc),
	.w5(32'h3c411c4e),
	.w6(32'h39bcd0d5),
	.w7(32'hbc0517db),
	.w8(32'hbb4f6295),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4b7b),
	.w1(32'hbaaba9e0),
	.w2(32'hbac22f34),
	.w3(32'hbb62eab9),
	.w4(32'h3c701086),
	.w5(32'h3a74c90c),
	.w6(32'h3ba26dc3),
	.w7(32'h3bc18fe7),
	.w8(32'hbba5ecf4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe61834),
	.w1(32'hbbb8dceb),
	.w2(32'h3ba5cef9),
	.w3(32'h3b892014),
	.w4(32'hbb166e03),
	.w5(32'h3c037070),
	.w6(32'hbb6896ef),
	.w7(32'h3af10fa5),
	.w8(32'hbc0b0129),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6108c0),
	.w1(32'hbcb532d2),
	.w2(32'hbacd2c5f),
	.w3(32'hbb87a083),
	.w4(32'hbb850dd5),
	.w5(32'h39214e71),
	.w6(32'hbc1e2a2c),
	.w7(32'hbb4954e8),
	.w8(32'hbb12638e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce53b7),
	.w1(32'hbbcfa02f),
	.w2(32'h3b5dad84),
	.w3(32'h3b0f516c),
	.w4(32'h39c1c376),
	.w5(32'hbb89ec96),
	.w6(32'h3c27863c),
	.w7(32'hbc046024),
	.w8(32'h3b85e690),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a530d),
	.w1(32'h3b8887b3),
	.w2(32'hbceebafe),
	.w3(32'h3ba0da53),
	.w4(32'h3b888b2c),
	.w5(32'hba50d236),
	.w6(32'h3af71202),
	.w7(32'hbb8db013),
	.w8(32'hbbaf5c8f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004ce2),
	.w1(32'hb97efaa4),
	.w2(32'hbb7b7e26),
	.w3(32'hbbadaf74),
	.w4(32'h3aeb8e74),
	.w5(32'h3a7cda1f),
	.w6(32'h3b8a22e0),
	.w7(32'h3d546744),
	.w8(32'hbb7e5c11),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc51d),
	.w1(32'h3d390844),
	.w2(32'h3b08bd77),
	.w3(32'hbc948e97),
	.w4(32'hbc1b584b),
	.w5(32'hbb491e19),
	.w6(32'hbb07b238),
	.w7(32'h3b8f9c7e),
	.w8(32'hbb9450ff),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20914d),
	.w1(32'hbb5fb797),
	.w2(32'hbad23966),
	.w3(32'h3b7675a4),
	.w4(32'hbbae8470),
	.w5(32'h3c519287),
	.w6(32'hba251849),
	.w7(32'hbc5a267c),
	.w8(32'hbc2af96c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb091d),
	.w1(32'h3b038a6c),
	.w2(32'hba0bf6b0),
	.w3(32'hbc007e81),
	.w4(32'h3b84f0e4),
	.w5(32'h3b2feb21),
	.w6(32'hbb88b96c),
	.w7(32'hbb52da59),
	.w8(32'hbc2fe9c6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef5709),
	.w1(32'h3aad4b22),
	.w2(32'hbc05d242),
	.w3(32'h3bfc17aa),
	.w4(32'h3a36c187),
	.w5(32'hb9d07fc8),
	.w6(32'h3b7fbc3f),
	.w7(32'h3af53d92),
	.w8(32'hbbd5ee61),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4319d),
	.w1(32'hbb68903f),
	.w2(32'hbb58218b),
	.w3(32'hba90190f),
	.w4(32'hbafaee86),
	.w5(32'h3b8f078a),
	.w6(32'h3b92dec3),
	.w7(32'h3c20cc9b),
	.w8(32'h3b55b117),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030a7f),
	.w1(32'hbad039d4),
	.w2(32'hbb967aac),
	.w3(32'hbb2f7ae2),
	.w4(32'hbba8c238),
	.w5(32'hbbbc59ce),
	.w6(32'hbb5fe527),
	.w7(32'h3b075905),
	.w8(32'h3b8c5bfd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e651ce),
	.w1(32'h3b6311ff),
	.w2(32'hbb8306ef),
	.w3(32'h3bd28c52),
	.w4(32'hba9db1be),
	.w5(32'h3a171a34),
	.w6(32'hbc98208d),
	.w7(32'h3ab06139),
	.w8(32'hbb82cf7b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6e016),
	.w1(32'h3c4cb86d),
	.w2(32'hbc4c7b82),
	.w3(32'hbb53fb45),
	.w4(32'hbc44aec6),
	.w5(32'hbbb0d35c),
	.w6(32'hbbc3cabb),
	.w7(32'hbb017f10),
	.w8(32'hbb00e761),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21263b),
	.w1(32'h3c779ce4),
	.w2(32'h399f2394),
	.w3(32'h3bc51623),
	.w4(32'hb97efec0),
	.w5(32'h3bac5356),
	.w6(32'hb8df8bc7),
	.w7(32'h3bb490df),
	.w8(32'h3b1bb730),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59b3d),
	.w1(32'hbb9967ec),
	.w2(32'h3aea1023),
	.w3(32'h3b6536d8),
	.w4(32'hba4b9230),
	.w5(32'hbc8d6064),
	.w6(32'hbbc236ec),
	.w7(32'hbba553ef),
	.w8(32'hbbb77428),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a850c9f),
	.w1(32'h3d381348),
	.w2(32'h3a95348c),
	.w3(32'h3d4740fa),
	.w4(32'hbc0c4f58),
	.w5(32'h39e52f99),
	.w6(32'hb8ac7dc4),
	.w7(32'hbb21516d),
	.w8(32'h385b672b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d54dd),
	.w1(32'hbbfeb6d1),
	.w2(32'h3b81f20f),
	.w3(32'h39e969c9),
	.w4(32'hbae365d9),
	.w5(32'h3b0ec946),
	.w6(32'hbbd4e268),
	.w7(32'hbb3b8204),
	.w8(32'h3ac5af43),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba785c89),
	.w1(32'hbc03840c),
	.w2(32'hba9b328a),
	.w3(32'hbabf7bef),
	.w4(32'h3b66d32d),
	.w5(32'hbc7030ed),
	.w6(32'h3b4045ba),
	.w7(32'hbbf4b8e4),
	.w8(32'hbd292baf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05623b),
	.w1(32'h3b2b1bfe),
	.w2(32'hbaedc817),
	.w3(32'h3a07cdc5),
	.w4(32'h3b4c2e92),
	.w5(32'h3bbd2bc1),
	.w6(32'hbc183fe7),
	.w7(32'h3b56d497),
	.w8(32'h3b99c76b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aaa43),
	.w1(32'hbae8ca82),
	.w2(32'h3b2f1782),
	.w3(32'hbbb380c4),
	.w4(32'h3ba317e5),
	.w5(32'hbaaa1676),
	.w6(32'h3b0a4df4),
	.w7(32'hbb9e27d9),
	.w8(32'h3b74dde3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2dc65),
	.w1(32'hbb955c4e),
	.w2(32'hbcd244be),
	.w3(32'hba392bc8),
	.w4(32'hbaf42c4b),
	.w5(32'h3918647b),
	.w6(32'hbc56798a),
	.w7(32'h3a2b7053),
	.w8(32'hbbc35f0e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f827),
	.w1(32'h3b9692e4),
	.w2(32'h3d265186),
	.w3(32'h3c9e31e6),
	.w4(32'h3bcad623),
	.w5(32'hbab8230b),
	.w6(32'hbbad2685),
	.w7(32'hb9c3e220),
	.w8(32'h3c818262),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d36b888),
	.w1(32'hbbb38779),
	.w2(32'h3d023638),
	.w3(32'h39004eca),
	.w4(32'h3b0de0e6),
	.w5(32'h3a33696b),
	.w6(32'hbb01f114),
	.w7(32'hba5d6687),
	.w8(32'h3add5c70),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eeb26),
	.w1(32'h3d4a9541),
	.w2(32'h3a8eb80a),
	.w3(32'h3c15b08e),
	.w4(32'hbb300cf4),
	.w5(32'hbc7ce3b3),
	.w6(32'h3b56bd50),
	.w7(32'h3b345bce),
	.w8(32'h3ba908da),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c180),
	.w1(32'h3b127504),
	.w2(32'hbbeba6c2),
	.w3(32'hbba6e901),
	.w4(32'h3b1a7736),
	.w5(32'hbb1f7bf9),
	.w6(32'hbb4f3b44),
	.w7(32'h3c070a41),
	.w8(32'hb8637ad0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1466dc),
	.w1(32'hbbe611fd),
	.w2(32'h3b339b13),
	.w3(32'h3b973de2),
	.w4(32'hbaacd26f),
	.w5(32'hbab5f2d6),
	.w6(32'h3b8e42e8),
	.w7(32'hba0b8d70),
	.w8(32'h399f899f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3cb11),
	.w1(32'hbc1475b5),
	.w2(32'h37bed2c6),
	.w3(32'hbb2dc674),
	.w4(32'hbb02a805),
	.w5(32'hba859afe),
	.w6(32'h37833849),
	.w7(32'hbb7f7ecd),
	.w8(32'hbb5c66e5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b9b885),
	.w1(32'h3901c12e),
	.w2(32'h3bbc6041),
	.w3(32'h3c97c8e4),
	.w4(32'hbbb46bc5),
	.w5(32'h3a4f2084),
	.w6(32'h3aed17aa),
	.w7(32'hbb4de537),
	.w8(32'h3bd03f37),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1423c9),
	.w1(32'h3a25e874),
	.w2(32'hbc6a74d1),
	.w3(32'hbbb051ea),
	.w4(32'h3a53b3a6),
	.w5(32'h39114d50),
	.w6(32'hbabbe8c8),
	.w7(32'h3b682f25),
	.w8(32'hbb9a952d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f68e),
	.w1(32'hbbd41995),
	.w2(32'hbb09473a),
	.w3(32'hbb77e832),
	.w4(32'h3b308b83),
	.w5(32'h3c9ba228),
	.w6(32'hbb76bc3a),
	.w7(32'hbc676831),
	.w8(32'hbaeae943),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76c8b8),
	.w1(32'h3be302d1),
	.w2(32'hbb633328),
	.w3(32'hba7191bf),
	.w4(32'h3b95f3cf),
	.w5(32'h3b80b863),
	.w6(32'h3bb31d02),
	.w7(32'hbb85bcc7),
	.w8(32'hbb6c4fde),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f448c),
	.w1(32'hbace5a8f),
	.w2(32'h3a460d0e),
	.w3(32'h3b19dd0f),
	.w4(32'h37e144fe),
	.w5(32'hbbc08b35),
	.w6(32'h3bd41b24),
	.w7(32'h3871aea2),
	.w8(32'hbbc0c18f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeac37),
	.w1(32'hbb1df67c),
	.w2(32'h3b615334),
	.w3(32'h3c2a7422),
	.w4(32'hbb2003ca),
	.w5(32'h37945af5),
	.w6(32'h3a4852ac),
	.w7(32'h3b502fdd),
	.w8(32'h3b2d8ba4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba110e86),
	.w1(32'hba5ac964),
	.w2(32'hba30cac7),
	.w3(32'h3b362273),
	.w4(32'h3b4eecdc),
	.w5(32'hbc01b6ce),
	.w6(32'h3aa8d2ea),
	.w7(32'hbae1defd),
	.w8(32'hbb83bbf5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c3c26),
	.w1(32'h3b3703f5),
	.w2(32'hbb32aea9),
	.w3(32'hbad013ca),
	.w4(32'h3aa29af9),
	.w5(32'hbb85d9d5),
	.w6(32'h3b2eca6f),
	.w7(32'h3b34804f),
	.w8(32'hbb8178ab),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f257),
	.w1(32'hbb395f8d),
	.w2(32'h3b50af69),
	.w3(32'h3a5b6c64),
	.w4(32'hbb96b753),
	.w5(32'hb9c25e94),
	.w6(32'h3b633e02),
	.w7(32'hbbb4750b),
	.w8(32'h3b9d8b1b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ce4e0),
	.w1(32'h3adb261c),
	.w2(32'h3b878fe1),
	.w3(32'h3b72e9aa),
	.w4(32'hbb0fb0fb),
	.w5(32'h3a15495d),
	.w6(32'h3acf1927),
	.w7(32'hbb7c5576),
	.w8(32'h3b125b5c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39940880),
	.w1(32'h3b26806f),
	.w2(32'h3b6c0897),
	.w3(32'h3ab31333),
	.w4(32'h3b0fa904),
	.w5(32'hba305167),
	.w6(32'hbb377e1d),
	.w7(32'h38dece17),
	.w8(32'hba2f6774),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a809c62),
	.w1(32'hbb111c5a),
	.w2(32'hba3bdfdf),
	.w3(32'hba874c82),
	.w4(32'hbaa332d8),
	.w5(32'h3ae393a1),
	.w6(32'h3a57c124),
	.w7(32'h3a9eef07),
	.w8(32'hbbf86dc5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e9ff9),
	.w1(32'h3aa056a5),
	.w2(32'h3afb2cb1),
	.w3(32'hbb9a5f8e),
	.w4(32'hbaaa607b),
	.w5(32'hbb9dd215),
	.w6(32'hbbbc83a5),
	.w7(32'h3c869f39),
	.w8(32'h3b637da1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b550b5e),
	.w1(32'hbaff6cfa),
	.w2(32'h3b72e95f),
	.w3(32'h39c4d0ed),
	.w4(32'hbb2870b2),
	.w5(32'hbb429503),
	.w6(32'h3a89a632),
	.w7(32'h3ac675d2),
	.w8(32'hbbd20d73),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f46f4),
	.w1(32'hbb99a403),
	.w2(32'h36d8211e),
	.w3(32'h3bfa2386),
	.w4(32'h3bcf28bf),
	.w5(32'h3c2e6c8e),
	.w6(32'h3a06865e),
	.w7(32'h3bd52d16),
	.w8(32'h38aa11c5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed9c6e),
	.w1(32'hbbee2ce5),
	.w2(32'hbb913d97),
	.w3(32'h384f2fe2),
	.w4(32'hbaf620c7),
	.w5(32'hbb577502),
	.w6(32'h3b1ce493),
	.w7(32'h3b80f452),
	.w8(32'hba565e88),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85453f),
	.w1(32'h3aac2e02),
	.w2(32'hbb1b5242),
	.w3(32'hba81fd1b),
	.w4(32'h3ab3f71c),
	.w5(32'hbaa9a91f),
	.w6(32'hbb571fb3),
	.w7(32'h3b46b577),
	.w8(32'hba4ab36c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a817cbd),
	.w1(32'hb30d7c4c),
	.w2(32'h3a13e36c),
	.w3(32'hbab8461e),
	.w4(32'h3c1db952),
	.w5(32'h3bad90ca),
	.w6(32'h3bfe3162),
	.w7(32'h38468549),
	.w8(32'h3adc0739),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a630bc3),
	.w1(32'hba9fa4de),
	.w2(32'h3aef6ae1),
	.w3(32'h3a7676b4),
	.w4(32'hbba1503c),
	.w5(32'h3cae03f8),
	.w6(32'hba874962),
	.w7(32'hba9e032a),
	.w8(32'h3b9e7cf3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875d47),
	.w1(32'h383c7d47),
	.w2(32'h3ba76e8f),
	.w3(32'h3b1edce2),
	.w4(32'hbb8d58f2),
	.w5(32'h3bd60d2e),
	.w6(32'hbc74e5f9),
	.w7(32'h3a8bd140),
	.w8(32'h3bbac4e8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf303),
	.w1(32'h3b52638e),
	.w2(32'h3ab11412),
	.w3(32'h3be9c3a3),
	.w4(32'hbb7a57a9),
	.w5(32'hb5b5bdfc),
	.w6(32'h3aa1691a),
	.w7(32'hbb716dd5),
	.w8(32'h3c403fde),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6569),
	.w1(32'h39e77c1c),
	.w2(32'h3c3f7636),
	.w3(32'h3976a511),
	.w4(32'hba992485),
	.w5(32'h39db61ec),
	.w6(32'hb995631e),
	.w7(32'hba1a6cfb),
	.w8(32'hba2dbf71),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb3b1),
	.w1(32'hbb33fc6a),
	.w2(32'hbabc8345),
	.w3(32'h3be6d4ed),
	.w4(32'h3ae476a0),
	.w5(32'hbb7798b0),
	.w6(32'h3794f177),
	.w7(32'hbc070dd7),
	.w8(32'h3ab9c82a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb741215),
	.w1(32'h3bb5a4a9),
	.w2(32'hbad7ea9c),
	.w3(32'hbb4eb9b3),
	.w4(32'h3aa1392f),
	.w5(32'h3c316be0),
	.w6(32'h3a076304),
	.w7(32'h39b1974a),
	.w8(32'h39d19c7a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2966b0),
	.w1(32'h3b099a16),
	.w2(32'hbb09a51f),
	.w3(32'h3ad9be63),
	.w4(32'h3b1ab247),
	.w5(32'h3b0448e4),
	.w6(32'hbb2def4a),
	.w7(32'h3a3d4747),
	.w8(32'h36a61a61),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9671d),
	.w1(32'hbaae29d0),
	.w2(32'hb9420cdb),
	.w3(32'hbb2587e2),
	.w4(32'hba50b3a3),
	.w5(32'hbb88a85c),
	.w6(32'h3b2b943a),
	.w7(32'h3aaff5ea),
	.w8(32'hbafd81a8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd332ea),
	.w1(32'h3a23e642),
	.w2(32'hbb28e86a),
	.w3(32'h3bde385f),
	.w4(32'hbba356ac),
	.w5(32'hb9e6f09d),
	.w6(32'hb8067f51),
	.w7(32'hb9ae27b6),
	.w8(32'hba2fd8b2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9adeb0),
	.w1(32'hb895ed75),
	.w2(32'h3ad1c7ac),
	.w3(32'hbb9d43ce),
	.w4(32'hbb750d97),
	.w5(32'h3983875e),
	.w6(32'hb9edf5cf),
	.w7(32'hb8359fae),
	.w8(32'h3bdef985),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4db2c5),
	.w1(32'h3a3a762d),
	.w2(32'h3bc4ed92),
	.w3(32'hb86453f5),
	.w4(32'hbbbf28fc),
	.w5(32'hbabaae47),
	.w6(32'h3a5058f0),
	.w7(32'hbc242a16),
	.w8(32'h3b35210e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9707b32),
	.w1(32'hb9b53d3a),
	.w2(32'h39e8a45c),
	.w3(32'hbb583490),
	.w4(32'h3a78d79e),
	.w5(32'h3a733013),
	.w6(32'hb9028f8b),
	.w7(32'h3b442a5e),
	.w8(32'h3b2435e9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98269c9),
	.w1(32'h3ac71a57),
	.w2(32'hbb8d2d70),
	.w3(32'h3ad49494),
	.w4(32'h3b7bb034),
	.w5(32'hb88cbedc),
	.w6(32'h3ba9c2e6),
	.w7(32'hbac82d0f),
	.w8(32'h3ba5b768),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9763e),
	.w1(32'hb9bbab29),
	.w2(32'hbadded93),
	.w3(32'h3ba0d8a9),
	.w4(32'hbbeef642),
	.w5(32'h3be18956),
	.w6(32'hbc09f4da),
	.w7(32'h3a899819),
	.w8(32'hba801a70),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacebfa5),
	.w1(32'hb99ab27d),
	.w2(32'h3b59cb62),
	.w3(32'h3b136a3c),
	.w4(32'hba876e7f),
	.w5(32'hbc1ecdd5),
	.w6(32'hb9e2b9f0),
	.w7(32'h3ba5a19b),
	.w8(32'h3b304325),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcfb5a),
	.w1(32'hbbc1339a),
	.w2(32'hba24fed2),
	.w3(32'hbb560e7d),
	.w4(32'hbc2b9c32),
	.w5(32'hbae2d268),
	.w6(32'hba686b4e),
	.w7(32'hbc5fc8d0),
	.w8(32'hb985c6e5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa56907),
	.w1(32'hbb1137e0),
	.w2(32'hb9a4c948),
	.w3(32'h3aee903c),
	.w4(32'h3cf2af76),
	.w5(32'h3c0971c6),
	.w6(32'h3b399f06),
	.w7(32'hbb88191f),
	.w8(32'hb6e218a4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfa689),
	.w1(32'h3a3a3c1b),
	.w2(32'hbba312b3),
	.w3(32'hb9ae117a),
	.w4(32'h388de10b),
	.w5(32'hbaad3df4),
	.w6(32'h3d0e0002),
	.w7(32'hbb40fcef),
	.w8(32'hba702e69),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf9620),
	.w1(32'hb9eed509),
	.w2(32'h3bac26a1),
	.w3(32'hb906d408),
	.w4(32'hbcc6e498),
	.w5(32'hbae1afff),
	.w6(32'hbb039f7f),
	.w7(32'hbba487f0),
	.w8(32'h3be44c34),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5111),
	.w1(32'hbb2d05aa),
	.w2(32'hb9190667),
	.w3(32'hbaa84d9f),
	.w4(32'hbb486586),
	.w5(32'hbb789890),
	.w6(32'h3c0474d0),
	.w7(32'h3bc4bac8),
	.w8(32'h3ad7d5e6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95ddf2),
	.w1(32'hbc24d4cf),
	.w2(32'hbacdb456),
	.w3(32'hbbc4c527),
	.w4(32'h39f22488),
	.w5(32'h3b873d4f),
	.w6(32'h3b07e5ce),
	.w7(32'hba642290),
	.w8(32'h3b9d93dd),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8efffb5),
	.w1(32'h3b7dea9e),
	.w2(32'h3b4b9e80),
	.w3(32'hbcc1b8d6),
	.w4(32'h3c0a6764),
	.w5(32'hbad9630b),
	.w6(32'h3bc622eb),
	.w7(32'hbb5a029d),
	.w8(32'h3a91e6ea),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44fe2d),
	.w1(32'hba9337b5),
	.w2(32'h3c15a0c7),
	.w3(32'hbaaeb990),
	.w4(32'hbb9ba5fb),
	.w5(32'hbb8803cc),
	.w6(32'hbaa425f1),
	.w7(32'h3a95bac2),
	.w8(32'h3b53d58d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39d1d6),
	.w1(32'hbaa80a46),
	.w2(32'hbafeba28),
	.w3(32'hbc3f6b5c),
	.w4(32'hba007132),
	.w5(32'hbb89cca6),
	.w6(32'hb93a94ff),
	.w7(32'h3ba18beb),
	.w8(32'h3b88c0f4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394cf34a),
	.w1(32'h3af4cacf),
	.w2(32'h3b4c8967),
	.w3(32'hbb55664d),
	.w4(32'hbb8d9ef5),
	.w5(32'hb9827630),
	.w6(32'h3c17aeb7),
	.w7(32'hbc2e29b8),
	.w8(32'h3b7bedcc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba042e63),
	.w1(32'hb8e66ce5),
	.w2(32'hbb18499e),
	.w3(32'hb62c4045),
	.w4(32'hbbf208e6),
	.w5(32'h3b3fdb78),
	.w6(32'h3cdbd6be),
	.w7(32'h3791d12b),
	.w8(32'hbb8280b2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d43b),
	.w1(32'h3b2cecff),
	.w2(32'hbccf20d5),
	.w3(32'h3b8d0dfb),
	.w4(32'h38952f6b),
	.w5(32'hbb36b6d7),
	.w6(32'hbb061f0b),
	.w7(32'hbb2fbd6a),
	.w8(32'h3b593b1a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce8c980),
	.w1(32'hba8a2106),
	.w2(32'h3bfd7c44),
	.w3(32'hba807dc1),
	.w4(32'hba88d561),
	.w5(32'h38356428),
	.w6(32'h3ced8e4e),
	.w7(32'hbaa62e9e),
	.w8(32'h3c7266bb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27b20),
	.w1(32'h3b2af0e0),
	.w2(32'h3b1925b6),
	.w3(32'hbac2f18f),
	.w4(32'hbb7e36d8),
	.w5(32'hbaf3c0ad),
	.w6(32'h3b983bbb),
	.w7(32'h3948a6a8),
	.w8(32'h3a119148),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbefd3),
	.w1(32'h392c5c18),
	.w2(32'hbca6d270),
	.w3(32'hba8531fc),
	.w4(32'hbbf17c12),
	.w5(32'hbd029715),
	.w6(32'hbb58d495),
	.w7(32'h3b35a2c9),
	.w8(32'h3a8f59c9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b41e61),
	.w1(32'hba17cb9c),
	.w2(32'h3a61d864),
	.w3(32'hbb547b9f),
	.w4(32'hba00e599),
	.w5(32'h3b636f5d),
	.w6(32'hbbad2daf),
	.w7(32'h3bde5527),
	.w8(32'h3b8ae8be),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11a0e),
	.w1(32'h3c165a8d),
	.w2(32'hbb79e05e),
	.w3(32'h3b15dbe3),
	.w4(32'hbbcd7baa),
	.w5(32'h39996442),
	.w6(32'hba9af672),
	.w7(32'h3b0c45c3),
	.w8(32'hbb9d78ad),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f61bb),
	.w1(32'h3abde983),
	.w2(32'hb74a7011),
	.w3(32'hbc9438a1),
	.w4(32'h3a1fe8af),
	.w5(32'h3a75a03a),
	.w6(32'h3ba3d5ef),
	.w7(32'hbc1432e3),
	.w8(32'hbb7382d5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe8950),
	.w1(32'h396846fc),
	.w2(32'h3b5761e3),
	.w3(32'hbb6a6617),
	.w4(32'h3b0f20be),
	.w5(32'hbc9a6b27),
	.w6(32'hbabec93e),
	.w7(32'h3d065c95),
	.w8(32'h3ca2d5c4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a331990),
	.w1(32'hbb7cc81d),
	.w2(32'hbb2d35c2),
	.w3(32'hbb9359b0),
	.w4(32'h3a909340),
	.w5(32'h3c11a983),
	.w6(32'h3afcf067),
	.w7(32'h3d182719),
	.w8(32'hbb06a2a0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00f099),
	.w1(32'hba8a8792),
	.w2(32'h3c40a367),
	.w3(32'hba4e3abf),
	.w4(32'hba664383),
	.w5(32'hbb813362),
	.w6(32'h3d0db595),
	.w7(32'h3c00337d),
	.w8(32'hbbcf09b8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399475e7),
	.w1(32'h3b95a08e),
	.w2(32'h3b1edbbb),
	.w3(32'hbb8b4e65),
	.w4(32'h3ba1df03),
	.w5(32'hbb0fcc22),
	.w6(32'hbaed1a1a),
	.w7(32'h3afd7c2b),
	.w8(32'h3c104312),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb393646),
	.w1(32'hba52d456),
	.w2(32'h3aeaeb9f),
	.w3(32'hbb89ce63),
	.w4(32'hb980cb17),
	.w5(32'h38d941a4),
	.w6(32'h3a93f57c),
	.w7(32'h3bc7b577),
	.w8(32'h3ad9f5ce),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9428480),
	.w1(32'h3a7ed2c7),
	.w2(32'hbae81430),
	.w3(32'hbb7d3fbf),
	.w4(32'hbb30b7f8),
	.w5(32'hbad08420),
	.w6(32'hb74a443c),
	.w7(32'hb9d2802f),
	.w8(32'hbc4463dc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0b007),
	.w1(32'h3b83629a),
	.w2(32'hba7c48f2),
	.w3(32'hbb28acb2),
	.w4(32'h3b423e0f),
	.w5(32'hba9ac187),
	.w6(32'hbbbc1c32),
	.w7(32'h3a787dc0),
	.w8(32'hbacbda10),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99df20),
	.w1(32'hb9a3a863),
	.w2(32'h3b0ad742),
	.w3(32'h3b073a51),
	.w4(32'h3a89eb7a),
	.w5(32'h3b09f27c),
	.w6(32'hb9d331c7),
	.w7(32'hbb9d2aa1),
	.w8(32'h3ba15374),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46789c),
	.w1(32'hbc02e1c7),
	.w2(32'h3bf9b429),
	.w3(32'hbb7c582b),
	.w4(32'hbc9f6bcb),
	.w5(32'h3adc1c64),
	.w6(32'h3b8fcdff),
	.w7(32'hbb55ff7a),
	.w8(32'h3bcaeae2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25cad9),
	.w1(32'h3b492f64),
	.w2(32'h3b01b532),
	.w3(32'hbb177bf4),
	.w4(32'hba9f1c40),
	.w5(32'h3ae59aa2),
	.w6(32'hbb026cff),
	.w7(32'hbb89d1ef),
	.w8(32'hbbbae8ac),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6e446),
	.w1(32'h3b2ab114),
	.w2(32'hbab10736),
	.w3(32'h3b6b143a),
	.w4(32'h39fa6927),
	.w5(32'h3c9bc552),
	.w6(32'hbbc6ba30),
	.w7(32'h3ad17d22),
	.w8(32'hbbae2de1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc847815),
	.w1(32'h3a80b73e),
	.w2(32'h3a1a2d78),
	.w3(32'hbad8e964),
	.w4(32'hbbcb1650),
	.w5(32'hbb829aae),
	.w6(32'hb890d558),
	.w7(32'h38dba2cc),
	.w8(32'h3ccb099f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b377dfb),
	.w1(32'h3afb5d96),
	.w2(32'h3d157274),
	.w3(32'h3b695767),
	.w4(32'h3b1e6409),
	.w5(32'h39e8b3bc),
	.w6(32'hbaa03744),
	.w7(32'h3b9191c3),
	.w8(32'hba860754),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32c04a),
	.w1(32'hbae7781e),
	.w2(32'h3b92e6ab),
	.w3(32'hbb351a54),
	.w4(32'hba01d273),
	.w5(32'h3b93cd61),
	.w6(32'hbb807bff),
	.w7(32'h3a71a6ec),
	.w8(32'h3b3a393f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a270777),
	.w1(32'hba810487),
	.w2(32'h3ae815a2),
	.w3(32'h3c3606dd),
	.w4(32'h3b8ab7f7),
	.w5(32'hbb1c0bed),
	.w6(32'hbb8853de),
	.w7(32'hbb6438c3),
	.w8(32'hbb217345),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f6e0),
	.w1(32'hbb8de19b),
	.w2(32'h39e34b8e),
	.w3(32'h3b522f08),
	.w4(32'hbb3bf5bc),
	.w5(32'hbb98d0ea),
	.w6(32'hba4b9b60),
	.w7(32'h3afaeed0),
	.w8(32'h3a9e3dbb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8a924),
	.w1(32'hbaef061f),
	.w2(32'hba631ba1),
	.w3(32'hb914d570),
	.w4(32'h3998b12e),
	.w5(32'hbb98c8c4),
	.w6(32'hbab4dece),
	.w7(32'h3a218340),
	.w8(32'h3c3e303d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa99f11),
	.w1(32'hb8601607),
	.w2(32'h3a3bad84),
	.w3(32'h3a0a03d4),
	.w4(32'h3b905cfc),
	.w5(32'h3aa5ee65),
	.w6(32'hba2a16e7),
	.w7(32'h38f1f3c6),
	.w8(32'h3bb56fe5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79348),
	.w1(32'hbbe545d0),
	.w2(32'h3bd86bea),
	.w3(32'hbaaa667c),
	.w4(32'hbbbd2100),
	.w5(32'h39a41f89),
	.w6(32'hbaafe66e),
	.w7(32'h3b3eea7d),
	.w8(32'hbbe3c66e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b21c5),
	.w1(32'h3c427815),
	.w2(32'h3c267233),
	.w3(32'hb994eda6),
	.w4(32'hbac65784),
	.w5(32'h3ba2f182),
	.w6(32'hbadadae0),
	.w7(32'hb8cdf477),
	.w8(32'hbbd9dd32),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc924b58),
	.w1(32'h3c3d056a),
	.w2(32'hbafae0bb),
	.w3(32'h3bdb758d),
	.w4(32'hb990689b),
	.w5(32'h3c000c02),
	.w6(32'hba401631),
	.w7(32'hb7f8bf81),
	.w8(32'hb9e7106d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3761a229),
	.w1(32'h3b3e3049),
	.w2(32'h3b9d1f5b),
	.w3(32'h3b01ce21),
	.w4(32'hbb9ea22c),
	.w5(32'h3b271f94),
	.w6(32'h3c0d2f68),
	.w7(32'h3c181bd8),
	.w8(32'h3b667662),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d09b8),
	.w1(32'hbba7f747),
	.w2(32'h3ca94281),
	.w3(32'hbabdfca4),
	.w4(32'h3c9a6ef2),
	.w5(32'h3b14c290),
	.w6(32'hba4f0d2c),
	.w7(32'hbb2dda92),
	.w8(32'h3a85c51e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c6af8),
	.w1(32'hbac18124),
	.w2(32'hbb2847f2),
	.w3(32'h39f4bea9),
	.w4(32'hb928325c),
	.w5(32'hba9c94c6),
	.w6(32'hb72671d8),
	.w7(32'h3ac6826a),
	.w8(32'hbb15e71d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587b73),
	.w1(32'h3ab7d2e9),
	.w2(32'hbce09a50),
	.w3(32'h382a112e),
	.w4(32'h3badd294),
	.w5(32'hbb980f57),
	.w6(32'h3bceef4e),
	.w7(32'hbb29154a),
	.w8(32'h3b6420b7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc841e8),
	.w1(32'h39cf1942),
	.w2(32'hbb64f95f),
	.w3(32'h3c321d18),
	.w4(32'hb9f6f40f),
	.w5(32'hbb1bdeb6),
	.w6(32'hbcbe38b2),
	.w7(32'h3b2be83e),
	.w8(32'h3bec8969),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4382b),
	.w1(32'h3b02626a),
	.w2(32'h3b0ec14d),
	.w3(32'h3b376c50),
	.w4(32'h38cad33b),
	.w5(32'hbca807e5),
	.w6(32'hbb6d09a2),
	.w7(32'hbbb319dc),
	.w8(32'h3b119bc8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf24864),
	.w1(32'h37935770),
	.w2(32'h3b214359),
	.w3(32'h3953f5b6),
	.w4(32'h3b0fb765),
	.w5(32'h3a9a11d5),
	.w6(32'hbb48522f),
	.w7(32'hbc9d300b),
	.w8(32'h37fe5a6c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87d87d),
	.w1(32'h3b13d4d9),
	.w2(32'hba945d78),
	.w3(32'hb8e7b522),
	.w4(32'h3c63965c),
	.w5(32'hbb67dc9e),
	.w6(32'h3a9554e7),
	.w7(32'hbb8887de),
	.w8(32'hba79ba1b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3a6e7),
	.w1(32'h3cab80e6),
	.w2(32'h3ba7d2f5),
	.w3(32'h3b0746dd),
	.w4(32'h39fd0a4e),
	.w5(32'hbba5bc21),
	.w6(32'hbbabe662),
	.w7(32'hbaa671aa),
	.w8(32'h3845ad82),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3abd2d),
	.w1(32'hba05c2db),
	.w2(32'h3c92d0fe),
	.w3(32'h3b4dd8d2),
	.w4(32'hbbcf182b),
	.w5(32'h3a31d00d),
	.w6(32'hbb81538d),
	.w7(32'hb902d0e9),
	.w8(32'hbac412c8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf00745),
	.w1(32'hb9ac3a7f),
	.w2(32'hbb339320),
	.w3(32'h3a3c784a),
	.w4(32'h3b1a360e),
	.w5(32'h39e9bc24),
	.w6(32'hbb2d8290),
	.w7(32'hba916376),
	.w8(32'hbc8502f9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cadd),
	.w1(32'hbb6dae7c),
	.w2(32'hbb1b3b65),
	.w3(32'hbadf3c72),
	.w4(32'hb8a512a4),
	.w5(32'h3a0a9f45),
	.w6(32'hba93e16e),
	.w7(32'hb9652517),
	.w8(32'h3a569006),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad09141),
	.w1(32'h3b2a65ff),
	.w2(32'hb9cb47d5),
	.w3(32'h3b247ffd),
	.w4(32'hbb030dbd),
	.w5(32'h3b8f53cc),
	.w6(32'h38f20518),
	.w7(32'hbb1b4c88),
	.w8(32'h3ad19597),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e81b7a),
	.w1(32'hba8ca0ef),
	.w2(32'h396fa4c5),
	.w3(32'hbb92a5bd),
	.w4(32'h38b75695),
	.w5(32'hba9a5517),
	.w6(32'h3a0135e2),
	.w7(32'hbabe78e5),
	.w8(32'hbbddd5b5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffc796),
	.w1(32'h3ab06d8d),
	.w2(32'hbace751e),
	.w3(32'h39d47d9b),
	.w4(32'hbb459537),
	.w5(32'hbaf921bc),
	.w6(32'h38c126ec),
	.w7(32'h3a37ca32),
	.w8(32'h384d0b4b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0096),
	.w1(32'h3bc2514a),
	.w2(32'h3c1c6e74),
	.w3(32'h3b85237b),
	.w4(32'hb9e439b1),
	.w5(32'h3a385e08),
	.w6(32'h3b1c309f),
	.w7(32'hb9c379eb),
	.w8(32'hbbb12f2d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33e088),
	.w1(32'h3b009ba4),
	.w2(32'hbac2404d),
	.w3(32'hbba4f3dc),
	.w4(32'h3b2e8930),
	.w5(32'h39efc8b5),
	.w6(32'h3b6d1b5e),
	.w7(32'hbb0e1ea3),
	.w8(32'h3bb4c46d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01260b),
	.w1(32'hba850ba3),
	.w2(32'hba4d6040),
	.w3(32'hba91e968),
	.w4(32'h3b221f2f),
	.w5(32'h3aac2a7d),
	.w6(32'hba8e1d7d),
	.w7(32'hbaa120b6),
	.w8(32'h3ae360fc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29dca),
	.w1(32'h3b1ac146),
	.w2(32'h3aaca6db),
	.w3(32'hbbb4f820),
	.w4(32'h3cb1594e),
	.w5(32'hbba94394),
	.w6(32'hbc495e5c),
	.w7(32'hbaaf13c3),
	.w8(32'h3acd3560),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86a7f8),
	.w1(32'hbc6c353f),
	.w2(32'h3b120b67),
	.w3(32'h3aa0d6ff),
	.w4(32'hb9097766),
	.w5(32'hbb1c198f),
	.w6(32'hbad390c1),
	.w7(32'h3b3ccb10),
	.w8(32'hb9d465dd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b457e67),
	.w1(32'hbaa32b39),
	.w2(32'hb89cb252),
	.w3(32'hbc22a852),
	.w4(32'hbaa648c5),
	.w5(32'h3b09e25f),
	.w6(32'h3b6fcd47),
	.w7(32'hbad3f9f7),
	.w8(32'h3ab71e29),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae2a1d),
	.w1(32'hbafee429),
	.w2(32'hb80f6156),
	.w3(32'h3a083282),
	.w4(32'h3aa30485),
	.w5(32'h3b8d8e06),
	.w6(32'h3936818a),
	.w7(32'h3b207844),
	.w8(32'h3a31b294),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba815eaf),
	.w1(32'h39b9c46e),
	.w2(32'h3b454870),
	.w3(32'hb9bf7284),
	.w4(32'h39b7871a),
	.w5(32'h3a1eec38),
	.w6(32'h3aa30596),
	.w7(32'h3adef059),
	.w8(32'h3a8ece64),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35def),
	.w1(32'h3a881996),
	.w2(32'hbbb22349),
	.w3(32'h3b2f9e65),
	.w4(32'h3b40b199),
	.w5(32'h3b905bc9),
	.w6(32'hb9f84dca),
	.w7(32'hbaae70d3),
	.w8(32'hb997905f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36622208),
	.w1(32'hbb33257b),
	.w2(32'hbae1cfd3),
	.w3(32'hbb05018e),
	.w4(32'hbb1fd1c1),
	.w5(32'h3b372b8b),
	.w6(32'h3b2ba1f9),
	.w7(32'h3a43d6e0),
	.w8(32'h3a1ea591),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac56752),
	.w1(32'hba9b6263),
	.w2(32'hbb9054bb),
	.w3(32'hb952139d),
	.w4(32'h399149b2),
	.w5(32'h39698957),
	.w6(32'h3b329d5c),
	.w7(32'hbc1291bd),
	.w8(32'h3cd85371),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986e2f9),
	.w1(32'h3ac95305),
	.w2(32'h3a8cfd29),
	.w3(32'hbbb9069b),
	.w4(32'hba1a422a),
	.w5(32'hbbd8edbd),
	.w6(32'h3b2bdd14),
	.w7(32'hbb5cc2de),
	.w8(32'h3a16d6ac),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72607d),
	.w1(32'hbb483d1a),
	.w2(32'hba6bd1fc),
	.w3(32'hbbb5abf9),
	.w4(32'h3cb585c9),
	.w5(32'hbb05b951),
	.w6(32'hb9eecb38),
	.w7(32'h3a898ab1),
	.w8(32'hbb10e7fd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36544240),
	.w1(32'h3a4fd62e),
	.w2(32'hbc6f6e39),
	.w3(32'h3b0c37c7),
	.w4(32'hb8369f21),
	.w5(32'h39fbc472),
	.w6(32'hbaea0f16),
	.w7(32'hba884db0),
	.w8(32'h3a8b9641),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab030d4),
	.w1(32'hba3413dc),
	.w2(32'h3b786766),
	.w3(32'h3b4ff856),
	.w4(32'h38a0d769),
	.w5(32'h3a7fe529),
	.w6(32'h3a10ebe2),
	.w7(32'hbb13e87f),
	.w8(32'hbc947e49),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90919c),
	.w1(32'h3ac9f911),
	.w2(32'h351eabef),
	.w3(32'hbc2979f8),
	.w4(32'hb9f7b253),
	.w5(32'h3b4208d7),
	.w6(32'hb981c46e),
	.w7(32'hbada7133),
	.w8(32'h38126e40),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33d09a),
	.w1(32'h39eb9321),
	.w2(32'h3b64a9f0),
	.w3(32'h3998dd5a),
	.w4(32'h3a9b2281),
	.w5(32'h3b414c01),
	.w6(32'h3a341081),
	.w7(32'hb955406c),
	.w8(32'h3b955b5f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dec24e),
	.w1(32'h3b786877),
	.w2(32'h3c1c414f),
	.w3(32'h3d090f5e),
	.w4(32'hbb19eadc),
	.w5(32'hbb35a85b),
	.w6(32'hbad2fc5a),
	.w7(32'hbbff2dfe),
	.w8(32'hb9b62f8e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b493b),
	.w1(32'hbae011ec),
	.w2(32'hba2115c5),
	.w3(32'hba6ddf51),
	.w4(32'h3a872caf),
	.w5(32'h3a95271a),
	.w6(32'hba88663a),
	.w7(32'h3ae2d57c),
	.w8(32'h3ba9480f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa10a),
	.w1(32'h3b03c702),
	.w2(32'hba1bb5ca),
	.w3(32'h3a45f39c),
	.w4(32'h3950af62),
	.w5(32'hba74e76e),
	.w6(32'h3ca431d8),
	.w7(32'h3a3b8d5b),
	.w8(32'h37a1fcb6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caea5dc),
	.w1(32'h3b55919b),
	.w2(32'h399528c1),
	.w3(32'h38a60d6d),
	.w4(32'h3cd7dc9d),
	.w5(32'h3a563885),
	.w6(32'hbad4d385),
	.w7(32'hb6487858),
	.w8(32'hbc820d24),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a675094),
	.w1(32'hbb143de0),
	.w2(32'hb92b5bb3),
	.w3(32'hbb1cdd29),
	.w4(32'hbc81d8f2),
	.w5(32'hbc3a3e09),
	.w6(32'h3aa4fac8),
	.w7(32'hbad2c213),
	.w8(32'h39abf81c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde919),
	.w1(32'hb9fbc4bd),
	.w2(32'hbb6c413a),
	.w3(32'h3b9562ff),
	.w4(32'hbbf47aa2),
	.w5(32'h3ac782b2),
	.w6(32'h3ae96e43),
	.w7(32'h39a8228b),
	.w8(32'h3babd94b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54d5fd),
	.w1(32'h3b4b59ad),
	.w2(32'h3a6ed57b),
	.w3(32'hbbd490c7),
	.w4(32'h3b12b331),
	.w5(32'hbb475526),
	.w6(32'h395a7ada),
	.w7(32'hbb521132),
	.w8(32'h3a67434c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae19c54),
	.w1(32'h3be60cb5),
	.w2(32'h3a4bc434),
	.w3(32'hba9c26da),
	.w4(32'h3a5a4c65),
	.w5(32'hb9a4ee4d),
	.w6(32'h3b21b963),
	.w7(32'hbadb9c43),
	.w8(32'hb9c7016f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1abe63),
	.w1(32'h39c2a03a),
	.w2(32'hb937a50a),
	.w3(32'hbbc5979c),
	.w4(32'h3b62aad9),
	.w5(32'h3af6a16f),
	.w6(32'h3a019c72),
	.w7(32'hbabe0cc9),
	.w8(32'hb9f899b4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8bc1),
	.w1(32'hbaabdb87),
	.w2(32'h3ac82fff),
	.w3(32'h3a3d0c2d),
	.w4(32'h388cd9fd),
	.w5(32'hbbe8495e),
	.w6(32'h3abbb082),
	.w7(32'hbad52d2e),
	.w8(32'hbc02c292),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20fc2c),
	.w1(32'h39f68d77),
	.w2(32'h3a16dba2),
	.w3(32'hbaf8f897),
	.w4(32'hbbb3e080),
	.w5(32'hbae66f53),
	.w6(32'h3ac8a92e),
	.w7(32'hb9392688),
	.w8(32'h3aaa935f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4632),
	.w1(32'hb9f73534),
	.w2(32'h3b3ebeb3),
	.w3(32'h3a60d80c),
	.w4(32'h391f3a86),
	.w5(32'h3aabdc14),
	.w6(32'h3aa41287),
	.w7(32'h3b079eb1),
	.w8(32'h3ad95a00),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5595f),
	.w1(32'hbb54d3a4),
	.w2(32'hbac7f07f),
	.w3(32'h398fd50c),
	.w4(32'hbbba1114),
	.w5(32'h3b5d76ff),
	.w6(32'h3b738c6a),
	.w7(32'hbc00decb),
	.w8(32'h3a83fc99),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7bc56),
	.w1(32'h3ae58635),
	.w2(32'hb888dee3),
	.w3(32'hbbd0fea9),
	.w4(32'h3ace92d2),
	.w5(32'h3a04d2b7),
	.w6(32'h3ba406eb),
	.w7(32'h3b756679),
	.w8(32'h3ad80e7c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2cd57),
	.w1(32'hba797a96),
	.w2(32'h3b0336f5),
	.w3(32'hbac3c753),
	.w4(32'hbb93b756),
	.w5(32'hbaa44e45),
	.w6(32'hb995901c),
	.w7(32'hbb5f3ed6),
	.w8(32'hbc1a46ef),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6951c),
	.w1(32'hbae86600),
	.w2(32'hba6dfe0a),
	.w3(32'hb8cbb33b),
	.w4(32'hb9e78c4a),
	.w5(32'h3c9bd26c),
	.w6(32'hbb3da789),
	.w7(32'h3b5e6176),
	.w8(32'hba3e9e9c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca7145),
	.w1(32'hba3a3f69),
	.w2(32'h3b8ff559),
	.w3(32'h3bc3250c),
	.w4(32'h3b16caab),
	.w5(32'h39f7a9fc),
	.w6(32'h3a6ecb8c),
	.w7(32'h3cb4af3a),
	.w8(32'h3b33a34e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fbfd1f),
	.w1(32'hbb5ce153),
	.w2(32'hb814155b),
	.w3(32'hbb2235df),
	.w4(32'h3abb6b96),
	.w5(32'hbb70a98d),
	.w6(32'hba41bc55),
	.w7(32'h39929e6f),
	.w8(32'hbae86158),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917bb75),
	.w1(32'hbb3d0c51),
	.w2(32'hbba0fb29),
	.w3(32'hba5da23e),
	.w4(32'hbb96ea26),
	.w5(32'hb80aaf0d),
	.w6(32'h3931bb87),
	.w7(32'h3ab1cf9b),
	.w8(32'h3b23e2a2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4dfcf),
	.w1(32'hb905c864),
	.w2(32'hbb3b3885),
	.w3(32'h3b63f43d),
	.w4(32'h3b08f687),
	.w5(32'h3aa27ecd),
	.w6(32'hb96b50b0),
	.w7(32'hbb04b0fe),
	.w8(32'hba9ac48f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d2fb),
	.w1(32'hba227619),
	.w2(32'h3b8d4bf4),
	.w3(32'hbbabee31),
	.w4(32'hbbde41eb),
	.w5(32'h3b0bd627),
	.w6(32'h3b1539e4),
	.w7(32'h3add2125),
	.w8(32'hbac17c6e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266840),
	.w1(32'h3ac3deef),
	.w2(32'h3b75b056),
	.w3(32'h39c73a95),
	.w4(32'hba9dc18e),
	.w5(32'h3a2aa352),
	.w6(32'hb9be0e1e),
	.w7(32'hb9c74bdc),
	.w8(32'h3b4455a2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5ac1e),
	.w1(32'hbabfe176),
	.w2(32'hbb8c7857),
	.w3(32'hbb78d963),
	.w4(32'hbbcbfbd0),
	.w5(32'hba1b87ba),
	.w6(32'hbb9e9e3d),
	.w7(32'hbb5350bc),
	.w8(32'h3b1a3d7f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa270),
	.w1(32'hbaa6afc3),
	.w2(32'hba232bed),
	.w3(32'hbb7b62f5),
	.w4(32'h3a5db197),
	.w5(32'hbb69c681),
	.w6(32'h3b9f42fa),
	.w7(32'h3ba4c661),
	.w8(32'hbbaed37c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93a36e),
	.w1(32'hba9c9da3),
	.w2(32'h39ccdeb1),
	.w3(32'hb8763f41),
	.w4(32'hb6cf9801),
	.w5(32'h3b1531bb),
	.w6(32'h3a170f84),
	.w7(32'h3b88fbd1),
	.w8(32'h38a4ca66),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a977af5),
	.w1(32'hbb1488e3),
	.w2(32'hbbedac64),
	.w3(32'h3b6c4c28),
	.w4(32'h39c628e7),
	.w5(32'hbaebf9a9),
	.w6(32'h3b8b64b3),
	.w7(32'h3bf57996),
	.w8(32'h3aa247a7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc345fd0),
	.w1(32'h3ca01e1f),
	.w2(32'hba85ba4b),
	.w3(32'hbaebc658),
	.w4(32'hba3b94f5),
	.w5(32'hba8df768),
	.w6(32'h3aa1da89),
	.w7(32'h3c655ede),
	.w8(32'h3b07d68a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa045),
	.w1(32'h38922e44),
	.w2(32'hbb68360b),
	.w3(32'hb85f30f2),
	.w4(32'hbb0ae292),
	.w5(32'hbb10ab5e),
	.w6(32'hbb432b09),
	.w7(32'h394d17ce),
	.w8(32'hbabe5034),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07798),
	.w1(32'h3b0aa3ba),
	.w2(32'h39d1fbdb),
	.w3(32'h3a99583f),
	.w4(32'hba215eae),
	.w5(32'h3af60766),
	.w6(32'h3b3a0ec1),
	.w7(32'hbc2da4ef),
	.w8(32'hbbc68571),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1e12f),
	.w1(32'h3b05a653),
	.w2(32'hbae87743),
	.w3(32'hbc933e35),
	.w4(32'h3aaa160f),
	.w5(32'h39ac1641),
	.w6(32'hbac7a83d),
	.w7(32'hbb5ef52b),
	.w8(32'hbb28f3d0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a35ed),
	.w1(32'hba0bd0f5),
	.w2(32'hbb7df939),
	.w3(32'hbb83c466),
	.w4(32'hb8db57ab),
	.w5(32'h3a1a270b),
	.w6(32'h3a2a02bf),
	.w7(32'hbb64825f),
	.w8(32'h398037d2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf3a75),
	.w1(32'h3b06937a),
	.w2(32'hb965f128),
	.w3(32'hbaba22e6),
	.w4(32'hbc69aacc),
	.w5(32'h3aaf752b),
	.w6(32'h3a654e15),
	.w7(32'h3a8e42f8),
	.w8(32'hbc125637),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7025d01),
	.w1(32'h3afb2e5d),
	.w2(32'hbb105cf1),
	.w3(32'hbabebf37),
	.w4(32'hba47854f),
	.w5(32'hbb1932ff),
	.w6(32'h3bc619d2),
	.w7(32'hbb0a92c4),
	.w8(32'h3cc7c1f1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1440ca),
	.w1(32'hb85f2f0d),
	.w2(32'hbb75075f),
	.w3(32'hbbc20c01),
	.w4(32'hb98c390d),
	.w5(32'hbad7c26e),
	.w6(32'h3c2cd880),
	.w7(32'hba932339),
	.w8(32'h3c364074),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba756c95),
	.w1(32'h3b984aed),
	.w2(32'h39897605),
	.w3(32'h39bd924a),
	.w4(32'hba407ee4),
	.w5(32'hbb0cf884),
	.w6(32'hb920e2a0),
	.w7(32'h3c9c19e2),
	.w8(32'h3ac9afa1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f3a1),
	.w1(32'hba6214dd),
	.w2(32'h3bab9610),
	.w3(32'h3a30d70b),
	.w4(32'hbb272df7),
	.w5(32'hbade560b),
	.w6(32'hbb5c2070),
	.w7(32'hbb5ebe51),
	.w8(32'h3ac9f866),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf64dbb),
	.w1(32'hbb320722),
	.w2(32'h376f1782),
	.w3(32'hbab0adfb),
	.w4(32'hba57ffbc),
	.w5(32'hba1c5116),
	.w6(32'h3bb79f42),
	.w7(32'hbb46f5f6),
	.w8(32'h3ab08fec),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f46f),
	.w1(32'hb94df33f),
	.w2(32'h3aa9598e),
	.w3(32'h389d370d),
	.w4(32'h3a0b533c),
	.w5(32'hba5c5ff1),
	.w6(32'h3a047f41),
	.w7(32'h3a1623ad),
	.w8(32'hb8c13902),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e25aa),
	.w1(32'hba226feb),
	.w2(32'h3a1acf98),
	.w3(32'hba068835),
	.w4(32'hbb233901),
	.w5(32'hb9072f25),
	.w6(32'hbac86270),
	.w7(32'hbb41cbc9),
	.w8(32'h39a21b07),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaecdc3),
	.w1(32'h3aa29dde),
	.w2(32'h3b32affd),
	.w3(32'h3ae82dba),
	.w4(32'hb99a653f),
	.w5(32'h3a8db43c),
	.w6(32'hbb4d34fc),
	.w7(32'hb836d4b4),
	.w8(32'hbb340394),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21784),
	.w1(32'hba48d4e5),
	.w2(32'h3a6b9147),
	.w3(32'h361e45cc),
	.w4(32'hbabea66e),
	.w5(32'hbbf79c4b),
	.w6(32'hba33d636),
	.w7(32'h3a5a272d),
	.w8(32'hbb78c145),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24eed1),
	.w1(32'hb9f49776),
	.w2(32'h3ae9f254),
	.w3(32'hba78b164),
	.w4(32'hba8db732),
	.w5(32'h3a0dc588),
	.w6(32'hba9ea9da),
	.w7(32'h3aa4c228),
	.w8(32'hbaa540d2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96a751),
	.w1(32'hbadb3089),
	.w2(32'hb93feaf0),
	.w3(32'h37f443eb),
	.w4(32'h3bcf5750),
	.w5(32'h3b158bb9),
	.w6(32'hb8de7f45),
	.w7(32'h3bb9e842),
	.w8(32'h3c83b402),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981648f),
	.w1(32'h3c2a2847),
	.w2(32'h3cd569e1),
	.w3(32'hbb49f428),
	.w4(32'h3bcaa7ed),
	.w5(32'h389f84eb),
	.w6(32'hbb2eb01d),
	.w7(32'hba4c760d),
	.w8(32'h3b53318b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule