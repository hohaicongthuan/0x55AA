module layer_10_featuremap_192(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf11540),
	.w1(32'hbb8d4e77),
	.w2(32'hbbc4b986),
	.w3(32'hbac22e37),
	.w4(32'hbad6a7f8),
	.w5(32'hbbac3827),
	.w6(32'hbbb1a6d8),
	.w7(32'hbbc45846),
	.w8(32'hbbd81db4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb689ca0),
	.w1(32'h3a82d6d1),
	.w2(32'h3bafa253),
	.w3(32'hbb9a70f3),
	.w4(32'hba60da97),
	.w5(32'h3afde4cd),
	.w6(32'h3abbab12),
	.w7(32'h3b9ea9c2),
	.w8(32'h3b0b6792),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac04e9),
	.w1(32'hbacf89ae),
	.w2(32'h3a668232),
	.w3(32'hbab7c8e9),
	.w4(32'hbb5b7d2b),
	.w5(32'hbb508b47),
	.w6(32'hbb0103cd),
	.w7(32'h3b323c59),
	.w8(32'h39b9c072),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade05e0),
	.w1(32'h3b3634f1),
	.w2(32'h3b8fe3cf),
	.w3(32'hbb871f18),
	.w4(32'h3b9ecadf),
	.w5(32'h3bfc9faf),
	.w6(32'hba333dd1),
	.w7(32'hbb2fda22),
	.w8(32'hbac0821e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cf6a2),
	.w1(32'h3ad69de3),
	.w2(32'h3bbf2a4d),
	.w3(32'h3c270430),
	.w4(32'hbb5b257a),
	.w5(32'h3b2ebdfe),
	.w6(32'h3af96d0b),
	.w7(32'h3ae48694),
	.w8(32'hbaf21f51),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec361),
	.w1(32'hbbaac6bb),
	.w2(32'hbbe52832),
	.w3(32'h392fa9ce),
	.w4(32'hbb8c4fc9),
	.w5(32'hbbb57304),
	.w6(32'hbbb1a098),
	.w7(32'hbbf38313),
	.w8(32'hbbd74805),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d6b5),
	.w1(32'h3b8fa8d9),
	.w2(32'h3c2f76c7),
	.w3(32'hbb702966),
	.w4(32'h39d6cdb9),
	.w5(32'h3b498782),
	.w6(32'h3b712375),
	.w7(32'h3c09577a),
	.w8(32'h3b107622),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2f310),
	.w1(32'h38bda054),
	.w2(32'hbb08d822),
	.w3(32'hb884dfa4),
	.w4(32'h390e270e),
	.w5(32'hba568ae0),
	.w6(32'h3b038ab1),
	.w7(32'h3a339ac7),
	.w8(32'h3b0b3f32),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad63328),
	.w1(32'hbb09ffbd),
	.w2(32'hbb4652d4),
	.w3(32'h3b18acf5),
	.w4(32'hbad3c3ba),
	.w5(32'hbb17d07c),
	.w6(32'hbb4ca62e),
	.w7(32'hbb3207c7),
	.w8(32'hbaf1c59f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd07f5e),
	.w1(32'hbade5502),
	.w2(32'hbad6c0ff),
	.w3(32'hbb952da8),
	.w4(32'hbad1334e),
	.w5(32'hbaacf391),
	.w6(32'hbb2bfd59),
	.w7(32'hba01451b),
	.w8(32'hbb0f3508),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17301d),
	.w1(32'hbac95e29),
	.w2(32'hbb4fcb9d),
	.w3(32'hbb1ce6c1),
	.w4(32'h3a56f2cd),
	.w5(32'h3a2fefe3),
	.w6(32'hbb1b39a0),
	.w7(32'hbb8cb484),
	.w8(32'hbb92f3fb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ba7a),
	.w1(32'h3bb7ae95),
	.w2(32'h3c03a830),
	.w3(32'hbad29326),
	.w4(32'h3b8a7e01),
	.w5(32'h3c177690),
	.w6(32'h39082aa1),
	.w7(32'h393856f6),
	.w8(32'h3b1fe30b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae64e8c),
	.w1(32'hbbbf6a57),
	.w2(32'hbc0d564b),
	.w3(32'h3baeb542),
	.w4(32'hbb9b1f38),
	.w5(32'hbbc605dc),
	.w6(32'hbbdc3a10),
	.w7(32'hbbe223cf),
	.w8(32'hbbcf2485),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b57d),
	.w1(32'h3ad418cc),
	.w2(32'hbb7b9445),
	.w3(32'h395a81d2),
	.w4(32'h3b950d03),
	.w5(32'hb96ae8e2),
	.w6(32'h3bda7fff),
	.w7(32'h3a2573b9),
	.w8(32'h3bb37697),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ea06),
	.w1(32'h39fa48d6),
	.w2(32'h3bf0efcb),
	.w3(32'h3b639fb0),
	.w4(32'hbbda26e2),
	.w5(32'h3bf3103d),
	.w6(32'hbaaedd16),
	.w7(32'hbb5c2027),
	.w8(32'hbaf7d494),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a9e3f),
	.w1(32'hbbe10be0),
	.w2(32'hbc191c44),
	.w3(32'h3ba1e752),
	.w4(32'hbbaf3e67),
	.w5(32'hbbf34b7e),
	.w6(32'hbbe68055),
	.w7(32'hbbd9664e),
	.w8(32'hbbe3e311),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b562a),
	.w1(32'h3b8fd230),
	.w2(32'h3b61585c),
	.w3(32'hbba5448f),
	.w4(32'h3ae19b8a),
	.w5(32'h3a253c8d),
	.w6(32'h3bb8e53c),
	.w7(32'h3bbf402f),
	.w8(32'h3b1c8ea5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176bd7),
	.w1(32'h3afe9bfb),
	.w2(32'h3b349651),
	.w3(32'hbb107c87),
	.w4(32'h3a82b89b),
	.w5(32'h3a5c68c1),
	.w6(32'h3a473e2d),
	.w7(32'h3bb2b5dd),
	.w8(32'h3a813453),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f9d0),
	.w1(32'hbb4eeef0),
	.w2(32'hbb8b4ea2),
	.w3(32'h3ac7a3ff),
	.w4(32'hbb4137d7),
	.w5(32'hbb58c681),
	.w6(32'hbac82cd0),
	.w7(32'hb9b98e07),
	.w8(32'hbb92aa3a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa17436),
	.w1(32'hba9c22a2),
	.w2(32'hbb2b28a5),
	.w3(32'hbabe763c),
	.w4(32'hba93c8a6),
	.w5(32'hbb167ee8),
	.w6(32'hbaad2d2d),
	.w7(32'hbb32fd88),
	.w8(32'hbb1ca58f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14558c),
	.w1(32'hba713c56),
	.w2(32'hba892861),
	.w3(32'hbb063ce9),
	.w4(32'hba029cbd),
	.w5(32'hba5c5076),
	.w6(32'hb9a4c6b7),
	.w7(32'hba1bb075),
	.w8(32'h3b099d23),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a609558),
	.w1(32'hbb4f9f1b),
	.w2(32'hbbc9d4ed),
	.w3(32'h3a4e1ddb),
	.w4(32'hbb106de9),
	.w5(32'hbb91a833),
	.w6(32'hbbbaf2fd),
	.w7(32'h3a3619cd),
	.w8(32'hbb88742a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2286ba),
	.w1(32'hbab3a9b3),
	.w2(32'hbacf1e6a),
	.w3(32'hbb228cfd),
	.w4(32'h3ac75b0b),
	.w5(32'h3b33abce),
	.w6(32'hba5dbebc),
	.w7(32'h38ed8723),
	.w8(32'h3b321ec2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0684),
	.w1(32'hba9c9bae),
	.w2(32'hbb3079ca),
	.w3(32'h3a117cc4),
	.w4(32'h3ad0f6c3),
	.w5(32'h3650754e),
	.w6(32'hba6afab6),
	.w7(32'hb86d8d18),
	.w8(32'h3aee457b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79004),
	.w1(32'hbbe319fa),
	.w2(32'hbbce38ed),
	.w3(32'hb9e66918),
	.w4(32'hbbaea889),
	.w5(32'hbb96a10c),
	.w6(32'hbc03d9b3),
	.w7(32'hbb93d69a),
	.w8(32'hbb8ae957),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd77e),
	.w1(32'hbaaa2235),
	.w2(32'hba812068),
	.w3(32'hbbd8f6a8),
	.w4(32'hbb6a3c7d),
	.w5(32'hbaf0a99d),
	.w6(32'h3b4a2f8e),
	.w7(32'h3a687311),
	.w8(32'h3a27b192),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f4074),
	.w1(32'hbad186a0),
	.w2(32'hbb2a9023),
	.w3(32'hba81027e),
	.w4(32'hbad36dec),
	.w5(32'hbb1dfb9f),
	.w6(32'hbab8da1e),
	.w7(32'hbb265b09),
	.w8(32'hba53579c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9594648),
	.w1(32'hbb378cf7),
	.w2(32'hbba866ec),
	.w3(32'hba8d7b7c),
	.w4(32'hbb5a44da),
	.w5(32'hbb7d1662),
	.w6(32'hbb87f369),
	.w7(32'hbba7b7ce),
	.w8(32'hbb8f4625),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a1e8),
	.w1(32'hbb6a3f5e),
	.w2(32'hbbd338fa),
	.w3(32'hbc08eef0),
	.w4(32'hbb00186e),
	.w5(32'hbb97d233),
	.w6(32'hbbe4f28d),
	.w7(32'hbbe2bb95),
	.w8(32'h38a546b7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba358d),
	.w1(32'h3acc1cd5),
	.w2(32'h3b04ec69),
	.w3(32'hbb317b0c),
	.w4(32'h3a588c1d),
	.w5(32'h3afeed24),
	.w6(32'h3a89a267),
	.w7(32'h3b26df8e),
	.w8(32'h3a29d3f9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22edba),
	.w1(32'hbab8e24f),
	.w2(32'hbade8753),
	.w3(32'h3a9fbd07),
	.w4(32'hba5728c0),
	.w5(32'hbaa776e0),
	.w6(32'hbaa59910),
	.w7(32'hbac2abb4),
	.w8(32'h3a270beb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14fb2f),
	.w1(32'hbb550a78),
	.w2(32'hbb6d5df8),
	.w3(32'h3a2a2d11),
	.w4(32'hbb41b729),
	.w5(32'hbb49ea03),
	.w6(32'hbb54a541),
	.w7(32'hbb6485cd),
	.w8(32'hbae8468e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cc425),
	.w1(32'h3974a05c),
	.w2(32'hba3cb4c5),
	.w3(32'hbac56d27),
	.w4(32'h3b27eb72),
	.w5(32'h3b034b05),
	.w6(32'h3a563c28),
	.w7(32'hb9394d69),
	.w8(32'h38c48f7c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8cad),
	.w1(32'hbb83c69b),
	.w2(32'hbbc67566),
	.w3(32'hbb9da779),
	.w4(32'hbb8b2504),
	.w5(32'hbb7e29a0),
	.w6(32'hbb7e8ee1),
	.w7(32'hbbb6f484),
	.w8(32'hbae1bc83),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44af2a),
	.w1(32'h3949dd63),
	.w2(32'h3b911d4b),
	.w3(32'hbb3b1d0d),
	.w4(32'hbb1308d6),
	.w5(32'h3a9b3b6e),
	.w6(32'hba62efdb),
	.w7(32'h3adcdbdb),
	.w8(32'h3a80c617),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac63a9c),
	.w1(32'hbb6c0566),
	.w2(32'hbb96f147),
	.w3(32'hba6e0e84),
	.w4(32'hbb6f4b5d),
	.w5(32'hbb9b3f5a),
	.w6(32'hbb1177d1),
	.w7(32'hbb439965),
	.w8(32'hbabf32df),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd33d85),
	.w1(32'h3abc92ed),
	.w2(32'h3bb9ef90),
	.w3(32'hbb8b3e16),
	.w4(32'hbb103edc),
	.w5(32'h3b4c3727),
	.w6(32'hbb53ecaa),
	.w7(32'h3b7c769e),
	.w8(32'h3a591d6b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc044a11),
	.w1(32'h3bad29af),
	.w2(32'h3c6e1b86),
	.w3(32'hbc096e3a),
	.w4(32'h3b4852c3),
	.w5(32'h3c383d5a),
	.w6(32'hbbc1bf5c),
	.w7(32'h3bc3f33d),
	.w8(32'h3c04defa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd6b67),
	.w1(32'h3a985f03),
	.w2(32'h3c0cc2ca),
	.w3(32'hbc1ab258),
	.w4(32'h3ad98c86),
	.w5(32'h3c04f33a),
	.w6(32'hbc25d1ef),
	.w7(32'hba6a95f5),
	.w8(32'h3bce2ee2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e15ed),
	.w1(32'h3a09a011),
	.w2(32'h3b8fee30),
	.w3(32'hba07a89e),
	.w4(32'hbb2278a8),
	.w5(32'h3a9003b4),
	.w6(32'hba25de10),
	.w7(32'h3b39ed67),
	.w8(32'h3a54cb9f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b8cf),
	.w1(32'h3aa86d73),
	.w2(32'h3b1c9ce8),
	.w3(32'hb93bae87),
	.w4(32'h3a6a7beb),
	.w5(32'h3b103c31),
	.w6(32'h3b020f5a),
	.w7(32'h3b32725a),
	.w8(32'h3a4b37fe),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5321b8),
	.w1(32'h3b873d30),
	.w2(32'h3c073fc6),
	.w3(32'h3a4bef40),
	.w4(32'hbb33547e),
	.w5(32'hb79caf9f),
	.w6(32'h3baf5b45),
	.w7(32'h3bcd2788),
	.w8(32'h3b44030e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59e5ff),
	.w1(32'hbb13c16a),
	.w2(32'hbb3a4c84),
	.w3(32'hbb6bd231),
	.w4(32'hbafbda15),
	.w5(32'hbb00931f),
	.w6(32'hbb34c170),
	.w7(32'hbb49e609),
	.w8(32'hba5d384b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4618f),
	.w1(32'h3b91f00e),
	.w2(32'h39e336fd),
	.w3(32'hbbaf824e),
	.w4(32'h3b5efb74),
	.w5(32'hba862d6f),
	.w6(32'h3b8dc442),
	.w7(32'h3ba06fce),
	.w8(32'h3a927148),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9281d2c),
	.w1(32'h3ab58b69),
	.w2(32'h3a256f24),
	.w3(32'hb9878239),
	.w4(32'h3b2f4751),
	.w5(32'hbadee91a),
	.w6(32'h3ac5fbc4),
	.w7(32'h3bc3acaa),
	.w8(32'h3bf89ce8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9a9e8),
	.w1(32'hbbdec03a),
	.w2(32'hbb64ad46),
	.w3(32'hbb953fb2),
	.w4(32'hbbe90a9d),
	.w5(32'hbbdd67d8),
	.w6(32'hbc203a59),
	.w7(32'hb98fd928),
	.w8(32'hbb88875e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124f63),
	.w1(32'h3bd1397f),
	.w2(32'h3c5f04f9),
	.w3(32'hbc04eed0),
	.w4(32'h3b88d5fd),
	.w5(32'h3c829096),
	.w6(32'h3a4dfc97),
	.w7(32'h3abaa29d),
	.w8(32'h3b3ad5d0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65429d),
	.w1(32'hbba90485),
	.w2(32'hbc4d5f00),
	.w3(32'h3c8e1fdc),
	.w4(32'hba920534),
	.w5(32'hbbd66e40),
	.w6(32'h3aa1b4a7),
	.w7(32'hbb84ab8e),
	.w8(32'hbbf779a4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f6df),
	.w1(32'hbb3e8e86),
	.w2(32'hbb748323),
	.w3(32'hb9db0f74),
	.w4(32'hbb18cf08),
	.w5(32'hbb337843),
	.w6(32'hbb349ee0),
	.w7(32'hbb6ad210),
	.w8(32'hbb19553c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a673),
	.w1(32'h3b237319),
	.w2(32'h3a78131c),
	.w3(32'hbaf508c4),
	.w4(32'h3b3f4f42),
	.w5(32'h3a9887d7),
	.w6(32'h3b5d3edc),
	.w7(32'h3b023bf4),
	.w8(32'h3b820481),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f911a),
	.w1(32'h3a0f4d29),
	.w2(32'h3b8efc54),
	.w3(32'h3b788133),
	.w4(32'hbb68a16d),
	.w5(32'hbb1b43cd),
	.w6(32'h398ee18e),
	.w7(32'h3b5ad7f8),
	.w8(32'h39f78da7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05555c),
	.w1(32'hbb872dc2),
	.w2(32'hbbe0d984),
	.w3(32'hbb87bebd),
	.w4(32'h3a973836),
	.w5(32'hbab97eeb),
	.w6(32'hbb6a9112),
	.w7(32'hbbec2fe7),
	.w8(32'hbb01c0fd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dbf82),
	.w1(32'hbbdd3193),
	.w2(32'hbbeefc9f),
	.w3(32'h3884e3b9),
	.w4(32'hbbc9021e),
	.w5(32'hbbe94da8),
	.w6(32'hbbd40ee3),
	.w7(32'hbbf1190f),
	.w8(32'hbbdfd6ec),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0ded),
	.w1(32'hbc0a3068),
	.w2(32'hbc459642),
	.w3(32'hbbfd20ab),
	.w4(32'hbc1ccbca),
	.w5(32'hbc241b77),
	.w6(32'hbc066512),
	.w7(32'hbbe240ba),
	.w8(32'hbc21e47c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0921ce),
	.w1(32'hbba020b0),
	.w2(32'hbb990e49),
	.w3(32'hbbf36c62),
	.w4(32'hbbb8eb55),
	.w5(32'hbb9a86c9),
	.w6(32'hbbb5c291),
	.w7(32'hbba84021),
	.w8(32'hbbc1d680),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe005),
	.w1(32'hba7d63b7),
	.w2(32'hbaaba814),
	.w3(32'hbbd20440),
	.w4(32'hba811da0),
	.w5(32'hbae82b62),
	.w6(32'hba1cae9a),
	.w7(32'hba24748e),
	.w8(32'hbaa2d995),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac934cd),
	.w1(32'h3c0d7e95),
	.w2(32'h3c4cbdf9),
	.w3(32'hba7bd037),
	.w4(32'h3b9830fa),
	.w5(32'h3bcf6934),
	.w6(32'h3bff0208),
	.w7(32'h3c40ddb9),
	.w8(32'h3c0bf62e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c182748),
	.w1(32'h3bb537d3),
	.w2(32'h3c16f27d),
	.w3(32'h3bc6b396),
	.w4(32'hbac48ce5),
	.w5(32'h3b7afd79),
	.w6(32'h3b410faa),
	.w7(32'h3bc2a867),
	.w8(32'hbae3ca37),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb738413),
	.w1(32'h3a3f2611),
	.w2(32'h3bbfaee7),
	.w3(32'h3a43ea71),
	.w4(32'hba923459),
	.w5(32'h3b032a58),
	.w6(32'hba788ff0),
	.w7(32'h3b30f416),
	.w8(32'h3af03b0d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed6c3d),
	.w1(32'hb8b1927f),
	.w2(32'hba3a1cb0),
	.w3(32'hba9f5a80),
	.w4(32'h3a33cb34),
	.w5(32'hb9d22842),
	.w6(32'h3801146c),
	.w7(32'hba1659ad),
	.w8(32'h3a92747a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f595b),
	.w1(32'hbbdee24a),
	.w2(32'hbb4aa263),
	.w3(32'hbb73dfc4),
	.w4(32'hbc0d1594),
	.w5(32'hbbb4c414),
	.w6(32'hbc13cad4),
	.w7(32'hbb3fb2dc),
	.w8(32'hbb28f28b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43250a),
	.w1(32'h3ad46f02),
	.w2(32'h39af51f0),
	.w3(32'hbbca3ad8),
	.w4(32'h3b223e34),
	.w5(32'h3a568760),
	.w6(32'h3acdaeaf),
	.w7(32'h3b0a796b),
	.w8(32'h3b8454fc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75b336),
	.w1(32'h3b03dffc),
	.w2(32'h3ad2ad0f),
	.w3(32'h3b596e56),
	.w4(32'h3b56ccf6),
	.w5(32'h3b94c155),
	.w6(32'h3b9cdd3a),
	.w7(32'h3afc9003),
	.w8(32'h3b9af289),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa5fe8),
	.w1(32'h3b77c336),
	.w2(32'h3b7fbde6),
	.w3(32'h3ae8262c),
	.w4(32'h3b08c4f3),
	.w5(32'h3a9b298c),
	.w6(32'h3b936e43),
	.w7(32'h3b864434),
	.w8(32'h3b02448e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8005a0),
	.w1(32'hbb011f8b),
	.w2(32'hba44893a),
	.w3(32'hb9a0bae0),
	.w4(32'hbad2bf77),
	.w5(32'hbab00e64),
	.w6(32'hbb26a67b),
	.w7(32'hba7ffaf9),
	.w8(32'hbacf85c8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30035e),
	.w1(32'hbaa7655c),
	.w2(32'hbaa481a3),
	.w3(32'hbb52f411),
	.w4(32'hbb9d4dcc),
	.w5(32'hbb90ea14),
	.w6(32'hbb6120ed),
	.w7(32'hbaeb1450),
	.w8(32'hbbb68f3d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe947fe),
	.w1(32'h3ad801e3),
	.w2(32'h3a0bbb8b),
	.w3(32'hbb4325c7),
	.w4(32'h3a2a4275),
	.w5(32'h3a9ed554),
	.w6(32'h3b59f338),
	.w7(32'h3b104f9f),
	.w8(32'hba94d70d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fa70),
	.w1(32'hbb0917f4),
	.w2(32'hbab64109),
	.w3(32'hba13fdb9),
	.w4(32'h3a9fa086),
	.w5(32'h3a997495),
	.w6(32'hbb1c1e21),
	.w7(32'h3a938045),
	.w8(32'h3b08c73c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f17c7),
	.w1(32'hbb817385),
	.w2(32'hbaf9136f),
	.w3(32'hba1ccdae),
	.w4(32'hbb2e757f),
	.w5(32'hbaa7491e),
	.w6(32'hbbdf5680),
	.w7(32'hbb5c10dc),
	.w8(32'hba5a15bb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18e83b),
	.w1(32'h390a9c25),
	.w2(32'h3b02a947),
	.w3(32'hbbf815a3),
	.w4(32'hbaf8896d),
	.w5(32'hba4299c1),
	.w6(32'hbb8623f1),
	.w7(32'h3ba409ac),
	.w8(32'h3b14b87b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254fe4),
	.w1(32'h3aebe8ec),
	.w2(32'h3bad1613),
	.w3(32'hba810d1b),
	.w4(32'hba3b6763),
	.w5(32'h3ab77783),
	.w6(32'h3a9a5b7b),
	.w7(32'h3b6c8fb8),
	.w8(32'h3afeb246),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c34df),
	.w1(32'hb9cd20f0),
	.w2(32'hba0d00d9),
	.w3(32'hb8bad24b),
	.w4(32'hb9ce2b4c),
	.w5(32'hba4d1f5f),
	.w6(32'hb98cdbf9),
	.w7(32'hba1f5b89),
	.w8(32'h3a5325bc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cbd29),
	.w1(32'hba9cc007),
	.w2(32'hbaf8d009),
	.w3(32'h3ab9ec37),
	.w4(32'hba5aa216),
	.w5(32'hbae1d0d1),
	.w6(32'hba6a573c),
	.w7(32'hbae254f3),
	.w8(32'hb98f07f7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc50b8),
	.w1(32'hbb8fdd40),
	.w2(32'hbbb9b225),
	.w3(32'hbab98762),
	.w4(32'hbb7c6283),
	.w5(32'hbb93a19c),
	.w6(32'hbb9be260),
	.w7(32'hbb8005a8),
	.w8(32'hbb0ec9e0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e4792),
	.w1(32'hbb88072e),
	.w2(32'hbac580f4),
	.w3(32'hbb147c3a),
	.w4(32'hbbbd7954),
	.w5(32'hbb989105),
	.w6(32'hbb6cf07a),
	.w7(32'hbb38d941),
	.w8(32'hbb5ba5a3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b0cf),
	.w1(32'h3c0cf2d9),
	.w2(32'h3bece8ac),
	.w3(32'hbbbe9201),
	.w4(32'h3c098d2f),
	.w5(32'h3c2c445b),
	.w6(32'h3c321087),
	.w7(32'h3b7b6416),
	.w8(32'h3bf9e7e5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49f37d),
	.w1(32'hba7c6e48),
	.w2(32'hbbea084f),
	.w3(32'h3bc38a06),
	.w4(32'h3b197312),
	.w5(32'hbb6832ef),
	.w6(32'h3a41f734),
	.w7(32'hbaf81126),
	.w8(32'h38f701d1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f03c),
	.w1(32'hba91e704),
	.w2(32'h39890a47),
	.w3(32'h3aefea58),
	.w4(32'h392c5dd8),
	.w5(32'h3ab95f97),
	.w6(32'h3a22f776),
	.w7(32'h3aae16c6),
	.w8(32'h3a47b28f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6499a1),
	.w1(32'h3b23cc03),
	.w2(32'hb9d201c7),
	.w3(32'hbb329e01),
	.w4(32'h3aec64cb),
	.w5(32'h397518d7),
	.w6(32'h3b2f3227),
	.w7(32'h3acdd35e),
	.w8(32'hbac6c5a5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba733b09),
	.w1(32'hbb2f951f),
	.w2(32'hbbb0e11f),
	.w3(32'hba43e903),
	.w4(32'hbaaeec6d),
	.w5(32'hbb53ad49),
	.w6(32'hba8e5639),
	.w7(32'hbb4d1a61),
	.w8(32'hb9b5e243),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedae68),
	.w1(32'hb914bbea),
	.w2(32'h398c391d),
	.w3(32'hba73795f),
	.w4(32'h3a414611),
	.w5(32'h3abfb6ff),
	.w6(32'hbaf89f2a),
	.w7(32'hb9149490),
	.w8(32'h3af547a1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9f9c),
	.w1(32'h3a13ef1a),
	.w2(32'h3bf14e9d),
	.w3(32'h3b1e81e4),
	.w4(32'hbb4c356e),
	.w5(32'h3905a196),
	.w6(32'h3ab0a1a7),
	.w7(32'h3be526c0),
	.w8(32'h3b2755ed),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3afcb),
	.w1(32'hbae472d9),
	.w2(32'hbb1b2036),
	.w3(32'hba866142),
	.w4(32'hbad9684a),
	.w5(32'hbb00f60a),
	.w6(32'hba30f9da),
	.w7(32'hbaadafa4),
	.w8(32'hbaa961c9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a50be),
	.w1(32'hbac0bb56),
	.w2(32'h3b02f002),
	.w3(32'hbb1bf244),
	.w4(32'hbad3e097),
	.w5(32'h39535c93),
	.w6(32'hbb26bcb8),
	.w7(32'h3a9d1cb1),
	.w8(32'h3a3fa72a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95968e),
	.w1(32'h3a6cf0ed),
	.w2(32'h3a9a3540),
	.w3(32'hbacc49dc),
	.w4(32'h3b282610),
	.w5(32'h3b1ba8a6),
	.w6(32'h38aba6d4),
	.w7(32'h3a14ca13),
	.w8(32'h3ad94814),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02e407),
	.w1(32'h3c78a0e8),
	.w2(32'h3c9b910f),
	.w3(32'h3b40b11e),
	.w4(32'h3c3a4bd2),
	.w5(32'h3c511aab),
	.w6(32'h3c5e35e6),
	.w7(32'h3c8c9ff3),
	.w8(32'h3c44e9d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ced1b),
	.w1(32'h3ab1edb5),
	.w2(32'h38ef3937),
	.w3(32'h3bbf4048),
	.w4(32'h3a80e60b),
	.w5(32'h3af0997e),
	.w6(32'hb9030b6a),
	.w7(32'hbb502deb),
	.w8(32'hbb28f7ea),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a09a60),
	.w1(32'hbb087a51),
	.w2(32'hbad59294),
	.w3(32'hbac8a3ff),
	.w4(32'hbab04f61),
	.w5(32'hbaa17eab),
	.w6(32'hba957415),
	.w7(32'hbaf043a5),
	.w8(32'h39b9f035),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7e21d),
	.w1(32'hbc11a6ca),
	.w2(32'hbc185caa),
	.w3(32'hb994dfa9),
	.w4(32'hbc06fa45),
	.w5(32'hbbfd8281),
	.w6(32'hbc0874bb),
	.w7(32'hbbe73ee1),
	.w8(32'hbc04677b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5eea),
	.w1(32'hbb7748a4),
	.w2(32'hbb9f836b),
	.w3(32'hbc158f52),
	.w4(32'hbb2e24a9),
	.w5(32'hbb5a1d75),
	.w6(32'hbb68506d),
	.w7(32'hbb61b0ab),
	.w8(32'hbaacb6d0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13b992),
	.w1(32'hbad7609d),
	.w2(32'hba36e9a7),
	.w3(32'hbb09f46e),
	.w4(32'hb99c4349),
	.w5(32'h3abc98c6),
	.w6(32'hbbaca7d7),
	.w7(32'hbb0a3953),
	.w8(32'h3a74f2c3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706ace),
	.w1(32'h3b8f4ef2),
	.w2(32'h3c06b110),
	.w3(32'hbb33f3b2),
	.w4(32'h3b44904c),
	.w5(32'h3bb9883d),
	.w6(32'h3b8ba746),
	.w7(32'h3c0c9eed),
	.w8(32'h3bc08651),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba011e6),
	.w1(32'hbb808f5f),
	.w2(32'hbac82dda),
	.w3(32'h3af12362),
	.w4(32'hbb8f87ca),
	.w5(32'hbb0bdd4a),
	.w6(32'hbbbcbddd),
	.w7(32'hbb2ea228),
	.w8(32'hbb4bd812),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5cbbc),
	.w1(32'hbb715489),
	.w2(32'hbbce704f),
	.w3(32'hbbed3d0d),
	.w4(32'hb981be88),
	.w5(32'hba99b102),
	.w6(32'hbb64aedb),
	.w7(32'hbb0fb197),
	.w8(32'h39043102),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70cb7),
	.w1(32'hbb7d09d0),
	.w2(32'hba7ff4e8),
	.w3(32'h3ac318a1),
	.w4(32'hbb7e8698),
	.w5(32'hba94b19b),
	.w6(32'hbb33feea),
	.w7(32'hba0c990e),
	.w8(32'hba959167),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974094),
	.w1(32'hbc085a2e),
	.w2(32'hbc3391fb),
	.w3(32'hbbb84098),
	.w4(32'hbbd0ac36),
	.w5(32'hbbf6a94d),
	.w6(32'hbc44fe54),
	.w7(32'hbc24f838),
	.w8(32'hbc2a8b07),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0645cc),
	.w1(32'h3aeca639),
	.w2(32'h3afb3c4a),
	.w3(32'hbbd97bce),
	.w4(32'h3a9a636d),
	.w5(32'h3961a19f),
	.w6(32'h3aaf0ca3),
	.w7(32'h3a8f93a3),
	.w8(32'h39e5fcec),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e8148),
	.w1(32'hbb55313a),
	.w2(32'hbba41dd5),
	.w3(32'hb8249d5f),
	.w4(32'hb9fa5cae),
	.w5(32'hb99087cd),
	.w6(32'hbb41aeb1),
	.w7(32'hbb5f2b4c),
	.w8(32'h3a313366),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770baf),
	.w1(32'h3a6f9619),
	.w2(32'h3c12c4e2),
	.w3(32'h3b32a02d),
	.w4(32'hbad3e910),
	.w5(32'h3b9c229b),
	.w6(32'h39553aea),
	.w7(32'h3bae00c5),
	.w8(32'h3b7b5894),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9995ac),
	.w1(32'hbc0c9920),
	.w2(32'hbc0c4d5a),
	.w3(32'hbb7fbab9),
	.w4(32'hbbc00ccd),
	.w5(32'hbbec676c),
	.w6(32'hbc302144),
	.w7(32'hbba21d2a),
	.w8(32'hbbdde0dc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6d66),
	.w1(32'h3beeb0d6),
	.w2(32'h3c925c3a),
	.w3(32'hbc35761c),
	.w4(32'h3ac4e119),
	.w5(32'h3c871f55),
	.w6(32'hbb24d2a2),
	.w7(32'h3c04ea65),
	.w8(32'h3c2009cf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28eed0),
	.w1(32'hbae19981),
	.w2(32'h3aecb02a),
	.w3(32'hbb85cf45),
	.w4(32'hbb5cf6a2),
	.w5(32'hbb3f6b79),
	.w6(32'hbbc1e91b),
	.w7(32'h3bff80ec),
	.w8(32'hbbacac04),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2f3d),
	.w1(32'h3b35fff8),
	.w2(32'hbba2da90),
	.w3(32'hbab93279),
	.w4(32'h3c0b677d),
	.w5(32'h3b3080dc),
	.w6(32'h3bb7992c),
	.w7(32'h3a22c9f8),
	.w8(32'h3bbd5ab4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0678a1),
	.w1(32'hba40259e),
	.w2(32'hbac5ad4e),
	.w3(32'h3bc28355),
	.w4(32'hba362199),
	.w5(32'hbadcb778),
	.w6(32'hba459b44),
	.w7(32'hbaedfcf4),
	.w8(32'hb7c64f23),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b3d62),
	.w1(32'hbaa28a79),
	.w2(32'hbbb8f3ed),
	.w3(32'hbae38fff),
	.w4(32'h3b363748),
	.w5(32'hba849090),
	.w6(32'h3944f863),
	.w7(32'h3804358a),
	.w8(32'h3a98d4e0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873dc4),
	.w1(32'h395cfeec),
	.w2(32'hbab276a5),
	.w3(32'h3adf4a7b),
	.w4(32'hb9d295e5),
	.w5(32'hbad33d15),
	.w6(32'hba8bc208),
	.w7(32'hbae50128),
	.w8(32'hbac69fce),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8766f1),
	.w1(32'hbb57605e),
	.w2(32'hba9a1957),
	.w3(32'hba697497),
	.w4(32'hbb7270f9),
	.w5(32'hbb3c2bc8),
	.w6(32'hbb32c492),
	.w7(32'hba4ff71f),
	.w8(32'hba20dfb3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145c3e),
	.w1(32'hbb249a3a),
	.w2(32'hbb131b6b),
	.w3(32'hbb8797f3),
	.w4(32'hbac1c9aa),
	.w5(32'hbaad7fb4),
	.w6(32'hbb055059),
	.w7(32'hbac44f54),
	.w8(32'h3a1b1854),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d40f1),
	.w1(32'hbb0d807b),
	.w2(32'hbc0ee98b),
	.w3(32'h39a03741),
	.w4(32'h3a7cab78),
	.w5(32'hbb97d520),
	.w6(32'h3ad3a100),
	.w7(32'hbb287739),
	.w8(32'hbae0c5a1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96c7a2),
	.w1(32'h38f3764e),
	.w2(32'h3adf33fa),
	.w3(32'h3abaf663),
	.w4(32'hba97b8cc),
	.w5(32'hbb31186b),
	.w6(32'hba7d3d91),
	.w7(32'h3a8f76d8),
	.w8(32'h3af999b9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf13c5),
	.w1(32'hbb93765e),
	.w2(32'hbbaaa279),
	.w3(32'hbb19f107),
	.w4(32'hbb4ecefc),
	.w5(32'hbb27e40a),
	.w6(32'hbb872006),
	.w7(32'hbbaf5c98),
	.w8(32'hbb1c7385),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e0c6),
	.w1(32'hb92ea489),
	.w2(32'hbbd57966),
	.w3(32'hbb78872b),
	.w4(32'h3bb8aca5),
	.w5(32'h3a573b61),
	.w6(32'h3b18eac7),
	.w7(32'hbbb0ceb3),
	.w8(32'h3b12cfb6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e26be),
	.w1(32'hbbb46e34),
	.w2(32'hbbb6a8f8),
	.w3(32'hbaaa1796),
	.w4(32'hbba117bf),
	.w5(32'hbbb2fe51),
	.w6(32'hbc024cae),
	.w7(32'hbbc9dc46),
	.w8(32'hbb8d8b41),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac415),
	.w1(32'hbb287c1d),
	.w2(32'h39830a0c),
	.w3(32'hbbf8f27b),
	.w4(32'hbbec7099),
	.w5(32'hbba44f0d),
	.w6(32'hbaa3bd8e),
	.w7(32'hba67c5e2),
	.w8(32'hbb9240f0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9055b5),
	.w1(32'h3aa29824),
	.w2(32'hba2cec60),
	.w3(32'hbc0d32d7),
	.w4(32'h3b3e65bf),
	.w5(32'h3a86010e),
	.w6(32'h3ad3819d),
	.w7(32'hb932289b),
	.w8(32'h3b448ffc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894c89),
	.w1(32'h3b00aaf6),
	.w2(32'hbb5650fb),
	.w3(32'h3b56a4c8),
	.w4(32'h3b9a3571),
	.w5(32'hb918805e),
	.w6(32'h3b8295ee),
	.w7(32'hb9b97735),
	.w8(32'h3b6643a3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dfd6c),
	.w1(32'h3ad30a35),
	.w2(32'h3910e559),
	.w3(32'h3b81c50a),
	.w4(32'h3b2adaf1),
	.w5(32'h3a9e1ab9),
	.w6(32'h3b0bc989),
	.w7(32'h3a959df0),
	.w8(32'h3b12a757),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031c1b),
	.w1(32'h3acaf96e),
	.w2(32'hba1810b7),
	.w3(32'h3b30908f),
	.w4(32'h3b35aa39),
	.w5(32'h3a48c578),
	.w6(32'h3ae1735c),
	.w7(32'h3978ffb4),
	.w8(32'h3acea362),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a939f8c),
	.w1(32'hbb0fef63),
	.w2(32'hbb5bb833),
	.w3(32'h3b1c244b),
	.w4(32'hbac41c49),
	.w5(32'hbb819732),
	.w6(32'hbb1294f7),
	.w7(32'h3b348fe7),
	.w8(32'h3a677582),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a1f2),
	.w1(32'hbb4e40c7),
	.w2(32'h3987e432),
	.w3(32'hbb7a7de6),
	.w4(32'hbb9f7b6a),
	.w5(32'hbb292b47),
	.w6(32'hbc0439ce),
	.w7(32'hba7d37ac),
	.w8(32'hbb6f4347),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3bd22),
	.w1(32'hbbca6867),
	.w2(32'hbbd0d7eb),
	.w3(32'hbb624628),
	.w4(32'hbbce024a),
	.w5(32'hbbce118e),
	.w6(32'hbbb43bff),
	.w7(32'hbbcadb27),
	.w8(32'hbb6c7beb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39219c),
	.w1(32'hbba1adc9),
	.w2(32'hbbe9856b),
	.w3(32'hbb354664),
	.w4(32'hbb758b4d),
	.w5(32'hbbb3fe7e),
	.w6(32'hbb6391c5),
	.w7(32'hbbb5ddb4),
	.w8(32'hbbec8b79),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc040493),
	.w1(32'h398504a0),
	.w2(32'hb9b853b0),
	.w3(32'hbbd937b7),
	.w4(32'h3ad8d7b8),
	.w5(32'h3a895a03),
	.w6(32'hba7ec46a),
	.w7(32'hb929c704),
	.w8(32'h3afa868d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d9d93),
	.w1(32'hbaac7d4e),
	.w2(32'hba38e865),
	.w3(32'h3b249c77),
	.w4(32'h3a526356),
	.w5(32'hbaad0ae4),
	.w6(32'hbb859850),
	.w7(32'h3bcc839e),
	.w8(32'h3ae6f5b6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bfe53),
	.w1(32'hbc16f68d),
	.w2(32'hbc1ce0a4),
	.w3(32'hb9f8eb90),
	.w4(32'hbc11ab67),
	.w5(32'hbc1a99d7),
	.w6(32'hbc1533b7),
	.w7(32'hbc2b59f9),
	.w8(32'hbc18583f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c4a0),
	.w1(32'hbb7ce90f),
	.w2(32'hbbb10480),
	.w3(32'hbc0619e7),
	.w4(32'hbb3c35ed),
	.w5(32'hbb8bba1f),
	.w6(32'hbb559bc4),
	.w7(32'hbb9d3ef1),
	.w8(32'hbad1f774),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6655),
	.w1(32'hba75da1f),
	.w2(32'hbab32a88),
	.w3(32'hbac4dcae),
	.w4(32'hb91bf037),
	.w5(32'h37faa31a),
	.w6(32'hb944f75e),
	.w7(32'hb94e6702),
	.w8(32'h391cdb6b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48c3c3),
	.w1(32'hba6cb13a),
	.w2(32'hba99b384),
	.w3(32'h3a88d63d),
	.w4(32'h3a536af2),
	.w5(32'hba553970),
	.w6(32'hba3f8849),
	.w7(32'hb913c054),
	.w8(32'hba396718),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eab8a),
	.w1(32'hbb0d87ef),
	.w2(32'hbba343cc),
	.w3(32'hba8b42ac),
	.w4(32'hba3a08d7),
	.w5(32'hbb0339f5),
	.w6(32'hbaf9a061),
	.w7(32'hba961612),
	.w8(32'hbae58ba9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8959a6e),
	.w1(32'h38121991),
	.w2(32'hb7203c20),
	.w3(32'hb78ffe9c),
	.w4(32'h38c0b62d),
	.w5(32'h38ab125a),
	.w6(32'hb8314b8d),
	.w7(32'h386f3c66),
	.w8(32'h37683f3d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53f56f),
	.w1(32'hb9bcbd1c),
	.w2(32'h36450a01),
	.w3(32'hba75a66a),
	.w4(32'hb9f3aee1),
	.w5(32'hb8ffbcee),
	.w6(32'hba8218bf),
	.w7(32'hb9ea9090),
	.w8(32'hb81f5e8d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e8969),
	.w1(32'hb8692102),
	.w2(32'h3895a31e),
	.w3(32'hba38369c),
	.w4(32'h3972c4bc),
	.w5(32'h3a1b7cc5),
	.w6(32'hba204be8),
	.w7(32'hb7697118),
	.w8(32'h39845b4b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98241b),
	.w1(32'hba3de271),
	.w2(32'hba463220),
	.w3(32'hba26eabc),
	.w4(32'hb9e36266),
	.w5(32'hb9925e74),
	.w6(32'hba9fa1b3),
	.w7(32'hba2959f8),
	.w8(32'hb9c37b1b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9afcc5),
	.w1(32'hb9d56f46),
	.w2(32'hba1bcd85),
	.w3(32'hb992760d),
	.w4(32'h3a867919),
	.w5(32'h3aeb0843),
	.w6(32'hb9c8197e),
	.w7(32'h3a419670),
	.w8(32'h3a9b6f7c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19d073),
	.w1(32'hbaed651b),
	.w2(32'hbb65a80f),
	.w3(32'h39c5d53d),
	.w4(32'hb9c4e8fb),
	.w5(32'hbaec5d5f),
	.w6(32'hba009cb2),
	.w7(32'hbac59dc1),
	.w8(32'hbb2d052f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac50fe),
	.w1(32'hba65a254),
	.w2(32'hbab87aa2),
	.w3(32'hba8602f9),
	.w4(32'hb9164487),
	.w5(32'hb8547676),
	.w6(32'hbaf7ee4e),
	.w7(32'hba7d13bd),
	.w8(32'hba2a1565),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122200),
	.w1(32'hbaba4eec),
	.w2(32'hbafc9455),
	.w3(32'h3a59e119),
	.w4(32'h3a96151a),
	.w5(32'h3af8271a),
	.w6(32'h3a92c4a5),
	.w7(32'h3a979eaf),
	.w8(32'h3a9a74db),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccda41),
	.w1(32'hba1a2961),
	.w2(32'hbaad05eb),
	.w3(32'h3978346b),
	.w4(32'h39b034f2),
	.w5(32'h382d4557),
	.w6(32'hba85ff92),
	.w7(32'hba9370fe),
	.w8(32'hba91c325),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedfe50),
	.w1(32'hba1e7cc9),
	.w2(32'hb9d0ef70),
	.w3(32'hba7f0fda),
	.w4(32'h392818c6),
	.w5(32'h39e87437),
	.w6(32'hbaceee52),
	.w7(32'hb90b131c),
	.w8(32'h381a7bbc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08f054),
	.w1(32'hbaebae2c),
	.w2(32'hbb52c589),
	.w3(32'h3a4f991b),
	.w4(32'hb91be8fa),
	.w5(32'hba893a0d),
	.w6(32'hb78b307c),
	.w7(32'hba52307c),
	.w8(32'hbaa2c4d5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bd94c),
	.w1(32'hb9f51d22),
	.w2(32'hba0550b2),
	.w3(32'hba0f0015),
	.w4(32'hb9315122),
	.w5(32'hb9387928),
	.w6(32'hba73597a),
	.w7(32'hb9e4fed4),
	.w8(32'hb9b3b885),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080d43),
	.w1(32'hb9e00ee5),
	.w2(32'hbaf6fb45),
	.w3(32'hbaab526e),
	.w4(32'h39606beb),
	.w5(32'h3a2916c2),
	.w6(32'hbaf34de6),
	.w7(32'hbaa5554d),
	.w8(32'hbabc433d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d512e8),
	.w1(32'h3a42fdd8),
	.w2(32'h3a93d782),
	.w3(32'hb8373d20),
	.w4(32'h3a7848f5),
	.w5(32'h3af3846c),
	.w6(32'hb9ab2faa),
	.w7(32'h39a8e7a0),
	.w8(32'h3a416d03),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3728f743),
	.w1(32'h37839722),
	.w2(32'hb74a6f2d),
	.w3(32'hb7618774),
	.w4(32'h36565bf0),
	.w5(32'hb781d2e3),
	.w6(32'hb6be27e7),
	.w7(32'h3670edb0),
	.w8(32'hb75079fe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59570c4),
	.w1(32'h3733f25a),
	.w2(32'hb7a6e870),
	.w3(32'hb8673f4f),
	.w4(32'hb7259614),
	.w5(32'hb8255933),
	.w6(32'hb77f0c45),
	.w7(32'h37b317cf),
	.w8(32'h3480a228),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e60b90),
	.w1(32'h398d9a70),
	.w2(32'h39296c40),
	.w3(32'hba32f988),
	.w4(32'h3966d332),
	.w5(32'h39a5104e),
	.w6(32'hba5d598b),
	.w7(32'hb9b3ce1d),
	.w8(32'hb988c09f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3178a7),
	.w1(32'hba0d725f),
	.w2(32'hbafdb20e),
	.w3(32'hba245c0a),
	.w4(32'h38aa642e),
	.w5(32'hba325df0),
	.w6(32'hba83263c),
	.w7(32'hbaa4b239),
	.w8(32'hbac2afa5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa1e83),
	.w1(32'hbb6c6a27),
	.w2(32'hbbaeb1d8),
	.w3(32'hbba72852),
	.w4(32'hbb34e9ed),
	.w5(32'hbb60fe77),
	.w6(32'hbbbce68a),
	.w7(32'hbb7ebac3),
	.w8(32'hbb834d49),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3744a115),
	.w1(32'h36baabd7),
	.w2(32'hb4b598a9),
	.w3(32'h372ac64f),
	.w4(32'hb60c8cd9),
	.w5(32'hb687418d),
	.w6(32'h3741b9e4),
	.w7(32'h34e7c6f9),
	.w8(32'hb49c4fbe),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ab047),
	.w1(32'hbb036b67),
	.w2(32'hbb82d817),
	.w3(32'hbab1441f),
	.w4(32'hba49fe3b),
	.w5(32'hbaf9340e),
	.w6(32'hbb1e38b9),
	.w7(32'hbaabd7d6),
	.w8(32'hbb043c76),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadca9f1),
	.w1(32'hbb04bde7),
	.w2(32'hbb47c81b),
	.w3(32'hba226f59),
	.w4(32'hbaa14ecc),
	.w5(32'hbadf12ab),
	.w6(32'hba9e8298),
	.w7(32'hbaba6b94),
	.w8(32'hbaefbfdc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af91a4),
	.w1(32'hbb918b02),
	.w2(32'hbbed232e),
	.w3(32'h3a4c9651),
	.w4(32'hbb13ffd6),
	.w5(32'hbb59b29d),
	.w6(32'h39c7d2f1),
	.w7(32'hbaec0be6),
	.w8(32'hbb1702f8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42f9ca),
	.w1(32'h39efd331),
	.w2(32'hb9d61be0),
	.w3(32'hb9c947f5),
	.w4(32'h3a87a4e4),
	.w5(32'h3a536d15),
	.w6(32'hba5d75a0),
	.w7(32'hb8d5dd4c),
	.w8(32'h397de0ef),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfae30),
	.w1(32'h3a41ac6c),
	.w2(32'h3b0a4ae1),
	.w3(32'h3a11819d),
	.w4(32'h3a694ba4),
	.w5(32'h3afb6504),
	.w6(32'h39ccf689),
	.w7(32'h39846a67),
	.w8(32'h3a189511),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb3e46),
	.w1(32'h39c22160),
	.w2(32'h39ba1bbd),
	.w3(32'h39eb30bc),
	.w4(32'h39c15fbd),
	.w5(32'h393e4f3c),
	.w6(32'h39e5f9d6),
	.w7(32'h39c11f03),
	.w8(32'h38f1c968),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4767e2),
	.w1(32'hb8582dee),
	.w2(32'h39a727de),
	.w3(32'hbb0840a2),
	.w4(32'h39cbca54),
	.w5(32'h3a1606fb),
	.w6(32'hbb4c2bce),
	.w7(32'hb9a8a7c9),
	.w8(32'h3839bc58),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91bee7),
	.w1(32'h3ac79f4e),
	.w2(32'h3b1bc391),
	.w3(32'h3948a546),
	.w4(32'h3b5e906c),
	.w5(32'h3ba7b7b4),
	.w6(32'h3aadc55d),
	.w7(32'h3b476a2a),
	.w8(32'h3b32868c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b047b),
	.w1(32'h3a3c875f),
	.w2(32'h3b05f748),
	.w3(32'hbb39c14e),
	.w4(32'h3a326d94),
	.w5(32'h3b0342bb),
	.w6(32'hbb50de20),
	.w7(32'h39bd16e3),
	.w8(32'h3aaddc24),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9334143),
	.w1(32'h380ab9e0),
	.w2(32'hb8c7801f),
	.w3(32'hb8ee6bdc),
	.w4(32'h388bde69),
	.w5(32'hb7d89c59),
	.w6(32'hb908aac4),
	.w7(32'h38821ad5),
	.w8(32'hb8a0ea12),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82391de),
	.w1(32'hb80293cb),
	.w2(32'hb85d3ac5),
	.w3(32'hb8513cd2),
	.w4(32'hb875a3f0),
	.w5(32'hb8abce07),
	.w6(32'hb8e4ac73),
	.w7(32'hb88b119a),
	.w8(32'hb8ce8f11),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba435a99),
	.w1(32'hbae1be9d),
	.w2(32'hbb0a99f7),
	.w3(32'hb88af0ea),
	.w4(32'hb93315d6),
	.w5(32'hb9f728eb),
	.w6(32'hba5ccb6f),
	.w7(32'hba0a26fd),
	.w8(32'hba149396),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959d90e),
	.w1(32'h386a3b99),
	.w2(32'hb9034364),
	.w3(32'h3937f446),
	.w4(32'h387101f8),
	.w5(32'h38462eea),
	.w6(32'h38be8675),
	.w7(32'hb7482f49),
	.w8(32'hb8daca63),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f0d5c),
	.w1(32'hb929d0eb),
	.w2(32'hb999719b),
	.w3(32'hb831efd6),
	.w4(32'h38f1c989),
	.w5(32'h3763698e),
	.w6(32'hba8b665e),
	.w7(32'hb9ca0ca1),
	.w8(32'hb9028e5b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cea561),
	.w1(32'hb40bf0dd),
	.w2(32'hb7b3967e),
	.w3(32'hb6485026),
	.w4(32'h379694ac),
	.w5(32'hb7c6c00a),
	.w6(32'h382a40db),
	.w7(32'hb7bd4cf7),
	.w8(32'h37b6c3f2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c060),
	.w1(32'hb9deffb4),
	.w2(32'h3b0867e9),
	.w3(32'hbb877a58),
	.w4(32'h39020b8f),
	.w5(32'h3aadb61e),
	.w6(32'hbbc05627),
	.w7(32'h39faf92c),
	.w8(32'h3ac426d7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383535d7),
	.w1(32'h385b90bc),
	.w2(32'h36a23df6),
	.w3(32'h388f0576),
	.w4(32'h388818dd),
	.w5(32'h3636c8e5),
	.w6(32'h38c1a27d),
	.w7(32'h3894825a),
	.w8(32'h37b2eca6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891fe94),
	.w1(32'hb8918c14),
	.w2(32'hb8e2eddc),
	.w3(32'h382f9642),
	.w4(32'hb7dc8770),
	.w5(32'hb8025f52),
	.w6(32'h3908a90f),
	.w7(32'h3913b9e2),
	.w8(32'h3780a1b9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3f436),
	.w1(32'hbab6a807),
	.w2(32'hbb04123a),
	.w3(32'h39e14edd),
	.w4(32'h3985fe8b),
	.w5(32'h39f64abc),
	.w6(32'hba19618d),
	.w7(32'hb9fc9d09),
	.w8(32'h360a5f2e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95142e),
	.w1(32'hbb130245),
	.w2(32'hbb6effeb),
	.w3(32'hbb24f730),
	.w4(32'hb99f6951),
	.w5(32'hbae6d1ef),
	.w6(32'hbb4f07f3),
	.w7(32'hb983eb98),
	.w8(32'hbaaec8ce),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb475e53),
	.w1(32'h3a5d824e),
	.w2(32'h3ae4d719),
	.w3(32'hbb256194),
	.w4(32'h3a829ef1),
	.w5(32'h3af8cf6b),
	.w6(32'hbb5e0dc9),
	.w7(32'h39abcdff),
	.w8(32'h3aa664c5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15cea0),
	.w1(32'hbb29d108),
	.w2(32'hbb5f3e4f),
	.w3(32'hbac52014),
	.w4(32'hbb070e1f),
	.w5(32'hbb026f4f),
	.w6(32'hbb239caf),
	.w7(32'hbb1babc0),
	.w8(32'hbb00fac4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dabfab),
	.w1(32'hb93e3831),
	.w2(32'hba0d3d8c),
	.w3(32'h377910da),
	.w4(32'h37c4b379),
	.w5(32'hb6fac42f),
	.w6(32'h39a7832d),
	.w7(32'h389935d5),
	.w8(32'h3706853a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb960f35),
	.w1(32'hbb8a6246),
	.w2(32'hbbe781b7),
	.w3(32'hbb42ac2f),
	.w4(32'hbacede09),
	.w5(32'hbb2a216d),
	.w6(32'hbb87a19c),
	.w7(32'hbb910cff),
	.w8(32'hbb8d5dce),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d7933),
	.w1(32'hba82181f),
	.w2(32'hba489493),
	.w3(32'hbabda250),
	.w4(32'hb8eea3ee),
	.w5(32'h3a490f8d),
	.w6(32'hbaf157d9),
	.w7(32'hb71e6ee2),
	.w8(32'h3a1b0da7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46e661),
	.w1(32'hbaf90146),
	.w2(32'hbb617d0b),
	.w3(32'hbaea3f3f),
	.w4(32'hba705000),
	.w5(32'hbb031d1c),
	.w6(32'hbb248071),
	.w7(32'hbaadc10e),
	.w8(32'hbb00b52f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883c9b3),
	.w1(32'h38167a33),
	.w2(32'hb7ae4aa7),
	.w3(32'h38d31154),
	.w4(32'h38b220e1),
	.w5(32'h382b9f1b),
	.w6(32'h38e4e569),
	.w7(32'h38bacfed),
	.w8(32'hb73381e4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9950f19),
	.w1(32'hb95dedcc),
	.w2(32'hbb10f53d),
	.w3(32'h39768284),
	.w4(32'h3a7b5203),
	.w5(32'h388c84cc),
	.w6(32'hb93366bc),
	.w7(32'h3918e796),
	.w8(32'hb9db4627),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885c2eb),
	.w1(32'h36bb1088),
	.w2(32'hb7e37855),
	.w3(32'h382f1cd3),
	.w4(32'hb5b6e1fc),
	.w5(32'hb819d172),
	.w6(32'h3823bc80),
	.w7(32'hb6a5634f),
	.w8(32'hb7dac16a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52a8bc),
	.w1(32'hba6539f4),
	.w2(32'hba9d22cb),
	.w3(32'hba0fb5ea),
	.w4(32'hba115b1f),
	.w5(32'hba6cf43a),
	.w6(32'hba174d5c),
	.w7(32'hba0af89c),
	.w8(32'hba1853f1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fb2a4),
	.w1(32'hb8404738),
	.w2(32'hb830083f),
	.w3(32'hb914f5ec),
	.w4(32'hb6b77c79),
	.w5(32'h37f74fc1),
	.w6(32'hb95c3113),
	.w7(32'h36a36303),
	.w8(32'h3869bcbf),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1685b1),
	.w1(32'hbadc9bb2),
	.w2(32'hbb6a2e5c),
	.w3(32'hba9aa14e),
	.w4(32'hb996d6d8),
	.w5(32'hba8bd259),
	.w6(32'hbac72e92),
	.w7(32'hba8866d2),
	.w8(32'hbaddba64),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37994ca9),
	.w1(32'h369c9998),
	.w2(32'hb7154829),
	.w3(32'h3748844e),
	.w4(32'hb5e8124e),
	.w5(32'hb7705dd5),
	.w6(32'h3789c70a),
	.w7(32'h36d38b81),
	.w8(32'hb6924485),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ce29f4),
	.w1(32'h38078827),
	.w2(32'h37947ef8),
	.w3(32'h38410f1d),
	.w4(32'h3766b096),
	.w5(32'hb7df5998),
	.w6(32'h3832cc5d),
	.w7(32'h3706dc3c),
	.w8(32'hb7eebf21),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacab6e1),
	.w1(32'h3986ff5e),
	.w2(32'h3a2c8a74),
	.w3(32'hba989156),
	.w4(32'h39ca6298),
	.w5(32'h3a30d444),
	.w6(32'hbacf5a4c),
	.w7(32'hb93e6e33),
	.w8(32'h39828c3e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb091a9c),
	.w1(32'h3a8117a3),
	.w2(32'h3add4ed8),
	.w3(32'hbae47ae6),
	.w4(32'h3aff6f89),
	.w5(32'h3b5b86d3),
	.w6(32'hbb23f744),
	.w7(32'hb904b1bd),
	.w8(32'h3a9d2180),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8accfc),
	.w1(32'h3906604b),
	.w2(32'hb9272a88),
	.w3(32'hba4be4e1),
	.w4(32'h3a0d674e),
	.w5(32'h39991075),
	.w6(32'hb94d72c2),
	.w7(32'h3a9f34a8),
	.w8(32'h37ce3e04),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953e85b),
	.w1(32'hb920aee1),
	.w2(32'hb87e0698),
	.w3(32'hb9af3899),
	.w4(32'hb8d1ff8f),
	.w5(32'hb928f623),
	.w6(32'hb8d907f0),
	.w7(32'hb7aa2c3c),
	.w8(32'hb90d4e66),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2a26),
	.w1(32'hbc0d5d18),
	.w2(32'hbc6935d6),
	.w3(32'hbc04b3fc),
	.w4(32'hbbe741ac),
	.w5(32'hbc44ef88),
	.w6(32'hbc0f5985),
	.w7(32'hbbf49a1c),
	.w8(32'hbc2d95b0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe570d),
	.w1(32'hb92df852),
	.w2(32'hbab02184),
	.w3(32'hbb7302d7),
	.w4(32'h3af5e77c),
	.w5(32'h3b64e0c8),
	.w6(32'hbb3ac7ad),
	.w7(32'h3ab495af),
	.w8(32'h3b0747a0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d9c0d),
	.w1(32'hb893feeb),
	.w2(32'hb969ced5),
	.w3(32'h3929b06e),
	.w4(32'hb8e01fd8),
	.w5(32'hb9202b2d),
	.w6(32'h397795d8),
	.w7(32'hb753f6ee),
	.w8(32'hb99d15ff),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379430f9),
	.w1(32'h348b11c4),
	.w2(32'hb64eb8f5),
	.w3(32'h37977e60),
	.w4(32'hb7536f3e),
	.w5(32'hb67eaa4f),
	.w6(32'h37d73bf9),
	.w7(32'hb65961b7),
	.w8(32'hb77e93e0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ecb28),
	.w1(32'h37e4fddd),
	.w2(32'h37c38e9d),
	.w3(32'hb78f3944),
	.w4(32'hb798e357),
	.w5(32'hb8298343),
	.w6(32'hb63edce1),
	.w7(32'hb7f32d76),
	.w8(32'hb801970c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384dfc93),
	.w1(32'h37166728),
	.w2(32'hb7722db4),
	.w3(32'h380562a9),
	.w4(32'hb573e30e),
	.w5(32'hb7953ef2),
	.w6(32'h38220776),
	.w7(32'h36e1a556),
	.w8(32'hb6f2a948),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3689a5),
	.w1(32'hb7c1c20d),
	.w2(32'hb90acd0d),
	.w3(32'h3a40e667),
	.w4(32'h396a4b38),
	.w5(32'h397fd349),
	.w6(32'h38bf0000),
	.w7(32'hb9aa22df),
	.w8(32'hb9297fc3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad44b46),
	.w1(32'hbab51102),
	.w2(32'hba09fc81),
	.w3(32'hb98ec5ce),
	.w4(32'h395c88f0),
	.w5(32'h3a909125),
	.w6(32'hbad88729),
	.w7(32'hbb0766a3),
	.w8(32'hbaf65f0a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3bce1),
	.w1(32'hbb91bf4b),
	.w2(32'hbbd302cb),
	.w3(32'hbb87e88d),
	.w4(32'hbb162669),
	.w5(32'hbb5dca8c),
	.w6(32'hbba830b3),
	.w7(32'hbb2e1687),
	.w8(32'hbb536e43),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79c1e9),
	.w1(32'hb9059b48),
	.w2(32'hb7edaefa),
	.w3(32'hba7917d8),
	.w4(32'hb915be9e),
	.w5(32'h3923e31e),
	.w6(32'hba9daf44),
	.w7(32'h3806ea25),
	.w8(32'h394ffc49),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadce923),
	.w1(32'hbb86c330),
	.w2(32'hbbba6059),
	.w3(32'hba0aed3c),
	.w4(32'hbb0f249b),
	.w5(32'hbb590e5b),
	.w6(32'hbb183126),
	.w7(32'hbb5a6d1f),
	.w8(32'hbb52ef0d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59321b),
	.w1(32'h38623a29),
	.w2(32'hb997b1c8),
	.w3(32'hba40f899),
	.w4(32'h358f2abc),
	.w5(32'hb8e018c7),
	.w6(32'hba51cda8),
	.w7(32'hb9acc95e),
	.w8(32'hb9beb7f4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385d90c8),
	.w1(32'h37c2349c),
	.w2(32'h36bca75d),
	.w3(32'h3828c617),
	.w4(32'h371efede),
	.w5(32'hb6f4205d),
	.w6(32'h38596dff),
	.w7(32'h37953186),
	.w8(32'h367d3d78),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e420ea),
	.w1(32'hb9a5d915),
	.w2(32'hb9672c25),
	.w3(32'hb97b09cc),
	.w4(32'hb885c95a),
	.w5(32'h38ad0079),
	.w6(32'hb890fcb5),
	.w7(32'h390303d2),
	.w8(32'h3952b9e2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c56d8f),
	.w1(32'h379fccce),
	.w2(32'hb7924c8b),
	.w3(32'h38751223),
	.w4(32'hb74544c5),
	.w5(32'hb845db29),
	.w6(32'h38a0b221),
	.w7(32'h378ca87c),
	.w8(32'hb75fcfbf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc03a),
	.w1(32'hba73093f),
	.w2(32'hba56c287),
	.w3(32'hbacadc91),
	.w4(32'hb99b9a49),
	.w5(32'h38eb05b9),
	.w6(32'hbb1c515c),
	.w7(32'hba66d4c9),
	.w8(32'hba165081),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6662a1),
	.w1(32'h39bbc62a),
	.w2(32'h3b75b361),
	.w3(32'hbb1e9340),
	.w4(32'h3ab29172),
	.w5(32'h3b96fe5f),
	.w6(32'hbb24877e),
	.w7(32'h3aca36a5),
	.w8(32'h3b685176),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf343ab),
	.w1(32'hbac5449c),
	.w2(32'hbaf6f191),
	.w3(32'hba36137d),
	.w4(32'hb8e890b8),
	.w5(32'hb7a43eaa),
	.w6(32'hbaaeb3fc),
	.w7(32'hb99ae6ab),
	.w8(32'hb8d52a25),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f2217),
	.w1(32'h3a5ccfb7),
	.w2(32'h3b05c308),
	.w3(32'hba4333c7),
	.w4(32'h3a041b74),
	.w5(32'h3ae33dd4),
	.w6(32'hba4f592e),
	.w7(32'h39a0f4b0),
	.w8(32'h3aab8099),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f792),
	.w1(32'hbb184e55),
	.w2(32'hbb3ff6a2),
	.w3(32'hba87a26b),
	.w4(32'hba103fbd),
	.w5(32'hb9129f5f),
	.w6(32'hbb0a1fa8),
	.w7(32'hbad2c2f6),
	.w8(32'hba6ecea3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ee0a),
	.w1(32'hbaac1998),
	.w2(32'hbb07c3b4),
	.w3(32'hba308ed0),
	.w4(32'hba7403b3),
	.w5(32'hba94e242),
	.w6(32'hbadd9ba3),
	.w7(32'hbaae3fe4),
	.w8(32'hba9c64f4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf22ed4),
	.w1(32'hbb4aee6a),
	.w2(32'hbb40516d),
	.w3(32'hbbcff44d),
	.w4(32'hbb2a7b45),
	.w5(32'hbb145973),
	.w6(32'hbbdf416e),
	.w7(32'hbb840cf7),
	.w8(32'hbb8e4022),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cab5f9),
	.w1(32'h362ee59b),
	.w2(32'hb6d928de),
	.w3(32'h375053df),
	.w4(32'hb5ff737e),
	.w5(32'hb775f2ec),
	.w6(32'h378face9),
	.w7(32'hb4d96ea0),
	.w8(32'hb749f8a9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a1c6aa),
	.w1(32'h383068bc),
	.w2(32'h37a02146),
	.w3(32'h378579d6),
	.w4(32'h37bce38f),
	.w5(32'h37575494),
	.w6(32'hb39a27d2),
	.w7(32'h3793bfea),
	.w8(32'h37b107bf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236708),
	.w1(32'hb608ee5a),
	.w2(32'h3ac9ba57),
	.w3(32'hba8a28c2),
	.w4(32'h3a9e6b83),
	.w5(32'h3b2f0772),
	.w6(32'hbadfd9a8),
	.w7(32'h3a3d7378),
	.w8(32'h3abe20ad),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817cfb),
	.w1(32'hbaefa0c5),
	.w2(32'hbb02929e),
	.w3(32'hbb0668ac),
	.w4(32'hb9da46a0),
	.w5(32'hba1ec385),
	.w6(32'hbb361cf0),
	.w7(32'hba16f702),
	.w8(32'hb9f3cd91),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f1791),
	.w1(32'hbae968ea),
	.w2(32'hbb30ddd4),
	.w3(32'hbad633ca),
	.w4(32'hb7e46470),
	.w5(32'hb9f4c2a4),
	.w6(32'hbb41032c),
	.w7(32'hba74ad08),
	.w8(32'hbaaf22e1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a483c5e),
	.w1(32'h391ad3b6),
	.w2(32'h387c3c24),
	.w3(32'h386199c8),
	.w4(32'hb8d484d1),
	.w5(32'h398071b1),
	.w6(32'h3a2dc35b),
	.w7(32'h3977c97e),
	.w8(32'hb9c24535),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386cfc1e),
	.w1(32'hb894001c),
	.w2(32'hb8b51a56),
	.w3(32'h386ece9b),
	.w4(32'hb8844d57),
	.w5(32'hb80d9391),
	.w6(32'hb80059e2),
	.w7(32'hb8cc4f1a),
	.w8(32'hb8075937),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d9b84),
	.w1(32'hb95809b7),
	.w2(32'hb96ddb9b),
	.w3(32'hb8152dab),
	.w4(32'hb844d9a5),
	.w5(32'hb8d742d0),
	.w6(32'hb7353f57),
	.w7(32'h3880b07e),
	.w8(32'hb86ecc23),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ed369),
	.w1(32'h397342de),
	.w2(32'hb9430b67),
	.w3(32'h39d22d06),
	.w4(32'h399839e6),
	.w5(32'hba4428f1),
	.w6(32'hb94983a0),
	.w7(32'h3996fe00),
	.w8(32'hba54f67e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00b46),
	.w1(32'hbba90d26),
	.w2(32'hbbbd0951),
	.w3(32'hbbb3cbcf),
	.w4(32'hbb890aba),
	.w5(32'hbbab2af7),
	.w6(32'hbbd39d36),
	.w7(32'hbb97aa03),
	.w8(32'hbbaa3a11),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37d67d),
	.w1(32'hbabe8168),
	.w2(32'hbbac52b1),
	.w3(32'h3aa043ba),
	.w4(32'h3a4c3234),
	.w5(32'hba75caa7),
	.w6(32'h3ac838f5),
	.w7(32'h3a3c343c),
	.w8(32'hbad54dd0),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a315),
	.w1(32'h3afb9fca),
	.w2(32'h3b322ebe),
	.w3(32'hbb097fa2),
	.w4(32'h3b0ebb47),
	.w5(32'h3b7112fc),
	.w6(32'hbb068fbb),
	.w7(32'h3a9b3355),
	.w8(32'h3b0bc1dc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9fbe),
	.w1(32'hbab289ba),
	.w2(32'hb9b2669b),
	.w3(32'hbb839ce0),
	.w4(32'hb9ee01f8),
	.w5(32'h3a635394),
	.w6(32'hbb8f1064),
	.w7(32'hba438658),
	.w8(32'h39db3a5e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ae6b69),
	.w1(32'h3726b05a),
	.w2(32'h363e26d0),
	.w3(32'h3776d3f7),
	.w4(32'h36ac488b),
	.w5(32'hb5cf4675),
	.w6(32'h379980c1),
	.w7(32'h3704c4f0),
	.w8(32'h3663b05d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f4fdc),
	.w1(32'h36c0d69b),
	.w2(32'h36890e20),
	.w3(32'h37304f9f),
	.w4(32'hb5960835),
	.w5(32'hb71220a7),
	.w6(32'h3798e699),
	.w7(32'h36a947ab),
	.w8(32'h34383402),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39647a60),
	.w1(32'h393c8f73),
	.w2(32'h38f40fed),
	.w3(32'h3a2dce63),
	.w4(32'h39900652),
	.w5(32'h38dabb11),
	.w6(32'h3884d7e9),
	.w7(32'hb8a55c7c),
	.w8(32'hb87ed2b8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382777b2),
	.w1(32'h365bec8b),
	.w2(32'hb80d9a85),
	.w3(32'h38105888),
	.w4(32'hb7098534),
	.w5(32'hb7dc7410),
	.w6(32'h3832d8e5),
	.w7(32'h363bb013),
	.w8(32'hb78b9f14),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996a081),
	.w1(32'hb9392d42),
	.w2(32'hb9533f1a),
	.w3(32'h38601092),
	.w4(32'hb4f890f8),
	.w5(32'h37e48bbe),
	.w6(32'hb8b6375d),
	.w7(32'hb92990dd),
	.w8(32'hb98901be),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a562b),
	.w1(32'hba9d90ec),
	.w2(32'hbac47995),
	.w3(32'hba8731c6),
	.w4(32'h395ae3d4),
	.w5(32'hb9a9ed89),
	.w6(32'hbaf3248f),
	.w7(32'hb99a6bcc),
	.w8(32'hb913011b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb55cf),
	.w1(32'hbaf14fca),
	.w2(32'hbb0ab414),
	.w3(32'hba8dbd55),
	.w4(32'hba57b107),
	.w5(32'hba5f53b0),
	.w6(32'hba987540),
	.w7(32'hba93f9cd),
	.w8(32'hba61df73),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eab415),
	.w1(32'h37396f1c),
	.w2(32'h36d32497),
	.w3(32'h37cbade0),
	.w4(32'h374c797e),
	.w5(32'h36202bbc),
	.w6(32'h37d5c422),
	.w7(32'h37767647),
	.w8(32'h369afa05),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845e3e),
	.w1(32'hbaf183b9),
	.w2(32'hbb675049),
	.w3(32'h3981d4cd),
	.w4(32'hb9944bb9),
	.w5(32'hba89f4ab),
	.w6(32'hba5ccc0b),
	.w7(32'hb9beb59e),
	.w8(32'hba0617f0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ea599),
	.w1(32'hb9f2d341),
	.w2(32'hba740373),
	.w3(32'hb7c40e8a),
	.w4(32'hb8b8bb2c),
	.w5(32'hba252628),
	.w6(32'hb9fcfbfb),
	.w7(32'hb9d9a07c),
	.w8(32'hba8e8edc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f6c3f),
	.w1(32'hb76b92a5),
	.w2(32'h395bf6e5),
	.w3(32'hb8d7dc41),
	.w4(32'h384b391b),
	.w5(32'h399f9670),
	.w6(32'hb8dff5b2),
	.w7(32'h3907c6a2),
	.w8(32'h39c2aa54),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9998395),
	.w1(32'hba098ae8),
	.w2(32'hba937933),
	.w3(32'h38fdb975),
	.w4(32'hb875c280),
	.w5(32'hb9c9017e),
	.w6(32'hba1a0e54),
	.w7(32'hba406373),
	.w8(32'hba76afc4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6ebfd),
	.w1(32'h387d66ce),
	.w2(32'h3819b567),
	.w3(32'h3896374c),
	.w4(32'h382d514d),
	.w5(32'h379c5147),
	.w6(32'h389698d1),
	.w7(32'h3815d743),
	.w8(32'h37eaf65c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dc9a17),
	.w1(32'h3874aef5),
	.w2(32'h38f2abfb),
	.w3(32'h385ae4b2),
	.w4(32'h3895b8ee),
	.w5(32'h38b8d5fa),
	.w6(32'hb822ef30),
	.w7(32'hb6b5a524),
	.w8(32'h379f0d52),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375abf73),
	.w1(32'h379ce6e1),
	.w2(32'h3808789e),
	.w3(32'h37129d7e),
	.w4(32'h38119c57),
	.w5(32'h381f2121),
	.w6(32'h38120867),
	.w7(32'h386302f2),
	.w8(32'h38041f12),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e32164),
	.w1(32'h3765e00e),
	.w2(32'h355910ed),
	.w3(32'h37ab2b61),
	.w4(32'h36e2ec5f),
	.w5(32'hb6da91b3),
	.w6(32'h37d84512),
	.w7(32'h36fb8042),
	.w8(32'hb5aae61d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948fc5),
	.w1(32'hb9ecb86c),
	.w2(32'h39086f9d),
	.w3(32'hba880807),
	.w4(32'hba0b82bd),
	.w5(32'h39a6193b),
	.w6(32'hbabb1b3d),
	.w7(32'hba466f7f),
	.w8(32'h38e94351),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb568),
	.w1(32'hbb0e3071),
	.w2(32'hbb6082f9),
	.w3(32'hba8d1c5b),
	.w4(32'hba69be6d),
	.w5(32'hba9840b8),
	.w6(32'hbb0e9e4e),
	.w7(32'hbb1242f6),
	.w8(32'hbafa43dd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec75e1),
	.w1(32'hba9bf0af),
	.w2(32'hbb161504),
	.w3(32'hba7c2ad2),
	.w4(32'hba06988f),
	.w5(32'hbaa2b26a),
	.w6(32'hbb0082d5),
	.w7(32'hba9be5da),
	.w8(32'hbab96758),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b7380),
	.w1(32'hbb6cd6b8),
	.w2(32'hbbd486dc),
	.w3(32'hbb0610f9),
	.w4(32'hbb13853c),
	.w5(32'hbb88bb86),
	.w6(32'hbb15e7e5),
	.w7(32'hbb325d83),
	.w8(32'hbb845b2a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2da97),
	.w1(32'hb8b453cb),
	.w2(32'h38895b4c),
	.w3(32'hb9005aac),
	.w4(32'hb8bc1e51),
	.w5(32'h38689423),
	.w6(32'hb8fedff1),
	.w7(32'hb8d2e792),
	.w8(32'hb791ac89),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e6cc61),
	.w1(32'hb8bfae22),
	.w2(32'hb8c12886),
	.w3(32'hb7a678bb),
	.w4(32'h3774e866),
	.w5(32'h37480b22),
	.w6(32'h37494342),
	.w7(32'h380d92a6),
	.w8(32'h37341631),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371b85ee),
	.w1(32'hb5680118),
	.w2(32'hb6900318),
	.w3(32'h3659ff35),
	.w4(32'hb6a18363),
	.w5(32'hb7110100),
	.w6(32'h372a82f8),
	.w7(32'hb637395e),
	.w8(32'hb68aab21),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e55d74),
	.w1(32'hb6cdaafb),
	.w2(32'h37835158),
	.w3(32'h38438e2f),
	.w4(32'h3821d08c),
	.w5(32'h38078fbd),
	.w6(32'hb65a46a9),
	.w7(32'h372eaded),
	.w8(32'h3827c683),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f378),
	.w1(32'hbaa59a58),
	.w2(32'hbb79412b),
	.w3(32'h38794618),
	.w4(32'h3745d9ee),
	.w5(32'hbab44322),
	.w6(32'hb9850670),
	.w7(32'hb9ccbbce),
	.w8(32'hbac18785),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89bf14f),
	.w1(32'hb7b2347f),
	.w2(32'h372d95c8),
	.w3(32'hb8cdcc6f),
	.w4(32'hb8902ca6),
	.w5(32'hb874553d),
	.w6(32'hb8821741),
	.w7(32'hb8a41287),
	.w8(32'hb881a0c0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6786b3),
	.w1(32'h3a3dacfd),
	.w2(32'h3a8444b1),
	.w3(32'hba4a5313),
	.w4(32'h3a181e9c),
	.w5(32'h3a79c496),
	.w6(32'hba5b3166),
	.w7(32'h39e4f006),
	.w8(32'h3a214d8b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf1350),
	.w1(32'hb78668e2),
	.w2(32'h39b56de7),
	.w3(32'hba998f73),
	.w4(32'h3833fc31),
	.w5(32'h3a143420),
	.w6(32'hba7349be),
	.w7(32'h37592737),
	.w8(32'h3999d311),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a4841),
	.w1(32'h36843497),
	.w2(32'hb6b2c674),
	.w3(32'h36e47016),
	.w4(32'hb6a3fbc7),
	.w5(32'hb7156684),
	.w6(32'h370f793f),
	.w7(32'hb70ff61e),
	.w8(32'hb6e59ead),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17128c),
	.w1(32'hba9ca92b),
	.w2(32'hbae12e9c),
	.w3(32'hba0f3dbc),
	.w4(32'hba400d52),
	.w5(32'hba93a4a1),
	.w6(32'hba495383),
	.w7(32'hba783581),
	.w8(32'hba9b78fb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d76ec6),
	.w1(32'hb80dbffa),
	.w2(32'hb80508e2),
	.w3(32'h3858e1c7),
	.w4(32'hb606a70d),
	.w5(32'hb781effa),
	.w6(32'h382429ce),
	.w7(32'h379443a2),
	.w8(32'hb8183627),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0cc3),
	.w1(32'hbb61e0f7),
	.w2(32'hbbbbbb50),
	.w3(32'hb970d32b),
	.w4(32'hba9e01aa),
	.w5(32'hbae233c1),
	.w6(32'hb9257e3f),
	.w7(32'hba663081),
	.w8(32'hba8a9658),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77a2061),
	.w1(32'hb7ef4f4f),
	.w2(32'hb8206186),
	.w3(32'h37823b67),
	.w4(32'hb692504f),
	.w5(32'hb7adf929),
	.w6(32'h37e033f4),
	.w7(32'hb5c03f82),
	.w8(32'hb800d423),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b20d7),
	.w1(32'h3a9261c9),
	.w2(32'h3b1d7428),
	.w3(32'hbaebf195),
	.w4(32'h3ae7140a),
	.w5(32'h3b9165c3),
	.w6(32'hbb42036a),
	.w7(32'h39ab75a0),
	.w8(32'h3b4a34bb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule