module layer_6_featuremap_13(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494e6a),
	.w1(32'h3a13b7bc),
	.w2(32'h3c974f4e),
	.w3(32'h3aad5633),
	.w4(32'hbba87122),
	.w5(32'hbb5ee190),
	.w6(32'hbc050635),
	.w7(32'h3c50ca41),
	.w8(32'hbbe8cb14),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf1b1a),
	.w1(32'h3b8ce6b4),
	.w2(32'h39b075aa),
	.w3(32'hbbd4488e),
	.w4(32'hbb89aa59),
	.w5(32'hbbc6b92d),
	.w6(32'hba4df33b),
	.w7(32'hbb8040ee),
	.w8(32'hb950ff5c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2cd2),
	.w1(32'h3bd5f6bb),
	.w2(32'hbb6b9cb8),
	.w3(32'hbb0b25de),
	.w4(32'h3bbae003),
	.w5(32'hbc0b6372),
	.w6(32'h3c467da0),
	.w7(32'h3ba4083d),
	.w8(32'hbc924434),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1ffc1),
	.w1(32'h3ba70f76),
	.w2(32'h3b978808),
	.w3(32'hbc9c1999),
	.w4(32'h3a188dae),
	.w5(32'h3aa906e4),
	.w6(32'hbb0eb987),
	.w7(32'hbbf25334),
	.w8(32'hbc2a56d6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37b35a),
	.w1(32'hb8d53032),
	.w2(32'h3b18431f),
	.w3(32'hbb21c0d6),
	.w4(32'h3b2adb3e),
	.w5(32'h3bbf6dcd),
	.w6(32'hb9642d4a),
	.w7(32'h3b0852a4),
	.w8(32'h3a8310bb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e89e31),
	.w1(32'h3ba2568a),
	.w2(32'hbca2b99e),
	.w3(32'h3b5df834),
	.w4(32'hbb9c5d47),
	.w5(32'hbc96ca01),
	.w6(32'h3bb035b5),
	.w7(32'hbc0798bb),
	.w8(32'h3a56a829),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b6e0),
	.w1(32'h3c3f4753),
	.w2(32'h3c82fdbb),
	.w3(32'hbb919ba8),
	.w4(32'h3c14ac47),
	.w5(32'h3c533a17),
	.w6(32'h3bea4fc8),
	.w7(32'h3c52a2dd),
	.w8(32'h3c0cb61c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52bcee),
	.w1(32'h3b456864),
	.w2(32'hbc758b4e),
	.w3(32'h3c328a80),
	.w4(32'hbac5ffce),
	.w5(32'hbc4c00db),
	.w6(32'h3abdb049),
	.w7(32'hbbf2c3d8),
	.w8(32'hbd1595aa),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd230724),
	.w1(32'hbc1af6d3),
	.w2(32'hbbd5a3d1),
	.w3(32'hbcd6b815),
	.w4(32'hbba5425d),
	.w5(32'hbb6a590f),
	.w6(32'hbbe630a5),
	.w7(32'hbb798b5a),
	.w8(32'hbb62b9bd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60034),
	.w1(32'h3c14f10e),
	.w2(32'h3c6198c3),
	.w3(32'hb93c3c28),
	.w4(32'h3bf5ab01),
	.w5(32'h3c3a6666),
	.w6(32'h3be6514d),
	.w7(32'h3c422776),
	.w8(32'h3b82f418),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7e02d),
	.w1(32'h3ba9adad),
	.w2(32'hbbdea2e1),
	.w3(32'h3b95adaa),
	.w4(32'h3baba4cb),
	.w5(32'h38d47ca0),
	.w6(32'h3bcc37b4),
	.w7(32'hbb16d9f9),
	.w8(32'h3b9422f2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e26f),
	.w1(32'h3be2c180),
	.w2(32'hbbd6228a),
	.w3(32'h3bbe0684),
	.w4(32'hba838fbe),
	.w5(32'hbc3e257b),
	.w6(32'h3bf6a7d7),
	.w7(32'hbc05e943),
	.w8(32'h3bac8ab0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9373e),
	.w1(32'h3bd62493),
	.w2(32'h3afb6765),
	.w3(32'hbb8aba2a),
	.w4(32'h3baa4527),
	.w5(32'h3bb66da8),
	.w6(32'h3c725d12),
	.w7(32'h3c908081),
	.w8(32'hbb409722),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca643c6),
	.w1(32'h3b8e2e66),
	.w2(32'h3b3a2c70),
	.w3(32'hbc3e78df),
	.w4(32'h3ba377b6),
	.w5(32'hbb81a1d7),
	.w6(32'h3b70aad1),
	.w7(32'hbb08521c),
	.w8(32'hbac0c387),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61938f),
	.w1(32'hba7a13f8),
	.w2(32'hbb62ad1a),
	.w3(32'hba9b37d0),
	.w4(32'h3a4ce581),
	.w5(32'hbae55289),
	.w6(32'h3c08ded8),
	.w7(32'h395c05e5),
	.w8(32'h3bbf57b6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b189),
	.w1(32'h3ae74cd3),
	.w2(32'hbccd71df),
	.w3(32'h3bb0048b),
	.w4(32'h3b438a8b),
	.w5(32'hbc5f0e87),
	.w6(32'h3c0ca748),
	.w7(32'hbc871d00),
	.w8(32'h3b99fb32),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dbb72),
	.w1(32'hbc00b4f4),
	.w2(32'h3c07d4bb),
	.w3(32'h3bfa337c),
	.w4(32'hbafaf810),
	.w5(32'h3c153afe),
	.w6(32'hbbb84def),
	.w7(32'h3c01a2e7),
	.w8(32'hbc995d12),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a74ad),
	.w1(32'hb9fa07e1),
	.w2(32'hbc4d7323),
	.w3(32'h3b4d07ae),
	.w4(32'h3ba28226),
	.w5(32'hb9c69039),
	.w6(32'h3b53de2a),
	.w7(32'hbb19a25d),
	.w8(32'hbb8dbc0c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c26f24),
	.w1(32'hbbbc849c),
	.w2(32'hbb1f4fab),
	.w3(32'h3b69f738),
	.w4(32'hbb3938a1),
	.w5(32'h391b683f),
	.w6(32'hbb9ae1ee),
	.w7(32'hbb29c187),
	.w8(32'hbc0358cb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea68b3),
	.w1(32'h3b4b421d),
	.w2(32'hbcd9f08a),
	.w3(32'hbba5d212),
	.w4(32'hbb7d0bd7),
	.w5(32'hbce2b4d1),
	.w6(32'h3ba777ba),
	.w7(32'hbc1f0b4a),
	.w8(32'h3c80f7d5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84980a),
	.w1(32'hbbf06ff7),
	.w2(32'hbc5747f1),
	.w3(32'hbc10749e),
	.w4(32'hbbc34475),
	.w5(32'hbb758c56),
	.w6(32'hbafb4740),
	.w7(32'hbb2e3c0b),
	.w8(32'h3c9bfda6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c044e),
	.w1(32'hbb9306a6),
	.w2(32'hbb129386),
	.w3(32'h3b5ae5fd),
	.w4(32'hba99fff8),
	.w5(32'h3b38aeb0),
	.w6(32'hbb85b0d9),
	.w7(32'hbb7feed9),
	.w8(32'h3bb215b5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2bf77),
	.w1(32'h3ae324a3),
	.w2(32'hbb50beb8),
	.w3(32'h3b373404),
	.w4(32'h3b817eb7),
	.w5(32'h371b5def),
	.w6(32'hba067a69),
	.w7(32'hbb9f3e5b),
	.w8(32'hbb2b9bb2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f9a3),
	.w1(32'h3c40bd9a),
	.w2(32'h3d0bdf94),
	.w3(32'h3b8f635c),
	.w4(32'hbc0163b6),
	.w5(32'h3b8034fa),
	.w6(32'h3bdcf6f7),
	.w7(32'h3d00dd64),
	.w8(32'h3d43b8cd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ad24f),
	.w1(32'hb95d29f8),
	.w2(32'h3c205046),
	.w3(32'h3c3809a2),
	.w4(32'hbbfa0f81),
	.w5(32'hbb295524),
	.w6(32'h3b5245c1),
	.w7(32'h3c05ff83),
	.w8(32'hbc001957),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0a162),
	.w1(32'h3a7c13c4),
	.w2(32'hbbd5f5b8),
	.w3(32'hbbf6d8fa),
	.w4(32'h3bfd4926),
	.w5(32'hbaa78ab0),
	.w6(32'h3b76780b),
	.w7(32'h3b18ec1c),
	.w8(32'hb90fb2b7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23b99a),
	.w1(32'hba306e0f),
	.w2(32'hbc144ade),
	.w3(32'hb9ef1838),
	.w4(32'hbbdf4baf),
	.w5(32'hbbf1a8cc),
	.w6(32'hbb21bb9e),
	.w7(32'hbc00224b),
	.w8(32'h3c961a88),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96fc46),
	.w1(32'h3a4ce080),
	.w2(32'hbc66522c),
	.w3(32'h3b02c3ab),
	.w4(32'h3b1cf702),
	.w5(32'hbc9b1c83),
	.w6(32'h3c45bf51),
	.w7(32'hbaa82cf3),
	.w8(32'h3c1b949a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bdae6),
	.w1(32'h3b2bc813),
	.w2(32'hbb651158),
	.w3(32'hbbb613a7),
	.w4(32'h3b47caa9),
	.w5(32'hbae12788),
	.w6(32'h3b9b557a),
	.w7(32'hb943854f),
	.w8(32'hbbc42155),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca10f19),
	.w1(32'h3c481835),
	.w2(32'h3d04ee28),
	.w3(32'hbbee1b0c),
	.w4(32'hbad4279a),
	.w5(32'h3c4c1d35),
	.w6(32'hb7d941df),
	.w7(32'h3cab9361),
	.w8(32'hbc0ee884),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109f7a),
	.w1(32'hbbb75744),
	.w2(32'h3ae8077e),
	.w3(32'hbb972f06),
	.w4(32'hba5c329e),
	.w5(32'hbbf22e81),
	.w6(32'hbc1526c6),
	.w7(32'hbb18c923),
	.w8(32'h3b639b04),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc206605),
	.w1(32'h3b149e33),
	.w2(32'hbc093d4d),
	.w3(32'hbba04138),
	.w4(32'h3b29e4a1),
	.w5(32'hbb974762),
	.w6(32'h3921356c),
	.w7(32'hbb38dc85),
	.w8(32'h3c0d7716),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dee2e),
	.w1(32'hb91e64f3),
	.w2(32'hbb9963ef),
	.w3(32'h3b1a7fcf),
	.w4(32'hbc566757),
	.w5(32'hbc30e624),
	.w6(32'h3bfe1b2a),
	.w7(32'h3c95665d),
	.w8(32'h3c9e36b7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbabb11),
	.w1(32'hbb2a31fe),
	.w2(32'hbba3da01),
	.w3(32'hba8628ba),
	.w4(32'hbc059fa8),
	.w5(32'hbc125331),
	.w6(32'hbb4c8fff),
	.w7(32'hbba48ba0),
	.w8(32'h39642a9c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36162c4f),
	.w1(32'hbb8df3e8),
	.w2(32'hbc07a51a),
	.w3(32'hba446e53),
	.w4(32'hbc14e8e7),
	.w5(32'hbbffc6e5),
	.w6(32'h3b5b5890),
	.w7(32'hbb29f6b2),
	.w8(32'h3b098a59),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b98d0d),
	.w1(32'h3acfebd0),
	.w2(32'hbbb68cca),
	.w3(32'hbb42c219),
	.w4(32'h3b8d905b),
	.w5(32'h3b578adb),
	.w6(32'h3b738517),
	.w7(32'h3c1e3133),
	.w8(32'hbc0444e6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46920b),
	.w1(32'h3b4b01dd),
	.w2(32'h3bc46465),
	.w3(32'hbc10ecca),
	.w4(32'h3ab8b956),
	.w5(32'h3b5f4bb1),
	.w6(32'h3910df01),
	.w7(32'h3b3de70c),
	.w8(32'h3b417c67),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43420),
	.w1(32'hbb2cc0f5),
	.w2(32'hbbbfb6ee),
	.w3(32'h3b8d4e7f),
	.w4(32'hba9cce2c),
	.w5(32'hbbe3ef1d),
	.w6(32'h3a3c80bf),
	.w7(32'hba6f360c),
	.w8(32'h3bcf54d8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e68c),
	.w1(32'h3d211131),
	.w2(32'h3d72319c),
	.w3(32'hbbd13729),
	.w4(32'h3cfc5c51),
	.w5(32'h3d44fc76),
	.w6(32'h3d01699f),
	.w7(32'h3d51c20d),
	.w8(32'h3d1f3be2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d451b5d),
	.w1(32'h3aa799ab),
	.w2(32'h3af35d1c),
	.w3(32'h3d166975),
	.w4(32'h3b95e2c9),
	.w5(32'hbab6ab2f),
	.w6(32'hbb58b395),
	.w7(32'hbb8e1acf),
	.w8(32'hba682068),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7a99),
	.w1(32'h3b01f7fa),
	.w2(32'h3b6239dd),
	.w3(32'hbb3f0433),
	.w4(32'hba2f82b3),
	.w5(32'hba766816),
	.w6(32'h3a580853),
	.w7(32'h3a00f7d6),
	.w8(32'h3a40536e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8174138),
	.w1(32'h3c9eac8f),
	.w2(32'h3cf89329),
	.w3(32'hbb085af9),
	.w4(32'h3c6d8c8b),
	.w5(32'h3cc4b325),
	.w6(32'h3c87c9e6),
	.w7(32'h3cda6d20),
	.w8(32'h3cbc84b1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd534e3),
	.w1(32'hbbd566b6),
	.w2(32'hbc84ca8b),
	.w3(32'h3ca2f2a4),
	.w4(32'hbb357cbb),
	.w5(32'hba86548c),
	.w6(32'h39e43a32),
	.w7(32'hbac2c84b),
	.w8(32'h39d9e7a6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00e2e8),
	.w1(32'hbca4bcfa),
	.w2(32'h3cc993cf),
	.w3(32'h3b917267),
	.w4(32'h3ad9f16e),
	.w5(32'hbb054252),
	.w6(32'h3ad6417d),
	.w7(32'hbcf1c736),
	.w8(32'h3c067813),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09ce72),
	.w1(32'h3c2dfd86),
	.w2(32'h3c8c6f92),
	.w3(32'hbc2fcd00),
	.w4(32'h3bc6eb8a),
	.w5(32'h3bbf2f4b),
	.w6(32'hbbd36664),
	.w7(32'hbb6e2453),
	.w8(32'h3b901a88),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6729ea),
	.w1(32'h3c151d4a),
	.w2(32'h3cc2d79e),
	.w3(32'h3ba75928),
	.w4(32'hbbb27884),
	.w5(32'hb9df803c),
	.w6(32'h3b6ac3b2),
	.w7(32'h3ced6f6b),
	.w8(32'h3cd2c73b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3af2d),
	.w1(32'hbb80658b),
	.w2(32'hbb56a0ec),
	.w3(32'hbb1601b1),
	.w4(32'h3a58f5b0),
	.w5(32'h3a890293),
	.w6(32'hbba52484),
	.w7(32'hbb9843ff),
	.w8(32'h3b9878eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1a9ab),
	.w1(32'h39eeac7a),
	.w2(32'h39fa9b9f),
	.w3(32'h3c2a54d7),
	.w4(32'hbbb98cff),
	.w5(32'hb9518cbe),
	.w6(32'hbb97fe37),
	.w7(32'h3b81dc5e),
	.w8(32'h3ba31e9b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ac3aa),
	.w1(32'hbb809ec6),
	.w2(32'h3b87881c),
	.w3(32'h3b454946),
	.w4(32'h3a8bb592),
	.w5(32'h3b366cb2),
	.w6(32'h3b3cae35),
	.w7(32'h3b91a072),
	.w8(32'hb9fe1426),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63cf7c),
	.w1(32'hbc2bb7ff),
	.w2(32'hbbb2393e),
	.w3(32'h3a33e27d),
	.w4(32'hbbcb94cc),
	.w5(32'h3b7b080f),
	.w6(32'hbc123df1),
	.w7(32'hbc2aa18e),
	.w8(32'h3c168e57),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7edd9a),
	.w1(32'hbb3b8991),
	.w2(32'h3a70e3c5),
	.w3(32'h3becf2b1),
	.w4(32'hbb18c93a),
	.w5(32'hbb146228),
	.w6(32'hbb26cfeb),
	.w7(32'hbb43ae09),
	.w8(32'hbb892021),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fae02),
	.w1(32'hbc193c38),
	.w2(32'hbb77c8d0),
	.w3(32'hbb82e052),
	.w4(32'hba60234c),
	.w5(32'hbc36a3ac),
	.w6(32'h3ba6d9e0),
	.w7(32'hbc1de26e),
	.w8(32'hbb51de7d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5780df),
	.w1(32'hbb1cd580),
	.w2(32'hbb96440e),
	.w3(32'h3b3ab71f),
	.w4(32'hbac345e0),
	.w5(32'hbb9c4056),
	.w6(32'h3b20db36),
	.w7(32'h3abf22d1),
	.w8(32'hba02ca0b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1064),
	.w1(32'hb98a2abf),
	.w2(32'h3bc40f55),
	.w3(32'hbb667474),
	.w4(32'hbb84d80a),
	.w5(32'hbb1325fc),
	.w6(32'hbb962552),
	.w7(32'hb9b5afaa),
	.w8(32'h390d3ab6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bcdf3),
	.w1(32'hbb0146ad),
	.w2(32'hbb2fc455),
	.w3(32'hbaa7d335),
	.w4(32'hbb8a4349),
	.w5(32'hbc18de63),
	.w6(32'h3c131bab),
	.w7(32'h3a533da3),
	.w8(32'h3c09ee1e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d895),
	.w1(32'hbc26ef01),
	.w2(32'hbc068201),
	.w3(32'h3ac1b334),
	.w4(32'h3bb6df03),
	.w5(32'h3b5ef364),
	.w6(32'hbb5a2174),
	.w7(32'hbbb3af6b),
	.w8(32'h3c02fd5f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a153772),
	.w1(32'hbbcc9a1f),
	.w2(32'hbb9d9996),
	.w3(32'h3c0360f9),
	.w4(32'hbbfee014),
	.w5(32'hbc251c32),
	.w6(32'h3c0a8e31),
	.w7(32'h3a7e1ab5),
	.w8(32'h39f35eb5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0744b1),
	.w1(32'hbc1765f5),
	.w2(32'h3bfbb5fc),
	.w3(32'hbba986ec),
	.w4(32'hbb99aecb),
	.w5(32'h3c20eeab),
	.w6(32'h3b8a57ad),
	.w7(32'hbbdb53b9),
	.w8(32'hba81fd06),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f371),
	.w1(32'hb9f6b89f),
	.w2(32'hbbf77430),
	.w3(32'h3b91fd06),
	.w4(32'h3b27421b),
	.w5(32'hb9b30ab4),
	.w6(32'hbabde14b),
	.w7(32'hbc1e443b),
	.w8(32'h3b56f48b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49392e),
	.w1(32'h3c1b1d32),
	.w2(32'h3c0eaf12),
	.w3(32'h3c3cd1a5),
	.w4(32'h3bef565b),
	.w5(32'hb62ef7ca),
	.w6(32'hbc2cd3d2),
	.w7(32'hbbd232b4),
	.w8(32'h3b8cc56e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afee218),
	.w1(32'hbb4078d0),
	.w2(32'h3c018c44),
	.w3(32'h3bfac88b),
	.w4(32'h3ba2e876),
	.w5(32'h3b68d9b2),
	.w6(32'h3a6caf7e),
	.w7(32'h3b947403),
	.w8(32'h3bd8c9bc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2826f9),
	.w1(32'hbc3ffdd1),
	.w2(32'hbcb71dec),
	.w3(32'h3b9cc6ba),
	.w4(32'hbb716236),
	.w5(32'hbc5bffc1),
	.w6(32'hbaa90fbd),
	.w7(32'hbc26688e),
	.w8(32'h399d0fa4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881c54),
	.w1(32'hbaf6c81a),
	.w2(32'hba10e883),
	.w3(32'h3b1f52b6),
	.w4(32'hba209003),
	.w5(32'hba1ca942),
	.w6(32'hba12592d),
	.w7(32'hba16d443),
	.w8(32'hba450f1d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53f5f8),
	.w1(32'h3b32a7f2),
	.w2(32'h3aa3c855),
	.w3(32'h3b673c0c),
	.w4(32'h3b504ec1),
	.w5(32'h3aea4503),
	.w6(32'h3b2fe34c),
	.w7(32'h3b34e202),
	.w8(32'h3b142bf3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule