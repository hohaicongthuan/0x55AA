module layer_10_featuremap_50(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2f0d),
	.w1(32'hba89e0ee),
	.w2(32'hbb9fde7b),
	.w3(32'h3c5e28a6),
	.w4(32'hbb5baf87),
	.w5(32'hbb8783c0),
	.w6(32'h3c154765),
	.w7(32'hbc66870e),
	.w8(32'hbc330423),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f6856),
	.w1(32'hbc86c61b),
	.w2(32'hbc9e7434),
	.w3(32'hbc2fb64b),
	.w4(32'hbc651531),
	.w5(32'hbc172864),
	.w6(32'hbc925c36),
	.w7(32'hbb950105),
	.w8(32'h3c0ccbfb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dd851),
	.w1(32'hbbce9541),
	.w2(32'hbc2004a0),
	.w3(32'h3ca0858a),
	.w4(32'h3c04ba7d),
	.w5(32'hbc5bc7e3),
	.w6(32'h3c7de403),
	.w7(32'hbab3d4dc),
	.w8(32'h3bcf07d0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b16d4),
	.w1(32'hbc0226cd),
	.w2(32'h3bd4648b),
	.w3(32'hba83cc36),
	.w4(32'hbb42084f),
	.w5(32'hbab38520),
	.w6(32'h3bbe55a7),
	.w7(32'h3b81e2c5),
	.w8(32'hbc93c025),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e7c8),
	.w1(32'hbae3eb60),
	.w2(32'hbc03f583),
	.w3(32'hbc3687de),
	.w4(32'hbbeef8c3),
	.w5(32'hbc68fe19),
	.w6(32'hbb64bad2),
	.w7(32'hbc01d7e6),
	.w8(32'h3b6d5f65),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d3879),
	.w1(32'hbbe3b178),
	.w2(32'hbc021432),
	.w3(32'h3c25991d),
	.w4(32'h3c2ee5e2),
	.w5(32'hbbe1dbe0),
	.w6(32'h3ccf07b8),
	.w7(32'h3c75d51e),
	.w8(32'hbb9385f5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ebac),
	.w1(32'hbb9e563f),
	.w2(32'h3c3cdc25),
	.w3(32'hbb0b6d09),
	.w4(32'h3aa496a0),
	.w5(32'h3bfd66fe),
	.w6(32'h3abddf70),
	.w7(32'hbb3b2e2f),
	.w8(32'hbc56616c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9104a7),
	.w1(32'h3adb814b),
	.w2(32'h3b5e0dad),
	.w3(32'hbb9dbfb8),
	.w4(32'hbc75b0c0),
	.w5(32'h3c25a53b),
	.w6(32'hbba8a4c7),
	.w7(32'h3b352142),
	.w8(32'h3be4f048),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1819d2),
	.w1(32'h3b2115ab),
	.w2(32'hbbab2b7a),
	.w3(32'h3ba43bae),
	.w4(32'h3bc43810),
	.w5(32'h3b678835),
	.w6(32'hbb7300da),
	.w7(32'hbb77f6c2),
	.w8(32'h3a6aae78),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03dc7b),
	.w1(32'hb9a27425),
	.w2(32'hba0a70ce),
	.w3(32'hbba3c7f9),
	.w4(32'h3bae687b),
	.w5(32'hba69de21),
	.w6(32'h3b2ed79f),
	.w7(32'h3c4ce439),
	.w8(32'hbaad8cb6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5495b9),
	.w1(32'hbb1fa216),
	.w2(32'hbc49d079),
	.w3(32'hbadbc592),
	.w4(32'hbadd5f06),
	.w5(32'hbc9f862b),
	.w6(32'hbb316d2d),
	.w7(32'hba0f780b),
	.w8(32'h3c32db9e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc863fac),
	.w1(32'hbbd27333),
	.w2(32'h3b111579),
	.w3(32'hbc3b5ada),
	.w4(32'hbbef6da1),
	.w5(32'h3b067138),
	.w6(32'h3c6ae5b3),
	.w7(32'h3b603d43),
	.w8(32'hbb013703),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3b926),
	.w1(32'h3b3b3518),
	.w2(32'h3c36c37e),
	.w3(32'hba0b0cc8),
	.w4(32'h3b2b9919),
	.w5(32'h3c1b866a),
	.w6(32'hba657643),
	.w7(32'hba3d9e51),
	.w8(32'h3b0bac56),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a5246),
	.w1(32'hbb988d2c),
	.w2(32'hbc1a52fd),
	.w3(32'h3bffa5e4),
	.w4(32'hbc227d66),
	.w5(32'hbbc95f9a),
	.w6(32'h3ad24024),
	.w7(32'hbb3099e9),
	.w8(32'hbc3e8113),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac62f30),
	.w1(32'h3b97b4df),
	.w2(32'hbb97bf80),
	.w3(32'hbc1707cf),
	.w4(32'hba5bc31e),
	.w5(32'hbb8a78e6),
	.w6(32'hbbbc6d70),
	.w7(32'hbbd0d7bf),
	.w8(32'hbae34a71),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882be16),
	.w1(32'hb9a9109f),
	.w2(32'hbab2c772),
	.w3(32'h3a16d9a0),
	.w4(32'hbbcdc3cc),
	.w5(32'hba63c8d5),
	.w6(32'hbac2aa86),
	.w7(32'hb8f049d9),
	.w8(32'hba2a4a2c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7df6),
	.w1(32'hbb0f7161),
	.w2(32'h39c88387),
	.w3(32'h39c035c4),
	.w4(32'hba22310c),
	.w5(32'hb9fa79a4),
	.w6(32'h38972fcd),
	.w7(32'hba354548),
	.w8(32'hbb3e4bd2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87eef4),
	.w1(32'h3c165488),
	.w2(32'h3c559a3b),
	.w3(32'h3ba3f09c),
	.w4(32'h3bbc5dfb),
	.w5(32'h3c83e256),
	.w6(32'h3beee36d),
	.w7(32'h3b7244c9),
	.w8(32'h3c6959cc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a50cd),
	.w1(32'h3bafd0f9),
	.w2(32'h3b660b4b),
	.w3(32'h3bb53aab),
	.w4(32'h3b1ce26e),
	.w5(32'h3bde5324),
	.w6(32'h3c4b799f),
	.w7(32'h3be51164),
	.w8(32'h3c287d5f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba124d6),
	.w1(32'hbbb98c2a),
	.w2(32'h3b09335c),
	.w3(32'hbae612ad),
	.w4(32'hbbb98abc),
	.w5(32'hbbf85c80),
	.w6(32'hbc353a80),
	.w7(32'hbbf4f489),
	.w8(32'hbc23addc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf97d6a),
	.w1(32'hbbc85fbc),
	.w2(32'hbbfa726c),
	.w3(32'hbc5141aa),
	.w4(32'hbbbaacf6),
	.w5(32'hbc370d9f),
	.w6(32'hbbd61b9c),
	.w7(32'h3b0df426),
	.w8(32'hbb61eb0b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25a341),
	.w1(32'hbc164388),
	.w2(32'hbbdf2983),
	.w3(32'hbc17fccf),
	.w4(32'hbc0423b5),
	.w5(32'hbbd3eedd),
	.w6(32'hbc95f8c4),
	.w7(32'hbcc2c0e4),
	.w8(32'h3baf7614),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ae412),
	.w1(32'h3c2f1670),
	.w2(32'h3c37650b),
	.w3(32'h3cab0361),
	.w4(32'h3c307519),
	.w5(32'h3c1b57e2),
	.w6(32'h3c9f2f48),
	.w7(32'h3bb360c2),
	.w8(32'h3c8f9654),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce284c),
	.w1(32'h3b500f69),
	.w2(32'h3bdbd9e9),
	.w3(32'h398ce48d),
	.w4(32'h3b37429c),
	.w5(32'h3a9ba830),
	.w6(32'hbaa75397),
	.w7(32'h39b3fdaf),
	.w8(32'hbbbc5462),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c216de8),
	.w1(32'hbc1c042b),
	.w2(32'hbcd27cca),
	.w3(32'hb9a2ec71),
	.w4(32'hbc45fda0),
	.w5(32'h3c3db2d4),
	.w6(32'hb86f4382),
	.w7(32'hbc104ecf),
	.w8(32'hbb4f397f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d3b93),
	.w1(32'h3b9d9359),
	.w2(32'h3c672c94),
	.w3(32'h3ca62504),
	.w4(32'h3a53f39d),
	.w5(32'h3cd156ed),
	.w6(32'h3b935510),
	.w7(32'hba5f923a),
	.w8(32'hbbcb698e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb57b6),
	.w1(32'h3c5942c0),
	.w2(32'hb9c5ccec),
	.w3(32'h3c4ba049),
	.w4(32'hbc45aa4e),
	.w5(32'hb92041c8),
	.w6(32'hbc5a3198),
	.w7(32'hbc344b40),
	.w8(32'hb91ac1cf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00332f),
	.w1(32'hba74282f),
	.w2(32'hbb36929b),
	.w3(32'h3b91ec85),
	.w4(32'h399debc7),
	.w5(32'hbbe0ce23),
	.w6(32'hbb5cb3b7),
	.w7(32'hba00fdac),
	.w8(32'hbb901848),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46c48),
	.w1(32'hbb90499b),
	.w2(32'hbc032d9a),
	.w3(32'hbb0546f5),
	.w4(32'h3b06b1ce),
	.w5(32'h3c2d9215),
	.w6(32'hbba49f25),
	.w7(32'hba8cb04e),
	.w8(32'hbbb39126),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc679980),
	.w1(32'hbc1d602b),
	.w2(32'hbc08fa4a),
	.w3(32'h3d117807),
	.w4(32'h3d262c5a),
	.w5(32'hbbccbcf1),
	.w6(32'h3d70e0ee),
	.w7(32'h3d6ead83),
	.w8(32'hbc47aeb9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb680885),
	.w1(32'hbb968915),
	.w2(32'h3b4a7b43),
	.w3(32'h3b29353b),
	.w4(32'h3b2c3392),
	.w5(32'h3b11425a),
	.w6(32'hbb847a37),
	.w7(32'hbb91cfa6),
	.w8(32'hbb2368ad),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c6a12),
	.w1(32'h3bfb7844),
	.w2(32'hbba95408),
	.w3(32'h3ba64671),
	.w4(32'h3c98e2f8),
	.w5(32'h39b4e4bc),
	.w6(32'h3c0478a4),
	.w7(32'h3b88d06e),
	.w8(32'hbb2728fe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a3a9),
	.w1(32'hbbcfa77f),
	.w2(32'h3b09537d),
	.w3(32'h3bf7489e),
	.w4(32'h3bceacf1),
	.w5(32'h3a21f642),
	.w6(32'h3b3d8d47),
	.w7(32'h3c4f8add),
	.w8(32'hbb94f132),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c9563),
	.w1(32'hbbcc55fb),
	.w2(32'hbc0d416d),
	.w3(32'h3adb01e9),
	.w4(32'hbb0de37e),
	.w5(32'hbbb18c25),
	.w6(32'hbc22db9e),
	.w7(32'hbbd80ac9),
	.w8(32'h3ae74fb7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03c224),
	.w1(32'hbb10a878),
	.w2(32'hb92fe1ee),
	.w3(32'hbc875b01),
	.w4(32'hbc98a6d6),
	.w5(32'hbbb9ad0d),
	.w6(32'h3c746286),
	.w7(32'h3c111d9f),
	.w8(32'hba91ff75),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b187e),
	.w1(32'hbab1542e),
	.w2(32'hbc2e30a1),
	.w3(32'hbbe12065),
	.w4(32'hbbc38552),
	.w5(32'h3ba24d5b),
	.w6(32'hbaaea12c),
	.w7(32'hbac6fcef),
	.w8(32'h3cdf6f2d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc993cf1),
	.w1(32'hbc34dfaa),
	.w2(32'h3b88004b),
	.w3(32'h3c38756d),
	.w4(32'h3c81f5c1),
	.w5(32'h3bcb54fa),
	.w6(32'h3d08588b),
	.w7(32'hbb137fec),
	.w8(32'h3906a7f4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25bc6c),
	.w1(32'hbc08d946),
	.w2(32'hbc854597),
	.w3(32'h3c37cde9),
	.w4(32'h3a1840e8),
	.w5(32'hbc8b2c68),
	.w6(32'hbc3ba087),
	.w7(32'hbc379ee5),
	.w8(32'hbce7faae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb178b1),
	.w1(32'hbbd9ec85),
	.w2(32'hba827b3d),
	.w3(32'h3c8000c1),
	.w4(32'h3b9a1cdd),
	.w5(32'hbbc55856),
	.w6(32'hbd35a1ca),
	.w7(32'hbcf53170),
	.w8(32'hbbf5c873),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ebec),
	.w1(32'h3b3f3e47),
	.w2(32'h3b71a5e6),
	.w3(32'hbc1f0587),
	.w4(32'hba8d4ff6),
	.w5(32'h3a30ad63),
	.w6(32'hbaefde48),
	.w7(32'hbc07c6be),
	.w8(32'h3a9a0835),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9ef37),
	.w1(32'h3b7ce50c),
	.w2(32'h3b111e59),
	.w3(32'h3b019e6a),
	.w4(32'h3b6d36ca),
	.w5(32'hbc8ae07d),
	.w6(32'h3c903e9a),
	.w7(32'h3c81684f),
	.w8(32'hbc1fcd67),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1873f),
	.w1(32'hbba829d8),
	.w2(32'hbb290932),
	.w3(32'hbc83b9f5),
	.w4(32'hbc32d9de),
	.w5(32'h3ba5da35),
	.w6(32'hbc1aab7a),
	.w7(32'hbaf3855e),
	.w8(32'hbabc9981),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98157cd),
	.w1(32'hbb27fb56),
	.w2(32'hbb5a51e5),
	.w3(32'h3c3dae77),
	.w4(32'h3c53c9ec),
	.w5(32'hbba80d13),
	.w6(32'h3c2a563d),
	.w7(32'h3bef62c5),
	.w8(32'hbb67e1f5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7c49c),
	.w1(32'h3a529ed4),
	.w2(32'hbb4ab79a),
	.w3(32'hbb1f1a3e),
	.w4(32'h3b289266),
	.w5(32'hba07796b),
	.w6(32'h3ac13543),
	.w7(32'h3ace7b8a),
	.w8(32'hbc21136d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d84b),
	.w1(32'hbc80d593),
	.w2(32'h3bb0d123),
	.w3(32'hbca53d4e),
	.w4(32'hbca8f7d9),
	.w5(32'hbc87bf3d),
	.w6(32'h3ca99c12),
	.w7(32'h3c581c21),
	.w8(32'hbc2b0a3f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dc968),
	.w1(32'hbaa120e0),
	.w2(32'h3c476647),
	.w3(32'hbccc333a),
	.w4(32'hbcb52b9e),
	.w5(32'hbb4a4c92),
	.w6(32'h3c626c7b),
	.w7(32'h3c967b56),
	.w8(32'h3c0ca837),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93653a),
	.w1(32'h3ab5b2c8),
	.w2(32'h3ba09d69),
	.w3(32'hbbdd1b4a),
	.w4(32'h3b611a08),
	.w5(32'hbc2cb570),
	.w6(32'h3cc0a5f5),
	.w7(32'h3cf9c92e),
	.w8(32'hba46c625),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2e737),
	.w1(32'h3c15baca),
	.w2(32'h3caa2afa),
	.w3(32'hbc7930d2),
	.w4(32'hba701b08),
	.w5(32'h3c923fd3),
	.w6(32'h3ccf3f00),
	.w7(32'h3d2f4537),
	.w8(32'h3c899c11),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66d14e),
	.w1(32'hba1f56fd),
	.w2(32'h3c04fac8),
	.w3(32'hbae6b6be),
	.w4(32'hbba1593a),
	.w5(32'hba226316),
	.w6(32'h3b10386f),
	.w7(32'hba942efb),
	.w8(32'hbc1258aa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f56c9),
	.w1(32'h3b9544b0),
	.w2(32'hbb870426),
	.w3(32'h3b1c4263),
	.w4(32'hbbc20d5f),
	.w5(32'hbbc2c186),
	.w6(32'hbc3c9755),
	.w7(32'hbca832ba),
	.w8(32'hbaa2f296),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28539a),
	.w1(32'hbb8d9c59),
	.w2(32'h3b7cea01),
	.w3(32'hbc8755c4),
	.w4(32'hbc971671),
	.w5(32'hbb935d53),
	.w6(32'h3b9a938c),
	.w7(32'h3b38548a),
	.w8(32'hbaf2993e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de560),
	.w1(32'hbc73ccae),
	.w2(32'hb991c0e8),
	.w3(32'hbbeec652),
	.w4(32'hbc2ef138),
	.w5(32'h3b249202),
	.w6(32'h3c7ac221),
	.w7(32'h3abe4e81),
	.w8(32'h3b1be891),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d243f),
	.w1(32'hba02eb12),
	.w2(32'h3c7e1e42),
	.w3(32'hb9c0a844),
	.w4(32'hbb4f3fcf),
	.w5(32'h3a9231cf),
	.w6(32'h3b8a7bef),
	.w7(32'h3b54b576),
	.w8(32'hbb658436),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1370ae),
	.w1(32'h3cc26963),
	.w2(32'h3c48d2f5),
	.w3(32'hb9ea7148),
	.w4(32'hbb307680),
	.w5(32'h3c7ff4e5),
	.w6(32'hbbbc3d43),
	.w7(32'h3a42efc4),
	.w8(32'h3c9c478a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5213ce),
	.w1(32'h3b11d40f),
	.w2(32'hbbf63dba),
	.w3(32'h3ce10068),
	.w4(32'h3c79b2a0),
	.w5(32'hbb5916ff),
	.w6(32'hbc18196a),
	.w7(32'hbc22108b),
	.w8(32'hbcb15d55),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b9144),
	.w1(32'hba9a7019),
	.w2(32'h3badb9d8),
	.w3(32'hbc4f1ccf),
	.w4(32'hbc6d0c0f),
	.w5(32'hbc84879e),
	.w6(32'hbc8b00fc),
	.w7(32'hbc948e5d),
	.w8(32'hbb6010e7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b44e2),
	.w1(32'hbbc7cc00),
	.w2(32'h399ed174),
	.w3(32'hbc8a6e16),
	.w4(32'h3aa299cb),
	.w5(32'hbb71d623),
	.w6(32'hbb757b7b),
	.w7(32'hbb939522),
	.w8(32'hbbced024),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e1918),
	.w1(32'h3c36059e),
	.w2(32'hb9ef0a0d),
	.w3(32'hbb08530a),
	.w4(32'h3bb11480),
	.w5(32'hbba43c8d),
	.w6(32'hbb075a94),
	.w7(32'h3ac00456),
	.w8(32'hb98a7eb5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c6047),
	.w1(32'hb7074538),
	.w2(32'h3b11a2c9),
	.w3(32'h3adf90fb),
	.w4(32'h3b1f11f7),
	.w5(32'hb9648ecd),
	.w6(32'h3b6c799e),
	.w7(32'h3c535b23),
	.w8(32'h3be48faa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222080),
	.w1(32'h3b17c339),
	.w2(32'h3c839d70),
	.w3(32'hba5cd72f),
	.w4(32'hbc01b3de),
	.w5(32'hba82c5c7),
	.w6(32'h3c600fd5),
	.w7(32'h3aa77378),
	.w8(32'h3b26c27d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32b43b),
	.w1(32'h3c2a8ba5),
	.w2(32'h3c273aa1),
	.w3(32'hbbf2a773),
	.w4(32'hbc080f46),
	.w5(32'hbc6cbdab),
	.w6(32'h3bd5a869),
	.w7(32'h3b296647),
	.w8(32'hbc22823b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1abdf4),
	.w1(32'hbc1ebf81),
	.w2(32'h3c5a26bd),
	.w3(32'hbc1ea1c2),
	.w4(32'h39b2a546),
	.w5(32'h3b3bda4b),
	.w6(32'hbb057079),
	.w7(32'h3bb4eae8),
	.w8(32'h3c2f991d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c133b9d),
	.w1(32'hbb678312),
	.w2(32'hbbe7a93e),
	.w3(32'hbbba83d0),
	.w4(32'hbc032ac6),
	.w5(32'hbabc063b),
	.w6(32'h3b6dce23),
	.w7(32'hbac02592),
	.w8(32'hbbc8a380),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c5f1),
	.w1(32'hbb7f5ea7),
	.w2(32'hb96027ea),
	.w3(32'h3b3b97b0),
	.w4(32'h3afbec72),
	.w5(32'hbb3b8611),
	.w6(32'hbc130378),
	.w7(32'hbb91cfb0),
	.w8(32'hbb33fc07),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b9d97),
	.w1(32'hbbb7037c),
	.w2(32'hb964b850),
	.w3(32'h3b8df633),
	.w4(32'h3bb3721b),
	.w5(32'hbb1f0bab),
	.w6(32'hbbed45f6),
	.w7(32'hbbafdfdf),
	.w8(32'hba0fced8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2754ad),
	.w1(32'h3b780e75),
	.w2(32'hbab18020),
	.w3(32'hbbdfa580),
	.w4(32'hba2c8de8),
	.w5(32'hbb4cda62),
	.w6(32'hbbfcd8f3),
	.w7(32'hbb537f42),
	.w8(32'hbc1e32a1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88aee0),
	.w1(32'hbb992f4a),
	.w2(32'h3b3612f6),
	.w3(32'h3a85118e),
	.w4(32'h3ad3b6ca),
	.w5(32'hba992ab6),
	.w6(32'hbc37228c),
	.w7(32'hbb9dd9a7),
	.w8(32'h3b96817a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ede9b),
	.w1(32'h3b4af9b8),
	.w2(32'h3b8054ab),
	.w3(32'hbb8f9408),
	.w4(32'hbb725e36),
	.w5(32'hbb3e5f91),
	.w6(32'h3c1c0e6a),
	.w7(32'h3bd0300e),
	.w8(32'hbbb39c3d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1743b3),
	.w1(32'h3c49b02d),
	.w2(32'h3b72bac8),
	.w3(32'h3b9416e5),
	.w4(32'hba05342e),
	.w5(32'h3b623578),
	.w6(32'h3a7431d0),
	.w7(32'h3abc122d),
	.w8(32'h3b5757a7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5023a3),
	.w1(32'hbc2a8d16),
	.w2(32'hbb831efa),
	.w3(32'hbc47a526),
	.w4(32'hbc199e1c),
	.w5(32'hbc052157),
	.w6(32'hbc72a0e0),
	.w7(32'hbc289acb),
	.w8(32'hbb8221ae),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2394),
	.w1(32'h39c5f520),
	.w2(32'h3a544699),
	.w3(32'hbc3951af),
	.w4(32'hbc203a41),
	.w5(32'hbbee317a),
	.w6(32'hbbb3c2e9),
	.w7(32'hbbbbfba1),
	.w8(32'hbb4418aa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bbc19),
	.w1(32'h3b9030fc),
	.w2(32'h39800737),
	.w3(32'hbc40aa21),
	.w4(32'h3b5d88af),
	.w5(32'hbc513ff5),
	.w6(32'hbbdcc8d9),
	.w7(32'hbb8be20a),
	.w8(32'h3c476bff),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15efec),
	.w1(32'hbaee60bd),
	.w2(32'hbbfed3e8),
	.w3(32'hbbdcce48),
	.w4(32'hbb787bd1),
	.w5(32'h3bf68acc),
	.w6(32'h3cc42e01),
	.w7(32'h3c6c9a5d),
	.w8(32'hbc08f233),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8efe78),
	.w1(32'hbc64b625),
	.w2(32'hbb3df525),
	.w3(32'h3cd1470b),
	.w4(32'h3ca6a92a),
	.w5(32'hbb20fbf6),
	.w6(32'hbc7f5872),
	.w7(32'hbb8c548b),
	.w8(32'hbb946efb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c4ba),
	.w1(32'hbb89e4ca),
	.w2(32'hbb348095),
	.w3(32'hbb389981),
	.w4(32'hbb197215),
	.w5(32'hbba7de82),
	.w6(32'hbb96550c),
	.w7(32'hbbbea206),
	.w8(32'hbb14d8eb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55708f),
	.w1(32'h3b34fb72),
	.w2(32'h3c103cf4),
	.w3(32'hbb5d9e3e),
	.w4(32'hbb819804),
	.w5(32'h3c7ab5c8),
	.w6(32'hba1014e5),
	.w7(32'hbacf0236),
	.w8(32'h3b16ea15),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec2ebc),
	.w1(32'h3bcae837),
	.w2(32'h3b84256f),
	.w3(32'h3c6ae204),
	.w4(32'h3c37ba21),
	.w5(32'h3c092c47),
	.w6(32'h3be0cbe8),
	.w7(32'h3bffef2d),
	.w8(32'h3c110d5d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc475042),
	.w1(32'hbc2087d1),
	.w2(32'hba5fe712),
	.w3(32'hbb1e9bdf),
	.w4(32'hbbbfadc2),
	.w5(32'hbc236b83),
	.w6(32'h3c2514ba),
	.w7(32'h3b9b6a40),
	.w8(32'h3c1e352e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a250501),
	.w1(32'h3a14a3df),
	.w2(32'h3ba395d9),
	.w3(32'hbbe75380),
	.w4(32'hbb7439b7),
	.w5(32'h3b90c93b),
	.w6(32'h3c223c3e),
	.w7(32'hbb2be5cd),
	.w8(32'h3ba80a3f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80746b),
	.w1(32'h3b568598),
	.w2(32'h3a56180a),
	.w3(32'h3c24ae7b),
	.w4(32'h3b6fec1f),
	.w5(32'h3a0a73f2),
	.w6(32'h3bb0d9fb),
	.w7(32'h3b44639f),
	.w8(32'hbb9cb23c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397bf7b6),
	.w1(32'hba8f418a),
	.w2(32'hbb0c2124),
	.w3(32'hbbfa1d58),
	.w4(32'hbc2a9f61),
	.w5(32'hbb314da5),
	.w6(32'h38ae58be),
	.w7(32'h3ab86620),
	.w8(32'hbb9a7fd0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7d4b1),
	.w1(32'h3b4a26c0),
	.w2(32'hbc085298),
	.w3(32'h3b86faf2),
	.w4(32'h3bd0514a),
	.w5(32'hbc2a90b6),
	.w6(32'hbb1481b5),
	.w7(32'h3a64596e),
	.w8(32'h3cd95221),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60f4c0),
	.w1(32'hbbe5e761),
	.w2(32'hba19a95c),
	.w3(32'hbc325388),
	.w4(32'h3b8b8907),
	.w5(32'hbbdf4693),
	.w6(32'h3d1795d1),
	.w7(32'h3cbe58db),
	.w8(32'h3a781a9b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2ac89),
	.w1(32'hbc6569d5),
	.w2(32'h3ba7b778),
	.w3(32'hbc4b862a),
	.w4(32'h3a97752d),
	.w5(32'hbbeaff4d),
	.w6(32'h3b07c89f),
	.w7(32'h3c3cc4a0),
	.w8(32'hbab73efd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a269d28),
	.w1(32'hbbda5ac5),
	.w2(32'hbc1c4623),
	.w3(32'hbc47f1c8),
	.w4(32'hba6219af),
	.w5(32'hbc7d2e8c),
	.w6(32'h3c15a3ac),
	.w7(32'h3b1e3e89),
	.w8(32'h3cf2f0d3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc913cce),
	.w1(32'hbb6e967c),
	.w2(32'h3af167de),
	.w3(32'hbb32b981),
	.w4(32'h39558182),
	.w5(32'h3b0af03e),
	.w6(32'h3d074c62),
	.w7(32'hb9b9d68d),
	.w8(32'h3b2987fd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6695f),
	.w1(32'h3b90e768),
	.w2(32'hbb82e6a5),
	.w3(32'hbb8fa50c),
	.w4(32'h3b819838),
	.w5(32'hbbf67e9f),
	.w6(32'hbb99e215),
	.w7(32'h3b128fb3),
	.w8(32'hbc0343fa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c6d96),
	.w1(32'h3b3542ec),
	.w2(32'hba945ac6),
	.w3(32'hbaae6393),
	.w4(32'hbacf4d4e),
	.w5(32'h3bf0127b),
	.w6(32'hbb8df685),
	.w7(32'h391ae19e),
	.w8(32'h3ab261b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93b5d3),
	.w1(32'h3b1c14c9),
	.w2(32'h3b925a6f),
	.w3(32'h3bfd0439),
	.w4(32'hbbde1148),
	.w5(32'h3a757f63),
	.w6(32'h3c70d917),
	.w7(32'h3c7e9902),
	.w8(32'hbc0d20a5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83283f),
	.w1(32'h3c3076a0),
	.w2(32'h3c4d3117),
	.w3(32'h3bfbf545),
	.w4(32'h3bcaa132),
	.w5(32'h3c197cdb),
	.w6(32'h3cb2cdff),
	.w7(32'h3c400a47),
	.w8(32'h3c6f613a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27d455),
	.w1(32'hb936e2b3),
	.w2(32'h3b94bf05),
	.w3(32'hbbc37f59),
	.w4(32'hbbe1d107),
	.w5(32'h3b2f030d),
	.w6(32'hbb690998),
	.w7(32'h3bf89870),
	.w8(32'h3b96f287),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9757a8),
	.w1(32'hbb8f45bc),
	.w2(32'h3b2c17fd),
	.w3(32'h3bd2af00),
	.w4(32'h39b3fd5f),
	.w5(32'h3bd31629),
	.w6(32'h3b994356),
	.w7(32'hbab177c6),
	.w8(32'h3bbe9bec),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8911af),
	.w1(32'h3b676d80),
	.w2(32'hbb06eb8a),
	.w3(32'h3c29a045),
	.w4(32'h3c060557),
	.w5(32'hbaf16f28),
	.w6(32'h3c2342eb),
	.w7(32'h3c163cfc),
	.w8(32'hbb09d66e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5958c),
	.w1(32'h3c121480),
	.w2(32'h3bf257b2),
	.w3(32'h3baa7e6d),
	.w4(32'h3bfe0ef7),
	.w5(32'h3a4b4d15),
	.w6(32'h3bdbff05),
	.w7(32'h3c112ebc),
	.w8(32'h3c0a6e90),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba0074),
	.w1(32'h3b9d3a2a),
	.w2(32'h3be77b7c),
	.w3(32'hbb873c47),
	.w4(32'hbbcf53c3),
	.w5(32'h3c869531),
	.w6(32'hbb83ca52),
	.w7(32'h3b2f32be),
	.w8(32'h3ccac31f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69cf48),
	.w1(32'h3afcfd77),
	.w2(32'h396ca22c),
	.w3(32'h3cbbc68e),
	.w4(32'h3cb13746),
	.w5(32'hbc10614f),
	.w6(32'h3dd483e9),
	.w7(32'h3dadfa73),
	.w8(32'hbcc5f82d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2080),
	.w1(32'h3b401106),
	.w2(32'h3bf9957c),
	.w3(32'hbc904deb),
	.w4(32'hbc00a853),
	.w5(32'hba616965),
	.w6(32'hbc9dadd0),
	.w7(32'hbc00bebd),
	.w8(32'h3c28fd99),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7638),
	.w1(32'hbb654522),
	.w2(32'h3c5498e2),
	.w3(32'h3beddeea),
	.w4(32'h3be29fe0),
	.w5(32'h38cc526e),
	.w6(32'h3c6b2a5a),
	.w7(32'h3c540ea1),
	.w8(32'h3b63c2f9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28d112),
	.w1(32'h3c0e6a96),
	.w2(32'h3a1c855c),
	.w3(32'hbc71e1e4),
	.w4(32'hbbabc0be),
	.w5(32'h3a70567a),
	.w6(32'hbb73e934),
	.w7(32'hbc18fc59),
	.w8(32'hbb97becf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0937e2),
	.w1(32'h3bd44e7f),
	.w2(32'h3c19d753),
	.w3(32'h3c1e1a3e),
	.w4(32'h3bec2bfe),
	.w5(32'h3ac351cc),
	.w6(32'h3c344a33),
	.w7(32'h3c09fe85),
	.w8(32'h3b697bec),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3829f),
	.w1(32'hbb924297),
	.w2(32'hbae42e54),
	.w3(32'hbbb2bde0),
	.w4(32'hbc85aff9),
	.w5(32'hbc09c3ad),
	.w6(32'h3b053a54),
	.w7(32'hbb57c91c),
	.w8(32'hbc8a6c5e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13ec33),
	.w1(32'hbc266697),
	.w2(32'hbbc7db2f),
	.w3(32'h39358cf5),
	.w4(32'hb9fa0310),
	.w5(32'hbc357b89),
	.w6(32'h3c032ade),
	.w7(32'h3c2acc07),
	.w8(32'hbbbadd91),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1432d),
	.w1(32'h3b7abc3e),
	.w2(32'h3ca95e92),
	.w3(32'hb9a1c3e0),
	.w4(32'hbc19de2f),
	.w5(32'h3b34ff94),
	.w6(32'h3b92d389),
	.w7(32'hbbf4a19c),
	.w8(32'hbc19122a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffd909),
	.w1(32'hbb23dee9),
	.w2(32'hbb9c3cfa),
	.w3(32'hbca961c9),
	.w4(32'hbcb1a1de),
	.w5(32'hbc4d4fcd),
	.w6(32'hbc83e674),
	.w7(32'hbb88561d),
	.w8(32'h3c0a0ee9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c714),
	.w1(32'h3b941fb3),
	.w2(32'h3c8494d0),
	.w3(32'hbc819e48),
	.w4(32'hbb58e043),
	.w5(32'h3c26594f),
	.w6(32'h3cc617f6),
	.w7(32'h3c8a9dcb),
	.w8(32'h3c228dc2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacca693),
	.w1(32'h3b058ac5),
	.w2(32'h3a947b04),
	.w3(32'hbc17abef),
	.w4(32'hbba7a05b),
	.w5(32'hbacc1022),
	.w6(32'hbbc3e561),
	.w7(32'hbb858328),
	.w8(32'hb9bb7fb2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831269),
	.w1(32'hba9d0689),
	.w2(32'hb9d3dc24),
	.w3(32'hbb444872),
	.w4(32'h3953731f),
	.w5(32'hbc204ce3),
	.w6(32'hbacea604),
	.w7(32'hbaa915f3),
	.w8(32'hbafac54d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406fa6),
	.w1(32'hbaf6afcc),
	.w2(32'h3b24680c),
	.w3(32'hbbe1f41f),
	.w4(32'h3b41dacb),
	.w5(32'hbc9a8f84),
	.w6(32'h38e1bdb7),
	.w7(32'hba191347),
	.w8(32'hbbcc8850),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42fae0),
	.w1(32'hbbf6d8f4),
	.w2(32'h3b03dbdf),
	.w3(32'hbcd87ea8),
	.w4(32'hbb6da1ef),
	.w5(32'hbc1e9e21),
	.w6(32'hbaedb991),
	.w7(32'hbb090fd2),
	.w8(32'hbcd72122),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2a4f),
	.w1(32'h3abdfa96),
	.w2(32'h3b640b70),
	.w3(32'hbbdaa4bd),
	.w4(32'hbbea43a6),
	.w5(32'hbc7ccac4),
	.w6(32'hbcc53468),
	.w7(32'hbcf0422b),
	.w8(32'hbba7b6cc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868215f),
	.w1(32'hbba17fb4),
	.w2(32'h3c2e6c66),
	.w3(32'hbbe3642f),
	.w4(32'hb992803f),
	.w5(32'h3b83002d),
	.w6(32'hbb0040d5),
	.w7(32'hbc2fb76b),
	.w8(32'h3c46e1db),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91ed1),
	.w1(32'h3b51fde8),
	.w2(32'h3bd3f9f7),
	.w3(32'hbbe43d7c),
	.w4(32'hbc753789),
	.w5(32'hbbc79f25),
	.w6(32'h3c831109),
	.w7(32'h3c2f441d),
	.w8(32'hbb691c7d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c829e31),
	.w1(32'h3c09b92c),
	.w2(32'h3ba2bcde),
	.w3(32'hbc5ce568),
	.w4(32'hbcb424d8),
	.w5(32'hbbee7eba),
	.w6(32'hbc6a3ed1),
	.w7(32'hbcb7d9bd),
	.w8(32'hbb06bb29),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239958),
	.w1(32'hbbda672b),
	.w2(32'h3ba3d118),
	.w3(32'hbc537f06),
	.w4(32'hba9199b3),
	.w5(32'h3b714008),
	.w6(32'h3c2e1880),
	.w7(32'h3bf43a89),
	.w8(32'h3c00099f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b254e23),
	.w1(32'hbbdd1787),
	.w2(32'h3b41b3a8),
	.w3(32'hbb01dda8),
	.w4(32'h3a5ac6e0),
	.w5(32'h399c1de0),
	.w6(32'h3bfd8ca0),
	.w7(32'h3c4db1b6),
	.w8(32'hbbc00a36),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22f0ed),
	.w1(32'h3b53fc23),
	.w2(32'hbbcbe944),
	.w3(32'h3ba64c2b),
	.w4(32'h3bd55125),
	.w5(32'hbc061d00),
	.w6(32'hbb900f4d),
	.w7(32'hba00cde2),
	.w8(32'h3b594c9f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba113794),
	.w1(32'hbba69541),
	.w2(32'h3ae71142),
	.w3(32'hbbf9f920),
	.w4(32'hbbd3d92b),
	.w5(32'h3b7a3ada),
	.w6(32'hbb096826),
	.w7(32'h3b6011c4),
	.w8(32'hbb39390f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab92ef),
	.w1(32'h3ab9affa),
	.w2(32'hba800dd3),
	.w3(32'h3c01e88f),
	.w4(32'h3b04136b),
	.w5(32'h3bd373e9),
	.w6(32'h3b0d9ffc),
	.w7(32'h3acab667),
	.w8(32'hb9240a4c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ebd7),
	.w1(32'hbb3b4364),
	.w2(32'hbb115432),
	.w3(32'h3c745c7e),
	.w4(32'h3c0cdfc1),
	.w5(32'hbb65515f),
	.w6(32'h3c416c7b),
	.w7(32'h3c3522a7),
	.w8(32'hbc31442e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb6f1c),
	.w1(32'hbc0a2802),
	.w2(32'h3bf99906),
	.w3(32'hbb4ee085),
	.w4(32'hbacb9a84),
	.w5(32'hbb6c7dd5),
	.w6(32'hbb853abc),
	.w7(32'hbc1e8167),
	.w8(32'hbbc64c93),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951841),
	.w1(32'hb9daedff),
	.w2(32'h3ba971c8),
	.w3(32'hbc27c32a),
	.w4(32'hbc11a391),
	.w5(32'h3ae841d0),
	.w6(32'h3b5157a9),
	.w7(32'h3a2e1485),
	.w8(32'h3ab890f1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eefe1),
	.w1(32'h3b35f106),
	.w2(32'hbacffba8),
	.w3(32'h3a8ed0b9),
	.w4(32'hbac41910),
	.w5(32'hbad69001),
	.w6(32'h3b03e3f8),
	.w7(32'hbb10f344),
	.w8(32'hbac534ac),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0002),
	.w1(32'hbb6f9598),
	.w2(32'hbb629d5a),
	.w3(32'hbc0c1485),
	.w4(32'hbb71c6a5),
	.w5(32'h3a2a5bb4),
	.w6(32'hbbafce09),
	.w7(32'hbbaea899),
	.w8(32'hbafda5ea),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93a03d),
	.w1(32'hbb89ada1),
	.w2(32'hba986bc6),
	.w3(32'h3b5b98a4),
	.w4(32'h399ada47),
	.w5(32'hba5b95ee),
	.w6(32'h3bbe331d),
	.w7(32'h3ba31b5a),
	.w8(32'h38fb7c1d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88444f5),
	.w1(32'h3b329ab8),
	.w2(32'h3b9a2b28),
	.w3(32'hbb478c65),
	.w4(32'hbad36437),
	.w5(32'h3ba67420),
	.w6(32'hbb8c45bb),
	.w7(32'hb9b42027),
	.w8(32'hbc2c6107),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacaeb),
	.w1(32'h3c58f0b7),
	.w2(32'hbb2b6262),
	.w3(32'hbc18d16c),
	.w4(32'hbca5bd5c),
	.w5(32'h3aa9e570),
	.w6(32'h3b6a08cc),
	.w7(32'h3bc3842c),
	.w8(32'h3c1d9677),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6586),
	.w1(32'hba202cea),
	.w2(32'hbba38227),
	.w3(32'hbc3312dd),
	.w4(32'hbbdf3f24),
	.w5(32'hbc028007),
	.w6(32'h3cb8c966),
	.w7(32'h3c9c4c48),
	.w8(32'h3c13bc9f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8c75),
	.w1(32'h3b48bf28),
	.w2(32'h3b9076a9),
	.w3(32'hbc2733a0),
	.w4(32'hbc065b21),
	.w5(32'hbcddf74d),
	.w6(32'h3cbdb03c),
	.w7(32'h3c516bf4),
	.w8(32'hbb189baf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63633),
	.w1(32'h3bb6977c),
	.w2(32'h3c0a973c),
	.w3(32'hbcc6bc24),
	.w4(32'hbc68a60a),
	.w5(32'hbc40b01a),
	.w6(32'h3c1cb494),
	.w7(32'hbb497cfe),
	.w8(32'h3b1419cf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc270da),
	.w1(32'h3b6fc17c),
	.w2(32'hbc446146),
	.w3(32'hbcb6b804),
	.w4(32'hbbb38599),
	.w5(32'h3b703aa9),
	.w6(32'h3b459f4b),
	.w7(32'hbc9d3dcc),
	.w8(32'hbab72ea4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c7458),
	.w1(32'hbb673e56),
	.w2(32'h3a2d1362),
	.w3(32'h3cb3799c),
	.w4(32'h3c89279b),
	.w5(32'h3b26d784),
	.w6(32'hbb3c18ef),
	.w7(32'hbb39b37b),
	.w8(32'hbb95314b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb335f1),
	.w1(32'h39d28e3d),
	.w2(32'hbacfcac7),
	.w3(32'hbc114375),
	.w4(32'hbbc389d2),
	.w5(32'h3c9c3729),
	.w6(32'h3c0b8e82),
	.w7(32'hbab22dc4),
	.w8(32'hbcab8efa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39565),
	.w1(32'hbbcf2d25),
	.w2(32'h3b5c9e8c),
	.w3(32'h3ce14eb4),
	.w4(32'h3b812d02),
	.w5(32'hb999412f),
	.w6(32'hb9c54f52),
	.w7(32'h3b46b1b4),
	.w8(32'h3c9e4245),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30fb06),
	.w1(32'h3bacd137),
	.w2(32'hbab0f691),
	.w3(32'hbc5b8074),
	.w4(32'hb9970072),
	.w5(32'hbb71ec5c),
	.w6(32'h3c97fe2a),
	.w7(32'h3cb5cb55),
	.w8(32'hbaef3f66),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a511c15),
	.w1(32'h3bbadcb0),
	.w2(32'h3bc299e0),
	.w3(32'h3af2f15b),
	.w4(32'h3bdb1625),
	.w5(32'h3c633504),
	.w6(32'h3bb4f4d2),
	.w7(32'h3c12fce1),
	.w8(32'h3ba25e18),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd288),
	.w1(32'hbb9cc269),
	.w2(32'hbb0671f6),
	.w3(32'h3c33e6d4),
	.w4(32'hbb972f45),
	.w5(32'hbc80b14b),
	.w6(32'hbab4322f),
	.w7(32'hbc3c1f2c),
	.w8(32'hbabea74a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dd5ac),
	.w1(32'h3b04a449),
	.w2(32'h3b256db3),
	.w3(32'hbc8b08e2),
	.w4(32'hbbc6eeb4),
	.w5(32'h3ab33324),
	.w6(32'hbad554be),
	.w7(32'hbc15a404),
	.w8(32'hbb047b58),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0fedd),
	.w1(32'h3b9f6737),
	.w2(32'h3b8cfe7a),
	.w3(32'h3ba400cd),
	.w4(32'h3b44a382),
	.w5(32'h3bae8b8a),
	.w6(32'h3a9e1a10),
	.w7(32'hbab9b7da),
	.w8(32'h3b194796),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f62f),
	.w1(32'hbb0039fd),
	.w2(32'h3a55c1a2),
	.w3(32'h3a2b439c),
	.w4(32'h3a4b21b3),
	.w5(32'h3ba514c7),
	.w6(32'hbb4e3b8b),
	.w7(32'h38127a04),
	.w8(32'hbb612fee),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf48baf),
	.w1(32'hbaaf2ce2),
	.w2(32'hbace4fe4),
	.w3(32'h3bcacc0d),
	.w4(32'hbba581f3),
	.w5(32'h3947a352),
	.w6(32'h3bca45a6),
	.w7(32'h3c8b0a59),
	.w8(32'hba4f6566),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba945156),
	.w1(32'hbadec5a4),
	.w2(32'h3c1bf268),
	.w3(32'hba824283),
	.w4(32'hbab8f817),
	.w5(32'h3bce01c6),
	.w6(32'h3af1a9b3),
	.w7(32'hbae51e88),
	.w8(32'hbac70b40),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5416b7),
	.w1(32'hba53e913),
	.w2(32'h3c1355bd),
	.w3(32'h3ba52987),
	.w4(32'hbb89830d),
	.w5(32'hbca4b325),
	.w6(32'h3ace3a5f),
	.w7(32'hbbfe77c7),
	.w8(32'hbc20f0bb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42d462),
	.w1(32'h3ac87201),
	.w2(32'h3ba291ed),
	.w3(32'hbc76fae4),
	.w4(32'hbca094a2),
	.w5(32'h3b5d6911),
	.w6(32'h3b282232),
	.w7(32'h3b9457f6),
	.w8(32'h3b3980ca),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5246f),
	.w1(32'hba9b14ff),
	.w2(32'hba7b0821),
	.w3(32'hba39c40a),
	.w4(32'hb75943ed),
	.w5(32'h3ae27240),
	.w6(32'h3baae3fc),
	.w7(32'h3acadda9),
	.w8(32'h3a91770f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00f75a),
	.w1(32'h3ae3c713),
	.w2(32'h3bb81805),
	.w3(32'h3b504754),
	.w4(32'h3b9c3336),
	.w5(32'hbb58e5cd),
	.w6(32'h3ace50d1),
	.w7(32'h3b5bf0e4),
	.w8(32'hbb60e74d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30c0cb),
	.w1(32'hba9662b3),
	.w2(32'h3b455f8d),
	.w3(32'hbc628a1d),
	.w4(32'hbbd06593),
	.w5(32'h3b35a59b),
	.w6(32'hbc3f8a30),
	.w7(32'hbb65ddf8),
	.w8(32'h3b0ea62c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e375),
	.w1(32'hb9a8b513),
	.w2(32'hbc05fc1e),
	.w3(32'h3bb9fa36),
	.w4(32'h3b9b9621),
	.w5(32'hbcc8e745),
	.w6(32'h3bf4efcb),
	.w7(32'hbae45a64),
	.w8(32'hbc6d2683),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c7bb2),
	.w1(32'hbbe8e2cd),
	.w2(32'h3bd9ab5f),
	.w3(32'hbc477280),
	.w4(32'hbc2aabf0),
	.w5(32'h3bf9b645),
	.w6(32'h3bc31a81),
	.w7(32'h39b06a6c),
	.w8(32'hbbbc4c89),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1e85),
	.w1(32'hbb09f03d),
	.w2(32'h3ac828c5),
	.w3(32'hbb6c773c),
	.w4(32'hbbf824c9),
	.w5(32'hbc144b9c),
	.w6(32'hbbcdc28f),
	.w7(32'h3a623f5c),
	.w8(32'hbad37658),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836a41),
	.w1(32'hbb82d2bf),
	.w2(32'h3a33b710),
	.w3(32'hbcadc9a2),
	.w4(32'hbb283c7c),
	.w5(32'hbb20731d),
	.w6(32'h3a749787),
	.w7(32'hbbb31086),
	.w8(32'h3b31cffc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae383),
	.w1(32'hbbf2276e),
	.w2(32'hbb515adb),
	.w3(32'hbb1748ee),
	.w4(32'hbafcb6de),
	.w5(32'hbb836a8b),
	.w6(32'h3c2b58c6),
	.w7(32'h3c6db141),
	.w8(32'hbb3f62fc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0874ad),
	.w1(32'h39c6ffa1),
	.w2(32'h3b95b6ee),
	.w3(32'h3adf0f76),
	.w4(32'h3b780286),
	.w5(32'h3b86280c),
	.w6(32'h3b5ebe73),
	.w7(32'h38244313),
	.w8(32'h3bbb0525),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24c2c),
	.w1(32'hba6bf78f),
	.w2(32'h3c0510a7),
	.w3(32'h3bb7c018),
	.w4(32'h3af12a5c),
	.w5(32'hbc1193c2),
	.w6(32'h3aabe788),
	.w7(32'hbac807f2),
	.w8(32'h3cedf442),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd8138),
	.w1(32'h3b98cd88),
	.w2(32'hbc09c0b1),
	.w3(32'h3cc2c6f8),
	.w4(32'h3cbaacc6),
	.w5(32'hb9b7dc77),
	.w6(32'h3d4ac408),
	.w7(32'h3cfdfd2e),
	.w8(32'hbbfb3c13),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb416674),
	.w1(32'h3b7b56be),
	.w2(32'hba78d8df),
	.w3(32'hbbb61263),
	.w4(32'hbcb669f5),
	.w5(32'hbb2380ae),
	.w6(32'h3b2ace12),
	.w7(32'h3b3e0d55),
	.w8(32'hba420fac),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9272d4),
	.w1(32'h3a26f708),
	.w2(32'h3c24a53a),
	.w3(32'hbb068649),
	.w4(32'hbae79538),
	.w5(32'h3ae0016f),
	.w6(32'h388c2f62),
	.w7(32'h39617484),
	.w8(32'hb94bae70),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaca9c),
	.w1(32'h3b0bb570),
	.w2(32'hbb357412),
	.w3(32'h39f75c79),
	.w4(32'hb9962f9f),
	.w5(32'h3abf49a9),
	.w6(32'hbaa52b71),
	.w7(32'hbb5ff252),
	.w8(32'hbbbe1c0d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa58d1),
	.w1(32'h3b1583f7),
	.w2(32'hbaf7ab8c),
	.w3(32'h3bd5d2c1),
	.w4(32'h3b2c5682),
	.w5(32'hbba502e8),
	.w6(32'hbb36be3a),
	.w7(32'hba0bbfd7),
	.w8(32'hbb4c6578),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608756),
	.w1(32'hb9ae245a),
	.w2(32'h3b9feb7e),
	.w3(32'hbbb57f8d),
	.w4(32'hbaef69fd),
	.w5(32'h3ccb2172),
	.w6(32'hbab84bde),
	.w7(32'h3b3a54c3),
	.w8(32'h3bd2123e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b1274),
	.w1(32'h3b7d4757),
	.w2(32'h3c5a56eb),
	.w3(32'h3cb5a727),
	.w4(32'h3ca594dc),
	.w5(32'h3c426fe6),
	.w6(32'h3c52f1a0),
	.w7(32'h3c095b4f),
	.w8(32'hbb941984),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0b24c),
	.w1(32'h3bdde16d),
	.w2(32'h3af51b6b),
	.w3(32'h3c9c58cb),
	.w4(32'h3c9bf1b6),
	.w5(32'hbb0052f4),
	.w6(32'h3b78e2fa),
	.w7(32'h39d99694),
	.w8(32'hbb0f36ec),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b20a3),
	.w1(32'h3a2ee20e),
	.w2(32'hbb04955e),
	.w3(32'hbb63b110),
	.w4(32'h3b5c95e6),
	.w5(32'hbaa99fda),
	.w6(32'hbb9788d0),
	.w7(32'h3b353ad3),
	.w8(32'hba27a890),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc9c4c),
	.w1(32'hbb44b0cb),
	.w2(32'hbb8be15c),
	.w3(32'hbc5043f4),
	.w4(32'hbb37b673),
	.w5(32'hbbc57579),
	.w6(32'hbaec25e7),
	.w7(32'hb9fc444d),
	.w8(32'hbb9aa17c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354e9e),
	.w1(32'hbbaf8460),
	.w2(32'h3bed3948),
	.w3(32'hbbbcd4da),
	.w4(32'hbba18e65),
	.w5(32'h3c1ee422),
	.w6(32'hbbc3c3ea),
	.w7(32'hbbd77476),
	.w8(32'hbb14657b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842383),
	.w1(32'hbb15a032),
	.w2(32'h3b1e5bf9),
	.w3(32'h3c077c28),
	.w4(32'h3bcf16f0),
	.w5(32'hbba5cd07),
	.w6(32'hbaca828d),
	.w7(32'h3b998b07),
	.w8(32'hbbe5a357),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2f2da),
	.w1(32'hba83ef60),
	.w2(32'h3c6c0b02),
	.w3(32'hbbbafcc6),
	.w4(32'hba8fb132),
	.w5(32'hbc18a8dd),
	.w6(32'hbc20cf4a),
	.w7(32'hbb63e770),
	.w8(32'hbc8efa82),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccceea4),
	.w1(32'h3caf20b8),
	.w2(32'hbb615b4b),
	.w3(32'hbbc64936),
	.w4(32'hb8c13e19),
	.w5(32'h3afb1148),
	.w6(32'hbcccd073),
	.w7(32'hbc8702ab),
	.w8(32'h3c080f32),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067e0a),
	.w1(32'hbc0e0eb2),
	.w2(32'h3ab808fa),
	.w3(32'hbbce0b66),
	.w4(32'hbc58a904),
	.w5(32'hbb877fd7),
	.w6(32'h3b78f66b),
	.w7(32'h384467a7),
	.w8(32'hbbbdf4a3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01180d),
	.w1(32'hb9799ffc),
	.w2(32'h3c98b6d3),
	.w3(32'hbb6a5962),
	.w4(32'hbad22ab7),
	.w5(32'h3cb65188),
	.w6(32'h3bedcecf),
	.w7(32'h3bc954b9),
	.w8(32'h3c003616),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3923e9),
	.w1(32'hbb2a066a),
	.w2(32'h3bffff24),
	.w3(32'h3cc41976),
	.w4(32'h3c354d04),
	.w5(32'h3c160491),
	.w6(32'hba74e477),
	.w7(32'hba0b98f2),
	.w8(32'hbba7c974),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0a8b),
	.w1(32'h3b9f897a),
	.w2(32'h3b94cc31),
	.w3(32'h3c053e2b),
	.w4(32'h3bc3a7b6),
	.w5(32'h3ae9b7e8),
	.w6(32'hbafb46af),
	.w7(32'h3a3b9be9),
	.w8(32'h3aa58e79),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3fe0),
	.w1(32'h38d80d13),
	.w2(32'hbba8d1cd),
	.w3(32'hba2b3c65),
	.w4(32'h3a164464),
	.w5(32'h3aeb0ed8),
	.w6(32'hbb0fb6a3),
	.w7(32'hbb6b7b22),
	.w8(32'hba31eab8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d56a6),
	.w1(32'h387f15f4),
	.w2(32'h3b793184),
	.w3(32'h3b8f9f43),
	.w4(32'h3a190133),
	.w5(32'h3b84a12b),
	.w6(32'h3bc89d75),
	.w7(32'h3b811bcd),
	.w8(32'h3b6ca99d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4104e),
	.w1(32'hbbda0ba9),
	.w2(32'hbb94ec76),
	.w3(32'h3aa303db),
	.w4(32'hbbdd5fdf),
	.w5(32'hbb913eec),
	.w6(32'hbb8d4df4),
	.w7(32'hbaa51674),
	.w8(32'hbbb472ac),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9c4b),
	.w1(32'h3b38590b),
	.w2(32'h3c0654cf),
	.w3(32'hbb2bb24a),
	.w4(32'hb9947a99),
	.w5(32'h3c2433f4),
	.w6(32'h3bf22531),
	.w7(32'h3975b509),
	.w8(32'h3c0fe0de),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd486f4),
	.w1(32'hbb8e100d),
	.w2(32'hba26d405),
	.w3(32'h3b869a2c),
	.w4(32'h3b40edd8),
	.w5(32'h3a0d2f21),
	.w6(32'hbbac16bf),
	.w7(32'h3b2c8406),
	.w8(32'hba3f1638),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c1a4f),
	.w1(32'hbaf6e1f7),
	.w2(32'hbb678fd4),
	.w3(32'h3910937c),
	.w4(32'hbad614bf),
	.w5(32'hbbb86bff),
	.w6(32'hb9354c16),
	.w7(32'hbb869b55),
	.w8(32'h3b6c97b7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee5197),
	.w1(32'hbb276f22),
	.w2(32'h3b40942d),
	.w3(32'hbbe92d80),
	.w4(32'hbb528ca5),
	.w5(32'hba7d441b),
	.w6(32'h3a83684c),
	.w7(32'hb998ac8f),
	.w8(32'hbbeb7a90),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09ab49),
	.w1(32'h3a884c7d),
	.w2(32'h3b05690b),
	.w3(32'hbb982b3d),
	.w4(32'h3b0da074),
	.w5(32'hbbea3985),
	.w6(32'hbad7cb23),
	.w7(32'h3bb21642),
	.w8(32'hbbfec36f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beacd2c),
	.w1(32'h3c0185e3),
	.w2(32'h3baff17c),
	.w3(32'hbb0e6730),
	.w4(32'h39d93b88),
	.w5(32'h3be743ef),
	.w6(32'hbb7d7a89),
	.w7(32'hbaaab9f1),
	.w8(32'h3b10e331),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3dec3f),
	.w1(32'h3b9bb089),
	.w2(32'hbab8c810),
	.w3(32'h3904f439),
	.w4(32'h3b5df03b),
	.w5(32'h3a9771aa),
	.w6(32'h3b6a4eb5),
	.w7(32'h3a9f2ed4),
	.w8(32'h3b5fbdd0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80105b),
	.w1(32'hbb73b3e5),
	.w2(32'h3b3dd003),
	.w3(32'h3b919ac6),
	.w4(32'hbb263279),
	.w5(32'h3c308133),
	.w6(32'h3b83c3c2),
	.w7(32'h3bded616),
	.w8(32'h383808c8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b655606),
	.w1(32'hbb0e7a2a),
	.w2(32'hbc0c4589),
	.w3(32'h3c12ab2d),
	.w4(32'h3bb086a2),
	.w5(32'hbc82cffc),
	.w6(32'h3b6fd90e),
	.w7(32'h3c41810d),
	.w8(32'hbc6413e0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1a5f),
	.w1(32'h3b2edd00),
	.w2(32'h3b622979),
	.w3(32'hbca251c8),
	.w4(32'hbc50a2f8),
	.w5(32'hbba0071d),
	.w6(32'hbca05e6d),
	.w7(32'hbca6c238),
	.w8(32'hbacd4a15),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c222005),
	.w1(32'h3b61c081),
	.w2(32'h3b3a1dc9),
	.w3(32'h3af69716),
	.w4(32'h3b5f962e),
	.w5(32'hba82df8e),
	.w6(32'hbc265e61),
	.w7(32'hbc00761f),
	.w8(32'hbaad1195),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87fc95),
	.w1(32'hba9a3059),
	.w2(32'hb9a1c201),
	.w3(32'h3a7e4da5),
	.w4(32'hbb3f0afc),
	.w5(32'hba27fc0a),
	.w6(32'h3b9705fb),
	.w7(32'hb9bed805),
	.w8(32'hbb373890),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c6b3),
	.w1(32'h3bee2898),
	.w2(32'h3c35cc56),
	.w3(32'hbaf14ce4),
	.w4(32'h3b95772b),
	.w5(32'h3c0382c0),
	.w6(32'hbc01109d),
	.w7(32'h3add8966),
	.w8(32'hbb40ca97),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c289a47),
	.w1(32'h3c23f9bc),
	.w2(32'h3be19598),
	.w3(32'h3caa5523),
	.w4(32'h3c94a875),
	.w5(32'h3d01bd61),
	.w6(32'h3be9fa20),
	.w7(32'h3c7631ca),
	.w8(32'h3d0354a9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928868),
	.w1(32'hbcac2ab6),
	.w2(32'hbc087ab7),
	.w3(32'h3c2253c1),
	.w4(32'h380fabac),
	.w5(32'hbca1cb71),
	.w6(32'h3c98e18e),
	.w7(32'h3c876f76),
	.w8(32'hbc45bd3a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c3cb),
	.w1(32'h3b6e4915),
	.w2(32'h3bf4f595),
	.w3(32'hbca55390),
	.w4(32'hbbac2c39),
	.w5(32'h3b91f10c),
	.w6(32'hbc642bb3),
	.w7(32'hbc8f349b),
	.w8(32'h3b62db4a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b847066),
	.w1(32'hba2c1817),
	.w2(32'h3bcb89d4),
	.w3(32'h3a30d4f0),
	.w4(32'h3974ca3b),
	.w5(32'h3a3f8f66),
	.w6(32'h3b8f5156),
	.w7(32'h3b4231de),
	.w8(32'hbbe090e3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babca12),
	.w1(32'h3a990a35),
	.w2(32'hbbfa0678),
	.w3(32'h3c41a79d),
	.w4(32'h3c0b947e),
	.w5(32'h3b2cf704),
	.w6(32'hbb504cae),
	.w7(32'hbb3e483d),
	.w8(32'hbb34d0f1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01455c),
	.w1(32'hbb967ba3),
	.w2(32'hbbe64f90),
	.w3(32'hbc03ae1f),
	.w4(32'hbbd6b9d5),
	.w5(32'hbbbb4e07),
	.w6(32'hbaa4985d),
	.w7(32'hb9e3f244),
	.w8(32'hb945d413),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1924ed),
	.w1(32'hbbe70069),
	.w2(32'h3b14027c),
	.w3(32'hbc231619),
	.w4(32'hbc13b22f),
	.w5(32'hbb1bc2e2),
	.w6(32'hbb4fd62a),
	.w7(32'hbba6a55b),
	.w8(32'hbb7c18cf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf27d8d),
	.w1(32'h3ba8de48),
	.w2(32'h3b03c5ff),
	.w3(32'hb885b05c),
	.w4(32'h3b354852),
	.w5(32'h3bcd1a42),
	.w6(32'hba9c6a3d),
	.w7(32'hbad3c99f),
	.w8(32'h3b478aa7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c85529),
	.w1(32'hbb34b1b0),
	.w2(32'h3b9b7550),
	.w3(32'h39a57fa0),
	.w4(32'hbb877dd7),
	.w5(32'hb9489ef3),
	.w6(32'h38d8d48e),
	.w7(32'h3b192490),
	.w8(32'h3b388b3b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56ed35),
	.w1(32'h3b6ac535),
	.w2(32'hb9c23de4),
	.w3(32'hba286856),
	.w4(32'h3b60f56c),
	.w5(32'h392522c9),
	.w6(32'h3bb82ce2),
	.w7(32'h3ad8507e),
	.w8(32'hb9f2e203),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d43de),
	.w1(32'hba456c4d),
	.w2(32'h3c26b98a),
	.w3(32'h3b6c21f8),
	.w4(32'h3b1016b8),
	.w5(32'h3c0d1110),
	.w6(32'h3be0a884),
	.w7(32'h3b758754),
	.w8(32'h3b477cd4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a81b),
	.w1(32'h3b1bf044),
	.w2(32'hbb41638b),
	.w3(32'h3bc9bcf8),
	.w4(32'hb814f7c7),
	.w5(32'hbc15376e),
	.w6(32'h396b8f93),
	.w7(32'hbb28a61e),
	.w8(32'hbbba9acc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7cf58),
	.w1(32'h3a90de81),
	.w2(32'h3b672e2b),
	.w3(32'hbc1dd0c1),
	.w4(32'hbbb90450),
	.w5(32'h3b9187b4),
	.w6(32'hbbaf8c76),
	.w7(32'hb874ad0f),
	.w8(32'h3be0078e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba33497),
	.w1(32'h3c066534),
	.w2(32'h3b4bbf83),
	.w3(32'h3b9b3b48),
	.w4(32'h3c195380),
	.w5(32'hba55a9e6),
	.w6(32'h3c092e56),
	.w7(32'h3c2f57d7),
	.w8(32'hba14b289),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc332c),
	.w1(32'h3a32a558),
	.w2(32'hb965f063),
	.w3(32'hbab8759a),
	.w4(32'hbb8aa8c9),
	.w5(32'hbaac6433),
	.w6(32'hbbc0cd9d),
	.w7(32'hbb323c7c),
	.w8(32'h3985af14),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4630b2),
	.w1(32'hbb5d4c7f),
	.w2(32'hbb99dcb1),
	.w3(32'hbb4ede75),
	.w4(32'hbae28ab0),
	.w5(32'h3be83819),
	.w6(32'hbab9cbc6),
	.w7(32'hbb184ce8),
	.w8(32'h3c87d73b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670a03),
	.w1(32'hbc7b7a8c),
	.w2(32'hbb99a2d5),
	.w3(32'hbbb28012),
	.w4(32'hbbb823d0),
	.w5(32'hbc0e413a),
	.w6(32'h3badb1a7),
	.w7(32'h3b9503fd),
	.w8(32'hbba06c5f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd691a),
	.w1(32'hbaf241e1),
	.w2(32'hbb8fb187),
	.w3(32'hbbe8cd74),
	.w4(32'hbbdec54b),
	.w5(32'hbc27fd50),
	.w6(32'hba693f35),
	.w7(32'hbaaa980d),
	.w8(32'hbc28d65e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc416445),
	.w1(32'hbc0d436e),
	.w2(32'h3bdf8516),
	.w3(32'hbc8b76e5),
	.w4(32'hbc1115cb),
	.w5(32'h3c440e5a),
	.w6(32'hbc351f32),
	.w7(32'hbb4d873d),
	.w8(32'h398afb0b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91f025),
	.w1(32'hbb82a79a),
	.w2(32'hbae0f509),
	.w3(32'h3c2934fd),
	.w4(32'h3b077714),
	.w5(32'hbc2be686),
	.w6(32'hbb6bf915),
	.w7(32'hbadf1a55),
	.w8(32'hbbc4feed),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb55e8),
	.w1(32'h3a535cd0),
	.w2(32'h3c056fce),
	.w3(32'hbb397e61),
	.w4(32'hbb9331cc),
	.w5(32'h3bfe9fee),
	.w6(32'h3bbee8b4),
	.w7(32'h3ae701e7),
	.w8(32'h3af21fe5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee47e),
	.w1(32'h3b0302b6),
	.w2(32'h3b2170ea),
	.w3(32'h3bad2ff0),
	.w4(32'h3bf9c61d),
	.w5(32'hbb52b10c),
	.w6(32'hbb0f5b76),
	.w7(32'h3a2e1c10),
	.w8(32'hba17a6f8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa0207),
	.w1(32'h3a93d6c0),
	.w2(32'hb9cd6fc0),
	.w3(32'hbbee6764),
	.w4(32'hbb31bd63),
	.w5(32'hba1ecb8d),
	.w6(32'hbb3c47a8),
	.w7(32'h3a7acf49),
	.w8(32'hb8aedfdb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90cba),
	.w1(32'hbaef7a3a),
	.w2(32'hbb0b4186),
	.w3(32'h3b1686da),
	.w4(32'h3b435d09),
	.w5(32'hbc67e8fd),
	.w6(32'h3bbec74c),
	.w7(32'h3aec93fa),
	.w8(32'hbbba52d7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016522),
	.w1(32'h3adf6566),
	.w2(32'hbbd0c965),
	.w3(32'hbcbcb075),
	.w4(32'hbc3a2e47),
	.w5(32'hbb962cb5),
	.w6(32'hbc9b5c1e),
	.w7(32'hbc4178d2),
	.w8(32'h3bd7d667),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c6eff),
	.w1(32'h3c4662ef),
	.w2(32'h3b212f47),
	.w3(32'h3af12a82),
	.w4(32'hbacde104),
	.w5(32'h3b11e99b),
	.w6(32'h3c2a0aa1),
	.w7(32'h3bc8dd82),
	.w8(32'h3c1a0dc3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07bdbb),
	.w1(32'hba3e503c),
	.w2(32'hbb49538e),
	.w3(32'hbbe44003),
	.w4(32'hbabba725),
	.w5(32'hbb840f2a),
	.w6(32'hb91a93e9),
	.w7(32'h3b0f0a54),
	.w8(32'hbb10a085),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ee63),
	.w1(32'hbb885dcf),
	.w2(32'hb829467a),
	.w3(32'hbc14beab),
	.w4(32'hbb0658fb),
	.w5(32'h394ad01a),
	.w6(32'hbbaadcc1),
	.w7(32'h3aded433),
	.w8(32'h3910528c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4417a7),
	.w1(32'hb9eedc8f),
	.w2(32'h3bdf2195),
	.w3(32'hba942610),
	.w4(32'hbaa7edd3),
	.w5(32'hbafbcf9b),
	.w6(32'hba838908),
	.w7(32'hba3ffac8),
	.w8(32'hb9fd810b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7b55),
	.w1(32'h3bc878a3),
	.w2(32'hbbffd016),
	.w3(32'hbb0f43e5),
	.w4(32'h3b328dac),
	.w5(32'hbcba33e3),
	.w6(32'h3bd75c24),
	.w7(32'h39f20b46),
	.w8(32'hbb35ff26),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0555),
	.w1(32'hbb3dcfa5),
	.w2(32'hbc4b6500),
	.w3(32'hbcb93910),
	.w4(32'hbc9c6d57),
	.w5(32'hbc1a5936),
	.w6(32'hbbc82c5e),
	.w7(32'hbc1d0f99),
	.w8(32'h3bfc8318),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39545e),
	.w1(32'hbc037fcb),
	.w2(32'h3c67582f),
	.w3(32'hbc35695f),
	.w4(32'hbc067399),
	.w5(32'h3c136676),
	.w6(32'h3c547751),
	.w7(32'h3bef5e4d),
	.w8(32'h3a248c71),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2adc66),
	.w1(32'h3c228cfa),
	.w2(32'h3bf6cbe4),
	.w3(32'h3c1cefb2),
	.w4(32'h3b921e38),
	.w5(32'h3b2fdda7),
	.w6(32'h3a4a6792),
	.w7(32'hbb61fd3b),
	.w8(32'hba52734f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf1236),
	.w1(32'h3af79c5f),
	.w2(32'hbb3740a5),
	.w3(32'hbb3b1d54),
	.w4(32'hbac5f18c),
	.w5(32'hbb0dae49),
	.w6(32'hbb7d5afb),
	.w7(32'hb9dec03f),
	.w8(32'hba978cc7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009b74),
	.w1(32'hbb04c142),
	.w2(32'h3b86e863),
	.w3(32'h3ab68736),
	.w4(32'hbae73005),
	.w5(32'hbb31b1d0),
	.w6(32'h3b622c99),
	.w7(32'h3ae41c2e),
	.w8(32'h3ac9003d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfacd3e),
	.w1(32'h3b97d507),
	.w2(32'h38b611d4),
	.w3(32'hbb369ccd),
	.w4(32'h3b95e4bc),
	.w5(32'hbc1d6cb2),
	.w6(32'h3ac21805),
	.w7(32'h3befcfd5),
	.w8(32'hbc2b0661),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54ee97),
	.w1(32'hba341d97),
	.w2(32'h3ac4f272),
	.w3(32'hbc311e4d),
	.w4(32'hbc0bb284),
	.w5(32'h3b034302),
	.w6(32'hbc4b4f3c),
	.w7(32'hbc58f467),
	.w8(32'h3bdb0008),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24f925),
	.w1(32'hbc322250),
	.w2(32'hbb09a4b3),
	.w3(32'hbacbf3b3),
	.w4(32'hbb4c75d3),
	.w5(32'hbbe936e8),
	.w6(32'h3bf61da4),
	.w7(32'h3bd5b62f),
	.w8(32'h3af50e78),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0efba),
	.w1(32'h3b84aff2),
	.w2(32'hbbf5ca21),
	.w3(32'hbbcbe2fa),
	.w4(32'hbba75df4),
	.w5(32'hbbc5a1f9),
	.w6(32'h39b811aa),
	.w7(32'hbb762957),
	.w8(32'hbc121d2d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb6d8),
	.w1(32'hbc1f9e99),
	.w2(32'h3beebcde),
	.w3(32'hbbb05000),
	.w4(32'hbbfd224f),
	.w5(32'h3b9bfcb9),
	.w6(32'hbb92a124),
	.w7(32'hbb5d6e26),
	.w8(32'h3b9387c3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be062),
	.w1(32'h3c6bde73),
	.w2(32'h3abae135),
	.w3(32'h3bbc746b),
	.w4(32'h3c54b1c7),
	.w5(32'h3c2a67b5),
	.w6(32'h3b33a6c8),
	.w7(32'h3c1f6b2a),
	.w8(32'h3b83c1b8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a356c57),
	.w1(32'hba26ad18),
	.w2(32'hbbc8f89c),
	.w3(32'h3b09c135),
	.w4(32'h3c0fae7e),
	.w5(32'hbb0affe1),
	.w6(32'h3a3b8a6a),
	.w7(32'h3ad6d32c),
	.w8(32'hbbe55759),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66d21),
	.w1(32'hb8cdc4ab),
	.w2(32'h3b6beaf7),
	.w3(32'hbc28ac1f),
	.w4(32'h39c30582),
	.w5(32'h3b090872),
	.w6(32'hbb9330c0),
	.w7(32'hbb9aebf7),
	.w8(32'h39825fe2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0db987),
	.w1(32'h3c33b544),
	.w2(32'hbbd4cb24),
	.w3(32'h3bc29663),
	.w4(32'h3c1c6327),
	.w5(32'hbb5093e4),
	.w6(32'h3a24e33e),
	.w7(32'h3b2daea4),
	.w8(32'h3bbacf11),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5273da),
	.w1(32'hbab7fb36),
	.w2(32'hbba6a835),
	.w3(32'hbc5e2d1d),
	.w4(32'hbc08367f),
	.w5(32'hbc1adcad),
	.w6(32'hbb02a4e8),
	.w7(32'h3a954599),
	.w8(32'hbc512edb),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2415ea),
	.w1(32'h3b96520d),
	.w2(32'hbb86b642),
	.w3(32'hbbf0b811),
	.w4(32'hbbcaaaf8),
	.w5(32'hbbdf2d79),
	.w6(32'hbc56a67b),
	.w7(32'hbb8fee82),
	.w8(32'hbb1b22ca),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa4e6),
	.w1(32'hb840437a),
	.w2(32'hbb7ccd06),
	.w3(32'hbbd1b517),
	.w4(32'h3a250568),
	.w5(32'hbb5555c1),
	.w6(32'hbaf54367),
	.w7(32'h3a8aee14),
	.w8(32'h39865bcc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc422cf2),
	.w1(32'hbbb81e13),
	.w2(32'h3c230271),
	.w3(32'hbc350796),
	.w4(32'hbb375fb5),
	.w5(32'h3add4a54),
	.w6(32'hbbca7992),
	.w7(32'hbb6c03af),
	.w8(32'h3b809335),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd496d0),
	.w1(32'h3b34cc40),
	.w2(32'h3b63a871),
	.w3(32'h3c0e1ab8),
	.w4(32'h3c2c8e25),
	.w5(32'hbc009926),
	.w6(32'hba0fc642),
	.w7(32'h3b98dd77),
	.w8(32'hbbe15546),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf49f42),
	.w1(32'h3b87c14a),
	.w2(32'h3bf3c4b9),
	.w3(32'hbb4cde4e),
	.w4(32'hbb4e4837),
	.w5(32'h3bd4bbd9),
	.w6(32'hbb3d17a3),
	.w7(32'hba0ad14d),
	.w8(32'h3bac6261),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c022f42),
	.w1(32'hbab79a95),
	.w2(32'h3b0d6703),
	.w3(32'h3bc01426),
	.w4(32'h3c21e7ad),
	.w5(32'h3aa2ecbc),
	.w6(32'h3c0c8990),
	.w7(32'h3b85c569),
	.w8(32'hba8057a5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912bfd5),
	.w1(32'h3b763b2b),
	.w2(32'hb9f94bac),
	.w3(32'hbbceccbc),
	.w4(32'hbb943d16),
	.w5(32'hbc384fc8),
	.w6(32'hbbd5522d),
	.w7(32'hbc2ae2f9),
	.w8(32'hbc3fa00a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba146116),
	.w1(32'hbaac44b4),
	.w2(32'h3b94e63a),
	.w3(32'hbb8be209),
	.w4(32'hb9edf922),
	.w5(32'h3bf61e42),
	.w6(32'hbc2a7861),
	.w7(32'h3b09e003),
	.w8(32'h3b2e2bd1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac69d1),
	.w1(32'h39c427f9),
	.w2(32'h3c28b7a9),
	.w3(32'h3bfc98bb),
	.w4(32'h3bbf546b),
	.w5(32'h3c37a6e8),
	.w6(32'h3b965627),
	.w7(32'h3c37e932),
	.w8(32'h3aa13704),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1863e8),
	.w1(32'hbac9876b),
	.w2(32'h3bc1403a),
	.w3(32'h3c8341a7),
	.w4(32'h3c5d2740),
	.w5(32'h3bcc9e7c),
	.w6(32'h3bb6b633),
	.w7(32'h3bb09a80),
	.w8(32'h3b07e93e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba320503),
	.w1(32'h3a0a81ea),
	.w2(32'h3c033cc4),
	.w3(32'h3bbc27d6),
	.w4(32'h3b969436),
	.w5(32'h3bcd655e),
	.w6(32'h3b79b9a4),
	.w7(32'h3b0b1b45),
	.w8(32'hbb936f46),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ada0e),
	.w1(32'h3c0fc24b),
	.w2(32'hbc18d7ef),
	.w3(32'h3c4e0406),
	.w4(32'h3c2d8cdd),
	.w5(32'hbb10fe37),
	.w6(32'hb8ae155e),
	.w7(32'h3b20ebd2),
	.w8(32'h3c62f420),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaf311),
	.w1(32'hbae60eb3),
	.w2(32'h3c3789ea),
	.w3(32'hbbdfdd2b),
	.w4(32'hbbb899f0),
	.w5(32'h3c3abe19),
	.w6(32'h3c17339f),
	.w7(32'h3b7834e4),
	.w8(32'h3b05a905),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46944c),
	.w1(32'h3c1bdf51),
	.w2(32'h3bf43ea5),
	.w3(32'h3ca01053),
	.w4(32'h3c9bf04e),
	.w5(32'hbba32922),
	.w6(32'h3b621771),
	.w7(32'h3bd24c70),
	.w8(32'hbc2a4c24),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6d163),
	.w1(32'h3bcdc19b),
	.w2(32'h3b477c65),
	.w3(32'h3bd6f096),
	.w4(32'h3ba9a3ae),
	.w5(32'h3b6c55a3),
	.w6(32'hbaaaea40),
	.w7(32'hbbfc8d75),
	.w8(32'h39612fda),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb47ee5),
	.w1(32'hbb33ef3f),
	.w2(32'h3b0948ae),
	.w3(32'h3ad16984),
	.w4(32'hbba9888d),
	.w5(32'h3b2186e9),
	.w6(32'hbafb2320),
	.w7(32'h3b40b0bf),
	.w8(32'h3bbb8e36),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac18b2b),
	.w1(32'h3a64e5b5),
	.w2(32'hbadd83a4),
	.w3(32'hbb940ef0),
	.w4(32'hbb9c9bbc),
	.w5(32'hba3f0989),
	.w6(32'h3b5ffa44),
	.w7(32'h3aba80fa),
	.w8(32'h390b57ff),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf6dfd),
	.w1(32'hbb0eadac),
	.w2(32'hbb97df64),
	.w3(32'hbb1933d7),
	.w4(32'hba8a5ec2),
	.w5(32'hbb1a2561),
	.w6(32'hba323675),
	.w7(32'h3aa57fa3),
	.w8(32'h3ac9c95a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09b265),
	.w1(32'hbbee2c79),
	.w2(32'h3ab0a001),
	.w3(32'hbbb417eb),
	.w4(32'hbb9e110a),
	.w5(32'hbb79301e),
	.w6(32'hba441f22),
	.w7(32'h3989bddf),
	.w8(32'hbb8f8848),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee0e3),
	.w1(32'h3b24f80e),
	.w2(32'h3be090da),
	.w3(32'hbc4882ff),
	.w4(32'hbb9fb4b5),
	.w5(32'h3bcfe0df),
	.w6(32'hbb3b2f62),
	.w7(32'hba33d9d8),
	.w8(32'h3b874c0a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9631cc),
	.w1(32'h3b4a0fb8),
	.w2(32'hbb4432ba),
	.w3(32'h3beb4d6e),
	.w4(32'h3bcc8f12),
	.w5(32'hbb2808b0),
	.w6(32'h3bae870e),
	.w7(32'h3b8e94de),
	.w8(32'hbc0a05e3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285314),
	.w1(32'hbb10fa46),
	.w2(32'h3c1e620a),
	.w3(32'hbb622eb4),
	.w4(32'hbc12d8b9),
	.w5(32'h3c24a0d6),
	.w6(32'hbc184947),
	.w7(32'hbae17a6a),
	.w8(32'h3bb7334a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39be4),
	.w1(32'h3c051365),
	.w2(32'h3a672a81),
	.w3(32'h3a91a575),
	.w4(32'h3b2aa9bb),
	.w5(32'h3b96efa9),
	.w6(32'h3b11af8e),
	.w7(32'h3979fa6f),
	.w8(32'h3be42e94),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc78e37),
	.w1(32'h3bd7dffc),
	.w2(32'hbba9e21b),
	.w3(32'h3c5a614d),
	.w4(32'h3bea6353),
	.w5(32'hbc2b9358),
	.w6(32'h3c68ea08),
	.w7(32'h3bf2cc41),
	.w8(32'hbb6cb4b5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule