module layer_10_featuremap_346(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1a09a),
	.w1(32'hbbbf4de4),
	.w2(32'hbbe79a10),
	.w3(32'hbc02d682),
	.w4(32'hbc073162),
	.w5(32'hbb615a55),
	.w6(32'hbbfc0677),
	.w7(32'hbc18a396),
	.w8(32'hb9f42a06),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a0ada),
	.w1(32'h3b604c3f),
	.w2(32'h3ba5da0b),
	.w3(32'h3b032570),
	.w4(32'hbaf47170),
	.w5(32'hbb99ac5a),
	.w6(32'h39569884),
	.w7(32'hbb11c0b5),
	.w8(32'hbc3bbee5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae2d73),
	.w1(32'h3a61a4b2),
	.w2(32'hb902d329),
	.w3(32'h3a730d79),
	.w4(32'h3b92a54d),
	.w5(32'hbad62566),
	.w6(32'hbbe77b38),
	.w7(32'hb9d2cb0d),
	.w8(32'hbb849ef5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa896b6),
	.w1(32'hbb086b3d),
	.w2(32'h3a1b615c),
	.w3(32'h3aad8936),
	.w4(32'h3b6aa675),
	.w5(32'hbacacb9c),
	.w6(32'hba1bef05),
	.w7(32'h3b52d75e),
	.w8(32'h3b1e1ae1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61a52d),
	.w1(32'hb997e09f),
	.w2(32'h3b874ad7),
	.w3(32'hbb04bbe9),
	.w4(32'hbbc093c2),
	.w5(32'hb77fe463),
	.w6(32'h3bd307b5),
	.w7(32'h3b825945),
	.w8(32'h39afcc74),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b512f),
	.w1(32'h3aa285ad),
	.w2(32'h3ad156f3),
	.w3(32'h3b300d01),
	.w4(32'h3ba6ad32),
	.w5(32'hb9c94fc9),
	.w6(32'h3ab78b16),
	.w7(32'h3ba12150),
	.w8(32'h39e35779),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a8aea),
	.w1(32'h3c101dff),
	.w2(32'hbb65e4ec),
	.w3(32'h3a5eb310),
	.w4(32'h3b8c82fd),
	.w5(32'hbc1dcd5b),
	.w6(32'h3c71cd60),
	.w7(32'h3b932111),
	.w8(32'hbca097ba),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30c83),
	.w1(32'hbc404278),
	.w2(32'hbc540e21),
	.w3(32'hbc715102),
	.w4(32'h3a932060),
	.w5(32'hbb63b582),
	.w6(32'h3b7fa366),
	.w7(32'hbc09fc6b),
	.w8(32'h3b4b7d84),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e2ed6),
	.w1(32'hb9748ed6),
	.w2(32'hbaaef74a),
	.w3(32'h3aab2740),
	.w4(32'hb95ee249),
	.w5(32'h3939419d),
	.w6(32'hbafa3f8b),
	.w7(32'h3a5dcede),
	.w8(32'h3a220250),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31d4bf),
	.w1(32'h3b7533fa),
	.w2(32'hbbdcfc37),
	.w3(32'h3b90311b),
	.w4(32'h3bec705e),
	.w5(32'hbbaa2d0e),
	.w6(32'h3a16cf5a),
	.w7(32'h3b7d6657),
	.w8(32'hbbfa1e9d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f019a6),
	.w1(32'hbb157e98),
	.w2(32'h3abe3e81),
	.w3(32'h39bbc584),
	.w4(32'h3b6a452a),
	.w5(32'h3a12dff3),
	.w6(32'h3b7e07dd),
	.w7(32'h3c012498),
	.w8(32'h3b6a5cd8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4138),
	.w1(32'h3b657571),
	.w2(32'hbc09e2f2),
	.w3(32'hba88e206),
	.w4(32'h3b90f135),
	.w5(32'h3b25eb7d),
	.w6(32'h3b7635a4),
	.w7(32'h3c3a2f63),
	.w8(32'hbb76811a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f61e),
	.w1(32'hbb093920),
	.w2(32'hbc1fe16a),
	.w3(32'h3bcdbc40),
	.w4(32'h3bb41cc2),
	.w5(32'hbc8282f3),
	.w6(32'h3b9667fa),
	.w7(32'h3acfddce),
	.w8(32'hbc21e710),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0d4e),
	.w1(32'hbbb167dd),
	.w2(32'hbc62c92d),
	.w3(32'hbb1a97cc),
	.w4(32'hbc6ec2fa),
	.w5(32'hbbd18878),
	.w6(32'hbb74b3b4),
	.w7(32'hbc343d05),
	.w8(32'hba3017d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bf91),
	.w1(32'h3c0ade69),
	.w2(32'h3bf57882),
	.w3(32'h3a4808bf),
	.w4(32'h3c1663b8),
	.w5(32'h3b2b6c14),
	.w6(32'hba266389),
	.w7(32'h3ba2b8ff),
	.w8(32'h3c0f620d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183d64),
	.w1(32'hbbeffb31),
	.w2(32'hbc524a91),
	.w3(32'hba03b4e5),
	.w4(32'h3ababcc5),
	.w5(32'hbbae9b40),
	.w6(32'hbc3778cf),
	.w7(32'h3b4d6578),
	.w8(32'hbbe3c644),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7e02f),
	.w1(32'hb8c43e01),
	.w2(32'h3a692458),
	.w3(32'hb964f228),
	.w4(32'h3ac5c4b6),
	.w5(32'hbaeebcf8),
	.w6(32'h39814719),
	.w7(32'h3b0029ed),
	.w8(32'hbb0f4484),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14049d),
	.w1(32'hbc066f53),
	.w2(32'hbcefcc41),
	.w3(32'hbb33d722),
	.w4(32'hbb673062),
	.w5(32'hbc7421f4),
	.w6(32'hbb01a468),
	.w7(32'hbbbc424e),
	.w8(32'hbc75580e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99a70e),
	.w1(32'hbb8ec203),
	.w2(32'hbbf75e57),
	.w3(32'hbb33556c),
	.w4(32'hba7713f3),
	.w5(32'h3b8d60e0),
	.w6(32'hb9419405),
	.w7(32'h3aa529da),
	.w8(32'h3c62987e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c140b22),
	.w1(32'h3c9567df),
	.w2(32'h3cd1ded5),
	.w3(32'h3d1845e2),
	.w4(32'h3cbb14cf),
	.w5(32'hbb40debd),
	.w6(32'h3cc62423),
	.w7(32'h3d225c05),
	.w8(32'hb9f78dfc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e063e),
	.w1(32'h3aeac733),
	.w2(32'h3b6ba530),
	.w3(32'h3b930c49),
	.w4(32'h398f5890),
	.w5(32'hbb21d9ea),
	.w6(32'h3c06432c),
	.w7(32'h3b3046e6),
	.w8(32'hbadea23e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa622f2),
	.w1(32'hba714b3f),
	.w2(32'h3b3f60e1),
	.w3(32'hbad8a737),
	.w4(32'h3baa359f),
	.w5(32'h3c1af43c),
	.w6(32'hbb36f29a),
	.w7(32'h3b22e45e),
	.w8(32'h3c7910ac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf89581),
	.w1(32'hbc004eb4),
	.w2(32'hbcb62b52),
	.w3(32'hbc1151fd),
	.w4(32'hbc21e1ea),
	.w5(32'hbac83e55),
	.w6(32'h3bd4a3e4),
	.w7(32'h3b9b3a04),
	.w8(32'hbba4c7a3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0421c),
	.w1(32'h3a2e6e4f),
	.w2(32'h3b1d50b6),
	.w3(32'h3adfc06e),
	.w4(32'hba46f48f),
	.w5(32'hba06dd71),
	.w6(32'h3b431f11),
	.w7(32'h3b134d1c),
	.w8(32'hbc2246e8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054dd1),
	.w1(32'hbadc3fe6),
	.w2(32'h3c58533e),
	.w3(32'h3c336696),
	.w4(32'h3c3487e6),
	.w5(32'h3c508d25),
	.w6(32'hbc2b4b41),
	.w7(32'hbc0e972c),
	.w8(32'h3c019188),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3858),
	.w1(32'h39bde8a8),
	.w2(32'hb9a1e08c),
	.w3(32'hbade82d0),
	.w4(32'h3be19639),
	.w5(32'h3b060aae),
	.w6(32'hbb1eb357),
	.w7(32'h3b08c59f),
	.w8(32'hbac4ffc4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e77f7),
	.w1(32'hbb5cbc13),
	.w2(32'h3af9f99d),
	.w3(32'h3abf47b1),
	.w4(32'h3a221337),
	.w5(32'hba56c779),
	.w6(32'h39ffa3eb),
	.w7(32'h3a4c70b8),
	.w8(32'hbb2b0f7d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec68b8),
	.w1(32'hbbc73fc5),
	.w2(32'hbb98271e),
	.w3(32'h3b24005f),
	.w4(32'hbbfb1f1d),
	.w5(32'hbcba2012),
	.w6(32'hbc697751),
	.w7(32'hbc8c4cf7),
	.w8(32'hbc365f00),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556bd5),
	.w1(32'hbb849445),
	.w2(32'hbbed58dd),
	.w3(32'h3b5bbfdb),
	.w4(32'hbb6cf9fb),
	.w5(32'h3b7b57c0),
	.w6(32'h3c24e1d8),
	.w7(32'h3bade3c3),
	.w8(32'h3bd91c96),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd051b0),
	.w1(32'h3c4ea671),
	.w2(32'h3ca4c25a),
	.w3(32'h3b344947),
	.w4(32'hbbe265f9),
	.w5(32'h3b869c4c),
	.w6(32'h3bf87ad5),
	.w7(32'h3a540603),
	.w8(32'hbb87ca83),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6cd5),
	.w1(32'h3ac5af39),
	.w2(32'h39d3f3ca),
	.w3(32'h3b8c98e4),
	.w4(32'h3aab8bef),
	.w5(32'hbb759c6f),
	.w6(32'hbbb00603),
	.w7(32'h3c0f32fe),
	.w8(32'hbb3a77bb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae36d78),
	.w1(32'h3bf61207),
	.w2(32'h3b69ace3),
	.w3(32'hbbc3ba2a),
	.w4(32'hbb2b379d),
	.w5(32'hbacd5d49),
	.w6(32'h3b956ff2),
	.w7(32'hbbb112d5),
	.w8(32'h3b17b426),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021712),
	.w1(32'hbbcf405a),
	.w2(32'hbc1a6a3e),
	.w3(32'h3b0faf1d),
	.w4(32'h3b5eef89),
	.w5(32'hbb4bd8d0),
	.w6(32'hbbde868b),
	.w7(32'hbbaf2aaa),
	.w8(32'h39a35b93),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69ab6),
	.w1(32'hbb50218d),
	.w2(32'hbb064a02),
	.w3(32'hbc161563),
	.w4(32'h3ad452d3),
	.w5(32'hb968b3c5),
	.w6(32'hbc64bd4f),
	.w7(32'h391787e4),
	.w8(32'hbbe7d344),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a05fb),
	.w1(32'hb9dee249),
	.w2(32'hbb6ae90e),
	.w3(32'hbb093b79),
	.w4(32'h3c5da80d),
	.w5(32'hbb081825),
	.w6(32'hbc0e7638),
	.w7(32'hbc2407f4),
	.w8(32'hbbca891c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80b573),
	.w1(32'h3bf16a09),
	.w2(32'hbc151713),
	.w3(32'h3b04f7a0),
	.w4(32'h3acc9741),
	.w5(32'h3bbd78f6),
	.w6(32'h3b2c62f3),
	.w7(32'hbbdda2e8),
	.w8(32'hba83b461),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ad0a4),
	.w1(32'h3ce03b55),
	.w2(32'hb9ddbb4f),
	.w3(32'h39b6c5d1),
	.w4(32'h3c79871b),
	.w5(32'h3c83fe10),
	.w6(32'h3acd5d75),
	.w7(32'h3c77b0b2),
	.w8(32'h3bd91176),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dcd47),
	.w1(32'hbaa75af7),
	.w2(32'h3ceedd03),
	.w3(32'hba87c65a),
	.w4(32'h3c02b026),
	.w5(32'h3c4a0302),
	.w6(32'h38fdc78c),
	.w7(32'h3bd550c3),
	.w8(32'h3c332771),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56ba65),
	.w1(32'hbbeba193),
	.w2(32'h3c4f9e58),
	.w3(32'hbb1c1237),
	.w4(32'hbc63c630),
	.w5(32'h3b2e0bd2),
	.w6(32'h3c14d1e6),
	.w7(32'h3a84d60e),
	.w8(32'hba337fea),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be70c70),
	.w1(32'hb9bfd16d),
	.w2(32'h3b0963ac),
	.w3(32'h398ff273),
	.w4(32'h3ba3bd62),
	.w5(32'hba40ac11),
	.w6(32'hbc1fb468),
	.w7(32'h3ad29219),
	.w8(32'h3c0852f0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db64d),
	.w1(32'hbc2dfee9),
	.w2(32'hbbac59f3),
	.w3(32'hbc487c0a),
	.w4(32'h3b84b26b),
	.w5(32'h39e3c97f),
	.w6(32'hbc5f3c9f),
	.w7(32'h3b93f728),
	.w8(32'hbac79a81),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3349f),
	.w1(32'hbb090e2d),
	.w2(32'h3b205b29),
	.w3(32'hbac40840),
	.w4(32'h3bd91988),
	.w5(32'h3b03dacf),
	.w6(32'hba98dfce),
	.w7(32'h3b707bde),
	.w8(32'h3b762be0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf06e4a),
	.w1(32'h3ab53cbb),
	.w2(32'h3b9f723d),
	.w3(32'hba4bcd6e),
	.w4(32'h3bee0019),
	.w5(32'hbbdcf3b3),
	.w6(32'hbaac845f),
	.w7(32'h3bf339b4),
	.w8(32'hbb52a8c4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21893),
	.w1(32'hbbe9fb6b),
	.w2(32'hbc8278cb),
	.w3(32'hbc2017a7),
	.w4(32'hbb884605),
	.w5(32'hbcbfb711),
	.w6(32'hbc31a83f),
	.w7(32'hba733ff8),
	.w8(32'hbc6fddaf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb331159),
	.w1(32'h3b995470),
	.w2(32'h3b468cfc),
	.w3(32'hba2876b3),
	.w4(32'h3c0c023c),
	.w5(32'h3b86c104),
	.w6(32'h3aa5973e),
	.w7(32'h3afacf44),
	.w8(32'hba8854fa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ecc3),
	.w1(32'h3bb9d51b),
	.w2(32'h3a8ec19a),
	.w3(32'h3bf3cdd3),
	.w4(32'h3b565fb7),
	.w5(32'h3b8d02f2),
	.w6(32'h3ba997b3),
	.w7(32'h3bcca969),
	.w8(32'h3b525c1d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a994a42),
	.w1(32'hbb03543a),
	.w2(32'hbb8bcf77),
	.w3(32'h3c1f6535),
	.w4(32'h3b7b7a73),
	.w5(32'hbb0d57a0),
	.w6(32'hbb762fa3),
	.w7(32'hb97bf15c),
	.w8(32'hb9d246eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813a40),
	.w1(32'hbb5b7988),
	.w2(32'hbce256a8),
	.w3(32'hbab33383),
	.w4(32'hb9f2db18),
	.w5(32'hbc72b061),
	.w6(32'hbb6c618a),
	.w7(32'hbb8f6b9e),
	.w8(32'hbc77ea16),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9897e74),
	.w1(32'h3a97e52d),
	.w2(32'hb7fc18fc),
	.w3(32'h3b15669a),
	.w4(32'h3a9f78f6),
	.w5(32'hbbc4d96d),
	.w6(32'h3acdf614),
	.w7(32'h3b074582),
	.w8(32'hbba598ba),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f790),
	.w1(32'hbb48793c),
	.w2(32'hbaf2f982),
	.w3(32'hbbcf374a),
	.w4(32'h3b0c260a),
	.w5(32'hbad4e2aa),
	.w6(32'hbbe8e09f),
	.w7(32'hbb4ca1bd),
	.w8(32'h3b4523ae),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4ba75),
	.w1(32'h3bc3cd18),
	.w2(32'h3b951da7),
	.w3(32'h3b40beff),
	.w4(32'hb9a5f985),
	.w5(32'hbb59e8f4),
	.w6(32'hbb533fc3),
	.w7(32'hbba25f16),
	.w8(32'h3a7a51e9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1749e0),
	.w1(32'hbad839e8),
	.w2(32'h3b143949),
	.w3(32'hbb30394f),
	.w4(32'hbb7bb5d5),
	.w5(32'hbc3b3684),
	.w6(32'h3c2c2170),
	.w7(32'h3c0023ac),
	.w8(32'hbc154c08),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7d3c),
	.w1(32'hbc7bc9f6),
	.w2(32'hbc5e6b35),
	.w3(32'hbc6c3d5f),
	.w4(32'hbc1efa6b),
	.w5(32'hbaae4e76),
	.w6(32'hbc61cb71),
	.w7(32'hbbad9f02),
	.w8(32'h3a331163),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31d8dd),
	.w1(32'hbc2f6da7),
	.w2(32'hbce43412),
	.w3(32'hbb9b97f7),
	.w4(32'hbb2ea970),
	.w5(32'hbc1950ce),
	.w6(32'hbae6c185),
	.w7(32'hbb1105f9),
	.w8(32'hbb4fa101),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1dd0),
	.w1(32'h3c2f32f5),
	.w2(32'h3a936721),
	.w3(32'h3c03e5ac),
	.w4(32'hba959189),
	.w5(32'hbbf05776),
	.w6(32'h3ccb1fad),
	.w7(32'h3c0e8915),
	.w8(32'hbc31d2bc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c360247),
	.w1(32'hbc33ddba),
	.w2(32'hbb13bab5),
	.w3(32'h3ba9c4e6),
	.w4(32'h3c881cb7),
	.w5(32'h3b44cac3),
	.w6(32'hbc861857),
	.w7(32'h39dfd4fd),
	.w8(32'h3c4ed697),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d9167),
	.w1(32'hbb1c88cb),
	.w2(32'hba11bb3a),
	.w3(32'h3af036e9),
	.w4(32'h3c97bd6d),
	.w5(32'h3ac13955),
	.w6(32'hbc258424),
	.w7(32'h3ba7d90b),
	.w8(32'h3acb9000),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45e43b),
	.w1(32'h3babf67c),
	.w2(32'h3c058f9b),
	.w3(32'h3c6430a0),
	.w4(32'h3c12905f),
	.w5(32'hbb588174),
	.w6(32'h3c153557),
	.w7(32'h3c581fbb),
	.w8(32'hbaee91f4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89a123),
	.w1(32'h3a90e763),
	.w2(32'h3af8c84a),
	.w3(32'hbbaebb72),
	.w4(32'h3b275bc3),
	.w5(32'h399cdc97),
	.w6(32'hb9e6bf59),
	.w7(32'hba984f99),
	.w8(32'hba37fbd0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8f5f),
	.w1(32'hbb89c95f),
	.w2(32'h38c5e648),
	.w3(32'hbb58f747),
	.w4(32'h3b6a5874),
	.w5(32'h3b3e0868),
	.w6(32'hbc1602bc),
	.w7(32'hbb3b64af),
	.w8(32'hba0c5b9b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2c60a),
	.w1(32'hbb8e12e1),
	.w2(32'hbc39390c),
	.w3(32'h3ba87d80),
	.w4(32'hbb2429c7),
	.w5(32'hbc1d5613),
	.w6(32'h3b55a18d),
	.w7(32'h3b1e31ac),
	.w8(32'hbbced1c6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25f36d),
	.w1(32'hbc603a9c),
	.w2(32'hbc428d15),
	.w3(32'hbc1b8470),
	.w4(32'hbbb97fa8),
	.w5(32'hbc444277),
	.w6(32'hbbe54695),
	.w7(32'hbbbef711),
	.w8(32'hbca3b070),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14e9b3),
	.w1(32'hbbd95e99),
	.w2(32'h3ae1d5ea),
	.w3(32'hbbee5742),
	.w4(32'hbb816cd4),
	.w5(32'h3b1c480d),
	.w6(32'hba29866c),
	.w7(32'hbc5bd183),
	.w8(32'h3ba37071),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e1f10),
	.w1(32'hbb5d5987),
	.w2(32'hbb8a765e),
	.w3(32'hbbcaafe6),
	.w4(32'h3c9ab3c2),
	.w5(32'hbbc5a70c),
	.w6(32'hbbd171e1),
	.w7(32'hbb24bd8d),
	.w8(32'hbc1091bb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38de9b),
	.w1(32'hb99a8071),
	.w2(32'hbbe53d0a),
	.w3(32'hbbd484ac),
	.w4(32'hbb155698),
	.w5(32'hbbfdd974),
	.w6(32'h3c36db4a),
	.w7(32'hbc288e08),
	.w8(32'h3be4ff48),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc369ab3),
	.w1(32'hbb85f1c8),
	.w2(32'hbae30ac5),
	.w3(32'hbc3b7f00),
	.w4(32'hbbd0b9f3),
	.w5(32'hbb47ae4b),
	.w6(32'h3b33b526),
	.w7(32'h3b48f4db),
	.w8(32'hbba99a6c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b747c),
	.w1(32'hbbbd81d8),
	.w2(32'hbcaf4fd8),
	.w3(32'h3bf8761c),
	.w4(32'h3c1e6038),
	.w5(32'hbb6c6204),
	.w6(32'hbb7e2c96),
	.w7(32'hbb2f3773),
	.w8(32'hbca219d7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b8269),
	.w1(32'hbb2e95b0),
	.w2(32'hbc3ee173),
	.w3(32'h3c5b158f),
	.w4(32'h3c432a26),
	.w5(32'hbb4157b0),
	.w6(32'h3c7dd33c),
	.w7(32'h3c2dad4c),
	.w8(32'h3a310d36),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db160),
	.w1(32'hbbe1704d),
	.w2(32'hbcbc42a1),
	.w3(32'hb8b6df66),
	.w4(32'hbba341d6),
	.w5(32'hbbc16dfc),
	.w6(32'h3b112d09),
	.w7(32'hbc0f5e7a),
	.w8(32'hbc410fe7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ee34),
	.w1(32'h3bf0f4d4),
	.w2(32'h3c89de61),
	.w3(32'hbae17851),
	.w4(32'h3bd5691c),
	.w5(32'h3c0f8199),
	.w6(32'hbc7a110e),
	.w7(32'hba7b1e0c),
	.w8(32'h39fcc997),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f23f),
	.w1(32'h3a8bbe8b),
	.w2(32'h3b90ee65),
	.w3(32'hbba17b5a),
	.w4(32'h3af48470),
	.w5(32'h3b6045fc),
	.w6(32'hbb9bac99),
	.w7(32'h3b063c27),
	.w8(32'h3a0a23bf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f9ad),
	.w1(32'hbb5ad2f0),
	.w2(32'h3af96a47),
	.w3(32'hbb117722),
	.w4(32'hbb5939d7),
	.w5(32'hbb31f5f1),
	.w6(32'hbb13d8dd),
	.w7(32'hbb7fc4f9),
	.w8(32'h3bc12765),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce2138),
	.w1(32'hbb12fcb9),
	.w2(32'h3a17c54c),
	.w3(32'hbbcc8c14),
	.w4(32'hbbb82b08),
	.w5(32'h3a3bc9dd),
	.w6(32'h3b99ee6f),
	.w7(32'hbb600d38),
	.w8(32'h3b273c3a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b34b9),
	.w1(32'h3b2befa4),
	.w2(32'hbbb37b99),
	.w3(32'h3ba2f329),
	.w4(32'h3b60297c),
	.w5(32'hbb811d6a),
	.w6(32'h3b17b67a),
	.w7(32'h3b3fad68),
	.w8(32'hbbe3ae99),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0fdbd),
	.w1(32'hbbb1f221),
	.w2(32'h3aaeaf10),
	.w3(32'hba534936),
	.w4(32'h3b104d84),
	.w5(32'h395aed68),
	.w6(32'hbb8e547e),
	.w7(32'h3babf735),
	.w8(32'hba721d16),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d92d),
	.w1(32'hbb739192),
	.w2(32'hbc21982f),
	.w3(32'h3adeeac0),
	.w4(32'hba1b0843),
	.w5(32'hba196ac5),
	.w6(32'h3b286a79),
	.w7(32'h3b4bb105),
	.w8(32'hbb585d60),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c339077),
	.w1(32'hbba7b103),
	.w2(32'hbc4640d7),
	.w3(32'hbc083279),
	.w4(32'h3ac73c02),
	.w5(32'hbb9d7766),
	.w6(32'hbaa0ea5e),
	.w7(32'h3c8c6e43),
	.w8(32'hbc17183f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098212),
	.w1(32'h3b16fa71),
	.w2(32'h3bb25931),
	.w3(32'hbbd43b11),
	.w4(32'hbb6e1b91),
	.w5(32'h3af08d30),
	.w6(32'hbaa0061a),
	.w7(32'hba5a8902),
	.w8(32'hba0c4516),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f0a3),
	.w1(32'hbb95b48d),
	.w2(32'hbb9ac147),
	.w3(32'h3a781a9c),
	.w4(32'hb73379cc),
	.w5(32'hbb603fdb),
	.w6(32'hbb85e4af),
	.w7(32'h3aebf45e),
	.w8(32'hbb52a43d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d644),
	.w1(32'h3b6ed38f),
	.w2(32'hbc2437d8),
	.w3(32'h3b84930c),
	.w4(32'h3b5d3c7f),
	.w5(32'hbbcf1529),
	.w6(32'hbaf03a50),
	.w7(32'hbb994314),
	.w8(32'hbc2e5a3f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc8b6d),
	.w1(32'hbbdbd1d5),
	.w2(32'hbaa2600b),
	.w3(32'h3a8dbf58),
	.w4(32'h3ab53dd3),
	.w5(32'hbb8d40b5),
	.w6(32'hbbb18f46),
	.w7(32'hba950c64),
	.w8(32'hbaac74ac),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa09b),
	.w1(32'hbb3cc5e2),
	.w2(32'hbc139405),
	.w3(32'h37ca045b),
	.w4(32'h3af5e089),
	.w5(32'hbbd196e2),
	.w6(32'hbba5de21),
	.w7(32'h3aa0f522),
	.w8(32'hbc9c87bc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1748b0),
	.w1(32'hbc67923a),
	.w2(32'hbc6914ea),
	.w3(32'hbb66f818),
	.w4(32'hbbbf4296),
	.w5(32'hb9a31987),
	.w6(32'hbc0fe053),
	.w7(32'hbbd74e19),
	.w8(32'hbc01f0f1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2347c),
	.w1(32'hbc0560ba),
	.w2(32'hbb0690ea),
	.w3(32'h3babb829),
	.w4(32'hbacaccb6),
	.w5(32'hbbde61ec),
	.w6(32'h3b8f9895),
	.w7(32'hba138bbd),
	.w8(32'hbc1d0e9b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37875aad),
	.w1(32'hbbe8da44),
	.w2(32'hbbfa4acf),
	.w3(32'hbbc158cf),
	.w4(32'hbbe47d62),
	.w5(32'h3ae8b0d1),
	.w6(32'hbbf0edec),
	.w7(32'hbbb3dca0),
	.w8(32'h3a0c1eaa),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d50ca),
	.w1(32'hbb7ec345),
	.w2(32'hbb5b31c6),
	.w3(32'hbae0cda9),
	.w4(32'hbc059257),
	.w5(32'hbb08e33b),
	.w6(32'h380db630),
	.w7(32'hbb768a34),
	.w8(32'hba22c096),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b739f),
	.w1(32'h3a973021),
	.w2(32'h3c20590a),
	.w3(32'h3bcc8726),
	.w4(32'h3bb02ac8),
	.w5(32'h3c18bbfc),
	.w6(32'hbac53cd1),
	.w7(32'h3bd77bb0),
	.w8(32'h3cb40676),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f29fe),
	.w1(32'h3c078d2b),
	.w2(32'h3b9e7b80),
	.w3(32'h3c7807d6),
	.w4(32'h3c9b06e6),
	.w5(32'hbabd37da),
	.w6(32'h3c8fdd2a),
	.w7(32'h3cf04666),
	.w8(32'hbab49246),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5571),
	.w1(32'h3a221d9a),
	.w2(32'h3a86b5c4),
	.w3(32'h3ba87a7a),
	.w4(32'h3c13a127),
	.w5(32'hba0e8c3b),
	.w6(32'hbacaf634),
	.w7(32'h3c0491aa),
	.w8(32'hbb14996e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4606e2),
	.w1(32'hbc32d2ee),
	.w2(32'hbc97889f),
	.w3(32'hbc06f91d),
	.w4(32'hbc5ebfcb),
	.w5(32'hbbd22034),
	.w6(32'h3a2f1ebc),
	.w7(32'hbc377929),
	.w8(32'hbc489e3e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2929d0),
	.w1(32'hb99d4c83),
	.w2(32'h3b1c3215),
	.w3(32'h3908f214),
	.w4(32'hbbb4ae70),
	.w5(32'h3af77f82),
	.w6(32'h3b43bfaa),
	.w7(32'h3ac307b9),
	.w8(32'h3b2d7f32),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd3c3),
	.w1(32'hbb18b93a),
	.w2(32'hbc28dcd0),
	.w3(32'h3c4b3c5a),
	.w4(32'h3bc683fe),
	.w5(32'hbc16a585),
	.w6(32'h3c678698),
	.w7(32'h3c26918b),
	.w8(32'hbc56f95a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add675d),
	.w1(32'h3ab89d8e),
	.w2(32'h3c1e9113),
	.w3(32'hbbbef1d3),
	.w4(32'hbbc3a50a),
	.w5(32'h3bef44cb),
	.w6(32'h3b607072),
	.w7(32'hbbafe386),
	.w8(32'h3bd8df75),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e7af9a),
	.w1(32'hba0ea3ef),
	.w2(32'hbc19a8f1),
	.w3(32'h3c8a3d25),
	.w4(32'h3bd56ea5),
	.w5(32'hbb8aab7a),
	.w6(32'h3c32e2aa),
	.w7(32'h3a1ca1e5),
	.w8(32'hbb4ace3a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a66a9),
	.w1(32'hbbb713fa),
	.w2(32'hbb9a97fe),
	.w3(32'hb9c301f1),
	.w4(32'h3bb06f57),
	.w5(32'hbb3ec944),
	.w6(32'hbb40a95a),
	.w7(32'hb9d4f474),
	.w8(32'hbb302b4e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0715),
	.w1(32'hbb2406fa),
	.w2(32'h3c237b6c),
	.w3(32'hbbabcb2e),
	.w4(32'hbbbabdfa),
	.w5(32'h3b8d667e),
	.w6(32'hbb88496f),
	.w7(32'hbad7982a),
	.w8(32'hba010e46),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e9d7),
	.w1(32'h3b0b61b6),
	.w2(32'h3a4c95b6),
	.w3(32'h3b02ef0b),
	.w4(32'h3b0e2579),
	.w5(32'hbae0b17e),
	.w6(32'hbb80baad),
	.w7(32'h3b31e53e),
	.w8(32'hbb4089c7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99588a),
	.w1(32'hbc071a6a),
	.w2(32'hbc80e67b),
	.w3(32'hbc0f0a46),
	.w4(32'h3bad8973),
	.w5(32'hbbd440ca),
	.w6(32'hb9c51992),
	.w7(32'h3b7613b1),
	.w8(32'hbc0f35f8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a98f6),
	.w1(32'hbb965824),
	.w2(32'hbc857dc8),
	.w3(32'h3b8a53d2),
	.w4(32'h3bdd0d3f),
	.w5(32'h3901cc6f),
	.w6(32'h3ae0dcb8),
	.w7(32'h3ab93bc5),
	.w8(32'hbb9f6152),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb098d6),
	.w1(32'h3b983ef7),
	.w2(32'hbab51e5e),
	.w3(32'hbc5f9551),
	.w4(32'hbb17933b),
	.w5(32'h3c4fa3b9),
	.w6(32'hbb617fd7),
	.w7(32'h3c48884d),
	.w8(32'h3c176858),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed3f1),
	.w1(32'h3b9f6692),
	.w2(32'h3c99344e),
	.w3(32'h3ba772ab),
	.w4(32'h3c335815),
	.w5(32'h3cbe1257),
	.w6(32'hbb915fcf),
	.w7(32'h3bf660be),
	.w8(32'h3c21f8a9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724fd7),
	.w1(32'h3b611622),
	.w2(32'h3c0c682a),
	.w3(32'h3b994f0f),
	.w4(32'h3bad6029),
	.w5(32'h3a444f27),
	.w6(32'hbc06856c),
	.w7(32'hbb6d74ab),
	.w8(32'hba200326),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0815e),
	.w1(32'h3ba86311),
	.w2(32'hbc338be2),
	.w3(32'h3b08e6ca),
	.w4(32'h3bec9cf8),
	.w5(32'h3c00510f),
	.w6(32'h3aec6c13),
	.w7(32'h3c1343b4),
	.w8(32'hbb840671),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb423388),
	.w1(32'hbbd25574),
	.w2(32'hbb9c3b99),
	.w3(32'hbacb3e9f),
	.w4(32'h3adcd266),
	.w5(32'h3990d1ad),
	.w6(32'hbb6bc8a5),
	.w7(32'hbb31829d),
	.w8(32'hbb3a47bd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fce59),
	.w1(32'hbb74a68e),
	.w2(32'hbc01f3f5),
	.w3(32'hbc1f85a2),
	.w4(32'hbb5f110d),
	.w5(32'h3c326b9c),
	.w6(32'hbafef348),
	.w7(32'hb9fa28f1),
	.w8(32'h3c0b35ea),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a2b3),
	.w1(32'h3b31d592),
	.w2(32'hbb627158),
	.w3(32'hbadb9e41),
	.w4(32'h3ac2321c),
	.w5(32'hba9fbfa7),
	.w6(32'hbaf27e03),
	.w7(32'h3b7b7a7c),
	.w8(32'hbb482d1a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dd8da),
	.w1(32'hbb68bb54),
	.w2(32'hbb193057),
	.w3(32'hbb27cac4),
	.w4(32'h3b1c3f49),
	.w5(32'hbb0ca459),
	.w6(32'hbb9d6d6d),
	.w7(32'hba3ba3bf),
	.w8(32'hbadf3702),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aed27),
	.w1(32'hbba8cbf9),
	.w2(32'hbb981b13),
	.w3(32'hbb49ccce),
	.w4(32'hba733737),
	.w5(32'h3a83b19a),
	.w6(32'hbbe070ec),
	.w7(32'hbaf1e5a5),
	.w8(32'hb9e50f51),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37aaca),
	.w1(32'h3b88832b),
	.w2(32'hbab3a378),
	.w3(32'h3b534d90),
	.w4(32'h3b87910b),
	.w5(32'hbbfb56e3),
	.w6(32'h3ae8660b),
	.w7(32'h3b8a10b0),
	.w8(32'hbbeefb39),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9668a0),
	.w1(32'h3a5c6ea4),
	.w2(32'h3bc229b8),
	.w3(32'hba91d327),
	.w4(32'h3ad9f4df),
	.w5(32'h3ac1022a),
	.w6(32'hbaa4cb85),
	.w7(32'h3b18fbe9),
	.w8(32'h3a15645a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa4ec),
	.w1(32'hbc0cc37f),
	.w2(32'h3a67ab9f),
	.w3(32'hbadc5628),
	.w4(32'hbc1c92f2),
	.w5(32'h3ad632bf),
	.w6(32'hbb4a072b),
	.w7(32'hbc17958d),
	.w8(32'h3b932806),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b415b9e),
	.w1(32'h3b0be484),
	.w2(32'h3a7451f3),
	.w3(32'h3a0b0868),
	.w4(32'h3ab0bc3c),
	.w5(32'h3b4fa437),
	.w6(32'hba0c9f11),
	.w7(32'hbb3fca52),
	.w8(32'h3aa819c6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb330d8),
	.w1(32'h3c2ba76c),
	.w2(32'h3aa88790),
	.w3(32'h3b252d84),
	.w4(32'h3bd26681),
	.w5(32'h3b2f38ad),
	.w6(32'h3c019446),
	.w7(32'h3c2b3605),
	.w8(32'h3c0c585e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae60f3c),
	.w1(32'hbb67ed9d),
	.w2(32'hbbfed6e7),
	.w3(32'h3ab4d96d),
	.w4(32'hbb8ea52a),
	.w5(32'hbc0ae8bd),
	.w6(32'hbb7b0194),
	.w7(32'h3ad108e2),
	.w8(32'hbb9bc049),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f07d8),
	.w1(32'hb9d5756a),
	.w2(32'h3b699c68),
	.w3(32'h3b21e8da),
	.w4(32'h3bccc19f),
	.w5(32'h3bae9de9),
	.w6(32'hbb361c67),
	.w7(32'h3bfaba86),
	.w8(32'h3b8f893a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa524f7),
	.w1(32'hbb222d76),
	.w2(32'hbb6ce6e6),
	.w3(32'h3a29b360),
	.w4(32'h397ad9db),
	.w5(32'h3bb4fa14),
	.w6(32'hbb06d7e2),
	.w7(32'hbb0d6b27),
	.w8(32'h3bd7e20a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a7bb),
	.w1(32'h3ba8c234),
	.w2(32'h39b92ba3),
	.w3(32'h3be96558),
	.w4(32'h3b72ec4e),
	.w5(32'hba890b0e),
	.w6(32'h3bf8ec5a),
	.w7(32'h3b2bb898),
	.w8(32'hbb75638a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0979ca),
	.w1(32'hbb65a57c),
	.w2(32'hbb3a1f89),
	.w3(32'hb99dd305),
	.w4(32'h3b105c4a),
	.w5(32'hba551253),
	.w6(32'hbb8b9080),
	.w7(32'hbb10f5e6),
	.w8(32'hbb4b55f5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba586c52),
	.w1(32'hbb214336),
	.w2(32'hbaa12436),
	.w3(32'hbaaaf564),
	.w4(32'hba5e992d),
	.w5(32'h3c500d8b),
	.w6(32'hbb8eadfa),
	.w7(32'hbb76586c),
	.w8(32'h3c2bab8c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31ecb7),
	.w1(32'h3c1c7d56),
	.w2(32'h3c702f50),
	.w3(32'h3c62a881),
	.w4(32'h3c87b2bd),
	.w5(32'h3b166803),
	.w6(32'h3c2a991e),
	.w7(32'h3c79ca57),
	.w8(32'h3b98cae9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b5d05),
	.w1(32'hbb1a815a),
	.w2(32'hbbc4f443),
	.w3(32'h39801377),
	.w4(32'hbacb49fa),
	.w5(32'hba6bc602),
	.w6(32'h3bb50736),
	.w7(32'hbb39b304),
	.w8(32'hb951c668),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d61e),
	.w1(32'hb80259a6),
	.w2(32'hbbcb1e57),
	.w3(32'h3b820dbe),
	.w4(32'h3b2d6273),
	.w5(32'hbad2735a),
	.w6(32'h39f5a06a),
	.w7(32'h3abc0a4b),
	.w8(32'hbb5691f1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59e2c),
	.w1(32'h3b98db95),
	.w2(32'h3c4e7435),
	.w3(32'hbb3e4b93),
	.w4(32'hba2791a0),
	.w5(32'h3b1d5196),
	.w6(32'hbbb7b49b),
	.w7(32'hbbe9201f),
	.w8(32'h3ad665d1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6931),
	.w1(32'hba8decb3),
	.w2(32'hb9e7ea3a),
	.w3(32'hb9e35241),
	.w4(32'hbb0734ed),
	.w5(32'hbaf94e72),
	.w6(32'hb98876bc),
	.w7(32'h3a26a346),
	.w8(32'hba727a32),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb2d9d),
	.w1(32'hbb1b8a31),
	.w2(32'hbac22560),
	.w3(32'hb9aba2d1),
	.w4(32'hba9c91ee),
	.w5(32'h3a9ec140),
	.w6(32'hbaf23338),
	.w7(32'hba86dfc4),
	.w8(32'hbb0fa37c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2ad1),
	.w1(32'hb9c6dc7c),
	.w2(32'hbb231a32),
	.w3(32'hbac19e87),
	.w4(32'hbb1a14a1),
	.w5(32'hbb573d99),
	.w6(32'hbbbfbd52),
	.w7(32'hbbdaf231),
	.w8(32'hbb4a93a3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a794c),
	.w1(32'hbb91ee23),
	.w2(32'hbb87b76e),
	.w3(32'hbb2887e7),
	.w4(32'hb99e520d),
	.w5(32'h3a95bee7),
	.w6(32'hbbb44cee),
	.w7(32'hbb115e3c),
	.w8(32'h3b3686e9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ce64b),
	.w1(32'hbad3728b),
	.w2(32'hbbf92ae8),
	.w3(32'h3bd8eaf0),
	.w4(32'h3c022d7d),
	.w5(32'hbc616439),
	.w6(32'h3c5c7049),
	.w7(32'h3c01b91c),
	.w8(32'hbc290e20),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ec33f),
	.w1(32'hbb150397),
	.w2(32'hbc6b8508),
	.w3(32'hba9f9773),
	.w4(32'hbb2e6fd7),
	.w5(32'hbc2a7299),
	.w6(32'hba7baee7),
	.w7(32'hbb778d6e),
	.w8(32'hbc1c3e6a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a337370),
	.w1(32'hbb4e434d),
	.w2(32'hbbd6d45c),
	.w3(32'hb9f7b2c4),
	.w4(32'h399e922e),
	.w5(32'h3b3e6636),
	.w6(32'hbb08eb96),
	.w7(32'hb97d5106),
	.w8(32'h398b35e1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5bb7),
	.w1(32'hbb178f35),
	.w2(32'hbb6c2bfe),
	.w3(32'hbae445c4),
	.w4(32'h3a8732fb),
	.w5(32'hba1b10db),
	.w6(32'hbb07ffa6),
	.w7(32'hba5716b2),
	.w8(32'hba45b3a6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba030aa5),
	.w1(32'h3a3f7f6e),
	.w2(32'hb925cfef),
	.w3(32'h3ad7a4dd),
	.w4(32'hba653fa2),
	.w5(32'h3ac1aeef),
	.w6(32'h3a0a8906),
	.w7(32'hb93a5caf),
	.w8(32'hbb2dcec1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc3296),
	.w1(32'hbb06998b),
	.w2(32'hbaf15223),
	.w3(32'h3abe12e2),
	.w4(32'h3ad6a2b1),
	.w5(32'hb9d097bd),
	.w6(32'hbb5c4164),
	.w7(32'hbafd81ff),
	.w8(32'hb9e40817),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc517e0),
	.w1(32'hbb9b61cb),
	.w2(32'hb9ef2e77),
	.w3(32'h3b5773db),
	.w4(32'h3b4cd071),
	.w5(32'h3b5dd64a),
	.w6(32'hba54f978),
	.w7(32'h3ade9bc3),
	.w8(32'h3b8210de),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80e1f2),
	.w1(32'hb99cb095),
	.w2(32'hbcb7a749),
	.w3(32'h3c117ba0),
	.w4(32'h3bca559f),
	.w5(32'hbbcc3a52),
	.w6(32'hb9d62b21),
	.w7(32'hbb2e2acb),
	.w8(32'hbc426b8d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895248),
	.w1(32'h3bbe32c5),
	.w2(32'h3bf6971f),
	.w3(32'h3abca0d8),
	.w4(32'h3a871f0a),
	.w5(32'h3bd19bd5),
	.w6(32'h3a8b1ede),
	.w7(32'h3a283972),
	.w8(32'h3bdac798),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b749),
	.w1(32'h3ac1655e),
	.w2(32'hbbac7003),
	.w3(32'h3c31762c),
	.w4(32'h3ba563bb),
	.w5(32'hba098797),
	.w6(32'h3bc928dc),
	.w7(32'h3b7af48c),
	.w8(32'hbb2d4025),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9653f),
	.w1(32'hbb8549ce),
	.w2(32'hbc816bba),
	.w3(32'h3b8e2051),
	.w4(32'h3b2ba6ee),
	.w5(32'h3a87e017),
	.w6(32'h3b891c81),
	.w7(32'h3b4a48fa),
	.w8(32'hbb684c6c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a683792),
	.w1(32'h3bd9cb74),
	.w2(32'h3bd067d2),
	.w3(32'h3baf71af),
	.w4(32'h3be33066),
	.w5(32'h3c0c8480),
	.w6(32'h3a162b01),
	.w7(32'h3b89431e),
	.w8(32'h3c03f441),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc635f8),
	.w1(32'hba82ebd3),
	.w2(32'hbc0a6f0f),
	.w3(32'h3bd2d74a),
	.w4(32'h3b65842b),
	.w5(32'hbbd9d137),
	.w6(32'hb870836f),
	.w7(32'hb8d72094),
	.w8(32'hbc0db296),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952461),
	.w1(32'hbb9649a6),
	.w2(32'hbb95dbee),
	.w3(32'hbb9915fa),
	.w4(32'hbb3f715e),
	.w5(32'hbad0f676),
	.w6(32'hbb9b1e4b),
	.w7(32'hbb3c94c7),
	.w8(32'hb91d0ec9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54ee30),
	.w1(32'hbaab22e5),
	.w2(32'h3c569e4e),
	.w3(32'h3b13b138),
	.w4(32'h3a3aeaf1),
	.w5(32'h3c29f8c9),
	.w6(32'h3ad76c40),
	.w7(32'hbb9fe4a6),
	.w8(32'h3b8c8776),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab304a7),
	.w1(32'h3b13957b),
	.w2(32'h3b12b01a),
	.w3(32'h3ba91aec),
	.w4(32'h3a679969),
	.w5(32'hbb3cbdac),
	.w6(32'h3af9e03d),
	.w7(32'h3ab597be),
	.w8(32'hbb4b3f91),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c7c3),
	.w1(32'hb9859271),
	.w2(32'hba8a48ff),
	.w3(32'hbb1414b0),
	.w4(32'hba2666d9),
	.w5(32'hb97ad26b),
	.w6(32'hbab118c1),
	.w7(32'h3919d961),
	.w8(32'h3ac70ba0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa57c2),
	.w1(32'h3aece6f6),
	.w2(32'h3a027ba5),
	.w3(32'hba5b774f),
	.w4(32'h3afbe32d),
	.w5(32'h3a604e40),
	.w6(32'hba21eb1c),
	.w7(32'h3ad32b90),
	.w8(32'hba6a58bb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dce46),
	.w1(32'hba482207),
	.w2(32'hb96058be),
	.w3(32'h3b08c69f),
	.w4(32'h3ae413ab),
	.w5(32'h3ba02e06),
	.w6(32'hbb66589d),
	.w7(32'hba1b4cba),
	.w8(32'h399d442f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abef714),
	.w1(32'h3bd2fcdc),
	.w2(32'h3c23e946),
	.w3(32'h3bf11da1),
	.w4(32'h3bfc59f6),
	.w5(32'h3be0c169),
	.w6(32'hbb21ee09),
	.w7(32'h3aaf2bd1),
	.w8(32'h3b8c248e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80dc8),
	.w1(32'h3b2e1061),
	.w2(32'hbb475320),
	.w3(32'hbb3adfc5),
	.w4(32'hbb307987),
	.w5(32'hbbe8a2aa),
	.w6(32'hbb40c067),
	.w7(32'hbaf8bd77),
	.w8(32'hbbd844fc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e02b),
	.w1(32'hbb311b55),
	.w2(32'hbb49cab7),
	.w3(32'hbae52345),
	.w4(32'hba40ccff),
	.w5(32'h3a93fae7),
	.w6(32'hbb2b623e),
	.w7(32'hbb1857a4),
	.w8(32'h3af6c71b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa1781),
	.w1(32'h3aa329a2),
	.w2(32'hbc138fa1),
	.w3(32'h3bc38e64),
	.w4(32'h3aeb2e48),
	.w5(32'hbbff2f0f),
	.w6(32'h3b3f7198),
	.w7(32'hbb152801),
	.w8(32'hbc0b0d47),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8b876),
	.w1(32'h3b9434ee),
	.w2(32'h3b87d572),
	.w3(32'h3a54ddf4),
	.w4(32'h392cf92d),
	.w5(32'hbb648eee),
	.w6(32'hbb43219f),
	.w7(32'h3b090f4b),
	.w8(32'hbb92c6a9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb301e7),
	.w1(32'hbb6c90d1),
	.w2(32'hbc8ce944),
	.w3(32'h3c08bc2f),
	.w4(32'h3b0dc1fd),
	.w5(32'hb96b02c0),
	.w6(32'hba5754e7),
	.w7(32'hba7a03d3),
	.w8(32'hbbb8fbf8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0a12f),
	.w1(32'hbc37b90c),
	.w2(32'hb9ef5d59),
	.w3(32'h3b4379cb),
	.w4(32'hbaa91e8d),
	.w5(32'hbb9b73e2),
	.w6(32'hbb8fb9cc),
	.w7(32'hbc151816),
	.w8(32'hbc257e55),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd7e80),
	.w1(32'hb9a70bd4),
	.w2(32'h3b85e178),
	.w3(32'h3ad2e4ed),
	.w4(32'h3a290149),
	.w5(32'h3b185ec1),
	.w6(32'hbb70243b),
	.w7(32'hba213fbb),
	.w8(32'h3aab7612),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ea1e7),
	.w1(32'hb9886a69),
	.w2(32'h38ee3132),
	.w3(32'h3b04d0c6),
	.w4(32'h3aecf18b),
	.w5(32'hb9d348bb),
	.w6(32'h3ae3d71f),
	.w7(32'h3b1d38e3),
	.w8(32'h39a28e91),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b39a),
	.w1(32'h3a9cd2a5),
	.w2(32'h3b5c60ef),
	.w3(32'h3918d4a2),
	.w4(32'h3b44d8ec),
	.w5(32'h3b238916),
	.w6(32'h3a806d8a),
	.w7(32'h3b50c383),
	.w8(32'h3a990aaa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947261),
	.w1(32'hbb23e733),
	.w2(32'h3b9a6d2f),
	.w3(32'h3ad9c411),
	.w4(32'h3b158405),
	.w5(32'h3b3268d2),
	.w6(32'hbb3823f7),
	.w7(32'hbad09cd9),
	.w8(32'h3b6dd600),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8442),
	.w1(32'h3a6346ec),
	.w2(32'h3bc8a894),
	.w3(32'hbadd5f91),
	.w4(32'hba4a68ea),
	.w5(32'h3acdc3d5),
	.w6(32'hbb0a6c13),
	.w7(32'h39d0b317),
	.w8(32'hbab63126),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad85943),
	.w1(32'hbbf19118),
	.w2(32'hbb9e70a7),
	.w3(32'hbb855eb0),
	.w4(32'hbb9cea35),
	.w5(32'hbb6a9d5e),
	.w6(32'hbbe5811d),
	.w7(32'hbb6593be),
	.w8(32'hbac4dbc3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031ba9),
	.w1(32'hb9da06cd),
	.w2(32'hba9281a3),
	.w3(32'h3ab3d121),
	.w4(32'h3b95cfaa),
	.w5(32'hba760907),
	.w6(32'h3b0506f2),
	.w7(32'h3be05610),
	.w8(32'hbae25be9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9c319),
	.w1(32'h3964dc2a),
	.w2(32'hbbdac77f),
	.w3(32'h3b85de13),
	.w4(32'hb8a90e06),
	.w5(32'hbb92d14b),
	.w6(32'h3b8c3ce0),
	.w7(32'h3b6883f6),
	.w8(32'hbba5860b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abde9ac),
	.w1(32'hbbc1e309),
	.w2(32'hbb9a3f43),
	.w3(32'hbb2e9809),
	.w4(32'hba447093),
	.w5(32'hbb49d0c9),
	.w6(32'hbb824d24),
	.w7(32'hbb85b914),
	.w8(32'hbb13aac7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6b15c),
	.w1(32'hb9fa5283),
	.w2(32'h3af465fa),
	.w3(32'hbb317532),
	.w4(32'h3ad48ac4),
	.w5(32'h3a8fbc03),
	.w6(32'h3a38de02),
	.w7(32'h3ab82c3d),
	.w8(32'h3af51fa9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d8b64),
	.w1(32'hb9f98dc9),
	.w2(32'h3a0b7792),
	.w3(32'h3a81383f),
	.w4(32'h3aa20a35),
	.w5(32'hba4121ba),
	.w6(32'hbb3bf32e),
	.w7(32'h3a868dbb),
	.w8(32'h39ce8d42),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e5cda),
	.w1(32'h3bbd1c41),
	.w2(32'hbab9cc43),
	.w3(32'h3b91e75e),
	.w4(32'hbb028bcd),
	.w5(32'hbb0664d3),
	.w6(32'h3bdebd4b),
	.w7(32'hbb0e34a3),
	.w8(32'hbc2d8bdc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1554f2),
	.w1(32'hba5210a3),
	.w2(32'hba8e30d5),
	.w3(32'h3b400b86),
	.w4(32'h3abc4f00),
	.w5(32'h3a05119c),
	.w6(32'hbb877888),
	.w7(32'hbb52b2a9),
	.w8(32'h3a86fb69),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba815799),
	.w1(32'hbb1342cc),
	.w2(32'hbb3a644c),
	.w3(32'h3a1a3c7f),
	.w4(32'hb970f5de),
	.w5(32'h3b45a1f4),
	.w6(32'h39e9c063),
	.w7(32'h3a05cc0d),
	.w8(32'h3a871183),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7af74f),
	.w1(32'h3b3a85c2),
	.w2(32'h3bee498e),
	.w3(32'h3b3f6223),
	.w4(32'h3c0aacb8),
	.w5(32'h3a9547bf),
	.w6(32'hb9545a70),
	.w7(32'h3b8f8312),
	.w8(32'h3b381e91),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40c4ce),
	.w1(32'h3b53bf0f),
	.w2(32'hbc22868d),
	.w3(32'h3b97ae14),
	.w4(32'h3a6146ef),
	.w5(32'h3a99cd70),
	.w6(32'h3ac3d5cb),
	.w7(32'hbb0b029b),
	.w8(32'hbb8d6aa3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9c623),
	.w1(32'hba650825),
	.w2(32'h39cc7686),
	.w3(32'hba0220bf),
	.w4(32'h3aaffe9d),
	.w5(32'h3ba76a39),
	.w6(32'hbb1eb39b),
	.w7(32'h3a88f2f2),
	.w8(32'h3ae2337d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f765eb),
	.w1(32'h3b825dcd),
	.w2(32'h3b6e10a2),
	.w3(32'h3b3b5217),
	.w4(32'h3ae763f7),
	.w5(32'hbaac46c0),
	.w6(32'hbb6ee73b),
	.w7(32'hbb401513),
	.w8(32'hbb0f05d6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa48a89),
	.w1(32'hbba34724),
	.w2(32'hbbb348f5),
	.w3(32'hba967e92),
	.w4(32'h3a36e7e4),
	.w5(32'h3ba3d46e),
	.w6(32'hbc514262),
	.w7(32'hbb8d3b5b),
	.w8(32'h3b3c6740),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be15f79),
	.w1(32'hbb1bd3ac),
	.w2(32'hbbc27244),
	.w3(32'h3c48e067),
	.w4(32'h3c0d9920),
	.w5(32'hbc20c1fc),
	.w6(32'h3acbcce7),
	.w7(32'h3c3019f9),
	.w8(32'hbb8e17d3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b6b7),
	.w1(32'hbc091146),
	.w2(32'hbc4e0c7e),
	.w3(32'hb999d487),
	.w4(32'hbafb4367),
	.w5(32'hba2efc51),
	.w6(32'h3aae25f0),
	.w7(32'hbacadd93),
	.w8(32'h3b13ff6f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba205ec),
	.w1(32'hbbb29810),
	.w2(32'hbc63d0ff),
	.w3(32'hba2e89ad),
	.w4(32'h39a0ea28),
	.w5(32'hbc1a69c2),
	.w6(32'hbaf53441),
	.w7(32'hbb410c0a),
	.w8(32'hbc2b9451),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba938c0e),
	.w1(32'h3a8d66bb),
	.w2(32'hbb788af5),
	.w3(32'h3a925479),
	.w4(32'hbb199adc),
	.w5(32'hbae38b34),
	.w6(32'h3b6ef1ad),
	.w7(32'hbabcc4a1),
	.w8(32'hbb0749c6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82fb39),
	.w1(32'hbc0a597a),
	.w2(32'hbc10331b),
	.w3(32'h398cf99d),
	.w4(32'hb9e10763),
	.w5(32'hbb0704ea),
	.w6(32'hbb4b42fe),
	.w7(32'hba0595ac),
	.w8(32'hbaef3089),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0a78),
	.w1(32'hbab0ee29),
	.w2(32'hbb546954),
	.w3(32'h3a219314),
	.w4(32'hbb14a735),
	.w5(32'hb9727e65),
	.w6(32'h39d1e382),
	.w7(32'hbad2aa6b),
	.w8(32'hba4d31b7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f2581),
	.w1(32'hbb7a342c),
	.w2(32'h3b0d5191),
	.w3(32'hbb232f11),
	.w4(32'h3b682024),
	.w5(32'h3b6c5dad),
	.w6(32'hba887ae4),
	.w7(32'hb9f79af2),
	.w8(32'hba9a193b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b346ce8),
	.w1(32'h39e58dce),
	.w2(32'h3aacb55f),
	.w3(32'h3b64d725),
	.w4(32'h3b7e28f9),
	.w5(32'h3af9660d),
	.w6(32'hba2acaca),
	.w7(32'h39526c00),
	.w8(32'h3b019236),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaebf12),
	.w1(32'hbbbc0e54),
	.w2(32'hbc12fa2f),
	.w3(32'h39c1f016),
	.w4(32'hbab754c2),
	.w5(32'h3a1d32a0),
	.w6(32'hbb5df13b),
	.w7(32'hb93129a8),
	.w8(32'h3b5ba601),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b355c40),
	.w1(32'hbb5623a5),
	.w2(32'hbb40bf5b),
	.w3(32'hbb021b53),
	.w4(32'hbb969450),
	.w5(32'hba9a82e9),
	.w6(32'hbba5ef44),
	.w7(32'hbb5f457b),
	.w8(32'hbab0b10a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c63d9),
	.w1(32'hbabbc490),
	.w2(32'hbaea1321),
	.w3(32'hbb4d7ce9),
	.w4(32'hbb929d94),
	.w5(32'hbab92a18),
	.w6(32'hbb2b0744),
	.w7(32'hbb1608b3),
	.w8(32'hbb8a3fe0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66df3),
	.w1(32'hbba26d91),
	.w2(32'h3aac5f11),
	.w3(32'hbb04dc34),
	.w4(32'h3ac5b1d8),
	.w5(32'hbb0e0f02),
	.w6(32'hbc049354),
	.w7(32'hbba956b3),
	.w8(32'hbafeaad2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb3c02),
	.w1(32'hbbe5b3a1),
	.w2(32'hbc5657a8),
	.w3(32'hbabdb264),
	.w4(32'hba42256e),
	.w5(32'h3bbe92ca),
	.w6(32'hba787346),
	.w7(32'hbab1345e),
	.w8(32'h3aa837d3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa246),
	.w1(32'h3b8ab9fb),
	.w2(32'hbb6cfba0),
	.w3(32'hbbd8de91),
	.w4(32'hbb525250),
	.w5(32'h3bb551e1),
	.w6(32'hbc0f1328),
	.w7(32'hba37b880),
	.w8(32'h3bf8b508),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b9caf),
	.w1(32'hba4768e5),
	.w2(32'hbac8a874),
	.w3(32'h3b031fb3),
	.w4(32'hba3d5a2e),
	.w5(32'hbaf6ebca),
	.w6(32'h3aa837ef),
	.w7(32'hba12c172),
	.w8(32'hbb8a6b56),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d90b),
	.w1(32'hbbd990ac),
	.w2(32'hbcb893f6),
	.w3(32'h3af4673b),
	.w4(32'h3b31d883),
	.w5(32'hbc3aabaa),
	.w6(32'h3bb54e39),
	.w7(32'h3b3cc233),
	.w8(32'hbc41b247),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db3373),
	.w1(32'hbbdc3abb),
	.w2(32'h3b819378),
	.w3(32'h3c180064),
	.w4(32'h3b55580f),
	.w5(32'hbba044c9),
	.w6(32'hbb817217),
	.w7(32'h39176d68),
	.w8(32'hbb9d2b7c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28ac0f),
	.w1(32'hba07f6e5),
	.w2(32'hbbbd961d),
	.w3(32'hbb1b7ab9),
	.w4(32'hbb1d91ee),
	.w5(32'hbb06ff3c),
	.w6(32'hbb2f06ad),
	.w7(32'hbb17ec6c),
	.w8(32'hbbfb5b78),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99c081),
	.w1(32'hbb948040),
	.w2(32'hbb60bcf1),
	.w3(32'h39b14dcf),
	.w4(32'h3a234e58),
	.w5(32'hbb60d6a0),
	.w6(32'hbb99d5c1),
	.w7(32'hbbaa3646),
	.w8(32'hbb473825),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c1ab),
	.w1(32'hbb1dfa8b),
	.w2(32'h39f741c5),
	.w3(32'hbb48d975),
	.w4(32'hb91acbbf),
	.w5(32'hbb4b31a9),
	.w6(32'hbb80f668),
	.w7(32'h39eb95ef),
	.w8(32'hbb6a4c82),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5296),
	.w1(32'hbb870a35),
	.w2(32'hbb472b69),
	.w3(32'hbb9df137),
	.w4(32'hbbce0eb8),
	.w5(32'hbade8663),
	.w6(32'hbb8ed2cc),
	.w7(32'hbb674e03),
	.w8(32'hbb5ada66),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd49c5),
	.w1(32'h3b8c689a),
	.w2(32'hbbb9e103),
	.w3(32'hbb1f39d9),
	.w4(32'hba6abe39),
	.w5(32'h3b537888),
	.w6(32'hb8eefe62),
	.w7(32'hbac01da7),
	.w8(32'hba4b4703),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db503),
	.w1(32'h3ae3d7cf),
	.w2(32'h3ab0054a),
	.w3(32'h3be6e1fb),
	.w4(32'h3b1aca04),
	.w5(32'hbb00c824),
	.w6(32'h3b95a58d),
	.w7(32'h3ac4ae6e),
	.w8(32'hbb96e97b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022bdd),
	.w1(32'hbb279b33),
	.w2(32'h3b0bfb2e),
	.w3(32'hbc198bfd),
	.w4(32'hbb3bc3c7),
	.w5(32'h3bba315f),
	.w6(32'hbc249bec),
	.w7(32'hbb3571ad),
	.w8(32'h3c046d59),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27c75f),
	.w1(32'hb90a02e6),
	.w2(32'h3b2b6524),
	.w3(32'h3a8074f7),
	.w4(32'hbb31ed98),
	.w5(32'hbaa9bebc),
	.w6(32'hbb57f2cf),
	.w7(32'h3a0ec5e0),
	.w8(32'hbb01af2b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdef812),
	.w1(32'h39f50b25),
	.w2(32'hbc046cfd),
	.w3(32'hb94e4494),
	.w4(32'h3accfb14),
	.w5(32'hbb9dc861),
	.w6(32'h3a768558),
	.w7(32'h39ee475e),
	.w8(32'hbc087ba8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cbd9b),
	.w1(32'hba51a0cd),
	.w2(32'hbb62eb95),
	.w3(32'hbb26e44f),
	.w4(32'hbb5d82e8),
	.w5(32'hbb47d1a0),
	.w6(32'hbba50b78),
	.w7(32'hba53562f),
	.w8(32'hba9929f9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7a2e),
	.w1(32'hbb61a905),
	.w2(32'hbaa3c588),
	.w3(32'hbb76946d),
	.w4(32'hbaf07a25),
	.w5(32'h3acabef7),
	.w6(32'hbb641f64),
	.w7(32'hba9c487a),
	.w8(32'h3a289523),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd6aa),
	.w1(32'hbb744579),
	.w2(32'hbb120ae0),
	.w3(32'hbba84dc6),
	.w4(32'hbb29a87c),
	.w5(32'h39e7406a),
	.w6(32'h3a886f47),
	.w7(32'h3b8b7352),
	.w8(32'h3b2c7234),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae921c3),
	.w1(32'hbaa145a6),
	.w2(32'hb94ba213),
	.w3(32'hba1c1c40),
	.w4(32'h39d452c1),
	.w5(32'hbaa2fa88),
	.w6(32'hbb571be1),
	.w7(32'hbabc3013),
	.w8(32'hbb11ba84),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e541d),
	.w1(32'h3b6502a7),
	.w2(32'hbab6d18d),
	.w3(32'hbabbcaf5),
	.w4(32'h3ad956e3),
	.w5(32'hbb49b124),
	.w6(32'hba70e1eb),
	.w7(32'h3b26576b),
	.w8(32'hbb4323a0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd47e),
	.w1(32'hbba173d5),
	.w2(32'h3bcc27fe),
	.w3(32'h3a8a84f6),
	.w4(32'h3b224ec7),
	.w5(32'h3b99cd71),
	.w6(32'hbb97fd91),
	.w7(32'hbaffa7a2),
	.w8(32'h39a891c3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d1fcd),
	.w1(32'h3af80a8b),
	.w2(32'h3b57a889),
	.w3(32'h3aa6be8a),
	.w4(32'h3b20bc5e),
	.w5(32'h3b42816d),
	.w6(32'hba61ba71),
	.w7(32'h3b23b284),
	.w8(32'h3accb0d2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b47429),
	.w1(32'hba4eb46c),
	.w2(32'hba1e8874),
	.w3(32'h3a6f2383),
	.w4(32'h3b39bede),
	.w5(32'hbaa5302e),
	.w6(32'hbab3582d),
	.w7(32'h3aba6270),
	.w8(32'hbb4ede10),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb835df1),
	.w1(32'hbb4e2153),
	.w2(32'h3bce61bf),
	.w3(32'hba700097),
	.w4(32'h3b34326d),
	.w5(32'h3bbd0284),
	.w6(32'hbb5b6744),
	.w7(32'h39de56a3),
	.w8(32'h3bdca51f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4445f3),
	.w1(32'h3a1d85fd),
	.w2(32'hbb82a50d),
	.w3(32'h3ba9387f),
	.w4(32'h3b9e703c),
	.w5(32'hbbf53845),
	.w6(32'h3b12cc1a),
	.w7(32'h3b2e143e),
	.w8(32'hbc0ce1e8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202e66),
	.w1(32'hbc0e7848),
	.w2(32'hbc0f1719),
	.w3(32'hbc0245af),
	.w4(32'hbbf1380e),
	.w5(32'hbb9907cc),
	.w6(32'hbbdd5230),
	.w7(32'hbbcb53aa),
	.w8(32'hbbe2f691),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1e093),
	.w1(32'hbb184d43),
	.w2(32'h3990712e),
	.w3(32'hbaed1380),
	.w4(32'hb9e3742d),
	.w5(32'hbad2e803),
	.w6(32'hbba72170),
	.w7(32'hbb29473c),
	.w8(32'hba0ba301),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba932e09),
	.w1(32'hbb1f3845),
	.w2(32'hbb43cc6d),
	.w3(32'hbabd6f9d),
	.w4(32'hbb6ab1f8),
	.w5(32'hbbc5b305),
	.w6(32'hbb91aea7),
	.w7(32'hbb750205),
	.w8(32'hbbef20c7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c426),
	.w1(32'hbc0a7148),
	.w2(32'hbc271a88),
	.w3(32'hbb8c3a7a),
	.w4(32'hbbba6616),
	.w5(32'hbbd1e56f),
	.w6(32'h3ba28841),
	.w7(32'h3958a7e9),
	.w8(32'hbb473282),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8672e2),
	.w1(32'hbb23e0d0),
	.w2(32'hbc156658),
	.w3(32'hba00dfc5),
	.w4(32'hba5ff67c),
	.w5(32'hbb85709f),
	.w6(32'hbb8cbf7e),
	.w7(32'hba808d61),
	.w8(32'hbbf53e1b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba488037),
	.w1(32'hbb6fa570),
	.w2(32'hb8c64723),
	.w3(32'hbb233375),
	.w4(32'hbad1ff57),
	.w5(32'h3bc3f575),
	.w6(32'hbb8cbfc8),
	.w7(32'h3a59a525),
	.w8(32'h3b8f552b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c567e2f),
	.w1(32'hba37e108),
	.w2(32'hbc8b8e9d),
	.w3(32'h3ab30cb8),
	.w4(32'h3ba629e4),
	.w5(32'h3b47c531),
	.w6(32'hbba043bc),
	.w7(32'hbb2924b9),
	.w8(32'hbc38ca10),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ae9bc5),
	.w1(32'hba22af9f),
	.w2(32'hbad6857f),
	.w3(32'hb907725c),
	.w4(32'hba414bbe),
	.w5(32'h3b8c72c2),
	.w6(32'hbb9df095),
	.w7(32'hbb96dea6),
	.w8(32'h3b828902),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b725739),
	.w1(32'h3b1b76c3),
	.w2(32'h3aa9e726),
	.w3(32'h3bd1de9b),
	.w4(32'h3b920084),
	.w5(32'hbb572335),
	.w6(32'h3bb8e90f),
	.w7(32'h3b600e50),
	.w8(32'h3907cbd9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2d98),
	.w1(32'h3c4fba45),
	.w2(32'hbc2261b5),
	.w3(32'hbb8b4fb1),
	.w4(32'h3b8d8c8d),
	.w5(32'hbac801d3),
	.w6(32'h3b4273f0),
	.w7(32'h3c170ac0),
	.w8(32'hbbafb3fe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07cbf9),
	.w1(32'hbbc2bdae),
	.w2(32'hbc849790),
	.w3(32'h3b2b4f9c),
	.w4(32'h3b2281e9),
	.w5(32'hbb0c9e52),
	.w6(32'h3bc6e7cf),
	.w7(32'h3b4a88fb),
	.w8(32'hbbd20591),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4445df),
	.w1(32'h3b99fb18),
	.w2(32'hbbe3d110),
	.w3(32'h3b8084e0),
	.w4(32'hba9232ca),
	.w5(32'h3a88804f),
	.w6(32'hbafb9c5d),
	.w7(32'h3aa8d155),
	.w8(32'h3b1fdf04),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea73f),
	.w1(32'h3b7614d3),
	.w2(32'h3c4f7bbf),
	.w3(32'hb9889368),
	.w4(32'h3b90ef50),
	.w5(32'h3c0f0f8c),
	.w6(32'hbaca731d),
	.w7(32'h3c0f9076),
	.w8(32'h3bb10104),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90eeed),
	.w1(32'hba806dfb),
	.w2(32'h3be45620),
	.w3(32'hbb455ea4),
	.w4(32'h392e2914),
	.w5(32'hba61dfd0),
	.w6(32'hbbd3d724),
	.w7(32'hbbc22f53),
	.w8(32'hbb75e65a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba634e8),
	.w1(32'hbb9f199f),
	.w2(32'hbb45e3bf),
	.w3(32'hbb6d8bfb),
	.w4(32'hbb09e794),
	.w5(32'h3b0e8650),
	.w6(32'hbbd23cdb),
	.w7(32'hbb67e783),
	.w8(32'hbaed83e3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a211a),
	.w1(32'hba072a73),
	.w2(32'hbb184ea4),
	.w3(32'hb9208f1e),
	.w4(32'h3aee1b0c),
	.w5(32'hbba30e06),
	.w6(32'hbb6fe900),
	.w7(32'hbb0cb18d),
	.w8(32'hbbc3ca4b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c93918),
	.w1(32'hbc04c89c),
	.w2(32'hbba721ea),
	.w3(32'hbb634976),
	.w4(32'hb8ad787a),
	.w5(32'hbbaec3f1),
	.w6(32'hbb6b8aa9),
	.w7(32'hbb851d6b),
	.w8(32'hbbb58d63),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfef389),
	.w1(32'hbbb664c1),
	.w2(32'h3a44dc70),
	.w3(32'hbaff7eac),
	.w4(32'h3af718cb),
	.w5(32'hba64b961),
	.w6(32'hbbd6e89f),
	.w7(32'h38cea9d9),
	.w8(32'hbac7e24b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b78fc),
	.w1(32'hbb154be8),
	.w2(32'hbbbb8e82),
	.w3(32'hbad66dc6),
	.w4(32'hbb257cb5),
	.w5(32'hbb424e54),
	.w6(32'hb856086a),
	.w7(32'hbb7d0952),
	.w8(32'hbadf7de6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47cc91),
	.w1(32'hbbb8eb5d),
	.w2(32'hbc1a6e24),
	.w3(32'h3b1d1d28),
	.w4(32'h3b8efb0e),
	.w5(32'h3bac1cc4),
	.w6(32'h3b809ce7),
	.w7(32'h3afbaa0e),
	.w8(32'hb8336f99),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1e071),
	.w1(32'h3aa55237),
	.w2(32'h3b88f45c),
	.w3(32'h3c06e692),
	.w4(32'h3b8b2d6a),
	.w5(32'h3b514a6f),
	.w6(32'h39666f49),
	.w7(32'h3a86603a),
	.w8(32'hbb5e1e73),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39790856),
	.w1(32'hba175697),
	.w2(32'h39171a42),
	.w3(32'hb604aba1),
	.w4(32'hbaff4e03),
	.w5(32'hb77571e2),
	.w6(32'hbb0ce7c2),
	.w7(32'hbb28e348),
	.w8(32'h3a9315fa),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c721eb8),
	.w1(32'h3b819303),
	.w2(32'hbc2dfd6c),
	.w3(32'h3b038c0c),
	.w4(32'h3baca017),
	.w5(32'h3bd68774),
	.w6(32'h3a77d561),
	.w7(32'h3acc8ebc),
	.w8(32'h3b746669),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be66e62),
	.w1(32'h3afd3766),
	.w2(32'hbb5182bf),
	.w3(32'h3bf16244),
	.w4(32'h3b876174),
	.w5(32'h3a93122d),
	.w6(32'h3ba01bbe),
	.w7(32'h3a7f6b4d),
	.w8(32'hbb588556),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b192a),
	.w1(32'hb96c632f),
	.w2(32'hba613a2d),
	.w3(32'h3a8d503a),
	.w4(32'hba63533b),
	.w5(32'hbb089cbd),
	.w6(32'h39e83a17),
	.w7(32'h3b045b0e),
	.w8(32'h3981be33),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f0353),
	.w1(32'h3b04d4ec),
	.w2(32'hbc2e901e),
	.w3(32'h3b572476),
	.w4(32'h3bc51ff9),
	.w5(32'hbbe11d6f),
	.w6(32'h3c30f8b3),
	.w7(32'h3b3ae0f2),
	.w8(32'hbc13ae60),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25795a),
	.w1(32'h3bace59d),
	.w2(32'hba102976),
	.w3(32'hbb0c6f44),
	.w4(32'h3aa9e526),
	.w5(32'h3a95d33c),
	.w6(32'h3b10e9be),
	.w7(32'h3b3276f9),
	.w8(32'h3ade91d1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7614b),
	.w1(32'hb92d8f46),
	.w2(32'h3a33b77a),
	.w3(32'h3ab764f6),
	.w4(32'h3a5367c6),
	.w5(32'hb9c00868),
	.w6(32'h3aa7bc13),
	.w7(32'hb9f36f9e),
	.w8(32'hbb3be844),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109187),
	.w1(32'hbb13f8a7),
	.w2(32'hbb03c97a),
	.w3(32'hbb1733be),
	.w4(32'hbb05c01a),
	.w5(32'hba46a72c),
	.w6(32'hbb695e41),
	.w7(32'hbb746a34),
	.w8(32'hba89103d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d0a23),
	.w1(32'hbaccc15d),
	.w2(32'hba79376f),
	.w3(32'hbb1db284),
	.w4(32'hbb1465c3),
	.w5(32'h3aec02bc),
	.w6(32'hbb15d0b0),
	.w7(32'hbb14ca4c),
	.w8(32'h3a75a765),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4447),
	.w1(32'h3b292197),
	.w2(32'h3b9a8f11),
	.w3(32'hbafba17c),
	.w4(32'h3b226863),
	.w5(32'h3b7eeece),
	.w6(32'hbb0bd4f7),
	.w7(32'h3a421c0b),
	.w8(32'h3b1680b1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde20ca),
	.w1(32'hba1d7e5a),
	.w2(32'hbc39782f),
	.w3(32'h3bd3f802),
	.w4(32'h3a271ef8),
	.w5(32'hbc22a6b3),
	.w6(32'hbb852f0f),
	.w7(32'h3b04aa40),
	.w8(32'hbc45d9e2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65ca86),
	.w1(32'hbb53a909),
	.w2(32'hbc464f2e),
	.w3(32'h3b106559),
	.w4(32'h39bd5aa8),
	.w5(32'hbbc3e56e),
	.w6(32'h3b6fae29),
	.w7(32'h3ad1d47b),
	.w8(32'hbb17ec60),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ec1b),
	.w1(32'hbb3f0cf8),
	.w2(32'hbc3a0113),
	.w3(32'h3a2b487b),
	.w4(32'h3b10367c),
	.w5(32'hbbac5b93),
	.w6(32'h3892407a),
	.w7(32'hbabb256a),
	.w8(32'hbbe3e6f8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac28844),
	.w1(32'hba318571),
	.w2(32'h38eaa01f),
	.w3(32'h3b940cfe),
	.w4(32'h3b3f1cfe),
	.w5(32'h3b4a9c66),
	.w6(32'h3a39e34b),
	.w7(32'h3a17ef5e),
	.w8(32'hb9a49a08),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf4316),
	.w1(32'h3b28e232),
	.w2(32'h3b1c3777),
	.w3(32'h3a4e7f0a),
	.w4(32'hba72689a),
	.w5(32'hbb83fd9c),
	.w6(32'hb7d81a73),
	.w7(32'h3a6b46ac),
	.w8(32'hbb1a6cc5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1973f3),
	.w1(32'hbb27090f),
	.w2(32'hbb625560),
	.w3(32'hbb5ae334),
	.w4(32'hbb3798b4),
	.w5(32'hbb4d3ee4),
	.w6(32'hbb1c59cf),
	.w7(32'hbb313627),
	.w8(32'hbb3fe98d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8044),
	.w1(32'hbb6863c7),
	.w2(32'h3a284ce4),
	.w3(32'hbb109c51),
	.w4(32'hbb6ab308),
	.w5(32'h3b3f1ef1),
	.w6(32'hba71fe33),
	.w7(32'hbab50040),
	.w8(32'h3b3cb447),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43fce2),
	.w1(32'hbbc73229),
	.w2(32'hbc149adc),
	.w3(32'h3baba775),
	.w4(32'h3ab27269),
	.w5(32'hbbe10934),
	.w6(32'h3bb096a4),
	.w7(32'hb93dcbc9),
	.w8(32'hbbd21224),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd92d),
	.w1(32'hbb7ce30a),
	.w2(32'hba5f6bbc),
	.w3(32'hbb00a8a8),
	.w4(32'hbac8e208),
	.w5(32'h39b06b40),
	.w6(32'hbbe45b03),
	.w7(32'hbb5c6030),
	.w8(32'hb9d4a72f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a22b5),
	.w1(32'h3b7e61c8),
	.w2(32'h3bafb1de),
	.w3(32'h39068a20),
	.w4(32'hbaa224db),
	.w5(32'h3a6da7bb),
	.w6(32'h3b12e317),
	.w7(32'h3b1b110d),
	.w8(32'hba365aa1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdc2ac),
	.w1(32'hbac0694a),
	.w2(32'hbb69514d),
	.w3(32'hba5a807d),
	.w4(32'hbb06702e),
	.w5(32'h3a7da87a),
	.w6(32'hbac7ff0c),
	.w7(32'hba1a019a),
	.w8(32'h3b4fc0a5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba03611),
	.w1(32'h3b2a3dc4),
	.w2(32'h3b2213c0),
	.w3(32'h3b018229),
	.w4(32'h3b5913a7),
	.w5(32'hba1f0b75),
	.w6(32'h3c08b2cf),
	.w7(32'h3be15357),
	.w8(32'hbac8d160),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a939131),
	.w1(32'h39aa5ca1),
	.w2(32'hbb9f3e6a),
	.w3(32'hb8f1debf),
	.w4(32'hb9a1af8f),
	.w5(32'hb9cc785e),
	.w6(32'hbb000a86),
	.w7(32'hbad39674),
	.w8(32'hbaa97813),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b003bf5),
	.w1(32'h3addcbf2),
	.w2(32'h393ed5be),
	.w3(32'h39f5439f),
	.w4(32'h3a283610),
	.w5(32'hb89c1591),
	.w6(32'h3ad030a8),
	.w7(32'h3b07847f),
	.w8(32'hbb2df660),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a85c),
	.w1(32'hbc8471c9),
	.w2(32'hbc8bc587),
	.w3(32'h3b9c30e8),
	.w4(32'hbb9edde5),
	.w5(32'hbc4db316),
	.w6(32'hbbd9f1d4),
	.w7(32'hbba1cdcb),
	.w8(32'hbc0ad8b6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae26175),
	.w1(32'hb95160d3),
	.w2(32'hba8d5424),
	.w3(32'hba798c4a),
	.w4(32'hbaf382c9),
	.w5(32'hba5bf0ac),
	.w6(32'h3904a6e1),
	.w7(32'hba8c02dd),
	.w8(32'h39bebf54),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2520),
	.w1(32'h3aeb0348),
	.w2(32'h3b9c3639),
	.w3(32'hbb93f719),
	.w4(32'h3b2c2ed6),
	.w5(32'h3bd18c73),
	.w6(32'hbb465ca6),
	.w7(32'h3b90f8b1),
	.w8(32'h3bdd4f0b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule