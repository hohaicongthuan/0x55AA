module layer_10_featuremap_386(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba644237),
	.w1(32'h3a9d75c4),
	.w2(32'hbac6886f),
	.w3(32'hb9229a1a),
	.w4(32'h3b0667ce),
	.w5(32'hbbf8bb82),
	.w6(32'hbb942500),
	.w7(32'h39b3922d),
	.w8(32'hb8cfe291),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf1208),
	.w1(32'hbac67a41),
	.w2(32'hbb2de161),
	.w3(32'hbb622185),
	.w4(32'hbb87cebb),
	.w5(32'hbb61fdd2),
	.w6(32'h3a4d4b9c),
	.w7(32'hbb3206d1),
	.w8(32'h39d64627),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381155cb),
	.w1(32'hbb125b92),
	.w2(32'hbb61ae94),
	.w3(32'h39bd1d35),
	.w4(32'hbb60714f),
	.w5(32'h3a4854b9),
	.w6(32'h3a561cbd),
	.w7(32'hbb9e38ea),
	.w8(32'hbb4d7d98),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d42d0),
	.w1(32'hbb8c40f5),
	.w2(32'h3a0ab194),
	.w3(32'h394f1b65),
	.w4(32'hb9c381b2),
	.w5(32'hbb492538),
	.w6(32'hbac40d52),
	.w7(32'hba942121),
	.w8(32'h3b02d7b2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d16767),
	.w1(32'h38cb02fc),
	.w2(32'h3a9e7437),
	.w3(32'h3ba85883),
	.w4(32'hb99bd049),
	.w5(32'h3ae2aec6),
	.w6(32'h3bba12e8),
	.w7(32'h3a141965),
	.w8(32'h3a9113a5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce2d0),
	.w1(32'h3b507db2),
	.w2(32'h3b86af58),
	.w3(32'hba594334),
	.w4(32'hb98a1be1),
	.w5(32'h3c16e3d8),
	.w6(32'h3b3df32e),
	.w7(32'hba9b3295),
	.w8(32'h3bc4181a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5648),
	.w1(32'hbb5b503f),
	.w2(32'hbb3d9cfa),
	.w3(32'hb9fc1c56),
	.w4(32'h3a80f3b6),
	.w5(32'hba6944cb),
	.w6(32'hba2b05bf),
	.w7(32'h3a988094),
	.w8(32'h3b0c5128),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b3325),
	.w1(32'h3b8aebcd),
	.w2(32'h3bf615a1),
	.w3(32'h3b699c01),
	.w4(32'h3bcdbdbb),
	.w5(32'h3b5886ec),
	.w6(32'hba950091),
	.w7(32'h3b98bf0d),
	.w8(32'h3b2228f9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8795f7),
	.w1(32'hbaeedad9),
	.w2(32'hbb85a19a),
	.w3(32'h3b4e37e5),
	.w4(32'h3a024ab4),
	.w5(32'hbb9458c1),
	.w6(32'h3bc61dfe),
	.w7(32'hba204679),
	.w8(32'hb8acccd6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad67e),
	.w1(32'h3bcd5648),
	.w2(32'h3b9c57e9),
	.w3(32'hbb3a4b61),
	.w4(32'h3bdb8469),
	.w5(32'hbae728f2),
	.w6(32'h3b5f7f43),
	.w7(32'h3b1bc13b),
	.w8(32'hbac6b1af),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa251e5),
	.w1(32'hba393141),
	.w2(32'hbb5093fc),
	.w3(32'hbb6450c6),
	.w4(32'h394ee6f2),
	.w5(32'hbafdd015),
	.w6(32'h3b0b33be),
	.w7(32'hb9cb061c),
	.w8(32'h3b113acc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9404c64),
	.w1(32'hbb28bd89),
	.w2(32'hbc07492a),
	.w3(32'h3b2fbdc9),
	.w4(32'hbb183785),
	.w5(32'hbbb45517),
	.w6(32'h3a89d7c8),
	.w7(32'hbbd4c25f),
	.w8(32'hbc1ed6c7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3155b),
	.w1(32'hba571c81),
	.w2(32'hbb1d1c1e),
	.w3(32'hbb0aa56d),
	.w4(32'h399dcf01),
	.w5(32'h3bf08a6d),
	.w6(32'hbb5a63e8),
	.w7(32'h39b943fd),
	.w8(32'h3b1987e8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31ad26),
	.w1(32'hbab68098),
	.w2(32'hba04f56f),
	.w3(32'h3b398729),
	.w4(32'hbb1e40f5),
	.w5(32'h3a7f0331),
	.w6(32'hbb829c8e),
	.w7(32'hbbc59b2d),
	.w8(32'h3a594908),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd8af0),
	.w1(32'h3895faf0),
	.w2(32'h3ba83887),
	.w3(32'hba0e27d9),
	.w4(32'hbb0c31f0),
	.w5(32'h3c25d077),
	.w6(32'hba974617),
	.w7(32'hb9f899b0),
	.w8(32'hba6ba6eb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb370cee),
	.w1(32'h3b273d34),
	.w2(32'h3b401323),
	.w3(32'h3a79a117),
	.w4(32'h3b17ba84),
	.w5(32'h3c3d331c),
	.w6(32'h3aa111ad),
	.w7(32'h3b4eb8b2),
	.w8(32'h3b79c5c0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe34c),
	.w1(32'hbb877650),
	.w2(32'h3a63c88e),
	.w3(32'hb9aefd6d),
	.w4(32'hbb7d29ac),
	.w5(32'hbb2d05eb),
	.w6(32'hbaeccb5b),
	.w7(32'hbbb01059),
	.w8(32'hbb2f9576),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b283d),
	.w1(32'h3b169e3b),
	.w2(32'hbbabdb48),
	.w3(32'h3b7171de),
	.w4(32'hbb14d0a3),
	.w5(32'hbbe27718),
	.w6(32'h3ad23570),
	.w7(32'hbb78aebe),
	.w8(32'hbbadf4cf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74992b),
	.w1(32'hbaccf37f),
	.w2(32'hbb2f6900),
	.w3(32'hbb8c492a),
	.w4(32'hbb140ae3),
	.w5(32'h3a5adbf9),
	.w6(32'hbadbbb91),
	.w7(32'h3a55f6bc),
	.w8(32'h3af08c59),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c5760),
	.w1(32'h3c31eafb),
	.w2(32'h3cfefdd3),
	.w3(32'h3b9caee8),
	.w4(32'h3bf9e124),
	.w5(32'h3c1435e6),
	.w6(32'h3b16f3c3),
	.w7(32'h3c08f9e8),
	.w8(32'h3c4e64c2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccf5be),
	.w1(32'h3b8b5c03),
	.w2(32'h3b0abc62),
	.w3(32'h3cca4308),
	.w4(32'h39414421),
	.w5(32'h3b9ff311),
	.w6(32'h3ccba753),
	.w7(32'h3ad26c1c),
	.w8(32'h3a5cbedb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39de6),
	.w1(32'hb979e4f4),
	.w2(32'h38b1b7ef),
	.w3(32'hbad03b0f),
	.w4(32'hba86c629),
	.w5(32'h3b2f810f),
	.w6(32'hbb3d4118),
	.w7(32'h3b201a27),
	.w8(32'h3b63614f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda3a3d),
	.w1(32'hbb0296e7),
	.w2(32'h3b132775),
	.w3(32'h3afa4b0b),
	.w4(32'h39efc327),
	.w5(32'h3ad5aa1f),
	.w6(32'hbbbef578),
	.w7(32'h39ddb765),
	.w8(32'h3ae0195a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7f184),
	.w1(32'h3b6b5816),
	.w2(32'h3aec5608),
	.w3(32'hbad81eea),
	.w4(32'h383723e1),
	.w5(32'hb95c6fbd),
	.w6(32'h38a08f8a),
	.w7(32'h3b243a22),
	.w8(32'h39969895),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8e935),
	.w1(32'hbba2954a),
	.w2(32'h3aeef165),
	.w3(32'hbb328169),
	.w4(32'hbb84cf75),
	.w5(32'hbac756ae),
	.w6(32'hba8dc985),
	.w7(32'hbb5e3b72),
	.w8(32'h38b10f87),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c4348),
	.w1(32'hbba0b822),
	.w2(32'hb985cc3a),
	.w3(32'hbb21e481),
	.w4(32'hbbbf865c),
	.w5(32'hb88235ed),
	.w6(32'hba9827cc),
	.w7(32'hba04651f),
	.w8(32'hbbe292da),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4d3a),
	.w1(32'hbbb3e919),
	.w2(32'hbbe243b1),
	.w3(32'hbbf3fa10),
	.w4(32'hbba1dfff),
	.w5(32'hbab075c0),
	.w6(32'hbbcca011),
	.w7(32'h3a19fe44),
	.w8(32'h3b4632cd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12adda),
	.w1(32'h3b104497),
	.w2(32'h3ab11fc3),
	.w3(32'h3b9f5f57),
	.w4(32'h3b7a9e10),
	.w5(32'h3a85dda9),
	.w6(32'hba89e266),
	.w7(32'h3bbfffda),
	.w8(32'h3acc98a7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c829d),
	.w1(32'h39bd653f),
	.w2(32'h3b277bf0),
	.w3(32'h3b332099),
	.w4(32'h3a87d22c),
	.w5(32'h3a9a05de),
	.w6(32'h3ba5013c),
	.w7(32'h3a9391a7),
	.w8(32'h3b68be47),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80adc9),
	.w1(32'h39440f2c),
	.w2(32'h3a8143fd),
	.w3(32'h3affa754),
	.w4(32'hbace93be),
	.w5(32'hbb1e98e3),
	.w6(32'h3aebf97b),
	.w7(32'hbb0c3a25),
	.w8(32'hbbc68ec8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80206c),
	.w1(32'hbb13bd5e),
	.w2(32'h3a57ff2c),
	.w3(32'hbbe97e46),
	.w4(32'h3a8b7d39),
	.w5(32'hbab16695),
	.w6(32'hbb930669),
	.w7(32'h3b0db0f8),
	.w8(32'hbac4cafd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad913),
	.w1(32'hbab3300a),
	.w2(32'hbb1717b0),
	.w3(32'h3a908199),
	.w4(32'hbafede0e),
	.w5(32'hb9e24b59),
	.w6(32'hb9b84c39),
	.w7(32'hbae436ab),
	.w8(32'hba3093db),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d15b56),
	.w1(32'hbb8b9d10),
	.w2(32'hbb4f4a7f),
	.w3(32'h3b57b164),
	.w4(32'hba6e6ba0),
	.w5(32'hbb928aff),
	.w6(32'h3a1383d1),
	.w7(32'hbbc1a334),
	.w8(32'hb909530a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c3f0),
	.w1(32'hbab2d0a7),
	.w2(32'h3b3541af),
	.w3(32'hbb62df6c),
	.w4(32'hbad03543),
	.w5(32'hbb61f7e6),
	.w6(32'hba4ee57d),
	.w7(32'hb9fdd709),
	.w8(32'h3a3607aa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c42b8),
	.w1(32'h3b7c2ae1),
	.w2(32'h3b754135),
	.w3(32'hba0c6031),
	.w4(32'h3b10c186),
	.w5(32'h3a585775),
	.w6(32'h3b39b4dc),
	.w7(32'h3b2b6c6c),
	.w8(32'h3b392e55),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f3a4),
	.w1(32'hba054a5c),
	.w2(32'hbb50ec7b),
	.w3(32'hbae9762f),
	.w4(32'h3aaf50a0),
	.w5(32'hbb1dea00),
	.w6(32'h3ba43868),
	.w7(32'hbb67134a),
	.w8(32'h3a02ec2b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde8a73),
	.w1(32'hbad40ffa),
	.w2(32'hba5892ea),
	.w3(32'hbbc8e0a9),
	.w4(32'h39af1d1e),
	.w5(32'hba694b45),
	.w6(32'hbbaa3a02),
	.w7(32'hbb1f1f28),
	.w8(32'h3a6500ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabef2bb),
	.w1(32'hbb532794),
	.w2(32'hbaf07601),
	.w3(32'hba9d28f2),
	.w4(32'hbae77679),
	.w5(32'hbb3ff848),
	.w6(32'hbb5cd6af),
	.w7(32'hbbb9a94f),
	.w8(32'hbb3a2f90),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2d72b),
	.w1(32'hbb239654),
	.w2(32'h3983bdad),
	.w3(32'hba6cd04e),
	.w4(32'h3a1c2582),
	.w5(32'hbb78a65e),
	.w6(32'hbbc4030d),
	.w7(32'hbae302c5),
	.w8(32'hb992f4b7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a921122),
	.w1(32'h3a8a5ccb),
	.w2(32'h3b353915),
	.w3(32'hbadfa988),
	.w4(32'h3afd2d05),
	.w5(32'hbab9b98a),
	.w6(32'h3a716987),
	.w7(32'h39fc9ad7),
	.w8(32'h3a587fa9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71ac83),
	.w1(32'hbb921253),
	.w2(32'hba006507),
	.w3(32'h3bf6491b),
	.w4(32'hbb378a40),
	.w5(32'h3b17ada4),
	.w6(32'h3bd209fb),
	.w7(32'hba489a53),
	.w8(32'hbb959fba),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0201cf),
	.w1(32'hbb557597),
	.w2(32'hbb56afb4),
	.w3(32'h3b60a0ba),
	.w4(32'hbb3b91cc),
	.w5(32'h3aa716bc),
	.w6(32'hbb9b4fcf),
	.w7(32'hbaf0f574),
	.w8(32'hbb6931be),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac771ac),
	.w1(32'hbab2ec9b),
	.w2(32'hbbae7699),
	.w3(32'h3b12894f),
	.w4(32'hba747c68),
	.w5(32'hb93c6f8a),
	.w6(32'hbb10f87e),
	.w7(32'hbb6fde6c),
	.w8(32'hba86f2f5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfd480),
	.w1(32'h3bf1ec2e),
	.w2(32'h3c2b3914),
	.w3(32'h3a3d7cf9),
	.w4(32'h3c203e7e),
	.w5(32'hbb6565c0),
	.w6(32'h3b2272f3),
	.w7(32'h3c2c15da),
	.w8(32'h3b2ef319),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c315f94),
	.w1(32'h3889f395),
	.w2(32'h3b63c868),
	.w3(32'h3c4da3d1),
	.w4(32'hba9cf9f2),
	.w5(32'h3bbfba91),
	.w6(32'h3c533eab),
	.w7(32'hba305de2),
	.w8(32'h3ae308b7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9cbc7),
	.w1(32'h3b9d82a8),
	.w2(32'h3bd974ed),
	.w3(32'h3a81841e),
	.w4(32'h3a90f413),
	.w5(32'h3c619330),
	.w6(32'hba02d953),
	.w7(32'h3b10bf66),
	.w8(32'h3bbf333d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c15b6),
	.w1(32'h3b7771a0),
	.w2(32'hbb8cb71a),
	.w3(32'h3b0c5006),
	.w4(32'h3a0e2925),
	.w5(32'h3a3ed189),
	.w6(32'h3b9bb763),
	.w7(32'h3b14d1f5),
	.w8(32'hbad71e8b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696257),
	.w1(32'hba506b0b),
	.w2(32'h3b56cb50),
	.w3(32'h3bb528a4),
	.w4(32'hb9964c8c),
	.w5(32'h3a28320f),
	.w6(32'hbab5d01d),
	.w7(32'h3b28ed01),
	.w8(32'h3b1d3501),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61b063),
	.w1(32'h3b44dfb3),
	.w2(32'h3b41e0ad),
	.w3(32'hba52cb6b),
	.w4(32'h3b7512fd),
	.w5(32'hbb11bae9),
	.w6(32'h3a6e8d5d),
	.w7(32'h3afcea98),
	.w8(32'hb92af94c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2770d7),
	.w1(32'h3acc6d59),
	.w2(32'h38e7ab04),
	.w3(32'hbbe8925d),
	.w4(32'h3ae1c3b8),
	.w5(32'h3af6015a),
	.w6(32'hbbbb38f9),
	.w7(32'hba46e450),
	.w8(32'hba96c488),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae43311),
	.w1(32'hbb7089fa),
	.w2(32'hbb6e9b78),
	.w3(32'hbb4a9145),
	.w4(32'hbbe1425e),
	.w5(32'h3ae5ff24),
	.w6(32'hbb2cf7b9),
	.w7(32'hbadf2e89),
	.w8(32'h3a922885),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01c1d2),
	.w1(32'hbacc9e24),
	.w2(32'h3a9fe1f7),
	.w3(32'h3a8928aa),
	.w4(32'hbaf7681b),
	.w5(32'h3b10f7dc),
	.w6(32'hba895fdc),
	.w7(32'h3bb342b4),
	.w8(32'h3c0d71b2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd4cd),
	.w1(32'h3bda6bf4),
	.w2(32'h39eafaf4),
	.w3(32'h3af1a590),
	.w4(32'h3b540912),
	.w5(32'hb8ea75b9),
	.w6(32'h3a98a845),
	.w7(32'h3a1209e3),
	.w8(32'h3afbf3a7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac69c22),
	.w1(32'h3bdfbc3a),
	.w2(32'hba78cfed),
	.w3(32'hba08b7ed),
	.w4(32'h3be1f4fc),
	.w5(32'hbac97930),
	.w6(32'h3b1527b4),
	.w7(32'h3ac1ecef),
	.w8(32'h3af04581),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be037),
	.w1(32'h3b6115b7),
	.w2(32'h3bc8534f),
	.w3(32'h395d1db6),
	.w4(32'h3b9605f2),
	.w5(32'h3b1f2990),
	.w6(32'h3b481e6c),
	.w7(32'h3b23abf3),
	.w8(32'h3b4b78b7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f388),
	.w1(32'hb972f8ca),
	.w2(32'hba51b867),
	.w3(32'h3c3eacce),
	.w4(32'h3b1f95cc),
	.w5(32'hb9838bf9),
	.w6(32'h3c08d42d),
	.w7(32'hba812a04),
	.w8(32'hb9aa9ddd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e10e7),
	.w1(32'hbb46e36f),
	.w2(32'hbb85ce14),
	.w3(32'hbb837c4a),
	.w4(32'hbb2e236b),
	.w5(32'hba969f8e),
	.w6(32'hbb39c67e),
	.w7(32'hbb07ff1a),
	.w8(32'hbb3bda32),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c6e1),
	.w1(32'hba8aa3d5),
	.w2(32'h3be6eecb),
	.w3(32'hbb35e22e),
	.w4(32'hbbf586e9),
	.w5(32'h3c6b2156),
	.w6(32'hbb3abeee),
	.w7(32'hbba7af2b),
	.w8(32'hb93d999b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1413e4),
	.w1(32'h3ac1353e),
	.w2(32'hbb7eb0b1),
	.w3(32'hbbd93315),
	.w4(32'h398423a1),
	.w5(32'hbaa4046b),
	.w6(32'hbb9eadb4),
	.w7(32'hbabd1a35),
	.w8(32'h3ad76bc8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cd306),
	.w1(32'h3ad228d4),
	.w2(32'hbaa4f80d),
	.w3(32'hb74f798c),
	.w4(32'h3b00602b),
	.w5(32'h3a2065fd),
	.w6(32'hbb6360d4),
	.w7(32'h3ab27c22),
	.w8(32'hba7c7757),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68e429),
	.w1(32'hbba3f6d3),
	.w2(32'h3b656830),
	.w3(32'hba8a4ab6),
	.w4(32'h3a64426c),
	.w5(32'h3c0df3d7),
	.w6(32'h39f251a5),
	.w7(32'hb974e2d1),
	.w8(32'hbb4d8932),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13894a),
	.w1(32'h3b06b973),
	.w2(32'h3ab88030),
	.w3(32'hbb141bbc),
	.w4(32'h3afe5b96),
	.w5(32'hbaa27da6),
	.w6(32'hbae1be39),
	.w7(32'h3af814f8),
	.w8(32'h3b4c9de4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97279e),
	.w1(32'h3b3ac73e),
	.w2(32'hbb85fef5),
	.w3(32'h3c083acd),
	.w4(32'h3ad540da),
	.w5(32'hbb29f0c9),
	.w6(32'h3b8f1f68),
	.w7(32'h3ad2bd33),
	.w8(32'hbabf3df7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb6dfa),
	.w1(32'hb98dfb5b),
	.w2(32'hbabc0ce3),
	.w3(32'hbb61458c),
	.w4(32'h39d59721),
	.w5(32'h3b875939),
	.w6(32'hbb3ee5f6),
	.w7(32'h3b0e4d42),
	.w8(32'h3a32c2b0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fe433),
	.w1(32'h3a6ba652),
	.w2(32'h3aa80efd),
	.w3(32'h3adc1d4d),
	.w4(32'h3b7d305b),
	.w5(32'h38c73e38),
	.w6(32'hb99fbf56),
	.w7(32'h3b28b354),
	.w8(32'h3ae5b31a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f7b0b1),
	.w1(32'h3ab02c4c),
	.w2(32'hbb99ae06),
	.w3(32'h3b55c238),
	.w4(32'hba693ad4),
	.w5(32'hbb3b50c9),
	.w6(32'h3b3c0afb),
	.w7(32'hbaec93b4),
	.w8(32'hba99f99e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc2a84),
	.w1(32'hbb5582c4),
	.w2(32'hbaf305db),
	.w3(32'hba964d9a),
	.w4(32'hbb7d11f2),
	.w5(32'hbbe166dd),
	.w6(32'h3a8bedb6),
	.w7(32'h39b9e100),
	.w8(32'h3a802334),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed0a3),
	.w1(32'h3b2d8e8a),
	.w2(32'h3b9e4e63),
	.w3(32'hbb462ee9),
	.w4(32'h3adb0989),
	.w5(32'h3b007485),
	.w6(32'hbb3fb792),
	.w7(32'h3b88aa7f),
	.w8(32'hba0c914b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2941),
	.w1(32'h3bfa0171),
	.w2(32'h3a890ab5),
	.w3(32'hbbff86c3),
	.w4(32'h3c172488),
	.w5(32'hbb1c887c),
	.w6(32'hbbb13114),
	.w7(32'h3bbee51b),
	.w8(32'h3b6e5277),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a781b4f),
	.w1(32'h39da2066),
	.w2(32'h3a436b17),
	.w3(32'h3a89c892),
	.w4(32'hb98e3642),
	.w5(32'h38fecfd8),
	.w6(32'h3b384df2),
	.w7(32'hb8d5da18),
	.w8(32'hba6a0596),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a969d),
	.w1(32'hb69bb684),
	.w2(32'h36d2c8a4),
	.w3(32'hb587b86e),
	.w4(32'h3678a083),
	.w5(32'h372ee5e4),
	.w6(32'h37d74aae),
	.w7(32'h37d0ec5b),
	.w8(32'h3815fdd9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b9b809),
	.w1(32'hb7441318),
	.w2(32'h378260da),
	.w3(32'hb61b4abe),
	.w4(32'h37012b21),
	.w5(32'h3800c746),
	.w6(32'h3803b7c2),
	.w7(32'h381a9e66),
	.w8(32'h38690231),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84dbc06),
	.w1(32'hb8177dbc),
	.w2(32'hb7bd9184),
	.w3(32'hb73aa864),
	.w4(32'hb725e40a),
	.w5(32'hb69d5f15),
	.w6(32'h37a190e1),
	.w7(32'h378d2cd2),
	.w8(32'h381818e5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f85c26),
	.w1(32'h3981cd2f),
	.w2(32'hb968b524),
	.w3(32'h3919dc6b),
	.w4(32'h38e0267a),
	.w5(32'hb901e716),
	.w6(32'hb8580577),
	.w7(32'h3950d6c2),
	.w8(32'hb7f36b86),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78b1b16),
	.w1(32'hb6b13e01),
	.w2(32'h37108dde),
	.w3(32'hb76b7546),
	.w4(32'h36820a66),
	.w5(32'hb6d4513c),
	.w6(32'h37321b78),
	.w7(32'h37c95fad),
	.w8(32'h37162864),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b069fd),
	.w1(32'h39fadd9d),
	.w2(32'h39c6a9de),
	.w3(32'hb97859cb),
	.w4(32'h39f6cf8f),
	.w5(32'hb6f80c16),
	.w6(32'hb81b4b82),
	.w7(32'hb9238e0c),
	.w8(32'hb8b748f4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba770567),
	.w1(32'h3a79e9cc),
	.w2(32'h3ac28add),
	.w3(32'hb8c14994),
	.w4(32'h3a7dbe6b),
	.w5(32'h39c3a599),
	.w6(32'hba914043),
	.w7(32'h39f3dd2a),
	.w8(32'h3985e77a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c5020),
	.w1(32'hb8b98eac),
	.w2(32'h398c4de9),
	.w3(32'h391d937a),
	.w4(32'hb926a723),
	.w5(32'h394e9da3),
	.w6(32'h380d6de1),
	.w7(32'hb9aa7eed),
	.w8(32'hb9a5a322),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397092e0),
	.w1(32'h3a0de60a),
	.w2(32'h39dc710e),
	.w3(32'h3933a1b0),
	.w4(32'h39ac8357),
	.w5(32'h394b7dba),
	.w6(32'hb8c01b28),
	.w7(32'h38c1ac5b),
	.w8(32'h38ac7f06),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba277abe),
	.w1(32'h3a6597a8),
	.w2(32'h3a200907),
	.w3(32'hb9bcaaa1),
	.w4(32'h39aeeb06),
	.w5(32'hba41e18f),
	.w6(32'hb9beb679),
	.w7(32'h3987135c),
	.w8(32'hb9da34df),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c48b3),
	.w1(32'h382e3cf6),
	.w2(32'h3861ab79),
	.w3(32'h3a7a2cb3),
	.w4(32'h39b73d33),
	.w5(32'h399c9e68),
	.w6(32'h3a2f23e4),
	.w7(32'h3a052cf0),
	.w8(32'h37d6ab32),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e1b21),
	.w1(32'h3981f1d6),
	.w2(32'hb99c4ef4),
	.w3(32'h3891228e),
	.w4(32'h3810e922),
	.w5(32'hb98ad58c),
	.w6(32'hb9915a70),
	.w7(32'hb981236a),
	.w8(32'hb98f89d7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aa4490),
	.w1(32'h367b6bb2),
	.w2(32'h3741c37f),
	.w3(32'hb718a590),
	.w4(32'h3623871d),
	.w5(32'h3717cc0d),
	.w6(32'h368ea734),
	.w7(32'h379ab3b5),
	.w8(32'h3754decf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3650cb01),
	.w1(32'hb6e83a0c),
	.w2(32'hb5dda898),
	.w3(32'h3667e163),
	.w4(32'h351e823e),
	.w5(32'h35bbc81a),
	.w6(32'h369a2ffc),
	.w7(32'h3727f673),
	.w8(32'h3731e444),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628809f),
	.w1(32'hb5bb6c4f),
	.w2(32'h361683ce),
	.w3(32'hb5d29c8f),
	.w4(32'h35b7821b),
	.w5(32'h36b09cad),
	.w6(32'h365374a7),
	.w7(32'h36907071),
	.w8(32'h3715d502),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d62f62),
	.w1(32'hb9322cc9),
	.w2(32'hb9096b75),
	.w3(32'hb800babb),
	.w4(32'hb7872420),
	.w5(32'hb81858b9),
	.w6(32'hb6a16c6a),
	.w7(32'h36d68a38),
	.w8(32'h376e1e80),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a6560),
	.w1(32'hb976136e),
	.w2(32'h39c47b1c),
	.w3(32'h3962391b),
	.w4(32'hb918e125),
	.w5(32'h39f7dcea),
	.w6(32'h39106a2c),
	.w7(32'hb9280e7c),
	.w8(32'hb79f34d0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a86191),
	.w1(32'hb775585c),
	.w2(32'h38126106),
	.w3(32'hb8b5ba5d),
	.w4(32'hb7d53189),
	.w5(32'h36c2e596),
	.w6(32'hb8739672),
	.w7(32'hb88e4501),
	.w8(32'hb7b1f025),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a48311),
	.w1(32'h3942dc47),
	.w2(32'h394bf192),
	.w3(32'hb8aea250),
	.w4(32'h3877d567),
	.w5(32'h39627ba7),
	.w6(32'hb9db2e65),
	.w7(32'hb97b491c),
	.w8(32'hb9062081),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f3084),
	.w1(32'h3a4ebf99),
	.w2(32'h39bce712),
	.w3(32'h396d11e5),
	.w4(32'h39de9090),
	.w5(32'h370f503d),
	.w6(32'hb9f6eac0),
	.w7(32'h39822b9e),
	.w8(32'h389d7e48),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24ef2c),
	.w1(32'hba0a1930),
	.w2(32'hb8d5f7e1),
	.w3(32'hb8ed8614),
	.w4(32'hba182792),
	.w5(32'h3725fa3a),
	.w6(32'hb715d1a9),
	.w7(32'hba0e0d0b),
	.w8(32'hba3bb84d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29a82d),
	.w1(32'h3ac0990f),
	.w2(32'h3a39e574),
	.w3(32'hb893a5aa),
	.w4(32'h3a848f5c),
	.w5(32'hba1c08db),
	.w6(32'hb95a380f),
	.w7(32'hb8b6c401),
	.w8(32'hba378c6b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f7075),
	.w1(32'hba09ff59),
	.w2(32'hba334cae),
	.w3(32'h3866c40f),
	.w4(32'hb9e81793),
	.w5(32'hba5e511c),
	.w6(32'hba142b49),
	.w7(32'hbab4c39f),
	.w8(32'hbadcf052),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a705376),
	.w1(32'h3b192f2d),
	.w2(32'h3b19565f),
	.w3(32'h3a5b779a),
	.w4(32'h3a934c6c),
	.w5(32'h3a5372c1),
	.w6(32'h3a1c0033),
	.w7(32'h3ad0c68f),
	.w8(32'h3abd609a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994e6d8),
	.w1(32'h3a8886ef),
	.w2(32'h3ac97695),
	.w3(32'h39230cfa),
	.w4(32'h36910405),
	.w5(32'h3886ff41),
	.w6(32'h3a12b545),
	.w7(32'h3a2cfa8b),
	.w8(32'h3a40879f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dee753),
	.w1(32'hb9a438ff),
	.w2(32'h39267465),
	.w3(32'hb6be620e),
	.w4(32'hb97083d7),
	.w5(32'hb92a07d4),
	.w6(32'h3a02797e),
	.w7(32'h3a010df9),
	.w8(32'h38042f18),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5bd43),
	.w1(32'h39a5cdcf),
	.w2(32'hb78e1df0),
	.w3(32'hb9375f9e),
	.w4(32'hb9abe630),
	.w5(32'hb8ec10db),
	.w6(32'hb927914f),
	.w7(32'hb9a28b93),
	.w8(32'hba14157f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae98e),
	.w1(32'h3b1efb08),
	.w2(32'h3ac5ef15),
	.w3(32'hb8473f5e),
	.w4(32'h3a6a3f53),
	.w5(32'h3a34892e),
	.w6(32'h39622b33),
	.w7(32'h3a986476),
	.w8(32'h3a500314),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399684b1),
	.w1(32'h3aa02e90),
	.w2(32'h396606d7),
	.w3(32'h39dc6cd0),
	.w4(32'h391d4fe7),
	.w5(32'hbaab2568),
	.w6(32'hb9926f12),
	.w7(32'hba94fffd),
	.w8(32'hbb085ee1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb060784),
	.w1(32'h3b2cb2d8),
	.w2(32'h3b920067),
	.w3(32'hb97b0552),
	.w4(32'h3b3fa7da),
	.w5(32'h3b6af7d0),
	.w6(32'hbaf1249b),
	.w7(32'h39140a4b),
	.w8(32'h3ad21f0a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f302f),
	.w1(32'h3ac7cd7c),
	.w2(32'h3a8b6b07),
	.w3(32'h3aa32469),
	.w4(32'h3aabf20d),
	.w5(32'h3aa820b8),
	.w6(32'h3a90e244),
	.w7(32'h3a724a70),
	.w8(32'h38d84ad8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53b452),
	.w1(32'h3a879bcb),
	.w2(32'h3ad23b87),
	.w3(32'hb800dda9),
	.w4(32'h39e12ded),
	.w5(32'h3aa2674f),
	.w6(32'h39d0d634),
	.w7(32'h3a401af6),
	.w8(32'h3a51a94b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad68eff),
	.w1(32'h3ab139f4),
	.w2(32'h3a40e688),
	.w3(32'hb9a3116a),
	.w4(32'h3a09907c),
	.w5(32'hba9f1807),
	.w6(32'hbadea5ca),
	.w7(32'hbaafe68b),
	.w8(32'hbab0e897),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd09eb),
	.w1(32'hb95ff687),
	.w2(32'hba4fd72f),
	.w3(32'hb9d52451),
	.w4(32'hba21a890),
	.w5(32'hba8d1d82),
	.w6(32'hb9625f5f),
	.w7(32'hba5f7f97),
	.w8(32'hbaa75752),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7293d),
	.w1(32'h3b83b98a),
	.w2(32'h3b86aef0),
	.w3(32'hb9fbd271),
	.w4(32'h3b0818d1),
	.w5(32'h3b0e6d19),
	.w6(32'hba9986a9),
	.w7(32'hb8e3878b),
	.w8(32'h3ae23a0a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ee1ec),
	.w1(32'h3938978e),
	.w2(32'hba6b11a5),
	.w3(32'h3a11bb02),
	.w4(32'hb99240e7),
	.w5(32'hba0ceaf6),
	.w6(32'h39bc015a),
	.w7(32'hba4ea3a2),
	.w8(32'hba9cc07f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eca304),
	.w1(32'hb88193d5),
	.w2(32'hb908cb92),
	.w3(32'h37e62ddb),
	.w4(32'hb851c612),
	.w5(32'hb90b2cfe),
	.w6(32'hb912ed48),
	.w7(32'hb95bfc15),
	.w8(32'hb960275b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929f18a),
	.w1(32'h38d42d55),
	.w2(32'h3a5a6230),
	.w3(32'h3a214633),
	.w4(32'h3a0b4080),
	.w5(32'h3a12b4a0),
	.w6(32'h3952ad25),
	.w7(32'h3862c32e),
	.w8(32'h39fd33f3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54c131),
	.w1(32'h39c821c0),
	.w2(32'h38f6e508),
	.w3(32'hb945bd25),
	.w4(32'h3995e59c),
	.w5(32'h39120293),
	.w6(32'hb836f544),
	.w7(32'h3a15a051),
	.w8(32'h3a2ac1c2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fed9d),
	.w1(32'h3a42ca0a),
	.w2(32'h3acc5b22),
	.w3(32'hb8f58449),
	.w4(32'h3a25f93d),
	.w5(32'h3a8fccef),
	.w6(32'h3a0d7938),
	.w7(32'h3a97aa45),
	.w8(32'h3a967511),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ab732),
	.w1(32'hb9b46db9),
	.w2(32'hb9d8e725),
	.w3(32'h39cd947b),
	.w4(32'hb940d59c),
	.w5(32'hb9d13648),
	.w6(32'h39abca98),
	.w7(32'h392f20aa),
	.w8(32'hba48bd35),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c34a2b),
	.w1(32'h3998c12b),
	.w2(32'h395b9090),
	.w3(32'h39781cbb),
	.w4(32'h3846cb2e),
	.w5(32'h395f3a83),
	.w6(32'h3990ac7a),
	.w7(32'h39a59d6a),
	.w8(32'h38894165),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72e766),
	.w1(32'hba1d2544),
	.w2(32'hb62a9ad8),
	.w3(32'hba3489ee),
	.w4(32'hba4336d5),
	.w5(32'hb804f475),
	.w6(32'hbaa17b0a),
	.w7(32'hbaa4b395),
	.w8(32'hba4eddaa),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b070a85),
	.w1(32'h3afbe34c),
	.w2(32'h3b2a31cd),
	.w3(32'h3a655781),
	.w4(32'h3a52b32c),
	.w5(32'h3aa0a6ad),
	.w6(32'h3a031fb4),
	.w7(32'h39d9fbe8),
	.w8(32'h3a6eb81c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7d2e8),
	.w1(32'h399006fb),
	.w2(32'h3970f074),
	.w3(32'h39a3ae9a),
	.w4(32'h38a972b5),
	.w5(32'h3911e98e),
	.w6(32'h3948f06c),
	.w7(32'hb715987c),
	.w8(32'hb865426f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38816ac9),
	.w1(32'h37a968d8),
	.w2(32'h36bd5d66),
	.w3(32'h388c06e4),
	.w4(32'hb747a943),
	.w5(32'h37928d7e),
	.w6(32'h38db8e47),
	.w7(32'h3818e980),
	.w8(32'h385d2dac),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39426864),
	.w1(32'h398912e5),
	.w2(32'h39bc920d),
	.w3(32'h38b95b59),
	.w4(32'h394882f5),
	.w5(32'h3996b0f7),
	.w6(32'hb8f83cc4),
	.w7(32'h38e24427),
	.w8(32'h3721aea1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb581cacf),
	.w1(32'hb5a7637b),
	.w2(32'hb63f1d21),
	.w3(32'hb6a1a38d),
	.w4(32'hb5af8c7e),
	.w5(32'hb42d7c0f),
	.w6(32'h3702e2c4),
	.w7(32'h3730421f),
	.w8(32'h3722a73a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916400a),
	.w1(32'hb8a23a58),
	.w2(32'hb8ccba3c),
	.w3(32'hb86a8452),
	.w4(32'hb82db847),
	.w5(32'hb888694d),
	.w6(32'hb8fb7d37),
	.w7(32'hb8ead12d),
	.w8(32'hb91ba58a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8cc66),
	.w1(32'h38e30638),
	.w2(32'hb967fa65),
	.w3(32'h394fd189),
	.w4(32'hb9593f83),
	.w5(32'hb9fae99e),
	.w6(32'h3796ac22),
	.w7(32'hb9b66b22),
	.w8(32'hba60a8ad),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ec207),
	.w1(32'h38168b29),
	.w2(32'hb9ed2f6f),
	.w3(32'h39513eac),
	.w4(32'h38d165dc),
	.w5(32'hb9bf41a9),
	.w6(32'h39a781e6),
	.w7(32'h393fb49b),
	.w8(32'hb9d29aab),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f350c),
	.w1(32'h3a22c0ee),
	.w2(32'h3849a259),
	.w3(32'hb9054383),
	.w4(32'h39f1739d),
	.w5(32'hb8623f6b),
	.w6(32'hb8ddc009),
	.w7(32'h398cf7f2),
	.w8(32'h38e168c8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1331a6),
	.w1(32'hba034d72),
	.w2(32'h38be20d4),
	.w3(32'hba054cc0),
	.w4(32'hba06ec88),
	.w5(32'h38ca0b79),
	.w6(32'hb9d6a78e),
	.w7(32'hb9bceedd),
	.w8(32'hb978c323),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71830be),
	.w1(32'hb741bb94),
	.w2(32'hb4a58978),
	.w3(32'hb56f2485),
	.w4(32'hb64087e5),
	.w5(32'h3738a6db),
	.w6(32'h372b5ba0),
	.w7(32'h3707f5ed),
	.w8(32'h379ddb9e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389645db),
	.w1(32'h38df3a11),
	.w2(32'h3865f970),
	.w3(32'h38970f38),
	.w4(32'h38e16477),
	.w5(32'h387e1d1e),
	.w6(32'h386ebd7b),
	.w7(32'h38a938e4),
	.w8(32'h37449184),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8103f8b),
	.w1(32'h369733f2),
	.w2(32'h35f6d33c),
	.w3(32'hb707a86f),
	.w4(32'h37608fef),
	.w5(32'hb655a7cd),
	.w6(32'hb798e88e),
	.w7(32'h36e66beb),
	.w8(32'h3607ccc1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd45d5),
	.w1(32'h394dfabd),
	.w2(32'h397244ea),
	.w3(32'h384228ed),
	.w4(32'h38a01c0c),
	.w5(32'h390f94e3),
	.w6(32'hb86ae619),
	.w7(32'hb878750f),
	.w8(32'h36bf04f3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64210a),
	.w1(32'h3a4820fc),
	.w2(32'h3b08980f),
	.w3(32'hba315050),
	.w4(32'h3a6295df),
	.w5(32'h3a96c935),
	.w6(32'hbaa5da10),
	.w7(32'hba0e13c4),
	.w8(32'h39a3f834),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d09f9b),
	.w1(32'h3a595c06),
	.w2(32'h36c481c2),
	.w3(32'h3973b32b),
	.w4(32'h39602519),
	.w5(32'hb9b97344),
	.w6(32'hb9dcc4a1),
	.w7(32'hb8683ec2),
	.w8(32'hb9b8e142),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e4b29d),
	.w1(32'h38e2350c),
	.w2(32'h3716647f),
	.w3(32'h386c4539),
	.w4(32'h380d5243),
	.w5(32'h37d0faa0),
	.w6(32'h37fe3198),
	.w7(32'hb7b58d2b),
	.w8(32'hb7645e55),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbdd55),
	.w1(32'h39f6ee94),
	.w2(32'h3a1c1dd4),
	.w3(32'h39af7cbf),
	.w4(32'h3a099609),
	.w5(32'h39d580b2),
	.w6(32'hb8f6a640),
	.w7(32'h396d54bb),
	.w8(32'hb80ff1e9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3740d29d),
	.w1(32'hb8232293),
	.w2(32'h38837a40),
	.w3(32'h38af9fdd),
	.w4(32'h380f4bb7),
	.w5(32'hb75d2948),
	.w6(32'h38eda080),
	.w7(32'h3834e3f6),
	.w8(32'hb8ca4c5d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38795067),
	.w1(32'h39b27b80),
	.w2(32'h398680cc),
	.w3(32'h379a5c31),
	.w4(32'h3984ae75),
	.w5(32'h3972c900),
	.w6(32'hb79ec88e),
	.w7(32'h39a1ade9),
	.w8(32'h398fbadb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de0fe),
	.w1(32'h3a22fc33),
	.w2(32'h3aac2ef3),
	.w3(32'h3a1b0edf),
	.w4(32'h3a124d4d),
	.w5(32'h3a339112),
	.w6(32'hb682322a),
	.w7(32'h39cb0bcf),
	.w8(32'h39a07afb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6ab44),
	.w1(32'h3ab7753f),
	.w2(32'h380489a6),
	.w3(32'h3953bd4d),
	.w4(32'h39b362a7),
	.w5(32'hb9f38b5a),
	.w6(32'hb99c42fa),
	.w7(32'h39b0d1e4),
	.w8(32'h37fc0ec2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8efe206),
	.w1(32'hb7c9ca5e),
	.w2(32'h39a7dbd0),
	.w3(32'hb8f2ce98),
	.w4(32'hb8fd1da6),
	.w5(32'h38de2538),
	.w6(32'hb86d73cd),
	.w7(32'hb7692cda),
	.w8(32'hb84c3988),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc59d8),
	.w1(32'h3a910a42),
	.w2(32'h3a3d1c37),
	.w3(32'h3905022b),
	.w4(32'h3941ca58),
	.w5(32'h39271dd4),
	.w6(32'hb9969431),
	.w7(32'hb9c41f1d),
	.w8(32'h393d4f2b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39824269),
	.w1(32'h3a657261),
	.w2(32'h38bafcef),
	.w3(32'h39019a60),
	.w4(32'h38dda691),
	.w5(32'hb9f7faab),
	.w6(32'hb9edf6e0),
	.w7(32'hb961b000),
	.w8(32'hb880f6a8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d1b15b),
	.w1(32'h3786f205),
	.w2(32'h3a0c5032),
	.w3(32'hb79cda7b),
	.w4(32'hb9486d8f),
	.w5(32'h3a0bd713),
	.w6(32'hb88c6988),
	.w7(32'hb80dd818),
	.w8(32'h38c26d47),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e40e3),
	.w1(32'h3a66120c),
	.w2(32'h39794db3),
	.w3(32'h39e02ae4),
	.w4(32'h3a10163d),
	.w5(32'h38a5ab38),
	.w6(32'h39d8e57c),
	.w7(32'h3a0d4059),
	.w8(32'h393d5d50),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968287d),
	.w1(32'h3914576e),
	.w2(32'h3861e629),
	.w3(32'h38ec06f0),
	.w4(32'h38920f1d),
	.w5(32'hb780f082),
	.w6(32'h38b614e6),
	.w7(32'h37c88257),
	.w8(32'hb8dede3c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab71dd0),
	.w1(32'hba0c7068),
	.w2(32'h39daa0c2),
	.w3(32'hbaa99dce),
	.w4(32'hba0da105),
	.w5(32'h399515c2),
	.w6(32'h398d3b08),
	.w7(32'h3a55e9f0),
	.w8(32'h3a86b300),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7449194),
	.w1(32'h39478eea),
	.w2(32'hb7f143aa),
	.w3(32'h38c9e6cd),
	.w4(32'h389fac40),
	.w5(32'hb7cf81d3),
	.w6(32'hb88dc5be),
	.w7(32'h3986b219),
	.w8(32'h37b94608),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb607471c),
	.w1(32'h3795b344),
	.w2(32'h3718e4f0),
	.w3(32'h3761ef27),
	.w4(32'h37c0724b),
	.w5(32'h370eed45),
	.w6(32'hb78e4d3d),
	.w7(32'h372c8256),
	.w8(32'h36d52833),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37939f5f),
	.w1(32'h3816bda7),
	.w2(32'h37adf183),
	.w3(32'hb52ebf36),
	.w4(32'h37fddf92),
	.w5(32'h380442dc),
	.w6(32'h36eef956),
	.w7(32'h37759518),
	.w8(32'h3794e36c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987fa26),
	.w1(32'h38895239),
	.w2(32'h38ccda37),
	.w3(32'h388d5852),
	.w4(32'h37eae48c),
	.w5(32'hb8a31713),
	.w6(32'h3964a342),
	.w7(32'h397eae22),
	.w8(32'h3862835f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba069302),
	.w1(32'hb98f6617),
	.w2(32'h38c8d8dd),
	.w3(32'hb85e0a8a),
	.w4(32'hb809de8d),
	.w5(32'hb828e67f),
	.w6(32'hb85e3d9f),
	.w7(32'h39abc0c9),
	.w8(32'h397808cc),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39382467),
	.w1(32'h39d5ff7a),
	.w2(32'h385975f7),
	.w3(32'h3983dc28),
	.w4(32'h39ae4ccc),
	.w5(32'h38c77082),
	.w6(32'h395353c1),
	.w7(32'h39deaa06),
	.w8(32'h393b4f5f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e0fe74),
	.w1(32'hb663f55d),
	.w2(32'hb7073e9a),
	.w3(32'hb618afdd),
	.w4(32'h3611d06d),
	.w5(32'h35d8b41f),
	.w6(32'h367be393),
	.w7(32'h371f5184),
	.w8(32'h36db486d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6e1af),
	.w1(32'h3a589fe3),
	.w2(32'h38ebad45),
	.w3(32'h3a19a5c8),
	.w4(32'h3a1c1f25),
	.w5(32'hb9374e89),
	.w6(32'h3a07aefa),
	.w7(32'h3a3cb5d3),
	.w8(32'h38df3fea),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec5799),
	.w1(32'h39d43ac1),
	.w2(32'h3a3de2ca),
	.w3(32'hb9b90792),
	.w4(32'h38558e50),
	.w5(32'h39f3bb2d),
	.w6(32'hb8a1d753),
	.w7(32'h39aa90ff),
	.w8(32'h3a36ad07),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd98d),
	.w1(32'h3a98c45d),
	.w2(32'h3a4c8486),
	.w3(32'h3890ff77),
	.w4(32'h3a830930),
	.w5(32'h394e330a),
	.w6(32'hba197060),
	.w7(32'h39e74d7b),
	.w8(32'h37f84d3d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90caf3a),
	.w1(32'hba816c41),
	.w2(32'hba7ab2eb),
	.w3(32'h3afb4921),
	.w4(32'h391094b6),
	.w5(32'hb84b3205),
	.w6(32'h3a050a23),
	.w7(32'h3a05686e),
	.w8(32'hba966e92),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a1048),
	.w1(32'hb9522d2e),
	.w2(32'h3a38fc2e),
	.w3(32'hb9c6f996),
	.w4(32'hb980a341),
	.w5(32'h39f18b11),
	.w6(32'hba10cd75),
	.w7(32'hb9b8fbda),
	.w8(32'h39819c70),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a8f0b),
	.w1(32'hb998e53a),
	.w2(32'hb976d266),
	.w3(32'hba23cb6a),
	.w4(32'hba56e741),
	.w5(32'hba6e609d),
	.w6(32'hba7a8221),
	.w7(32'hbab8c1ba),
	.w8(32'hbac3a0a0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808313),
	.w1(32'h3a7c6dbb),
	.w2(32'h399ffd3c),
	.w3(32'h3a9d53f4),
	.w4(32'h3a51f5ab),
	.w5(32'h39b9d6dc),
	.w6(32'h3ac66800),
	.w7(32'h3aa691eb),
	.w8(32'h3a839acc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98593a6),
	.w1(32'hb81d51a0),
	.w2(32'h38635f61),
	.w3(32'h391037c6),
	.w4(32'h37834393),
	.w5(32'hb6a9d6ab),
	.w6(32'h39060606),
	.w7(32'hb7c3bc43),
	.w8(32'hb9cd7706),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf699),
	.w1(32'hb9f299d7),
	.w2(32'hb9619c5f),
	.w3(32'hb9e822c1),
	.w4(32'hb9cfad1c),
	.w5(32'hb94e6c35),
	.w6(32'hb9504723),
	.w7(32'hb94ef345),
	.w8(32'hb97e8a82),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943e31f),
	.w1(32'h383ffd81),
	.w2(32'hb8f4ace0),
	.w3(32'hb92e8b64),
	.w4(32'h38eec2df),
	.w5(32'hb89952d1),
	.w6(32'hb8e84c51),
	.w7(32'hb8cc7898),
	.w8(32'hb8b83d89),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84194af),
	.w1(32'hb7005a24),
	.w2(32'h385debe2),
	.w3(32'h3845eb92),
	.w4(32'h3628b9f4),
	.w5(32'h389ed54b),
	.w6(32'hb7586cb1),
	.w7(32'hb74484a5),
	.w8(32'h37cf3f1b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39929c68),
	.w1(32'h3aa06781),
	.w2(32'h3a108a4c),
	.w3(32'h38fab22c),
	.w4(32'h399edbeb),
	.w5(32'hb90e531e),
	.w6(32'hb9923e8a),
	.w7(32'h3944851f),
	.w8(32'h38a57050),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e03e21),
	.w1(32'hb95dffdf),
	.w2(32'hb99d2ee1),
	.w3(32'hb910b979),
	.w4(32'hb82346f7),
	.w5(32'hb9d49e48),
	.w6(32'hb90fb513),
	.w7(32'hb9525a7a),
	.w8(32'hb9b9abdc),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007a09),
	.w1(32'h38e71f6f),
	.w2(32'hb8c47aa6),
	.w3(32'h388c6559),
	.w4(32'hb912ed2d),
	.w5(32'hb6987c66),
	.w6(32'h396fd030),
	.w7(32'h39a2f7d3),
	.w8(32'hb8804480),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93189b1),
	.w1(32'hb9b59f75),
	.w2(32'hb9e94add),
	.w3(32'hb9046d1f),
	.w4(32'hb9542979),
	.w5(32'hb9a0b0ef),
	.w6(32'hb91afce5),
	.w7(32'hb8f8637a),
	.w8(32'hb95201ca),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b8c0),
	.w1(32'hb96e8db2),
	.w2(32'hba382e30),
	.w3(32'hba25b070),
	.w4(32'hb9d293cf),
	.w5(32'hba2b7f13),
	.w6(32'hba2da500),
	.w7(32'hb94ee431),
	.w8(32'hb8d6ab78),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79f4e6d),
	.w1(32'hb940b29a),
	.w2(32'hb9278df2),
	.w3(32'hb795ba89),
	.w4(32'hb92a3955),
	.w5(32'hb935315e),
	.w6(32'hb811d118),
	.w7(32'hb918b7ff),
	.w8(32'hb92fb20d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922c2d1),
	.w1(32'hb88c5952),
	.w2(32'hb906b250),
	.w3(32'hb8f9bf54),
	.w4(32'hb8dcfba0),
	.w5(32'hb918ff6f),
	.w6(32'hb947c954),
	.w7(32'hb984ddf7),
	.w8(32'hb9b1011b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2725d0),
	.w1(32'h398a6d23),
	.w2(32'h39a24910),
	.w3(32'h39662af7),
	.w4(32'h3891b768),
	.w5(32'hb93d3143),
	.w6(32'h39d451a5),
	.w7(32'h39225a3b),
	.w8(32'hb8ed7787),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9893f16),
	.w1(32'h3aa59fb5),
	.w2(32'h3a42ce90),
	.w3(32'h396f85a8),
	.w4(32'h3a76ad3e),
	.w5(32'h39bc85d4),
	.w6(32'h38657a36),
	.w7(32'h3a09d943),
	.w8(32'h3a123f91),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344f52),
	.w1(32'hb9f20b6c),
	.w2(32'hb88452be),
	.w3(32'hba377213),
	.w4(32'hb9ea9969),
	.w5(32'hb92c8cca),
	.w6(32'hba6655df),
	.w7(32'hba41a47d),
	.w8(32'hb9d44115),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39237e73),
	.w1(32'hb9ba5fe9),
	.w2(32'h39a3600a),
	.w3(32'hb89196f9),
	.w4(32'hba08c580),
	.w5(32'hb866f254),
	.w6(32'hb8e7f79e),
	.w7(32'hba0fe158),
	.w8(32'hb9e0b26c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d3f45),
	.w1(32'hba257c41),
	.w2(32'hb8e0520a),
	.w3(32'h3948ab9f),
	.w4(32'hba0bf673),
	.w5(32'hb9116297),
	.w6(32'h39e0bd99),
	.w7(32'hb8d3385a),
	.w8(32'hb9a58326),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ffe3c),
	.w1(32'h3a404558),
	.w2(32'h399d4b2f),
	.w3(32'h3afcfd2a),
	.w4(32'h396e72fb),
	.w5(32'hb93fad78),
	.w6(32'h3a8b0a6f),
	.w7(32'h3a17f833),
	.w8(32'hb86ff225),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b60ad),
	.w1(32'h3ad0f348),
	.w2(32'h3a9bd5ae),
	.w3(32'h3927a9b3),
	.w4(32'h3a22ace4),
	.w5(32'h39b6f422),
	.w6(32'hba2204da),
	.w7(32'hb95959cf),
	.w8(32'hba096cce),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4be64),
	.w1(32'h3ad221c5),
	.w2(32'h39dbd98c),
	.w3(32'h3ab2afc3),
	.w4(32'h3a701392),
	.w5(32'h387aa979),
	.w6(32'h3a4adf0e),
	.w7(32'h3a5f8524),
	.w8(32'h398d224f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f990e7),
	.w1(32'hb8d5f92e),
	.w2(32'hb9d326ec),
	.w3(32'hb98636b4),
	.w4(32'hb99063af),
	.w5(32'hb9ece4cb),
	.w6(32'hb9324083),
	.w7(32'hb985e406),
	.w8(32'hb9bbeb23),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ada191),
	.w1(32'h3a46966f),
	.w2(32'h3a383366),
	.w3(32'h39bb7b68),
	.w4(32'h39a5a3ca),
	.w5(32'h3971537e),
	.w6(32'h3a196821),
	.w7(32'h3a209efa),
	.w8(32'h3a26e119),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7124c97),
	.w1(32'hb690a099),
	.w2(32'h3649d761),
	.w3(32'hb72a7f6a),
	.w4(32'hb63afc8c),
	.w5(32'h36049c0d),
	.w6(32'hb4812bae),
	.w7(32'h36d417a7),
	.w8(32'h3734ff09),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b32df4),
	.w1(32'h395f5e9a),
	.w2(32'h391128b2),
	.w3(32'h38f817e2),
	.w4(32'h39354162),
	.w5(32'h388e2ce2),
	.w6(32'h389a7307),
	.w7(32'hb609bf8a),
	.w8(32'hb93ead8a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b9960),
	.w1(32'hb96d1118),
	.w2(32'hb936639b),
	.w3(32'hb942e6ed),
	.w4(32'hb9300af2),
	.w5(32'hb929715c),
	.w6(32'hb839a379),
	.w7(32'hb91e55eb),
	.w8(32'hb92675b5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ab0c2),
	.w1(32'h3a87d78a),
	.w2(32'h3ac5e112),
	.w3(32'h39b5e739),
	.w4(32'h39e309d8),
	.w5(32'h3a2436ef),
	.w6(32'h39a402fd),
	.w7(32'h3a080dd5),
	.w8(32'h3a02d622),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3d71f),
	.w1(32'hb72bea87),
	.w2(32'h3669d5c8),
	.w3(32'hb669ec11),
	.w4(32'hb6d41c36),
	.w5(32'h35de187b),
	.w6(32'h3609af69),
	.w7(32'hb6017da4),
	.w8(32'h36a8e65b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85cce16),
	.w1(32'h38802f76),
	.w2(32'h38c6f7ff),
	.w3(32'hb882ea57),
	.w4(32'h37fd2ef2),
	.w5(32'h383d9353),
	.w6(32'hb74189fd),
	.w7(32'h388ed833),
	.w8(32'h387bc206),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39039677),
	.w1(32'hb97edde9),
	.w2(32'hb89e8569),
	.w3(32'h39a396ee),
	.w4(32'h38a9169b),
	.w5(32'hb8deb170),
	.w6(32'hb9c979de),
	.w7(32'hb8280c65),
	.w8(32'hb9085c83),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a657288),
	.w1(32'h3abc831a),
	.w2(32'h3ab5b43a),
	.w3(32'h39eb9090),
	.w4(32'h39c93449),
	.w5(32'h3a775424),
	.w6(32'hba9c88e1),
	.w7(32'hba51e996),
	.w8(32'h388b7aa9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73c440),
	.w1(32'h3aba80f4),
	.w2(32'h3ab6d3e6),
	.w3(32'hb9081339),
	.w4(32'h3ac15cb8),
	.w5(32'h3a357e7b),
	.w6(32'hb9a30edd),
	.w7(32'h3a363476),
	.w8(32'h388b1f39),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9e277),
	.w1(32'hb88c05d8),
	.w2(32'hb8ee7de5),
	.w3(32'hb8dd9b4c),
	.w4(32'hb85b0572),
	.w5(32'hb8977329),
	.w6(32'hb98ae5e2),
	.w7(32'hb971f291),
	.w8(32'hb945cc1d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafcf28),
	.w1(32'h3b0bac76),
	.w2(32'h3a4579af),
	.w3(32'h3a332b2c),
	.w4(32'h3ad5ddf4),
	.w5(32'h3966e53c),
	.w6(32'h39c537a2),
	.w7(32'h3ad0c0dc),
	.w8(32'h3abb5cf2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874d81),
	.w1(32'hbad193a7),
	.w2(32'hba22f7e1),
	.w3(32'h3ad54df2),
	.w4(32'h3897e4d0),
	.w5(32'hba174ded),
	.w6(32'h3b28b03f),
	.w7(32'h3af53548),
	.w8(32'hba4acb33),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20fcd3),
	.w1(32'h385e5342),
	.w2(32'hb7af7ff2),
	.w3(32'hb9febbfd),
	.w4(32'h3907958a),
	.w5(32'h3784ca70),
	.w6(32'hb93123d8),
	.w7(32'h3903d614),
	.w8(32'h3832ba69),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da0bdc),
	.w1(32'h37a49814),
	.w2(32'h381c927f),
	.w3(32'hb642ac14),
	.w4(32'h37cd84d5),
	.w5(32'h381f14aa),
	.w6(32'h379eec38),
	.w7(32'h38130f70),
	.w8(32'h382ab6d2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928e57c),
	.w1(32'h39ebe986),
	.w2(32'h39d99e2a),
	.w3(32'h38a1926d),
	.w4(32'h399939ee),
	.w5(32'h3989d14f),
	.w6(32'h38dc14de),
	.w7(32'h39a9c609),
	.w8(32'h39b28fe2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be7bf2),
	.w1(32'hb787b3b8),
	.w2(32'h366bfa08),
	.w3(32'hb7fa1f2d),
	.w4(32'hb78cf5b7),
	.w5(32'h362e608f),
	.w6(32'hb7e25548),
	.w7(32'hb75e316e),
	.w8(32'hb6019b87),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba328f68),
	.w1(32'h38ebef49),
	.w2(32'h3933aac8),
	.w3(32'hb97ceab2),
	.w4(32'h3913a033),
	.w5(32'hb8e0fef6),
	.w6(32'hba2bf878),
	.w7(32'hb9afe920),
	.w8(32'h395de779),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927e674),
	.w1(32'h39ac9345),
	.w2(32'hb81f7ae3),
	.w3(32'hb9cb6581),
	.w4(32'hb89171cc),
	.w5(32'hb9183aa6),
	.w6(32'hba280c31),
	.w7(32'hb9c2768f),
	.w8(32'hba0a0fab),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c40926),
	.w1(32'h39c166e6),
	.w2(32'h3a990618),
	.w3(32'hb9952f17),
	.w4(32'h39b3336d),
	.w5(32'h3a51ce2d),
	.w6(32'hb8abd551),
	.w7(32'h39b696e5),
	.w8(32'h399b20b2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885a750),
	.w1(32'h389cf491),
	.w2(32'h38e7ecc9),
	.w3(32'hb8a33fad),
	.w4(32'hb8411f91),
	.w5(32'h38c306af),
	.w6(32'hb8c26aaa),
	.w7(32'hb8c2ac2f),
	.w8(32'hb9193fe1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a9ac8),
	.w1(32'hba4d18d7),
	.w2(32'h3b1c5379),
	.w3(32'hb9d14fe3),
	.w4(32'h3b8e3cdf),
	.w5(32'h3bcdc51b),
	.w6(32'hb95c6d48),
	.w7(32'hbbd82930),
	.w8(32'hbbb4d358),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4ae0),
	.w1(32'hbb50c27b),
	.w2(32'hbc455f7f),
	.w3(32'h3b78b3bc),
	.w4(32'hbb1428c0),
	.w5(32'hbc2d0b56),
	.w6(32'hbb9a5e36),
	.w7(32'h3bd47683),
	.w8(32'h3b505e12),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005dea),
	.w1(32'hbb22fddd),
	.w2(32'hbc2ef096),
	.w3(32'hba9d60a4),
	.w4(32'h3b4ebf4f),
	.w5(32'hbc531d09),
	.w6(32'h3c0551ec),
	.w7(32'h3c42719f),
	.w8(32'h3c8a962d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dde24),
	.w1(32'hbb4eba2a),
	.w2(32'hbac597f5),
	.w3(32'h3b8dd2fb),
	.w4(32'h3c3f6625),
	.w5(32'hba6cf416),
	.w6(32'h3bbf7b08),
	.w7(32'h3c09d3bf),
	.w8(32'h3b523d3b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb528038),
	.w1(32'h3a949827),
	.w2(32'h3b06d19d),
	.w3(32'hbbcb9dce),
	.w4(32'h3a4184c0),
	.w5(32'hbbb3f85b),
	.w6(32'hbaf3b183),
	.w7(32'hba05a1ab),
	.w8(32'h3b126723),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb851006),
	.w1(32'hb9a85d49),
	.w2(32'hbbde411d),
	.w3(32'hbbc264b3),
	.w4(32'h3a82580f),
	.w5(32'hbb9f6b9c),
	.w6(32'h3ab40977),
	.w7(32'hbbd2cf7e),
	.w8(32'hbb0dab42),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0db18d),
	.w1(32'h3bd16c33),
	.w2(32'h3b388e8d),
	.w3(32'hba58388a),
	.w4(32'h3c2e8df6),
	.w5(32'hbbd3f09a),
	.w6(32'hbb8cd287),
	.w7(32'h3c565602),
	.w8(32'h3c994b13),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8acae5),
	.w1(32'hbba0129c),
	.w2(32'hbba0df21),
	.w3(32'h3baeb2fe),
	.w4(32'hbb72d488),
	.w5(32'h3b2f35fc),
	.w6(32'h3bd4e92b),
	.w7(32'hbaeefd12),
	.w8(32'hbbb2c2bc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e7caf),
	.w1(32'hb9ee943f),
	.w2(32'h3b6872b3),
	.w3(32'hbc061790),
	.w4(32'h3c23a4e0),
	.w5(32'hbbd6071b),
	.w6(32'hbc21c716),
	.w7(32'h3c2f5765),
	.w8(32'h3c3d048c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ac30),
	.w1(32'hbab0b8fb),
	.w2(32'hba2bbe2a),
	.w3(32'hbb63ca1c),
	.w4(32'hbae29f3e),
	.w5(32'h3b30a7f4),
	.w6(32'h39b1644b),
	.w7(32'h3b512023),
	.w8(32'hb91dd0c7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b235f39),
	.w1(32'hbb16efba),
	.w2(32'h3ae83356),
	.w3(32'h3b597533),
	.w4(32'hbbaa79fd),
	.w5(32'hbb9aaf5e),
	.w6(32'hbb8e1ea9),
	.w7(32'h39c9c98f),
	.w8(32'hbb69962b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0ff0),
	.w1(32'h3c1ffa5f),
	.w2(32'h3babb419),
	.w3(32'hbbbb8176),
	.w4(32'hba7e6546),
	.w5(32'h39896be5),
	.w6(32'hbc13f6b7),
	.w7(32'hbc6e942e),
	.w8(32'hbc848992),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8561c7),
	.w1(32'hb9a6472f),
	.w2(32'hbb4fc56e),
	.w3(32'h3a6cbba6),
	.w4(32'h3b104459),
	.w5(32'hbb0956a4),
	.w6(32'hbbc6c26f),
	.w7(32'h3a662a6f),
	.w8(32'h3b3dc926),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920cbd),
	.w1(32'h3b9a63a9),
	.w2(32'h3b1906e4),
	.w3(32'hbae89524),
	.w4(32'h3b9c6d6b),
	.w5(32'hbb01496a),
	.w6(32'h3b19b4f8),
	.w7(32'hbaca8798),
	.w8(32'h3b599d94),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44d0e),
	.w1(32'h3a41f25b),
	.w2(32'hbb30b07b),
	.w3(32'h3bc3a9bf),
	.w4(32'h3b94a605),
	.w5(32'h3a2d6051),
	.w6(32'h3bb86c4e),
	.w7(32'hbbe1bd84),
	.w8(32'h3b793f4e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd8cc),
	.w1(32'hbafd22c1),
	.w2(32'hbbd8c736),
	.w3(32'hb9eb7a77),
	.w4(32'h3c84ea68),
	.w5(32'hbae94d60),
	.w6(32'hba75f8d3),
	.w7(32'hb87ed056),
	.w8(32'h3c58458d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03cc6a),
	.w1(32'h38c583b2),
	.w2(32'h3b33ff81),
	.w3(32'hbbd6ee51),
	.w4(32'hbb2638e9),
	.w5(32'hbb9a5ee7),
	.w6(32'h3b9fba89),
	.w7(32'hbacbcc4c),
	.w8(32'hbc0f649d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936357),
	.w1(32'hbbbd0b73),
	.w2(32'hbbb40e74),
	.w3(32'h3b43e994),
	.w4(32'hba7fd2a7),
	.w5(32'hbc2889d5),
	.w6(32'hba5c6454),
	.w7(32'h3c2d2347),
	.w8(32'hbb02aebb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ecd72),
	.w1(32'hbbb3c561),
	.w2(32'h3c224a17),
	.w3(32'h3b07fa8f),
	.w4(32'hbc138486),
	.w5(32'hbbd7b808),
	.w6(32'hb9b6c41a),
	.w7(32'hba4037c9),
	.w8(32'hbb9248ae),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3de9d),
	.w1(32'hbb5c49a0),
	.w2(32'hbb52feb5),
	.w3(32'hbbc0b00c),
	.w4(32'hbb5e933f),
	.w5(32'hbb8a85e8),
	.w6(32'hbb03d96a),
	.w7(32'hbb9db68d),
	.w8(32'hba715d48),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd74f30),
	.w1(32'hbb7ecfdb),
	.w2(32'hbafae333),
	.w3(32'hbc0fe887),
	.w4(32'hbb441410),
	.w5(32'h3b121803),
	.w6(32'hbb1eebde),
	.w7(32'h3b96730f),
	.w8(32'h3b135f97),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937f17),
	.w1(32'hbb6b4c5a),
	.w2(32'hbaafa4b0),
	.w3(32'hbafe351d),
	.w4(32'hbb239588),
	.w5(32'h3a6643ae),
	.w6(32'h3b1f973c),
	.w7(32'hbb756642),
	.w8(32'hba13c0f7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5e2d),
	.w1(32'h3bc6ca71),
	.w2(32'h3c031322),
	.w3(32'hbc07ac53),
	.w4(32'hbbdad409),
	.w5(32'h3b9a971e),
	.w6(32'h3aa79215),
	.w7(32'hbb574a8c),
	.w8(32'hbb9be530),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d8fa4),
	.w1(32'h3b1d30ef),
	.w2(32'h3c23bbd3),
	.w3(32'h3b8b8c3a),
	.w4(32'h3c08e750),
	.w5(32'h3bf8b637),
	.w6(32'hbc03d9e0),
	.w7(32'hbb94090e),
	.w8(32'hbbf527d1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2089),
	.w1(32'h3c0b0699),
	.w2(32'h3c8ddd40),
	.w3(32'h3c53acca),
	.w4(32'hbbd1dfe9),
	.w5(32'h38e7363a),
	.w6(32'hbafb2f35),
	.w7(32'hbc4383cc),
	.w8(32'hbc3e9d5d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10b7b3),
	.w1(32'hba8e2f2d),
	.w2(32'hba43f00f),
	.w3(32'h3a90ca35),
	.w4(32'hbc33b232),
	.w5(32'hbc0c9ae0),
	.w6(32'hbbfc9943),
	.w7(32'hbbc511df),
	.w8(32'h3b6bf6bc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a715a2b),
	.w1(32'h3b39045c),
	.w2(32'h3bdfd8e2),
	.w3(32'hbc2b1d2e),
	.w4(32'h3b840d27),
	.w5(32'hba180316),
	.w6(32'hbb537e74),
	.w7(32'hbb84ad1c),
	.w8(32'h3b66bfbe),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0ae9),
	.w1(32'hba12fd78),
	.w2(32'hba06c927),
	.w3(32'h3b165f66),
	.w4(32'hba3e6e6d),
	.w5(32'hbc1a67c6),
	.w6(32'h3b65e177),
	.w7(32'hbbd7be09),
	.w8(32'hbb1a7b1c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffab54),
	.w1(32'hbaf40896),
	.w2(32'hbba07a0d),
	.w3(32'hbbf358ea),
	.w4(32'hbb62dade),
	.w5(32'hbb71a0e7),
	.w6(32'h3a38fb4e),
	.w7(32'hbc191260),
	.w8(32'hbc087334),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfa181),
	.w1(32'hbba2af0f),
	.w2(32'hbae71525),
	.w3(32'h39eab9a8),
	.w4(32'hbb261c34),
	.w5(32'hba418749),
	.w6(32'hbb93a36e),
	.w7(32'hbbcd0cc4),
	.w8(32'hba848c5e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbaa32),
	.w1(32'hb7ba20e3),
	.w2(32'h3b9ab4e1),
	.w3(32'hba0410a6),
	.w4(32'h3b329093),
	.w5(32'hbbe80ea0),
	.w6(32'hbba1a473),
	.w7(32'h3c162182),
	.w8(32'h3c773f55),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf939b),
	.w1(32'hba2e7f94),
	.w2(32'h3b09d22e),
	.w3(32'hbafbb0b0),
	.w4(32'hbb578858),
	.w5(32'hbbd28bb7),
	.w6(32'h3bb7d5cf),
	.w7(32'hbb306ea3),
	.w8(32'h3adc3390),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00bbe0),
	.w1(32'hbb82260d),
	.w2(32'hbbd21867),
	.w3(32'hbb4ec87a),
	.w4(32'h3c55942e),
	.w5(32'hbc2c3e6a),
	.w6(32'h3ac3dde3),
	.w7(32'h3c048887),
	.w8(32'h3c00ca30),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35e61f),
	.w1(32'hba603f50),
	.w2(32'h3b67a9f6),
	.w3(32'hbbbaf202),
	.w4(32'hbb8e2c99),
	.w5(32'hbc4be3e6),
	.w6(32'h39c398b2),
	.w7(32'h3b258c5b),
	.w8(32'h3b8220cc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a59f),
	.w1(32'h3ac98cc3),
	.w2(32'hbc24d438),
	.w3(32'hbb91de4a),
	.w4(32'h3aa79398),
	.w5(32'hbc169be9),
	.w6(32'h3ab4e15c),
	.w7(32'h3bd443e5),
	.w8(32'h3b5b64e8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1936e),
	.w1(32'h3a868226),
	.w2(32'hba98a9c1),
	.w3(32'hbc130c1f),
	.w4(32'h3bb7f2b3),
	.w5(32'h386e1c2c),
	.w6(32'h3ae2f3c5),
	.w7(32'hbb8f1b2d),
	.w8(32'h3bb3455e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43c90),
	.w1(32'h3b647f4b),
	.w2(32'h3b2e720c),
	.w3(32'h3b928f0e),
	.w4(32'hba104f27),
	.w5(32'hbb835517),
	.w6(32'h3bf6af7f),
	.w7(32'hbb275922),
	.w8(32'hbb9d7586),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96747d),
	.w1(32'hb9d8c027),
	.w2(32'h3aa496e3),
	.w3(32'h3b67f32a),
	.w4(32'hbb169f51),
	.w5(32'hb89a289f),
	.w6(32'hba98acc5),
	.w7(32'h3b7c0d9e),
	.w8(32'h3b3f8e0a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a243683),
	.w1(32'hbb49964a),
	.w2(32'hbb67f629),
	.w3(32'h3bad47ff),
	.w4(32'h3bc00eb2),
	.w5(32'h3bce17c7),
	.w6(32'h3a699277),
	.w7(32'h3b918a57),
	.w8(32'h3bcd91f0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fe15d),
	.w1(32'hbbeb58a6),
	.w2(32'hbbcf57eb),
	.w3(32'hbb2c6719),
	.w4(32'h3b8a49ec),
	.w5(32'hbc7d4424),
	.w6(32'hbb3a6ff5),
	.w7(32'h3b208658),
	.w8(32'h3c1b1e1f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90182),
	.w1(32'h3b41e104),
	.w2(32'hbb742056),
	.w3(32'hbb6f41a4),
	.w4(32'h3c547f4e),
	.w5(32'hbc18bb1f),
	.w6(32'h3bb8c5e7),
	.w7(32'h3bbd25c2),
	.w8(32'h3c82bfb9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9152f8),
	.w1(32'hbbaa76b2),
	.w2(32'hbc18fd99),
	.w3(32'hbc183842),
	.w4(32'hbb5e489b),
	.w5(32'h39f1601e),
	.w6(32'h3bac5d34),
	.w7(32'h3b71e0f5),
	.w8(32'hb9b14877),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803dcb),
	.w1(32'h3ab7de88),
	.w2(32'hb9586299),
	.w3(32'hba5dd21b),
	.w4(32'h3c528448),
	.w5(32'hbb41bd8b),
	.w6(32'h3bda3d9c),
	.w7(32'h3b21e075),
	.w8(32'hbaf178a9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bd679),
	.w1(32'hbba8f103),
	.w2(32'hbb2d00c7),
	.w3(32'h3bc97c46),
	.w4(32'h3b827437),
	.w5(32'hbaff0c8f),
	.w6(32'h3ba93330),
	.w7(32'hbc24cd87),
	.w8(32'hbbbe71ec),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd67abd),
	.w1(32'h3b536316),
	.w2(32'h3b2d8b67),
	.w3(32'hbb701828),
	.w4(32'h3ae7e4be),
	.w5(32'hbb47b5b9),
	.w6(32'h3aab8283),
	.w7(32'h3c0b04a5),
	.w8(32'h39fbd2b8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8baf),
	.w1(32'h3b2326aa),
	.w2(32'h3b4a9b7a),
	.w3(32'hbb776a25),
	.w4(32'h3aa6477a),
	.w5(32'h3bc090b0),
	.w6(32'hbaf15da9),
	.w7(32'hbbb1a443),
	.w8(32'hbc179bad),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8fac),
	.w1(32'hbba19f9b),
	.w2(32'hbbdde6be),
	.w3(32'h3baaa99f),
	.w4(32'hbb0ff722),
	.w5(32'hbb1d239a),
	.w6(32'hbc2817c3),
	.w7(32'h3c1444eb),
	.w8(32'h3bb9770a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9192ca),
	.w1(32'h3a9f603a),
	.w2(32'h3a36ce12),
	.w3(32'h3b86855d),
	.w4(32'h3c03e657),
	.w5(32'h3b3a3ec6),
	.w6(32'h3bc58c11),
	.w7(32'hba8d1f3a),
	.w8(32'h3b4b8ea0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977f68),
	.w1(32'h3c0e2d1b),
	.w2(32'h3c8e9c7c),
	.w3(32'h3a2937cb),
	.w4(32'h3c5422a0),
	.w5(32'h3c4c70b3),
	.w6(32'h3b9010eb),
	.w7(32'hba1e8a9f),
	.w8(32'hbb8136ff),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5f8f0),
	.w1(32'hbbc62223),
	.w2(32'h3b66009e),
	.w3(32'h3c28bc34),
	.w4(32'hbba73a40),
	.w5(32'hbc35620c),
	.w6(32'hbad7a99e),
	.w7(32'h3b8ed49b),
	.w8(32'h3baa2fa8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06805),
	.w1(32'h3ab56bc0),
	.w2(32'hbb9ee209),
	.w3(32'hbbb69317),
	.w4(32'h3bf392ac),
	.w5(32'hbb48543b),
	.w6(32'h3aad85a7),
	.w7(32'h3c0dbd23),
	.w8(32'h3a310747),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07fb8),
	.w1(32'hbbb84f97),
	.w2(32'hbb47b044),
	.w3(32'hbb412eb0),
	.w4(32'hbc1ce681),
	.w5(32'hbae315c9),
	.w6(32'h3a6956df),
	.w7(32'hbbac2892),
	.w8(32'hbb6dec31),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bf272),
	.w1(32'h3b9da658),
	.w2(32'h3b8cbed5),
	.w3(32'hbbd0e7ae),
	.w4(32'h3b99061b),
	.w5(32'hbb1fdfc5),
	.w6(32'hbbb18242),
	.w7(32'hbb368b86),
	.w8(32'h3aa3453b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c98bf),
	.w1(32'hbbbd5db0),
	.w2(32'hbb16b9f4),
	.w3(32'h3bd0c364),
	.w4(32'hbb6d1db8),
	.w5(32'hbbccfbca),
	.w6(32'h3ba08b85),
	.w7(32'hbb29f9ab),
	.w8(32'hbbaaa3df),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2160f),
	.w1(32'h3b3698e2),
	.w2(32'h3b58b605),
	.w3(32'hbb6a2e42),
	.w4(32'h3c0651d2),
	.w5(32'h3afb6c8c),
	.w6(32'h3b48e8f1),
	.w7(32'hbbde0dd7),
	.w8(32'hbb8c1330),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecac88),
	.w1(32'hbbbf7836),
	.w2(32'hbbebb04e),
	.w3(32'h3be219ad),
	.w4(32'h3c49c888),
	.w5(32'hbca7120a),
	.w6(32'hbab0ed1d),
	.w7(32'h3bdfb996),
	.w8(32'h3c872087),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106eb0),
	.w1(32'hba2c6cfd),
	.w2(32'hbc100b6d),
	.w3(32'hba5441e9),
	.w4(32'h3b0f1c1a),
	.w5(32'hbc46d0a1),
	.w6(32'h394ffe8c),
	.w7(32'h3b3d53e7),
	.w8(32'h3c263281),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb350ef9),
	.w1(32'h3b0fb503),
	.w2(32'h3b51b47f),
	.w3(32'h3aa39279),
	.w4(32'h3940ffb5),
	.w5(32'h3ba243d7),
	.w6(32'h3bcc178d),
	.w7(32'hbc455ee7),
	.w8(32'hb9a5f8ab),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcde8cd),
	.w1(32'h3a702710),
	.w2(32'h3a9dad15),
	.w3(32'h3bea07dc),
	.w4(32'hbb7a9868),
	.w5(32'h3b0b203d),
	.w6(32'h3b27ed50),
	.w7(32'hbb2712e1),
	.w8(32'hbb9c9046),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule