module layer_10_featuremap_120(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba396c02),
	.w1(32'h392178a5),
	.w2(32'h38e8555d),
	.w3(32'h38f784f5),
	.w4(32'h3ba0cd87),
	.w5(32'h3ae3f0a7),
	.w6(32'h3a776fac),
	.w7(32'h39a496ab),
	.w8(32'hb9b640a3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b008),
	.w1(32'hbaa40c22),
	.w2(32'h39ddfaa1),
	.w3(32'hba5a0348),
	.w4(32'hb9f595f3),
	.w5(32'h3b21b81d),
	.w6(32'hbb02774a),
	.w7(32'h38fc6d35),
	.w8(32'h399f04ce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afcc3a),
	.w1(32'hb9262d18),
	.w2(32'h39372773),
	.w3(32'h3a9217f1),
	.w4(32'h39d2c18a),
	.w5(32'h38d8d46c),
	.w6(32'hba1cd088),
	.w7(32'h38925436),
	.w8(32'h3a3416b3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3d344),
	.w1(32'hbb6a8161),
	.w2(32'hbb7ba0d6),
	.w3(32'h3a1ff707),
	.w4(32'hbb8e7d4d),
	.w5(32'hbba2032b),
	.w6(32'h3ab0138b),
	.w7(32'h39e0b437),
	.w8(32'h3b19fbab),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121a44),
	.w1(32'hba84298f),
	.w2(32'h3a8f797d),
	.w3(32'hbb1c6a28),
	.w4(32'h38b07a5b),
	.w5(32'h38b54349),
	.w6(32'hb9d63740),
	.w7(32'h3a0a1f09),
	.w8(32'h394e810f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29f52a),
	.w1(32'h3af0ad5b),
	.w2(32'h39d19b42),
	.w3(32'h3a756743),
	.w4(32'h3b4f736d),
	.w5(32'h3b02f08a),
	.w6(32'h39e7668c),
	.w7(32'h3a7c9643),
	.w8(32'hbadda705),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b84894),
	.w1(32'hbabc7fdc),
	.w2(32'h3b3c2003),
	.w3(32'hba84bf36),
	.w4(32'h39473e3c),
	.w5(32'h3b27bab7),
	.w6(32'hb8603fe2),
	.w7(32'h3b19ea17),
	.w8(32'h3a8db588),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc855d),
	.w1(32'h38a38b95),
	.w2(32'hb91a848a),
	.w3(32'h3b1ce347),
	.w4(32'h3b0417c5),
	.w5(32'h39c61a60),
	.w6(32'h3999b612),
	.w7(32'h38a29a34),
	.w8(32'hb9f4b299),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5800ed),
	.w1(32'hbab41aa0),
	.w2(32'hba142f38),
	.w3(32'hba1c785b),
	.w4(32'hb9eddab5),
	.w5(32'hb9c68a46),
	.w6(32'h39945f07),
	.w7(32'hba4a21a6),
	.w8(32'hb9e09045),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9c4c),
	.w1(32'hbb08e7c5),
	.w2(32'h3a59e623),
	.w3(32'hbb4f54df),
	.w4(32'hb993181b),
	.w5(32'h3b5680f3),
	.w6(32'hbb07ed1e),
	.w7(32'h39f8108a),
	.w8(32'h3b2bbb8a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a0b28),
	.w1(32'h3b9fac96),
	.w2(32'h3b515785),
	.w3(32'h3a682a41),
	.w4(32'hbb1f373b),
	.w5(32'hbb264dce),
	.w6(32'hbb163051),
	.w7(32'hbb352ba2),
	.w8(32'hb9a082d4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc562fb),
	.w1(32'hba61fb7a),
	.w2(32'hb9d987ba),
	.w3(32'h3b184170),
	.w4(32'h3abe0a88),
	.w5(32'h3b3d3fad),
	.w6(32'hbac3853e),
	.w7(32'h3af4c001),
	.w8(32'hb9d08f01),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de36d),
	.w1(32'h3a93ce90),
	.w2(32'h3b17ab66),
	.w3(32'h3ac96d20),
	.w4(32'hb9bb48a8),
	.w5(32'h3a8e9327),
	.w6(32'hba6e0068),
	.w7(32'hba325119),
	.w8(32'h39b24abe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306f61),
	.w1(32'hbb28bd13),
	.w2(32'hba23a5e9),
	.w3(32'h39d56b57),
	.w4(32'h3a88dfb6),
	.w5(32'hb892176b),
	.w6(32'hbaee9112),
	.w7(32'hbad68d9b),
	.w8(32'hba02b4a4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6efeb),
	.w1(32'hb9687eee),
	.w2(32'h3a12484e),
	.w3(32'hba0c7e80),
	.w4(32'hbbaf6669),
	.w5(32'hbb12a4f5),
	.w6(32'h39bcca22),
	.w7(32'h3b3cdf2d),
	.w8(32'h3b1ad520),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae18e12),
	.w1(32'h3940620b),
	.w2(32'h3b24aad2),
	.w3(32'hbb4d6717),
	.w4(32'hb987a321),
	.w5(32'h3ac947f2),
	.w6(32'hba582474),
	.w7(32'hb86ec1bb),
	.w8(32'hb996878d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0553dc),
	.w1(32'hb9920643),
	.w2(32'h3bb1517a),
	.w3(32'hbaed627e),
	.w4(32'hbb90fc1e),
	.w5(32'h3b2b3d23),
	.w6(32'hbbffd863),
	.w7(32'h398bb61d),
	.w8(32'h39a25aff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76ca2),
	.w1(32'hbb41e0eb),
	.w2(32'h3a54eee5),
	.w3(32'hb9fa2f50),
	.w4(32'hba362fe6),
	.w5(32'h3ab97dd9),
	.w6(32'hba7b37db),
	.w7(32'h3a9a7dc5),
	.w8(32'hb78223eb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4a51),
	.w1(32'hbab1e093),
	.w2(32'h3acdad39),
	.w3(32'hba340ec2),
	.w4(32'hb9ddeda9),
	.w5(32'h3addf88f),
	.w6(32'hbb075728),
	.w7(32'h3a1f73de),
	.w8(32'h3b0c97e0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c7543),
	.w1(32'hbaecf04f),
	.w2(32'hba935ceb),
	.w3(32'h3aa0a12e),
	.w4(32'hba3ae8db),
	.w5(32'hbaa1217c),
	.w6(32'hb939cb37),
	.w7(32'hba253bca),
	.w8(32'hba81d459),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97cfec),
	.w1(32'h39ae02a6),
	.w2(32'h3b674c81),
	.w3(32'hba91c394),
	.w4(32'hb7a89a63),
	.w5(32'h3b07588d),
	.w6(32'hb816885b),
	.w7(32'h3b2b64ff),
	.w8(32'hbaed54aa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388aa13e),
	.w1(32'hb967ff3e),
	.w2(32'hbb48365b),
	.w3(32'hbb429c37),
	.w4(32'hbc14e796),
	.w5(32'hbbd87e0a),
	.w6(32'h3a128f61),
	.w7(32'h3b38510e),
	.w8(32'h3ace837f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad117b6),
	.w1(32'h3b758c98),
	.w2(32'h3c829dc9),
	.w3(32'hbb572f59),
	.w4(32'hbbc5af7d),
	.w5(32'h3c4bef4d),
	.w6(32'hba5a0b66),
	.w7(32'h3c94f805),
	.w8(32'h397379f0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be14103),
	.w1(32'hb989f442),
	.w2(32'h3b1df2c5),
	.w3(32'hbb850250),
	.w4(32'hb838997b),
	.w5(32'h3abffd31),
	.w6(32'hbad3eda8),
	.w7(32'hbaa01141),
	.w8(32'h39e99119),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bec86),
	.w1(32'hbaa7c4a3),
	.w2(32'h3b99dc35),
	.w3(32'hba8836e3),
	.w4(32'hb9de815e),
	.w5(32'h3badf53a),
	.w6(32'hbae3e75d),
	.w7(32'h3b122fc2),
	.w8(32'h3b370ecb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd14b3),
	.w1(32'hbb980d45),
	.w2(32'hbba68fef),
	.w3(32'h3a20301e),
	.w4(32'hbb699460),
	.w5(32'hbb696af0),
	.w6(32'hbbb022a3),
	.w7(32'hbbf7a4ca),
	.w8(32'hbbbba8d0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac156),
	.w1(32'hbac124d6),
	.w2(32'hbacd1018),
	.w3(32'hbbb81eae),
	.w4(32'hb9ea3235),
	.w5(32'hba8f3672),
	.w6(32'hb9022d7c),
	.w7(32'hba34ef3e),
	.w8(32'hbb072853),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4125ee),
	.w1(32'hb9d622b4),
	.w2(32'h3a86ec0d),
	.w3(32'hbb1b490d),
	.w4(32'h3abb8541),
	.w5(32'h3af89a96),
	.w6(32'h399d6563),
	.w7(32'hba276237),
	.w8(32'h3ab76672),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a931ace),
	.w1(32'hbb828945),
	.w2(32'h3bcb26b2),
	.w3(32'h3af45ecc),
	.w4(32'hbb58db0c),
	.w5(32'h3bfff9c8),
	.w6(32'hbb8eecde),
	.w7(32'h3c0550f7),
	.w8(32'h3b7eacf0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e6b72),
	.w1(32'hb9caf393),
	.w2(32'h3be94a88),
	.w3(32'h3b2358d9),
	.w4(32'hbb0c2c04),
	.w5(32'h3c0beebc),
	.w6(32'h3b951137),
	.w7(32'h3c2e828f),
	.w8(32'h3c3fc588),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfce5d1),
	.w1(32'h3a00716b),
	.w2(32'h3a999bec),
	.w3(32'hba88e5b8),
	.w4(32'h3835e5df),
	.w5(32'h3a0b6228),
	.w6(32'h3a378b8e),
	.w7(32'h3aebc1ec),
	.w8(32'hba849834),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d4f09),
	.w1(32'h39d3e2c5),
	.w2(32'h3a87f5af),
	.w3(32'hbadc0d91),
	.w4(32'h3a6b0cbd),
	.w5(32'h3aa7d521),
	.w6(32'hb9079958),
	.w7(32'hb64b53ef),
	.w8(32'hbb0b8a46),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b606bc),
	.w1(32'hbbb5dcda),
	.w2(32'hbb68eb80),
	.w3(32'hbad84a14),
	.w4(32'hbae202c1),
	.w5(32'hbac16f3d),
	.w6(32'hbba79dc0),
	.w7(32'hbabbc5ff),
	.w8(32'hb8341447),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c165fe),
	.w1(32'hbb6b477e),
	.w2(32'hbbc4fd54),
	.w3(32'hba7c28c1),
	.w4(32'hbbb686e5),
	.w5(32'hbbaff17a),
	.w6(32'h39ec2676),
	.w7(32'hbbd71cce),
	.w8(32'hbbbe0c8c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4644),
	.w1(32'h3a21373b),
	.w2(32'hb9ded57a),
	.w3(32'h3aadb31c),
	.w4(32'h3a482833),
	.w5(32'h39cc0199),
	.w6(32'h3a31aca1),
	.w7(32'h3a44767f),
	.w8(32'hba84ae26),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d34145),
	.w1(32'h3a51e07b),
	.w2(32'h3a13bef0),
	.w3(32'hba23eee3),
	.w4(32'h39ba8d5c),
	.w5(32'h3a4ef694),
	.w6(32'hb997d11e),
	.w7(32'h3aa2daa8),
	.w8(32'hba892652),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0395f7),
	.w1(32'hbabc0de4),
	.w2(32'h390811bc),
	.w3(32'hba6d4fc9),
	.w4(32'hbad578ba),
	.w5(32'h39965638),
	.w6(32'h39dabe1c),
	.w7(32'h3a23db6b),
	.w8(32'hbb43ee8e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431db7),
	.w1(32'hbaaa2146),
	.w2(32'h39ff0d93),
	.w3(32'h3b567af6),
	.w4(32'hbb21f40c),
	.w5(32'h3a77800d),
	.w6(32'h39f81cc8),
	.w7(32'hbaa05a78),
	.w8(32'h39e39d44),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ce5a7),
	.w1(32'h3b183480),
	.w2(32'h3b2308b4),
	.w3(32'h3b832534),
	.w4(32'h3b657319),
	.w5(32'h3b424589),
	.w6(32'h3b82ae75),
	.w7(32'h39341aad),
	.w8(32'h3ac45423),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73130f),
	.w1(32'hba72c072),
	.w2(32'h3a38b602),
	.w3(32'hba1d5167),
	.w4(32'hba5fac40),
	.w5(32'h39c6eaf1),
	.w6(32'hba0b26b2),
	.w7(32'hba09aa7c),
	.w8(32'hb9026256),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39987943),
	.w1(32'hbb66c8cd),
	.w2(32'h3a8263eb),
	.w3(32'h3a94a5e0),
	.w4(32'hbc371efc),
	.w5(32'h3b3bee50),
	.w6(32'h3bf118f7),
	.w7(32'h3c82f073),
	.w8(32'h3c52482b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4a379),
	.w1(32'h398d16fc),
	.w2(32'h39e38d69),
	.w3(32'hbc317159),
	.w4(32'hba049c8f),
	.w5(32'hb8522f6a),
	.w6(32'h393d6710),
	.w7(32'hb80c9600),
	.w8(32'hbb034c2b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953730a),
	.w1(32'hba0ed809),
	.w2(32'hba41ec18),
	.w3(32'hb9d189d5),
	.w4(32'hb995f93a),
	.w5(32'h39854e93),
	.w6(32'hba619a62),
	.w7(32'hbb215b6a),
	.w8(32'hbb81d703),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aec5a),
	.w1(32'hbb87375a),
	.w2(32'h3afa72f9),
	.w3(32'hbba1a52a),
	.w4(32'h38982c58),
	.w5(32'h3b906e4b),
	.w6(32'hbb3e6638),
	.w7(32'hbaeab9d6),
	.w8(32'h3af29ec7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae483b0),
	.w1(32'h3a628c63),
	.w2(32'h3b44a324),
	.w3(32'h3acfc352),
	.w4(32'h3a02fc0d),
	.w5(32'h3b1cdfe7),
	.w6(32'hb98076d2),
	.w7(32'h3a861dd4),
	.w8(32'h3b9b9fac),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc45a12),
	.w1(32'h39285031),
	.w2(32'h3b738052),
	.w3(32'h39e0f463),
	.w4(32'hb90558c3),
	.w5(32'h3b24d328),
	.w6(32'hb95bc77c),
	.w7(32'h3a725546),
	.w8(32'h3b09455c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b081a),
	.w1(32'hbb044a1e),
	.w2(32'h3aaadb4b),
	.w3(32'h3a9f3076),
	.w4(32'hbb18764a),
	.w5(32'h3b16e1ac),
	.w6(32'h3ab1605e),
	.w7(32'h3b6d5e7b),
	.w8(32'h3b4166fd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7f7e9),
	.w1(32'h3b768731),
	.w2(32'h3b4eef44),
	.w3(32'hbb1d5cb0),
	.w4(32'hba23beda),
	.w5(32'h3b118fc7),
	.w6(32'hbb893713),
	.w7(32'hbb5648c8),
	.w8(32'h3bf581b2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c908c7d),
	.w1(32'hbadd2393),
	.w2(32'hba7d0ccd),
	.w3(32'h3c1401c4),
	.w4(32'hba4a9794),
	.w5(32'h390689a1),
	.w6(32'hba2d54c1),
	.w7(32'hbaa6585a),
	.w8(32'hbb7702e9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c75b),
	.w1(32'h38cc5309),
	.w2(32'h3aaf80a8),
	.w3(32'hbb3325b0),
	.w4(32'h3afee019),
	.w5(32'h3ac78659),
	.w6(32'hb9b89e4c),
	.w7(32'hb973c105),
	.w8(32'hb98393ab),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba314989),
	.w1(32'hba6ee7a6),
	.w2(32'h3a944a23),
	.w3(32'h3924e393),
	.w4(32'h3a11504d),
	.w5(32'h3b17f551),
	.w6(32'hba9194a6),
	.w7(32'hba873b0f),
	.w8(32'hbb41ebc3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ade36),
	.w1(32'h3b57e850),
	.w2(32'h3b51a152),
	.w3(32'hbaa30af8),
	.w4(32'h3b4053bb),
	.w5(32'h3b846d3c),
	.w6(32'h3b5d2c61),
	.w7(32'h399b91a1),
	.w8(32'h3b09d39f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d7601),
	.w1(32'hba71095c),
	.w2(32'h39a2aa12),
	.w3(32'h3b844788),
	.w4(32'hb8fbd960),
	.w5(32'h3a7cb10d),
	.w6(32'hb7837180),
	.w7(32'h3aa5cc1f),
	.w8(32'hbb6fc56a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb740732),
	.w1(32'h3acba5c5),
	.w2(32'h3abb61b7),
	.w3(32'hbbe745b2),
	.w4(32'h3a2658bc),
	.w5(32'h3a83b4ff),
	.w6(32'hba6c691a),
	.w7(32'hbb101948),
	.w8(32'hb909964d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af94ef8),
	.w1(32'hbb6077c8),
	.w2(32'hbb57db39),
	.w3(32'h3abd6dfe),
	.w4(32'hbb13432b),
	.w5(32'hba0e7040),
	.w6(32'hbb5d2194),
	.w7(32'hbac7e262),
	.w8(32'hb93b6fe1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389bceaa),
	.w1(32'hbc38c1c4),
	.w2(32'h3b69fabe),
	.w3(32'hbb0296dc),
	.w4(32'hbc9c42cc),
	.w5(32'hbb39d10e),
	.w6(32'h3c22d15c),
	.w7(32'h3cd3ccc1),
	.w8(32'h3c8c1ede),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5f65),
	.w1(32'hba8bcf41),
	.w2(32'hbafce680),
	.w3(32'hbc6ce223),
	.w4(32'hbb943e48),
	.w5(32'hbad449c8),
	.w6(32'hb99036e3),
	.w7(32'hba2e512f),
	.w8(32'hbb290659),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d06dd),
	.w1(32'hba8d2b0e),
	.w2(32'hba9907c3),
	.w3(32'hbbc65351),
	.w4(32'h3a95efcd),
	.w5(32'hba2e1b4a),
	.w6(32'hbac08425),
	.w7(32'hbb67dfae),
	.w8(32'hbb35967e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cefbb),
	.w1(32'hbaef47e3),
	.w2(32'hba3e111d),
	.w3(32'h3a9b14e9),
	.w4(32'hba36391e),
	.w5(32'h39da19c6),
	.w6(32'hb810051f),
	.w7(32'h3a2e0b73),
	.w8(32'h39a500f6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a093396),
	.w1(32'hb9bb4b30),
	.w2(32'hb949e716),
	.w3(32'h3a88cc18),
	.w4(32'h3ad1fbff),
	.w5(32'h3a384827),
	.w6(32'h399f291c),
	.w7(32'hba187fb4),
	.w8(32'hba0f83b8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e393e3),
	.w1(32'h3aef83ee),
	.w2(32'h3ab7ccf6),
	.w3(32'h391df215),
	.w4(32'h3b2b066e),
	.w5(32'h3b32824f),
	.w6(32'h3a06af77),
	.w7(32'h3b00cee9),
	.w8(32'h39760d7b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391afd05),
	.w1(32'h39dd8b96),
	.w2(32'h3a950890),
	.w3(32'h3998c918),
	.w4(32'h3989968a),
	.w5(32'h3817aad2),
	.w6(32'h3b138e07),
	.w7(32'h3b0841fb),
	.w8(32'h3897cfc6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b021),
	.w1(32'hbb4fab01),
	.w2(32'hbac78ac4),
	.w3(32'hb9c3720a),
	.w4(32'hba4a3b14),
	.w5(32'hba013c45),
	.w6(32'hba9a887a),
	.w7(32'h3a91ca9b),
	.w8(32'hba9f4a2c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9135cef),
	.w1(32'hbab13913),
	.w2(32'hba27874a),
	.w3(32'hba8b9449),
	.w4(32'h3abf992c),
	.w5(32'h3b206ed7),
	.w6(32'hba5da106),
	.w7(32'hba04a049),
	.w8(32'h39e6c34d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5be2),
	.w1(32'hbb063982),
	.w2(32'hba9f50b2),
	.w3(32'h3b1a8a6b),
	.w4(32'h39800dcd),
	.w5(32'h3a0e9a05),
	.w6(32'hba1fe5bc),
	.w7(32'h3b026bfe),
	.w8(32'h3aa53d71),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39112dc1),
	.w1(32'hba30417e),
	.w2(32'hbb037a98),
	.w3(32'h3a8fdb34),
	.w4(32'h3977670e),
	.w5(32'hba81bbe6),
	.w6(32'hbb361365),
	.w7(32'hbbac48a9),
	.w8(32'hbb6a1251),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f05c),
	.w1(32'h3b44e323),
	.w2(32'h3bf52e97),
	.w3(32'h3a53ace0),
	.w4(32'hbb5e1f70),
	.w5(32'h3b0de07c),
	.w6(32'h3c809d53),
	.w7(32'h3c985fae),
	.w8(32'h3ca870f4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f93c),
	.w1(32'h3c17b63e),
	.w2(32'h3c60c0f5),
	.w3(32'hbb1d463f),
	.w4(32'hbbe6a9ec),
	.w5(32'h3c4a64d9),
	.w6(32'h3ab57b84),
	.w7(32'h3c52a502),
	.w8(32'h3baaef27),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64fa12),
	.w1(32'hb9518ed6),
	.w2(32'h3a6ec01b),
	.w3(32'hbb9765cf),
	.w4(32'h39f315c1),
	.w5(32'h398af342),
	.w6(32'h3a49cd23),
	.w7(32'h3910bf7b),
	.w8(32'hbb61ccc8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a0d23),
	.w1(32'h3a85814c),
	.w2(32'h3bb725bd),
	.w3(32'hbb823ea7),
	.w4(32'h3adcbdcb),
	.w5(32'h3b8b30d6),
	.w6(32'hbb39a0e1),
	.w7(32'hb9f01eec),
	.w8(32'h3b22466c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2b6a),
	.w1(32'hbaa34b58),
	.w2(32'hba473873),
	.w3(32'h39f9285c),
	.w4(32'hba4e7177),
	.w5(32'hb832e1b6),
	.w6(32'hb80b030c),
	.w7(32'h3a29a59c),
	.w8(32'h3a148ea9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ddec5),
	.w1(32'hba47be00),
	.w2(32'hba8271b3),
	.w3(32'h3a00c7eb),
	.w4(32'h39e7b669),
	.w5(32'hb9efb3e3),
	.w6(32'hba248b3a),
	.w7(32'hb9eb7184),
	.w8(32'hbab5723d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81896d),
	.w1(32'h39ccbf24),
	.w2(32'h39832c40),
	.w3(32'hb9fdfa37),
	.w4(32'h3aea1098),
	.w5(32'h3a56ac41),
	.w6(32'h3a276051),
	.w7(32'hb90b690f),
	.w8(32'hb9c86ce8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1db6e),
	.w1(32'h3b0be7be),
	.w2(32'h3b3b2957),
	.w3(32'h39ea35ce),
	.w4(32'h3a97940b),
	.w5(32'h3af281d5),
	.w6(32'hb99e2f4b),
	.w7(32'h3a2b7ccb),
	.w8(32'hbb05a07e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d6b78),
	.w1(32'h368ff383),
	.w2(32'h3a022315),
	.w3(32'hbace5efb),
	.w4(32'h3aa31271),
	.w5(32'h3ae7f4af),
	.w6(32'hb783b5d9),
	.w7(32'h3a5c23c7),
	.w8(32'h3a0ecd6a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb2f2),
	.w1(32'hbb2eb0d4),
	.w2(32'hbb304fe8),
	.w3(32'h3adbfac5),
	.w4(32'h3ab051b2),
	.w5(32'h3b0e61a9),
	.w6(32'hbb9e8a59),
	.w7(32'hbb286c7e),
	.w8(32'hbb706ee7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa5cc),
	.w1(32'hb9b2c36a),
	.w2(32'h3b03bc04),
	.w3(32'hbb0962a8),
	.w4(32'h3b49502c),
	.w5(32'h3b2cab34),
	.w6(32'hba07abf5),
	.w7(32'h3abeea9c),
	.w8(32'h3a8829bb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fda12d),
	.w1(32'h3a63ab71),
	.w2(32'h3ab8a25e),
	.w3(32'hbad081ff),
	.w4(32'h38d8b0a1),
	.w5(32'h3a2d61a4),
	.w6(32'hbaf2f0ba),
	.w7(32'h3a2361dc),
	.w8(32'h3a5cb439),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cb923),
	.w1(32'hbbb70fca),
	.w2(32'hbb41721f),
	.w3(32'hb9e6817c),
	.w4(32'hbb4baf09),
	.w5(32'h3b20ef62),
	.w6(32'hbc2e40f5),
	.w7(32'hbbc9001b),
	.w8(32'hbb8173eb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed8e0e),
	.w1(32'hba81c8d5),
	.w2(32'h3a354763),
	.w3(32'hbb93bf3d),
	.w4(32'hba8508ac),
	.w5(32'hba0d8de1),
	.w6(32'hba0dc9ae),
	.w7(32'h3aabca3a),
	.w8(32'hbab2a8fb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bfec),
	.w1(32'h3c08b294),
	.w2(32'h3c10bc5d),
	.w3(32'hbb4f762c),
	.w4(32'hbc1b6904),
	.w5(32'h3b6ab1c6),
	.w6(32'h3c215a4f),
	.w7(32'h3c5e9040),
	.w8(32'h3c3961b8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5851bd),
	.w1(32'h3a5db225),
	.w2(32'h3a00f6cf),
	.w3(32'hbba5fad1),
	.w4(32'h3a0d320c),
	.w5(32'h39ce4618),
	.w6(32'h39bcaacd),
	.w7(32'h3ac66fd3),
	.w8(32'hb9f11329),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39511bf5),
	.w1(32'h39f9d376),
	.w2(32'h3b2e5c5a),
	.w3(32'hb8c691cb),
	.w4(32'hbac553d2),
	.w5(32'h3aa4f0fc),
	.w6(32'h3aa2f3e4),
	.w7(32'h3b903ce7),
	.w8(32'h3b0fec02),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af794a9),
	.w1(32'hba9b6e7e),
	.w2(32'hbaa2205a),
	.w3(32'hbb35d9a7),
	.w4(32'h38013e37),
	.w5(32'h3a07ebad),
	.w6(32'hb98032bf),
	.w7(32'h3a5af462),
	.w8(32'h39d3bbb0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37881fe1),
	.w1(32'h3ca79148),
	.w2(32'h3c1c0c82),
	.w3(32'h398e6fbb),
	.w4(32'h3b83672e),
	.w5(32'h3be586fc),
	.w6(32'hbba9aa97),
	.w7(32'hbc17bf7f),
	.w8(32'hbac0f903),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4a423),
	.w1(32'hba78246e),
	.w2(32'h3a2c1aa8),
	.w3(32'h3c63ffcc),
	.w4(32'hba1a0069),
	.w5(32'h3ab09184),
	.w6(32'h3b1246ba),
	.w7(32'h3b7d5463),
	.w8(32'h3b29fa0c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb9389),
	.w1(32'h3ac5950a),
	.w2(32'hba20154c),
	.w3(32'hbade195d),
	.w4(32'h3b0c7309),
	.w5(32'h3a85ba75),
	.w6(32'h3a285b8e),
	.w7(32'hba41cec0),
	.w8(32'hbaaed73c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b6cc),
	.w1(32'h3a74557c),
	.w2(32'h3af0c685),
	.w3(32'hba316400),
	.w4(32'hb8c6da26),
	.w5(32'h3a27cfc2),
	.w6(32'h3968397d),
	.w7(32'h3acd0dd9),
	.w8(32'hba9000a3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fa0f3),
	.w1(32'hbb3bb6dd),
	.w2(32'hbaf3f119),
	.w3(32'hbb77702a),
	.w4(32'hbb5dae6b),
	.w5(32'hba4b3eb2),
	.w6(32'hbb641e53),
	.w7(32'hbb063b1c),
	.w8(32'hba9477a7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a230ca8),
	.w1(32'h3a8f8e26),
	.w2(32'h3b24fd8f),
	.w3(32'hbacbaa6d),
	.w4(32'h3acefa27),
	.w5(32'h3b036af7),
	.w6(32'h3b1755c7),
	.w7(32'h3b6e8f67),
	.w8(32'hba90aea4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4dcd),
	.w1(32'h3b759559),
	.w2(32'h3b9c88ee),
	.w3(32'hbb2f66f5),
	.w4(32'h3a8df649),
	.w5(32'h3b278c1b),
	.w6(32'h3a9f8756),
	.w7(32'h3818fe91),
	.w8(32'hbad6848a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78937e),
	.w1(32'hbb2c3900),
	.w2(32'h3a7a66db),
	.w3(32'h398345b1),
	.w4(32'hbb670835),
	.w5(32'h39584d72),
	.w6(32'hbaebd3a4),
	.w7(32'hb984e4f6),
	.w8(32'hb8cc9587),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad90360),
	.w1(32'h383ac1da),
	.w2(32'hb8924e54),
	.w3(32'hbb860ae5),
	.w4(32'hbaa77361),
	.w5(32'h37e6bd24),
	.w6(32'hbaa455fa),
	.w7(32'h3a38866d),
	.w8(32'hba4f4f6a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa16d9),
	.w1(32'h3b7d27b2),
	.w2(32'h3c89ad30),
	.w3(32'hbb8ab018),
	.w4(32'hbc591fe9),
	.w5(32'h3bf30980),
	.w6(32'h3b617854),
	.w7(32'h3ca15bee),
	.w8(32'h3c3e1697),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c395298),
	.w1(32'hba92f3c2),
	.w2(32'hb8f5728a),
	.w3(32'hbbf03636),
	.w4(32'hbb1f1c56),
	.w5(32'hb9d5dcce),
	.w6(32'hbaed168b),
	.w7(32'hbaaa9332),
	.w8(32'hbacf85d6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74f103),
	.w1(32'h3b126688),
	.w2(32'h3b0bc9ad),
	.w3(32'hbb1f6481),
	.w4(32'h3ad369fe),
	.w5(32'h3b01560d),
	.w6(32'h3ae5858b),
	.w7(32'h3a996cf3),
	.w8(32'h39ce665d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc205),
	.w1(32'hba0eec54),
	.w2(32'h3a5909cd),
	.w3(32'h3a8932ac),
	.w4(32'hba669296),
	.w5(32'h3c31b856),
	.w6(32'hbb19aa3e),
	.w7(32'h3c2cb58a),
	.w8(32'hbb3710fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ab9a),
	.w1(32'hbae634fb),
	.w2(32'hbafcb8f2),
	.w3(32'hbb955568),
	.w4(32'h3a0affe9),
	.w5(32'hbb37c9a3),
	.w6(32'hba1b42a7),
	.w7(32'hbb96d287),
	.w8(32'h39c1ff38),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2a617),
	.w1(32'h3a88def0),
	.w2(32'hb9b763da),
	.w3(32'h3a9e9fed),
	.w4(32'hb9cab6db),
	.w5(32'hb97ce654),
	.w6(32'h38855934),
	.w7(32'hb9ffb30f),
	.w8(32'hbb21eece),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8804b7),
	.w1(32'hba130985),
	.w2(32'h3b186938),
	.w3(32'h3abd3e5e),
	.w4(32'h3add8ff2),
	.w5(32'h3b738d7c),
	.w6(32'h3b618e67),
	.w7(32'h3bc9edc1),
	.w8(32'h3b30cb81),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc39a4),
	.w1(32'hbb463a4c),
	.w2(32'hbb3cd87c),
	.w3(32'h3a9fd975),
	.w4(32'hbb8a64ea),
	.w5(32'hbb655c55),
	.w6(32'hba8bea1f),
	.w7(32'hbbce23a6),
	.w8(32'hbc11732f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26fcd),
	.w1(32'hba9f149c),
	.w2(32'h3b038fe2),
	.w3(32'hbbabcf17),
	.w4(32'hbb87d630),
	.w5(32'hb9e51a1c),
	.w6(32'hbb880e7b),
	.w7(32'hbafbddee),
	.w8(32'hbab4ab63),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981b1b),
	.w1(32'hbae4c7d1),
	.w2(32'h3aafb67f),
	.w3(32'hbb9f6319),
	.w4(32'h3abdba1c),
	.w5(32'h3aab6d6d),
	.w6(32'hbad48d0f),
	.w7(32'hb9212651),
	.w8(32'hba8c7f62),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d895e),
	.w1(32'hbb0c4cc9),
	.w2(32'hbab7248f),
	.w3(32'hba1329e4),
	.w4(32'hb9fd016d),
	.w5(32'hba1a6c86),
	.w6(32'hba594755),
	.w7(32'hba9fc345),
	.w8(32'hbb3b1e87),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae630dd),
	.w1(32'h3a6893f7),
	.w2(32'h3ad21506),
	.w3(32'hbb320ab2),
	.w4(32'h3b5053fd),
	.w5(32'h3b077ad0),
	.w6(32'h3a82561d),
	.w7(32'h3b2e6524),
	.w8(32'h3add8597),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38faa109),
	.w1(32'hbb022676),
	.w2(32'hba3c8e47),
	.w3(32'hb9055cce),
	.w4(32'hba6acdb7),
	.w5(32'h395ad7b1),
	.w6(32'hba92b89f),
	.w7(32'hba22c49f),
	.w8(32'h392ddfab),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8f121),
	.w1(32'h3ad9e4b5),
	.w2(32'h3a807c5a),
	.w3(32'hbb09d2db),
	.w4(32'h3a5f11c7),
	.w5(32'h3961e001),
	.w6(32'h397d6680),
	.w7(32'h3a92bd67),
	.w8(32'h36e5a2da),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8052),
	.w1(32'h3b82452b),
	.w2(32'h3bd5fc6c),
	.w3(32'h3a0aad87),
	.w4(32'h3a68abed),
	.w5(32'h3b554114),
	.w6(32'h3934c078),
	.w7(32'h3b30aac0),
	.w8(32'hba9e6c68),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a279a54),
	.w1(32'hbaef1816),
	.w2(32'h3ae05b7d),
	.w3(32'hbbabc1fb),
	.w4(32'hb9c394e4),
	.w5(32'h3ac22ecb),
	.w6(32'hbb4b4784),
	.w7(32'hba3431e5),
	.w8(32'h3a3a9c56),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba4501),
	.w1(32'hbb0a86d1),
	.w2(32'h399f3985),
	.w3(32'hbb0b8863),
	.w4(32'hb90577bc),
	.w5(32'h3b067bc4),
	.w6(32'hbb3f9f24),
	.w7(32'hba3d3a3a),
	.w8(32'h3b89b451),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a41ed),
	.w1(32'h399eaa9f),
	.w2(32'h3a99e4ca),
	.w3(32'h3b2d9210),
	.w4(32'h3a78f5b9),
	.w5(32'h39f9565e),
	.w6(32'h3a9b7cfc),
	.w7(32'hba8a0edc),
	.w8(32'hbab784a2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cbb1c4),
	.w1(32'h3ab4885a),
	.w2(32'hb95ece91),
	.w3(32'hba84827f),
	.w4(32'h3b6a7415),
	.w5(32'h3b125b60),
	.w6(32'h3a907226),
	.w7(32'hbb27e181),
	.w8(32'h3a91ac5c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b414c52),
	.w1(32'h3b07d4b9),
	.w2(32'h3aa33a67),
	.w3(32'h3b3726c1),
	.w4(32'h3b1b0d3f),
	.w5(32'h3a6a86a3),
	.w6(32'h3b134472),
	.w7(32'h3755cb9f),
	.w8(32'hba38172c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48e85c),
	.w1(32'h3a95934a),
	.w2(32'h3b2f41b5),
	.w3(32'hbaac6f6a),
	.w4(32'hb7fa9a34),
	.w5(32'h3b38cbf4),
	.w6(32'hbaac4d46),
	.w7(32'hba05631b),
	.w8(32'hbabcb66c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85a6d3),
	.w1(32'hbabe5fc7),
	.w2(32'h3a9f90a5),
	.w3(32'hba8ed02e),
	.w4(32'hbb5ebdad),
	.w5(32'hba99dbd8),
	.w6(32'hbb1c362a),
	.w7(32'hbb7cbc83),
	.w8(32'hbb2ed842),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d1f9f),
	.w1(32'hb9856527),
	.w2(32'h3a8512ae),
	.w3(32'hbb282e88),
	.w4(32'h3b528940),
	.w5(32'h3b0ab1f9),
	.w6(32'hb98184ec),
	.w7(32'h3a77e057),
	.w8(32'h399eb6ae),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9f22b),
	.w1(32'h3a9268f4),
	.w2(32'h3a70a84b),
	.w3(32'h39768636),
	.w4(32'h3adfaf00),
	.w5(32'h3a7436cf),
	.w6(32'h38d94101),
	.w7(32'h39d419b0),
	.w8(32'hba214e56),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0197c9),
	.w1(32'h3ab2dc34),
	.w2(32'h3a212303),
	.w3(32'h399171b4),
	.w4(32'h3b2bd873),
	.w5(32'h3aa35b3a),
	.w6(32'h3953dc74),
	.w7(32'h39ace5b2),
	.w8(32'hb981278f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c0d9b),
	.w1(32'h3b489471),
	.w2(32'h3a184b59),
	.w3(32'h3a80721a),
	.w4(32'h3b0033d6),
	.w5(32'h3a7bdead),
	.w6(32'h3ac40984),
	.w7(32'h3b223fb0),
	.w8(32'h3addf602),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb952),
	.w1(32'hba30873a),
	.w2(32'h3a8527ed),
	.w3(32'h3aa169ea),
	.w4(32'h39b68622),
	.w5(32'h3a7bae58),
	.w6(32'h3a1bc4ba),
	.w7(32'hb9d43022),
	.w8(32'h3af66e6f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22ec13),
	.w1(32'h3a43c615),
	.w2(32'hbac976c7),
	.w3(32'h3b4ae05c),
	.w4(32'hba55f17f),
	.w5(32'hbb484208),
	.w6(32'h39b3b46a),
	.w7(32'hba732d66),
	.w8(32'hbb281285),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f37b),
	.w1(32'hb990d7de),
	.w2(32'hbafeb2f3),
	.w3(32'hbb8aeaa7),
	.w4(32'hb754ab04),
	.w5(32'hbb07a725),
	.w6(32'hb9a1cd3c),
	.w7(32'hbb1fa7d3),
	.w8(32'hba8ecb6c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56ec1c),
	.w1(32'h39169b12),
	.w2(32'h3af9332b),
	.w3(32'hba92b417),
	.w4(32'h39e6a9b5),
	.w5(32'h3af7bf88),
	.w6(32'h35a73ede),
	.w7(32'hba86a6ff),
	.w8(32'h3a94ffb6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b890a6),
	.w1(32'hba8bca81),
	.w2(32'hba0a7e19),
	.w3(32'h39a9040f),
	.w4(32'h3b337758),
	.w5(32'h3b36e6dc),
	.w6(32'h3ae13f42),
	.w7(32'h3b5edfd2),
	.w8(32'h3a628830),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ddc9),
	.w1(32'h3b60b346),
	.w2(32'h3acd6acc),
	.w3(32'h3ab869f9),
	.w4(32'h3b698352),
	.w5(32'h3b457069),
	.w6(32'h3b44b39e),
	.w7(32'h3b185497),
	.w8(32'hbb1c5ab4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8f685),
	.w1(32'h3ac5049e),
	.w2(32'h3a7824fa),
	.w3(32'hbb0b43a7),
	.w4(32'h3931ac43),
	.w5(32'hba4b0a38),
	.w6(32'h3a7e4fbf),
	.w7(32'hb9336ecc),
	.w8(32'hbb0ffa27),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a37625),
	.w1(32'hba0957fa),
	.w2(32'h393bb03c),
	.w3(32'hbb64d336),
	.w4(32'hba6205e0),
	.w5(32'hb9bcc24f),
	.w6(32'hba8286bc),
	.w7(32'hba89eaee),
	.w8(32'hb9931d49),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a9420),
	.w1(32'h38e82b01),
	.w2(32'h3a06ea0e),
	.w3(32'hba0c575b),
	.w4(32'hb982cfe3),
	.w5(32'h39978ba3),
	.w6(32'hb89fc0c4),
	.w7(32'h39ba6605),
	.w8(32'h39f10841),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba907e5f),
	.w1(32'hb95d069a),
	.w2(32'h3afaf396),
	.w3(32'hbb188415),
	.w4(32'hba840012),
	.w5(32'h3aa0def2),
	.w6(32'hbadb16f0),
	.w7(32'hba21167c),
	.w8(32'h3a8658ac),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f3586),
	.w1(32'hb74e9bd1),
	.w2(32'h37f83686),
	.w3(32'hb907d9ba),
	.w4(32'hb6ea4156),
	.w5(32'hb8302113),
	.w6(32'h3865dab5),
	.w7(32'h3847a75a),
	.w8(32'hb8f5f4ca),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bb3a6),
	.w1(32'h39480e8c),
	.w2(32'h396b8bc7),
	.w3(32'h396e200f),
	.w4(32'hb8fcf423),
	.w5(32'hb89e6050),
	.w6(32'h39cb743e),
	.w7(32'hb8f907c5),
	.w8(32'h384807fb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb48acc96),
	.w1(32'h37ed03d0),
	.w2(32'h390d228f),
	.w3(32'hb9afb374),
	.w4(32'hb9cabbb2),
	.w5(32'hb86587a9),
	.w6(32'hb6e72229),
	.w7(32'hb8ffcfdc),
	.w8(32'h390de5f3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c66b96),
	.w1(32'hb93a4111),
	.w2(32'h39f41c25),
	.w3(32'hba235cdf),
	.w4(32'hb9c273e0),
	.w5(32'h39200451),
	.w6(32'hb98e5688),
	.w7(32'hb86d79b6),
	.w8(32'h39ae8de5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09acd4),
	.w1(32'h3a908215),
	.w2(32'h3a93c996),
	.w3(32'hba2e53a0),
	.w4(32'hb962ce01),
	.w5(32'h397094e4),
	.w6(32'hba19c20e),
	.w7(32'hb92aed4e),
	.w8(32'h3a4d8532),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f8691),
	.w1(32'hba00e558),
	.w2(32'h3a91699b),
	.w3(32'hbab79756),
	.w4(32'hb9d62399),
	.w5(32'hb98d3e7d),
	.w6(32'hba912433),
	.w7(32'h3a0e61d6),
	.w8(32'h3938eac9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22d8e8),
	.w1(32'hb9ce12f0),
	.w2(32'h3a934a59),
	.w3(32'hbaec64b2),
	.w4(32'hbad1513e),
	.w5(32'h388ec346),
	.w6(32'hba7195b8),
	.w7(32'hba7a9ca3),
	.w8(32'h39bcd1e8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803aee1),
	.w1(32'h39257e32),
	.w2(32'h3a259e45),
	.w3(32'hbadb613f),
	.w4(32'hbb046e43),
	.w5(32'h38d2965c),
	.w6(32'hbad842ff),
	.w7(32'hba5403f5),
	.w8(32'h397fdf20),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5e3a0),
	.w1(32'hb9508da7),
	.w2(32'h39a0bd5a),
	.w3(32'hb94f94fc),
	.w4(32'h37adffb2),
	.w5(32'hba24eb19),
	.w6(32'h3a7e236e),
	.w7(32'h3a486868),
	.w8(32'hb8ce5ac0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f89b7),
	.w1(32'hb96f49d2),
	.w2(32'h3a460702),
	.w3(32'hba228bde),
	.w4(32'hba2d03d3),
	.w5(32'h3996d891),
	.w6(32'hba0be935),
	.w7(32'hb9d4b19c),
	.w8(32'h3a0eabca),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba495551),
	.w1(32'hba894b26),
	.w2(32'h3a189277),
	.w3(32'hbaf17a56),
	.w4(32'hbac12f5a),
	.w5(32'hb79f5b93),
	.w6(32'hbaded01f),
	.w7(32'hba9cebc3),
	.w8(32'hb9a17073),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9452f1f),
	.w1(32'hb931485a),
	.w2(32'h3946ac2b),
	.w3(32'hba011bd6),
	.w4(32'hb9b3d6f6),
	.w5(32'hb81062ec),
	.w6(32'hb9b2222d),
	.w7(32'hb943b4b9),
	.w8(32'h38ac8624),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf7b1f),
	.w1(32'h39c1f237),
	.w2(32'h3b122432),
	.w3(32'hbb04b61e),
	.w4(32'hbb02e325),
	.w5(32'h3a895bd1),
	.w6(32'hba7268c0),
	.w7(32'hba32e62b),
	.w8(32'h3af27e96),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cfb1c),
	.w1(32'hba34d16a),
	.w2(32'hb9325956),
	.w3(32'hba785cdc),
	.w4(32'hba967767),
	.w5(32'hba609a1f),
	.w6(32'hb92690b6),
	.w7(32'hb9f245f2),
	.w8(32'hba526fda),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb759d97b),
	.w1(32'hb7a7c9e4),
	.w2(32'h3533f48f),
	.w3(32'hb73cf43e),
	.w4(32'hb7147c58),
	.w5(32'hb6560f35),
	.w6(32'hb71a0922),
	.w7(32'hb6ed9932),
	.w8(32'hb741097a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f412d8),
	.w1(32'h372c285e),
	.w2(32'h37874698),
	.w3(32'hb71b9a2b),
	.w4(32'h37f9c3b1),
	.w5(32'h3802894c),
	.w6(32'h376441fe),
	.w7(32'h38542ddf),
	.w8(32'h37b3ec8c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec4975),
	.w1(32'h3929ac73),
	.w2(32'h3a1e776a),
	.w3(32'hb92ab5d1),
	.w4(32'hb822af7a),
	.w5(32'h3a1d88ad),
	.w6(32'hb90158ae),
	.w7(32'hb84984e7),
	.w8(32'h3a6b74ec),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24cbac),
	.w1(32'hba692974),
	.w2(32'h39ac2818),
	.w3(32'hbb085dbc),
	.w4(32'hbafba01e),
	.w5(32'hba6459b0),
	.w6(32'hba3db43d),
	.w7(32'hb9f472d1),
	.w8(32'h383c6209),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff84ac),
	.w1(32'h3a66bb36),
	.w2(32'h3b25f36c),
	.w3(32'hb9c41150),
	.w4(32'h3a44c982),
	.w5(32'h3aece51f),
	.w6(32'h3909e039),
	.w7(32'h3abc2ab8),
	.w8(32'h3b42b8a2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787667e),
	.w1(32'hb700e0c6),
	.w2(32'hb73880bb),
	.w3(32'hb76c79d7),
	.w4(32'h363eb977),
	.w5(32'h3685a664),
	.w6(32'hb7aebbde),
	.w7(32'hb6c62e8f),
	.w8(32'h3700b1ed),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c682ff),
	.w1(32'h390edd1c),
	.w2(32'h3ae2228a),
	.w3(32'hbabdd6f2),
	.w4(32'hba68bd25),
	.w5(32'h3a4df481),
	.w6(32'hba62902d),
	.w7(32'hb953218e),
	.w8(32'h3a7f00eb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29732),
	.w1(32'hba22a552),
	.w2(32'h3ac4d905),
	.w3(32'hbb32e5b0),
	.w4(32'hbae23b92),
	.w5(32'h3a0031cc),
	.w6(32'hbb185c65),
	.w7(32'hba816b94),
	.w8(32'h3a9b3839),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e6af9),
	.w1(32'h39b88958),
	.w2(32'h3ab977e9),
	.w3(32'hbaddaf6a),
	.w4(32'hb9e4be68),
	.w5(32'h3956c39d),
	.w6(32'hbabd2254),
	.w7(32'h3956c9f8),
	.w8(32'h3a516bf4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39832203),
	.w1(32'hb7b8493c),
	.w2(32'h3aab5649),
	.w3(32'hba6e8d5c),
	.w4(32'hba1d5a68),
	.w5(32'h3a851d5e),
	.w6(32'hba255358),
	.w7(32'hb8f5a7aa),
	.w8(32'h3aabca2f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4859),
	.w1(32'hba0e2512),
	.w2(32'hba016ae1),
	.w3(32'hb867319f),
	.w4(32'hb9a76673),
	.w5(32'hba0d1b5e),
	.w6(32'hba1f5f05),
	.w7(32'hba3b7b70),
	.w8(32'hba068c36),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2566ca),
	.w1(32'hb9b3b3a6),
	.w2(32'hb8b405b2),
	.w3(32'hba957e97),
	.w4(32'hb9bf2b81),
	.w5(32'hba340d4c),
	.w6(32'hbaa3bf65),
	.w7(32'hba84ffe8),
	.w8(32'hba50b825),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd96e),
	.w1(32'h39039e3b),
	.w2(32'h39fa1a2c),
	.w3(32'h3a511b99),
	.w4(32'hb9d76b55),
	.w5(32'hb85c96f9),
	.w6(32'h3aab1d7d),
	.w7(32'hb9502edd),
	.w8(32'h38ebd101),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516639),
	.w1(32'hba441851),
	.w2(32'hba8afe1c),
	.w3(32'hbaafe932),
	.w4(32'hbb08a55c),
	.w5(32'hbaaf5e1d),
	.w6(32'hb9fd71ce),
	.w7(32'hbaa83e4d),
	.w8(32'hb9dab424),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ff249),
	.w1(32'hb9272912),
	.w2(32'hb8edb673),
	.w3(32'h3a657037),
	.w4(32'h3843bee7),
	.w5(32'h3820310e),
	.w6(32'h3a72df87),
	.w7(32'h390077f9),
	.w8(32'h39998de7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5433e),
	.w1(32'h38839465),
	.w2(32'h38cbd9d4),
	.w3(32'hb92e6997),
	.w4(32'h38cbb084),
	.w5(32'h379797d6),
	.w6(32'h37b0d47b),
	.w7(32'h38be7b9e),
	.w8(32'hb83241e9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831fd51),
	.w1(32'hb698c3d5),
	.w2(32'h3834e588),
	.w3(32'h386bdf9b),
	.w4(32'hb80fad35),
	.w5(32'h383282f7),
	.w6(32'h3822151c),
	.w7(32'hb7a42ec7),
	.w8(32'h3846e8a8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df588b),
	.w1(32'hb9daf6e9),
	.w2(32'h3a1f81e6),
	.w3(32'hbaa996d0),
	.w4(32'hba7b5009),
	.w5(32'hb93d3090),
	.w6(32'hba803b8b),
	.w7(32'hba5a2c38),
	.w8(32'hb98439ed),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb827b0de),
	.w1(32'hb79bb3de),
	.w2(32'h37f65f93),
	.w3(32'hb84a3975),
	.w4(32'h368c6341),
	.w5(32'h3846a9b4),
	.w6(32'h36b8bdfa),
	.w7(32'h36f8677a),
	.w8(32'h37e476b8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bcc22a),
	.w1(32'hba1200df),
	.w2(32'h39a8ea46),
	.w3(32'hb9cb0a14),
	.w4(32'hba4f8632),
	.w5(32'h393ee6a7),
	.w6(32'hb9d842d1),
	.w7(32'hb9b1e7be),
	.w8(32'h39d0b679),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab9023),
	.w1(32'hb8106b83),
	.w2(32'hb8f745aa),
	.w3(32'h38d1ceb8),
	.w4(32'h38921c35),
	.w5(32'h372029d9),
	.w6(32'h3964bd56),
	.w7(32'h38dee71a),
	.w8(32'h39011120),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa1b3),
	.w1(32'h3a8a7936),
	.w2(32'h3a1efc8f),
	.w3(32'h3a354bdf),
	.w4(32'h3a575990),
	.w5(32'h3a4ed941),
	.w6(32'h39f75958),
	.w7(32'h3a3dc90d),
	.w8(32'h3a4f0fe0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d2145),
	.w1(32'hb968827d),
	.w2(32'hb8b513b3),
	.w3(32'hb93b8479),
	.w4(32'hb9164da7),
	.w5(32'hb858847b),
	.w6(32'hb984846e),
	.w7(32'hb920109c),
	.w8(32'hb956c8e3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382fcd96),
	.w1(32'h398923ba),
	.w2(32'h397f0c14),
	.w3(32'hb8c4d7de),
	.w4(32'h38b3c853),
	.w5(32'h38a03275),
	.w6(32'h373fe3cf),
	.w7(32'h392aba67),
	.w8(32'h38d54853),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53a5de),
	.w1(32'hbaeb080a),
	.w2(32'hb7cdd376),
	.w3(32'hbadb96f9),
	.w4(32'hbb2b3ad0),
	.w5(32'hba971cf1),
	.w6(32'hba71993c),
	.w7(32'hbaf828fe),
	.w8(32'hba9d64be),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b0b05),
	.w1(32'hba776e50),
	.w2(32'h3b07abd5),
	.w3(32'hbaf2cbcc),
	.w4(32'hbb0827fb),
	.w5(32'h3981dce7),
	.w6(32'hb8286ad3),
	.w7(32'hba4af7be),
	.w8(32'h3a404745),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33125b),
	.w1(32'hb89e4bde),
	.w2(32'h38b8667e),
	.w3(32'h3a8fd9bf),
	.w4(32'h39e6d4d6),
	.w5(32'h39f274e3),
	.w6(32'h3a4e3b05),
	.w7(32'h38c9029f),
	.w8(32'h3a10e69c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f514c),
	.w1(32'hba18da96),
	.w2(32'h3acd4f5c),
	.w3(32'hbb263eca),
	.w4(32'hbaf4200d),
	.w5(32'h3a01c5ce),
	.w6(32'hbb0ff3a1),
	.w7(32'hbabe0424),
	.w8(32'h3a84ec7c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a47e68),
	.w1(32'hb9812e0f),
	.w2(32'h38711c81),
	.w3(32'hba11509e),
	.w4(32'hb9f6134e),
	.w5(32'hb9049ec5),
	.w6(32'hb9ec83f2),
	.w7(32'hb9b5b196),
	.w8(32'hb8c1ad5e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae9c5),
	.w1(32'hbaa98bb4),
	.w2(32'h3a403b6c),
	.w3(32'hbab1f2f9),
	.w4(32'hbaa456a4),
	.w5(32'h39f9e830),
	.w6(32'h39662fdd),
	.w7(32'h39e27c24),
	.w8(32'h3ab7dfec),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20115a),
	.w1(32'h3a68150c),
	.w2(32'h3ab4e5d8),
	.w3(32'hb99b4aff),
	.w4(32'h38638aab),
	.w5(32'h3a070bcf),
	.w6(32'h3814ae2f),
	.w7(32'h3a2f0411),
	.w8(32'h3a6bb3bd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90dde88),
	.w1(32'h3670828d),
	.w2(32'h3aa8acf5),
	.w3(32'hba9e42a3),
	.w4(32'hb9f355fb),
	.w5(32'h39e66c05),
	.w6(32'hba503508),
	.w7(32'hb924c880),
	.w8(32'h3a56178b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bd3e1),
	.w1(32'hb9790193),
	.w2(32'hb85b6f33),
	.w3(32'hb919959a),
	.w4(32'hb91e2888),
	.w5(32'hb99c616e),
	.w6(32'hb8987a51),
	.w7(32'hb9db6e28),
	.w8(32'hba0808a3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63a421),
	.w1(32'hba500f07),
	.w2(32'h395ed431),
	.w3(32'hbace8d3b),
	.w4(32'hbaa7a769),
	.w5(32'hb972c77d),
	.w6(32'hba493f40),
	.w7(32'hba5476cb),
	.w8(32'hb9913249),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8042a88),
	.w1(32'hb7a21e8d),
	.w2(32'hb80e802f),
	.w3(32'hb7a93bc5),
	.w4(32'hb6ff4e8c),
	.w5(32'hb7d66ab6),
	.w6(32'hb774bc7b),
	.w7(32'hb7435352),
	.w8(32'hb79a419c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6d7a2),
	.w1(32'h3a4852df),
	.w2(32'h3a7af1ae),
	.w3(32'h377d56fa),
	.w4(32'h39f21b6a),
	.w5(32'h3a590568),
	.w6(32'h3910372a),
	.w7(32'h39d3f21b),
	.w8(32'h3a70ab29),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c100c2),
	.w1(32'h388e801c),
	.w2(32'hb80677f8),
	.w3(32'hb8c1d240),
	.w4(32'hb82a153d),
	.w5(32'h383ed277),
	.w6(32'hb886b1dc),
	.w7(32'hb8118202),
	.w8(32'hb6511eb4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980bdd0),
	.w1(32'h39e38f1f),
	.w2(32'h3a5b0eac),
	.w3(32'hba33c304),
	.w4(32'hba8003fd),
	.w5(32'h39bdb61e),
	.w6(32'hb99252be),
	.w7(32'h38fe2597),
	.w8(32'h3a806e8d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70ff77c),
	.w1(32'h36096465),
	.w2(32'hb6e40a07),
	.w3(32'hb6c7f658),
	.w4(32'h362ae2d3),
	.w5(32'hb6459b4c),
	.w6(32'hb74607a7),
	.w7(32'hb59c5820),
	.w8(32'hb5ed5ff3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379248d5),
	.w1(32'h387cc886),
	.w2(32'h38c02a6e),
	.w3(32'hb72273c2),
	.w4(32'h3865fb13),
	.w5(32'h387bc431),
	.w6(32'hb8989701),
	.w7(32'hb88f6e2d),
	.w8(32'hb7b78763),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a257a36),
	.w1(32'h39a20970),
	.w2(32'h399704cc),
	.w3(32'h3a1e6a93),
	.w4(32'h3910e352),
	.w5(32'h378e6fbc),
	.w6(32'h3a18763a),
	.w7(32'h39782fae),
	.w8(32'h397af791),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f01d7),
	.w1(32'hb86523f1),
	.w2(32'h3a2f6260),
	.w3(32'hb9e02114),
	.w4(32'hbaa389f6),
	.w5(32'hba4115e1),
	.w6(32'h380f9820),
	.w7(32'hb9a115df),
	.w8(32'hb88624fe),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f528ec),
	.w1(32'hb88d0f21),
	.w2(32'hb92016a0),
	.w3(32'h36f77a3b),
	.w4(32'hb74b48d6),
	.w5(32'hb91d4c84),
	.w6(32'h391d6a3c),
	.w7(32'hb80ba88f),
	.w8(32'hb906ae36),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390addc5),
	.w1(32'h3955fafa),
	.w2(32'h38c9cc90),
	.w3(32'h38fbc37a),
	.w4(32'h39310e08),
	.w5(32'hb741f343),
	.w6(32'h38f55510),
	.w7(32'hb7b871a8),
	.w8(32'hb8e38f32),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4c9aa),
	.w1(32'h3ad40e54),
	.w2(32'h3bae1972),
	.w3(32'hbb422db0),
	.w4(32'h3a8be396),
	.w5(32'h3b8b2251),
	.w6(32'hbb1f3b77),
	.w7(32'h3a4b3494),
	.w8(32'h3b8a1e8a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b15a0e),
	.w1(32'h38e0fcb7),
	.w2(32'h3afa330c),
	.w3(32'hbac96c73),
	.w4(32'hbb1aa5b8),
	.w5(32'h3a4e5779),
	.w6(32'hba95ac58),
	.w7(32'hbb095b75),
	.w8(32'h37f32a0c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffbe7f),
	.w1(32'hb97ee104),
	.w2(32'hb851d031),
	.w3(32'hb92e67b7),
	.w4(32'hb9335ffd),
	.w5(32'hb92f7cbd),
	.w6(32'hb930a952),
	.w7(32'hb96b5ee9),
	.w8(32'hb97785bb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a698d4),
	.w1(32'h37dd0470),
	.w2(32'hb78558aa),
	.w3(32'h37f438bf),
	.w4(32'h37d49d00),
	.w5(32'h36cbf2ff),
	.w6(32'h38278b12),
	.w7(32'h37deaf46),
	.w8(32'h36721b49),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870498f),
	.w1(32'h395427ab),
	.w2(32'h388dd308),
	.w3(32'h391a024d),
	.w4(32'h398d28ee),
	.w5(32'h3882ad81),
	.w6(32'h394ecda8),
	.w7(32'h3920a00d),
	.w8(32'h37635ddb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da85fb),
	.w1(32'h32bf7c84),
	.w2(32'hb6873de2),
	.w3(32'hb724a3e8),
	.w4(32'h3516018b),
	.w5(32'hb62a0a26),
	.w6(32'hb7870496),
	.w7(32'hb650a49a),
	.w8(32'hb7239496),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083712),
	.w1(32'hba2fa5bc),
	.w2(32'hb951148d),
	.w3(32'hba4cc054),
	.w4(32'hba537258),
	.w5(32'hba164c0a),
	.w6(32'hb9962b48),
	.w7(32'hba067c61),
	.w8(32'hba03988d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7587f3e),
	.w1(32'hb90053b3),
	.w2(32'h39a7c337),
	.w3(32'hba89e82a),
	.w4(32'hbab86ba5),
	.w5(32'hbacec109),
	.w6(32'hba0d1e42),
	.w7(32'hb9bd34e8),
	.w8(32'hb8c3b889),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d260d),
	.w1(32'h3880db9e),
	.w2(32'h3b062fee),
	.w3(32'hbaffd2f4),
	.w4(32'hba08c84c),
	.w5(32'h3a8cbf7a),
	.w6(32'hba93e250),
	.w7(32'h39506ab3),
	.w8(32'h3b0d2471),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d1696),
	.w1(32'h3a1c7894),
	.w2(32'h3a0d812a),
	.w3(32'h3960bce8),
	.w4(32'h38872879),
	.w5(32'h38de5f80),
	.w6(32'h38e22fed),
	.w7(32'h38878bdd),
	.w8(32'hb7f586f8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab76ca7),
	.w1(32'hba0d6471),
	.w2(32'h3b1d489a),
	.w3(32'hbb0f37ba),
	.w4(32'hba5e7772),
	.w5(32'h3ac3e0e6),
	.w6(32'hbae5f818),
	.w7(32'h39bf558e),
	.w8(32'h3b2526b3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37849f48),
	.w1(32'h399df712),
	.w2(32'h39cefd2c),
	.w3(32'hb9e3d882),
	.w4(32'hb7ff1306),
	.w5(32'h39f84618),
	.w6(32'hb9018b09),
	.w7(32'h3929fd3f),
	.w8(32'h3a6a97cd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77cb9e2),
	.w1(32'hb75cfb50),
	.w2(32'hb802b28e),
	.w3(32'h350283ab),
	.w4(32'hb559b4c0),
	.w5(32'hb79f36ab),
	.w6(32'hb6c02df1),
	.w7(32'hb6e5da37),
	.w8(32'hb7dde298),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83b282e),
	.w1(32'h371c53b1),
	.w2(32'hb8246002),
	.w3(32'hb8772050),
	.w4(32'h38d68f36),
	.w5(32'hb80784c8),
	.w6(32'h38811a54),
	.w7(32'h389d31cc),
	.w8(32'hb8d9f753),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72ffc75),
	.w1(32'h37495b90),
	.w2(32'hb80ec91a),
	.w3(32'h36ff32aa),
	.w4(32'h37cc4018),
	.w5(32'hb79bec9d),
	.w6(32'hb70660e8),
	.w7(32'h35acff7e),
	.w8(32'hb82f941b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82c88e),
	.w1(32'hba4864a9),
	.w2(32'h3aac9e5a),
	.w3(32'hbac39b51),
	.w4(32'hbadba8de),
	.w5(32'h3a0dfa44),
	.w6(32'hba81f288),
	.w7(32'hba352eab),
	.w8(32'h3ac6e70b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6bd8),
	.w1(32'h3a58825b),
	.w2(32'h38930dba),
	.w3(32'h371727d4),
	.w4(32'hba339fe8),
	.w5(32'hb9b1c31b),
	.w6(32'h39b21bbd),
	.w7(32'hb9b819b7),
	.w8(32'hb9e58c32),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba102963),
	.w1(32'hb9920d09),
	.w2(32'h3ac07fec),
	.w3(32'hbaf388fa),
	.w4(32'hbacbb96d),
	.w5(32'h39d6107a),
	.w6(32'hbabcf3bb),
	.w7(32'hba91c738),
	.w8(32'h3a44fb8b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b90bd3),
	.w1(32'hb9390ca4),
	.w2(32'hb899bf98),
	.w3(32'h397db028),
	.w4(32'hb90d80b5),
	.w5(32'hb879ec4f),
	.w6(32'h396d7f8d),
	.w7(32'hb915b062),
	.w8(32'h38b82145),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82f6d),
	.w1(32'hbacd6c29),
	.w2(32'h3aaf034c),
	.w3(32'hbb42bec8),
	.w4(32'hbb3abc30),
	.w5(32'hb7305846),
	.w6(32'hbb0db640),
	.w7(32'hbaf85c7a),
	.w8(32'h3a048c3b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af8e0b),
	.w1(32'hb99e61eb),
	.w2(32'h3ab0a6ca),
	.w3(32'hba83b48f),
	.w4(32'hba08283c),
	.w5(32'h3a5a9464),
	.w6(32'hba25bcbd),
	.w7(32'hb66a5a26),
	.w8(32'h3a5e776d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290414),
	.w1(32'h3ac4cc3f),
	.w2(32'h3b0a2c0c),
	.w3(32'h3a66bc93),
	.w4(32'h3aa5969a),
	.w5(32'h3aca2895),
	.w6(32'h3a7567a9),
	.w7(32'h3b0d619c),
	.w8(32'h3b28ad69),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8284c1e),
	.w1(32'hb6457ec5),
	.w2(32'hb8052fa1),
	.w3(32'hb7b4f22d),
	.w4(32'h373fcc37),
	.w5(32'hb6b31dbd),
	.w6(32'hb7b705ed),
	.w7(32'h376b360c),
	.w8(32'h351b6550),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5322b02),
	.w1(32'hb6ba39dd),
	.w2(32'hb7b1062a),
	.w3(32'h36e4daf3),
	.w4(32'h37567390),
	.w5(32'hb70b6ae2),
	.w6(32'h36cc2d21),
	.w7(32'h35f51113),
	.w8(32'hb73fc9f4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43ff08),
	.w1(32'h3a21e5d4),
	.w2(32'h3aa95956),
	.w3(32'hb98e501f),
	.w4(32'hb981f084),
	.w5(32'h39e9a87b),
	.w6(32'h395a8fdb),
	.w7(32'h395ba7c1),
	.w8(32'h3a830d7c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01cd81),
	.w1(32'h37c3e4c3),
	.w2(32'h3b03357c),
	.w3(32'hbaa8dced),
	.w4(32'hba905ab3),
	.w5(32'h39c8876b),
	.w6(32'hba217443),
	.w7(32'h387e8ccc),
	.w8(32'h3aab5938),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d82fad),
	.w1(32'hb7f49948),
	.w2(32'h3af13e12),
	.w3(32'hba8b0991),
	.w4(32'hba303324),
	.w5(32'h3aab3b92),
	.w6(32'hb9956b88),
	.w7(32'h3894a36f),
	.w8(32'h3af614f5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e396d7),
	.w1(32'hb8a1b296),
	.w2(32'hb6e55340),
	.w3(32'hb826f786),
	.w4(32'h3813017e),
	.w5(32'hb7f894bf),
	.w6(32'h38327b01),
	.w7(32'hb8652095),
	.w8(32'hb97a2b75),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ae02e),
	.w1(32'h37529122),
	.w2(32'hb4e90982),
	.w3(32'h36aa48d1),
	.w4(32'h380e310d),
	.w5(32'h377c1d11),
	.w6(32'h381b9bfb),
	.w7(32'h381e4ca1),
	.w8(32'h36c8938b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37549989),
	.w1(32'h39029105),
	.w2(32'h38589503),
	.w3(32'h380dc632),
	.w4(32'h38cef610),
	.w5(32'h389bee81),
	.w6(32'h37acb3c3),
	.w7(32'h37096569),
	.w8(32'h3742966b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eec791),
	.w1(32'hb906969f),
	.w2(32'h3890127f),
	.w3(32'hba08d4e9),
	.w4(32'h3880cf81),
	.w5(32'h387280fa),
	.w6(32'hb9227d91),
	.w7(32'h39ebb1dd),
	.w8(32'h3a0059b6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13e9a9),
	.w1(32'h3afa3514),
	.w2(32'h3b13de61),
	.w3(32'h3a794852),
	.w4(32'h3b41a1ad),
	.w5(32'h3ac60c9d),
	.w6(32'h3aeb2462),
	.w7(32'h3b794c50),
	.w8(32'h3b2593c5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394384),
	.w1(32'hba887a44),
	.w2(32'h39180c20),
	.w3(32'hbb4d5307),
	.w4(32'hbabbe6e7),
	.w5(32'hb9cd34da),
	.w6(32'hbaf005df),
	.w7(32'hba925a2e),
	.w8(32'hba5fdc90),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386e58a5),
	.w1(32'hba4fec1d),
	.w2(32'hba20c8b0),
	.w3(32'h399cf394),
	.w4(32'hba44ae9e),
	.w5(32'hba0a881b),
	.w6(32'h3a12b3ca),
	.w7(32'hb9ff0f32),
	.w8(32'hb9065dbb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1924e4),
	.w1(32'h3acd7bc8),
	.w2(32'h3b111782),
	.w3(32'h3ac1a448),
	.w4(32'h3a39f925),
	.w5(32'h3ac2ae16),
	.w6(32'h3abf82ba),
	.w7(32'h3a35f0d1),
	.w8(32'h3af98cb8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72245bb),
	.w1(32'hb6d0ca07),
	.w2(32'hb784bd20),
	.w3(32'hb5bde3e8),
	.w4(32'h34bf2fbe),
	.w5(32'hb7221387),
	.w6(32'hb71d14f6),
	.w7(32'hb688c223),
	.w8(32'hb743a717),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67c9647),
	.w1(32'hb4d4fa93),
	.w2(32'hb768363f),
	.w3(32'h36922b46),
	.w4(32'h3732d5e6),
	.w5(32'hb7014682),
	.w6(32'h35ff514d),
	.w7(32'h36a90f5b),
	.w8(32'hb6f5e648),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c2737f),
	.w1(32'hb6c58ce7),
	.w2(32'hb729aa3f),
	.w3(32'h369c7648),
	.w4(32'hb78ab47d),
	.w5(32'hb8479291),
	.w6(32'hb7d78afd),
	.w7(32'hb73df2bd),
	.w8(32'hb7e393f7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78411f5),
	.w1(32'hb794798b),
	.w2(32'hb7c86261),
	.w3(32'hb683e7f1),
	.w4(32'h35da5158),
	.w5(32'hb75176cd),
	.w6(32'hb7adef19),
	.w7(32'hb700ad1f),
	.w8(32'hb7d35966),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996e40a),
	.w1(32'h38b5342f),
	.w2(32'hb7653af9),
	.w3(32'h391361ce),
	.w4(32'hb888b1bc),
	.w5(32'h36ff55d8),
	.w6(32'h3912ea91),
	.w7(32'hb8b71389),
	.w8(32'hb702487c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f80f6),
	.w1(32'h392026c1),
	.w2(32'h3aa52d97),
	.w3(32'h37f017a4),
	.w4(32'hba4d0c97),
	.w5(32'h3a067ce7),
	.w6(32'h39939729),
	.w7(32'h394e620c),
	.w8(32'h3a8889bd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396dac8b),
	.w1(32'h37d9d803),
	.w2(32'h3ac99eff),
	.w3(32'hbad1651a),
	.w4(32'hbad61632),
	.w5(32'h39005d14),
	.w6(32'hbaa5a675),
	.w7(32'hba9a8221),
	.w8(32'h39bd3bc1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7966ecd),
	.w1(32'hb8062804),
	.w2(32'hb823ac03),
	.w3(32'hb6f113d6),
	.w4(32'hb7ae7c50),
	.w5(32'hb81257db),
	.w6(32'hb8001464),
	.w7(32'hb7c4c393),
	.w8(32'hb81e981d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca5e80),
	.w1(32'hb9a2f825),
	.w2(32'h3a34f04d),
	.w3(32'hbad8fbae),
	.w4(32'hb8908e74),
	.w5(32'hb9ebbcf4),
	.w6(32'hba6f61c0),
	.w7(32'h39ee5bfa),
	.w8(32'h392019bb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b51e5a),
	.w1(32'h3905b050),
	.w2(32'h398e693c),
	.w3(32'hba1a166d),
	.w4(32'hb5b8b43e),
	.w5(32'h370e3341),
	.w6(32'hb9d2c656),
	.w7(32'h392c31b0),
	.w8(32'h36e32ddd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c42f89),
	.w1(32'h38632196),
	.w2(32'h38ccfa76),
	.w3(32'hb851d5fa),
	.w4(32'h384f659c),
	.w5(32'h38bfde51),
	.w6(32'h37c851aa),
	.w7(32'h39196edd),
	.w8(32'h393b9a0c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e233b5),
	.w1(32'hb99da8c4),
	.w2(32'h3932f959),
	.w3(32'hba0a4417),
	.w4(32'hb98dc4dd),
	.w5(32'hb9192415),
	.w6(32'hb93f555a),
	.w7(32'h390950c4),
	.w8(32'h388721d6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb54b2c50),
	.w1(32'hb816414c),
	.w2(32'hb8cdcfe3),
	.w3(32'hb77d93b6),
	.w4(32'hb8ba7e5f),
	.w5(32'hb92be8c0),
	.w6(32'hb8db6b21),
	.w7(32'hb9207411),
	.w8(32'hb96aa2a3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c3918),
	.w1(32'hb98e1ae2),
	.w2(32'hb878d713),
	.w3(32'hb844d3f9),
	.w4(32'hb8b79002),
	.w5(32'h378a21a2),
	.w6(32'hb8d4a134),
	.w7(32'hb8f47ffe),
	.w8(32'hb83c651e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7301629),
	.w1(32'hb7061736),
	.w2(32'hb705e2b6),
	.w3(32'hb810a230),
	.w4(32'hb8218e71),
	.w5(32'hb7eabffc),
	.w6(32'hb7607743),
	.w7(32'hb7b1434f),
	.w8(32'hb7298b72),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d8332),
	.w1(32'hb789039a),
	.w2(32'hb810fcac),
	.w3(32'hb70f4a8b),
	.w4(32'hb6c737df),
	.w5(32'hb7dcf9db),
	.w6(32'hb7963fea),
	.w7(32'hb6cf428e),
	.w8(32'hb7dd078a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85ff19),
	.w1(32'h39c77faf),
	.w2(32'h390d1448),
	.w3(32'h3aaa7880),
	.w4(32'h39f8bbc8),
	.w5(32'h39823b2c),
	.w6(32'h3a87e265),
	.w7(32'h3a624b45),
	.w8(32'h3a20170d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d342c),
	.w1(32'hb827344e),
	.w2(32'h3acf0fbf),
	.w3(32'hbac07587),
	.w4(32'hba198c21),
	.w5(32'h3a6dbee4),
	.w6(32'hba0e80f4),
	.w7(32'h39e9959d),
	.w8(32'h3a96ab49),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb717d),
	.w1(32'hb8a336f5),
	.w2(32'h3a648964),
	.w3(32'hba98a6b4),
	.w4(32'hba757e31),
	.w5(32'hb90b70a0),
	.w6(32'hba27f89c),
	.w7(32'hb9b0f66b),
	.w8(32'h38a4fb9f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947be2c),
	.w1(32'h390c2a9b),
	.w2(32'h3aee067f),
	.w3(32'hba9c4030),
	.w4(32'hb9b52dbc),
	.w5(32'h3a9f3988),
	.w6(32'hba6612db),
	.w7(32'h382fe64a),
	.w8(32'h3ac3e1a7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b7490),
	.w1(32'hb88b078e),
	.w2(32'hb8c00740),
	.w3(32'hb8864e9f),
	.w4(32'hb89facc3),
	.w5(32'hb8bcd3b5),
	.w6(32'hb8871878),
	.w7(32'hb8847ed2),
	.w8(32'hb89a98df),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7312c23),
	.w1(32'hb57b1b86),
	.w2(32'h3629ec2f),
	.w3(32'hb54d1ef2),
	.w4(32'hb61570ad),
	.w5(32'hb4b18e66),
	.w6(32'hb6e8246c),
	.w7(32'hb7010622),
	.w8(32'hb6fa7674),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dea5b5),
	.w1(32'hb69ca739),
	.w2(32'h36ccc589),
	.w3(32'hb805f330),
	.w4(32'h382e0357),
	.w5(32'h37bc55b9),
	.w6(32'hb7d74b07),
	.w7(32'h37fa1171),
	.w8(32'h38052414),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62910c3),
	.w1(32'h370a17a4),
	.w2(32'h36fb862c),
	.w3(32'hb7c4f410),
	.w4(32'hb7abbac4),
	.w5(32'hb7c1e4e8),
	.w6(32'hb7a91484),
	.w7(32'hb80701e2),
	.w8(32'hb7ebb8c1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba702af1),
	.w1(32'hba21b1a8),
	.w2(32'h3a3e08e9),
	.w3(32'hbabc0189),
	.w4(32'hba879866),
	.w5(32'hb8a66bd6),
	.w6(32'hba82e12a),
	.w7(32'hba28db7d),
	.w8(32'h38960600),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959659e),
	.w1(32'h388db7b2),
	.w2(32'hb74fd347),
	.w3(32'h39875b1e),
	.w4(32'h39558d23),
	.w5(32'h3959a5b0),
	.w6(32'h3994e2ed),
	.w7(32'h39b08ea6),
	.w8(32'h397c10ef),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63260cc),
	.w1(32'h38d14b6e),
	.w2(32'h381dc09c),
	.w3(32'h3813bf0e),
	.w4(32'hb8e8f843),
	.w5(32'h3800388e),
	.w6(32'h38e53919),
	.w7(32'hb997f567),
	.w8(32'hb7c91a54),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39defea8),
	.w1(32'h394997e1),
	.w2(32'hb726f514),
	.w3(32'h399138e6),
	.w4(32'h3884981b),
	.w5(32'h388197df),
	.w6(32'h39c13332),
	.w7(32'h388a258b),
	.w8(32'h39176d4a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891c99b),
	.w1(32'hb6a79ab1),
	.w2(32'hb87072ff),
	.w3(32'h3880189b),
	.w4(32'h377313d5),
	.w5(32'hb82b0e36),
	.w6(32'h37d79bff),
	.w7(32'hb878c5a0),
	.w8(32'hb8e70a5f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b5378),
	.w1(32'hb79949a7),
	.w2(32'h3a609b2d),
	.w3(32'hba186383),
	.w4(32'hb9665d58),
	.w5(32'h3a156f4f),
	.w6(32'hba1c0acb),
	.w7(32'hb842196f),
	.w8(32'h3a0f3d8c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8020c5c),
	.w1(32'h3685e327),
	.w2(32'hb724f926),
	.w3(32'hb883b43c),
	.w4(32'hb7b64e1a),
	.w5(32'hb773b141),
	.w6(32'hb895277a),
	.w7(32'hb7fff690),
	.w8(32'hb69b13f4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dad855),
	.w1(32'h3a8700f0),
	.w2(32'h3adfc969),
	.w3(32'hbaa2e10b),
	.w4(32'hba639fb3),
	.w5(32'h3a491773),
	.w6(32'hba43ac4b),
	.w7(32'hb9b9d2aa),
	.w8(32'h398e1410),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374b0a55),
	.w1(32'hb8bb4303),
	.w2(32'hb966a7c5),
	.w3(32'h3713c579),
	.w4(32'h38747670),
	.w5(32'hb87a22e7),
	.w6(32'h39b4e7b4),
	.w7(32'h3990f94d),
	.w8(32'h39d2411d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45401c),
	.w1(32'h3b013a5b),
	.w2(32'h3a740d53),
	.w3(32'h3b0cff43),
	.w4(32'h3a21a56a),
	.w5(32'hb87a5cca),
	.w6(32'h3aedeae3),
	.w7(32'h392dc6f3),
	.w8(32'h39b1fdc4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule