module layer_10_featuremap_430(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eadc22),
	.w1(32'hbb6e63e6),
	.w2(32'hbb7825af),
	.w3(32'h3b96337d),
	.w4(32'hbb15647c),
	.w5(32'h3b9b512c),
	.w6(32'h3c3294da),
	.w7(32'hb99b762d),
	.w8(32'hb8b920be),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc917ef),
	.w1(32'h3b005c8a),
	.w2(32'hba5b6edb),
	.w3(32'hb9895144),
	.w4(32'h3acf1226),
	.w5(32'h3b7545d8),
	.w6(32'hb9521a7f),
	.w7(32'h3b81c545),
	.w8(32'h3b88c2b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8deb75),
	.w1(32'h3c3e48ea),
	.w2(32'h3c358c12),
	.w3(32'h3a140391),
	.w4(32'h3c282336),
	.w5(32'h3c514fc6),
	.w6(32'hbb5178c8),
	.w7(32'h3ba7d8a7),
	.w8(32'h3b885156),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f07be),
	.w1(32'hbb89cddc),
	.w2(32'hbb5aad98),
	.w3(32'h3c0cec79),
	.w4(32'hba398d9f),
	.w5(32'hbb149d96),
	.w6(32'h3c1e686c),
	.w7(32'hbb91e90d),
	.w8(32'hbbcf839b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0abc0a),
	.w1(32'hbb9541fb),
	.w2(32'hbb983aa1),
	.w3(32'hbc161275),
	.w4(32'hbbe614d6),
	.w5(32'hbc05c528),
	.w6(32'hbc22311d),
	.w7(32'hbb8cedfb),
	.w8(32'hbbf3112c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc72daf),
	.w1(32'h3bcccbc8),
	.w2(32'h3b8f40dd),
	.w3(32'hbbea034f),
	.w4(32'h3bd1e66d),
	.w5(32'h3b06b601),
	.w6(32'hbbb15e04),
	.w7(32'h3b59eb1e),
	.w8(32'h3b27f247),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07fbee),
	.w1(32'h3b8dcf98),
	.w2(32'h3b6d9457),
	.w3(32'h3b48f96f),
	.w4(32'h3a9e2e21),
	.w5(32'h3b775ff2),
	.w6(32'h3b6a7e67),
	.w7(32'h38cfa280),
	.w8(32'hba395e85),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03cdf),
	.w1(32'hbbbb69e8),
	.w2(32'hb98efc7c),
	.w3(32'h3b06b832),
	.w4(32'hbaebcef0),
	.w5(32'h3c09d607),
	.w6(32'hbb7e91c8),
	.w7(32'h3af80381),
	.w8(32'h3b86a24b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdf926),
	.w1(32'h3b1259f3),
	.w2(32'h3b73ce3b),
	.w3(32'h3c0ff206),
	.w4(32'h3ba760b8),
	.w5(32'h3bfb2265),
	.w6(32'h3be38b77),
	.w7(32'h3aa46279),
	.w8(32'h3b5cb97a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b2964),
	.w1(32'h3c1ecc8a),
	.w2(32'h3b97bf51),
	.w3(32'hbac7d604),
	.w4(32'h3b31a114),
	.w5(32'hbbe00e82),
	.w6(32'h3b0200ea),
	.w7(32'h3a5b1afd),
	.w8(32'hbbd5bb0c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b216827),
	.w1(32'h3bac7192),
	.w2(32'h3bf14a37),
	.w3(32'hbba2a393),
	.w4(32'h38b7a1b9),
	.w5(32'h3b0d747c),
	.w6(32'hbb366477),
	.w7(32'hbbc80b7d),
	.w8(32'hbbb3ac3c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12257b),
	.w1(32'h3b8f3331),
	.w2(32'h3bb22c7b),
	.w3(32'h3c19a095),
	.w4(32'h3b6e1549),
	.w5(32'h3bd970b8),
	.w6(32'h3a5e1b19),
	.w7(32'h3b52fb66),
	.w8(32'h3ba3938d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9ded8),
	.w1(32'h3b88fe52),
	.w2(32'h3aea734f),
	.w3(32'h3b22bbd1),
	.w4(32'h3bd9e1d2),
	.w5(32'h3b639682),
	.w6(32'h3b4476bd),
	.w7(32'h3bfcf769),
	.w8(32'h3bc2b5e7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a7d3f),
	.w1(32'hbb862a5b),
	.w2(32'h3af4fdef),
	.w3(32'h39efd970),
	.w4(32'hbb6c1059),
	.w5(32'h3ac1ab85),
	.w6(32'h3ac5fabc),
	.w7(32'hbabfdef7),
	.w8(32'h3b40d26b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880c956),
	.w1(32'hbc1f4afa),
	.w2(32'hbaeedde9),
	.w3(32'hba2ed30f),
	.w4(32'hbc6d5c7f),
	.w5(32'hbc319407),
	.w6(32'hba66bc28),
	.w7(32'hbc870cde),
	.w8(32'hbc4e47dd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39186cec),
	.w1(32'hbbd3af5f),
	.w2(32'hbb69030b),
	.w3(32'hbb1675ef),
	.w4(32'hbbc79398),
	.w5(32'hbaa93ace),
	.w6(32'hbbe0d28b),
	.w7(32'hbba0a445),
	.w8(32'hba50e2ef),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58795),
	.w1(32'h3af4dce4),
	.w2(32'h3afaf863),
	.w3(32'hbb3fe2d5),
	.w4(32'h3b679c81),
	.w5(32'h3bd21af4),
	.w6(32'hbb3d3e42),
	.w7(32'hbbc66768),
	.w8(32'hbb6c2c32),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22083b),
	.w1(32'hba73d317),
	.w2(32'hbb7fe973),
	.w3(32'h3bdd5617),
	.w4(32'h383fe018),
	.w5(32'h3a72e036),
	.w6(32'hbac05c75),
	.w7(32'h3a5adbdb),
	.w8(32'h3a803338),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0c3df),
	.w1(32'hb9303539),
	.w2(32'h3b38b4a8),
	.w3(32'hb94366a2),
	.w4(32'h3a8953a0),
	.w5(32'h3b720a5b),
	.w6(32'hbb25d889),
	.w7(32'hba69a8d8),
	.w8(32'h39f31448),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cdb36),
	.w1(32'hbaec7fb7),
	.w2(32'h3a785002),
	.w3(32'h3a441c33),
	.w4(32'hbb9c8f0e),
	.w5(32'hbacf5b41),
	.w6(32'hb94d3ca8),
	.w7(32'hbc1af878),
	.w8(32'h3b2ce4be),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6b398),
	.w1(32'h3be36679),
	.w2(32'hbab54286),
	.w3(32'h3b8175f0),
	.w4(32'h3c66d82f),
	.w5(32'hbad4809c),
	.w6(32'h3a7be177),
	.w7(32'h3bbf4c94),
	.w8(32'hbaf267cd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf943),
	.w1(32'hbb6535e6),
	.w2(32'hb8c131a1),
	.w3(32'hbb13dc82),
	.w4(32'h38cdac38),
	.w5(32'h3a8aac35),
	.w6(32'hba396722),
	.w7(32'hbb163c25),
	.w8(32'hb9d3717b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ad467),
	.w1(32'h3bbc00d5),
	.w2(32'h3b8c60c2),
	.w3(32'h3ae8d86e),
	.w4(32'hba707abc),
	.w5(32'hbb50cb00),
	.w6(32'hba313ef5),
	.w7(32'h3bcd2409),
	.w8(32'h3bc9ab7b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab53355),
	.w1(32'hba133ce2),
	.w2(32'h3bde6997),
	.w3(32'hbb5eb1fc),
	.w4(32'h3aec1221),
	.w5(32'h3c02978b),
	.w6(32'h3995d33e),
	.w7(32'hbb99b20f),
	.w8(32'h3a0de27e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4509ce),
	.w1(32'hbb3648b3),
	.w2(32'hbb96ebb9),
	.w3(32'h3b3a7673),
	.w4(32'h3b96629b),
	.w5(32'hbc1195bf),
	.w6(32'hbbd426a3),
	.w7(32'h3b3c3420),
	.w8(32'hbb02c1e8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21377d),
	.w1(32'h3c91ddc4),
	.w2(32'h3c3ee00b),
	.w3(32'hbc34222e),
	.w4(32'h3c8d0ccd),
	.w5(32'h3c24dd8b),
	.w6(32'hbbfe9efa),
	.w7(32'h3c1a221e),
	.w8(32'h3bc08715),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdcdca),
	.w1(32'hb8e0126e),
	.w2(32'h3abcacfc),
	.w3(32'h3b2fd116),
	.w4(32'h3abeb3d2),
	.w5(32'h3b42e2f0),
	.w6(32'hbac39337),
	.w7(32'h3b1fd956),
	.w8(32'h3ba9d093),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c909),
	.w1(32'h3b6fc9b9),
	.w2(32'h3bcab62f),
	.w3(32'h3bcb000f),
	.w4(32'h3ba2405c),
	.w5(32'h3bd34be2),
	.w6(32'h3b81b7d0),
	.w7(32'h3b585445),
	.w8(32'h3b0e3cea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f38c8),
	.w1(32'h3ca3be50),
	.w2(32'h3b6e5492),
	.w3(32'h3b00d1cd),
	.w4(32'h3bb2296a),
	.w5(32'h3a84f02b),
	.w6(32'h3986aa56),
	.w7(32'hbb80ba4c),
	.w8(32'hbbe75ff6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fa37b),
	.w1(32'hba2b349a),
	.w2(32'hbbb39061),
	.w3(32'hbb85e824),
	.w4(32'h3b8e8610),
	.w5(32'hbb967ee4),
	.w6(32'hbc8fb9fa),
	.w7(32'h3bb10237),
	.w8(32'h3b0b9193),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26d4e2),
	.w1(32'hbb8b705c),
	.w2(32'hbb07390b),
	.w3(32'hbc05c1be),
	.w4(32'hbaa31dee),
	.w5(32'h3bad09cb),
	.w6(32'hba6b6312),
	.w7(32'hbb7ef827),
	.w8(32'h3abee5aa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4ce6),
	.w1(32'hbb3ae73e),
	.w2(32'h3b8fbf5c),
	.w3(32'h3b1ca256),
	.w4(32'hbb1a68bc),
	.w5(32'h3c0491dd),
	.w6(32'h3b367e61),
	.w7(32'hbb0a9fac),
	.w8(32'h3b9521d1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb03c),
	.w1(32'hbbc7e756),
	.w2(32'hbb97d119),
	.w3(32'h3bc7d832),
	.w4(32'h3a77645e),
	.w5(32'h39e0c5bb),
	.w6(32'h3b690e85),
	.w7(32'h3bb728f3),
	.w8(32'h3b4eb7b0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba407c1c),
	.w1(32'h3a1a88af),
	.w2(32'h3bc686ef),
	.w3(32'h3a041778),
	.w4(32'h3ba28572),
	.w5(32'h3c4cf5d1),
	.w6(32'h3b5ea33b),
	.w7(32'h3b364fb5),
	.w8(32'h3c0b4c45),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094ddf),
	.w1(32'hbaa05cd2),
	.w2(32'h3b3cd378),
	.w3(32'h3c0202b6),
	.w4(32'h3b9342cf),
	.w5(32'h3bb4aba7),
	.w6(32'h3b1fb818),
	.w7(32'h3bef9d2e),
	.w8(32'h3bd6b7e9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd35d59),
	.w1(32'h3b1fef2d),
	.w2(32'hbac9238e),
	.w3(32'hbae5d31b),
	.w4(32'h3b7e1a71),
	.w5(32'hba0362ef),
	.w6(32'hba8e3659),
	.w7(32'h389a35d8),
	.w8(32'hbb1649d8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb666a19),
	.w1(32'hbb5baf26),
	.w2(32'hbb8a7f2a),
	.w3(32'hbbc8406a),
	.w4(32'hbbd18366),
	.w5(32'hbb5aa9f6),
	.w6(32'hbc06b2b6),
	.w7(32'hbb9eb70e),
	.w8(32'hba8b3a63),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c37cb9),
	.w1(32'h3b7ca02e),
	.w2(32'h3b4842e8),
	.w3(32'h3c050914),
	.w4(32'h3ae75008),
	.w5(32'h3af9f5fd),
	.w6(32'h3b7a96ea),
	.w7(32'h3af455d4),
	.w8(32'h39d0797b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f2976),
	.w1(32'h3bfe56e8),
	.w2(32'h3bece066),
	.w3(32'h3b00ce73),
	.w4(32'h3b75fc32),
	.w5(32'h3c0d1d29),
	.w6(32'hba5a89f4),
	.w7(32'h3b585bc3),
	.w8(32'h3b919bb6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba302d5),
	.w1(32'hbaf07375),
	.w2(32'hbad7393b),
	.w3(32'h3be63452),
	.w4(32'hbaaa6f7b),
	.w5(32'hbb6817a6),
	.w6(32'h3bd4ebb5),
	.w7(32'hbb095b60),
	.w8(32'hbb32e65c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457a1f),
	.w1(32'hbc14a86b),
	.w2(32'hbbc7af4b),
	.w3(32'hbc0b2d52),
	.w4(32'hbc16da7b),
	.w5(32'hbb222167),
	.w6(32'hbbfce966),
	.w7(32'hbbf54afa),
	.w8(32'hbb9f3e0e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd25aa7),
	.w1(32'hba8f650e),
	.w2(32'hbbf1d1cf),
	.w3(32'hbac39177),
	.w4(32'hbb25296b),
	.w5(32'hbc2b51a8),
	.w6(32'hbb81b8fb),
	.w7(32'hbb305281),
	.w8(32'hbc18c3e2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083e26),
	.w1(32'h3bb3a32b),
	.w2(32'h3b43cd1a),
	.w3(32'hbbafd79a),
	.w4(32'h3bf9e60c),
	.w5(32'h3b72eaad),
	.w6(32'hbbd55a75),
	.w7(32'h3bc7db6c),
	.w8(32'h3ba2f115),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2635e4),
	.w1(32'hbac16795),
	.w2(32'h37ee579c),
	.w3(32'hba4fb8d0),
	.w4(32'hb92c7e32),
	.w5(32'h3c3f7e9c),
	.w6(32'hba8fef25),
	.w7(32'hb9f8ca77),
	.w8(32'h3b801581),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca2991),
	.w1(32'hbb1d2ae4),
	.w2(32'hbb0219e1),
	.w3(32'hbc1a8934),
	.w4(32'hbb8687b9),
	.w5(32'hbaf5c624),
	.w6(32'hbc0dc431),
	.w7(32'hbb4ac858),
	.w8(32'hbab1c7a5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d1c14),
	.w1(32'hbbc4902a),
	.w2(32'hbbdac264),
	.w3(32'hbb1f1ae7),
	.w4(32'hbb9bbfc8),
	.w5(32'hbba73c6d),
	.w6(32'hba709d58),
	.w7(32'hbb9c46d9),
	.w8(32'hbbb217c8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebc844),
	.w1(32'h3bf97769),
	.w2(32'h3b9da6ee),
	.w3(32'hbbb11513),
	.w4(32'h3c0972d3),
	.w5(32'h3beb94e6),
	.w6(32'hbba8a5bf),
	.w7(32'hbb44858d),
	.w8(32'h3b7800b6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831ecf0),
	.w1(32'h3c315aab),
	.w2(32'hbb971a72),
	.w3(32'h3b2d9fd6),
	.w4(32'h3be9c389),
	.w5(32'hbba93a88),
	.w6(32'h3b92e33c),
	.w7(32'h3c03a669),
	.w8(32'hbb0fde29),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4df582),
	.w1(32'hbbe80751),
	.w2(32'hbb4e2b85),
	.w3(32'hbbd1e4f4),
	.w4(32'hbb0db691),
	.w5(32'h3b870962),
	.w6(32'hbc0ebc56),
	.w7(32'hbb505d9b),
	.w8(32'h3b3da83f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb055c),
	.w1(32'hbae545d1),
	.w2(32'h3af227e1),
	.w3(32'hbb92ba79),
	.w4(32'h3b1a1df1),
	.w5(32'h3c486e7a),
	.w6(32'hbb828aa9),
	.w7(32'h38e0e930),
	.w8(32'h3c03c413),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136880),
	.w1(32'h3b51d431),
	.w2(32'h3aec6acc),
	.w3(32'h3b8b5ccd),
	.w4(32'h3ad1b5fc),
	.w5(32'h3aa8582b),
	.w6(32'h3acf7616),
	.w7(32'h3abe0866),
	.w8(32'hba4c5668),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245ead),
	.w1(32'hba771fe0),
	.w2(32'hbb6d47af),
	.w3(32'h3aa1ee08),
	.w4(32'h3b0c0f1a),
	.w5(32'hbb44a610),
	.w6(32'hbb3391ee),
	.w7(32'h3aac42af),
	.w8(32'hbb2832a1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901e88),
	.w1(32'hb9bf4f01),
	.w2(32'hba7c5e8f),
	.w3(32'h3a8fdb51),
	.w4(32'h3b1161b2),
	.w5(32'h39c23589),
	.w6(32'hb985d1ec),
	.w7(32'h3b7938dd),
	.w8(32'h3b84f24a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0448d2),
	.w1(32'h38b46261),
	.w2(32'hba45d2ff),
	.w3(32'hbb912419),
	.w4(32'h3ab58871),
	.w5(32'hbb812c20),
	.w6(32'hbae7db75),
	.w7(32'h3adde95f),
	.w8(32'hb970b961),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43af20),
	.w1(32'h3bc95939),
	.w2(32'h3afbb6ed),
	.w3(32'hbbaaac23),
	.w4(32'h3c0647ac),
	.w5(32'h39169e65),
	.w6(32'hbba35175),
	.w7(32'h3bbf1f0f),
	.w8(32'h3b5296ee),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4cae6),
	.w1(32'h3c589ffb),
	.w2(32'h3c2f54d3),
	.w3(32'h3aaf8b49),
	.w4(32'h3cb30190),
	.w5(32'h3c827291),
	.w6(32'h3af85960),
	.w7(32'h3c9652d8),
	.w8(32'h3c51bec1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394dad88),
	.w1(32'hbae9e933),
	.w2(32'h3b3e4342),
	.w3(32'h3ab6d799),
	.w4(32'hbb665e5f),
	.w5(32'hbb2afd71),
	.w6(32'hbb1c525a),
	.w7(32'hbb69efcb),
	.w8(32'hbaf6c1d5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4890),
	.w1(32'h3a9a0eb7),
	.w2(32'hbbb3ef8e),
	.w3(32'h3b3813ca),
	.w4(32'h3add242f),
	.w5(32'hbb84219d),
	.w6(32'h398485ba),
	.w7(32'h3b22b425),
	.w8(32'hbbce174d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54589e),
	.w1(32'hbaa8066f),
	.w2(32'h3ab6dc1d),
	.w3(32'h3baf9303),
	.w4(32'hba7ced03),
	.w5(32'h3a52c814),
	.w6(32'h3bed147f),
	.w7(32'hbb9966cb),
	.w8(32'hbb255791),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed868),
	.w1(32'h3bef33df),
	.w2(32'hbbaa9a17),
	.w3(32'h3b450c3f),
	.w4(32'h3c702234),
	.w5(32'hbb0e86b0),
	.w6(32'hb9d54f60),
	.w7(32'h3bfcdfce),
	.w8(32'h3c411463),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc141693),
	.w1(32'h3c33d9bb),
	.w2(32'h3b804a9b),
	.w3(32'hbbf24dc4),
	.w4(32'h3c033779),
	.w5(32'h3aaa0047),
	.w6(32'hbac5463f),
	.w7(32'h3bceab34),
	.w8(32'h3bbcfd45),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98e3ff),
	.w1(32'hbaab4a67),
	.w2(32'h3b485e6a),
	.w3(32'h3b1fe625),
	.w4(32'h3a75971c),
	.w5(32'h3baeb990),
	.w6(32'h3be73306),
	.w7(32'h3aaac7e2),
	.w8(32'h3bbc0d3f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b577de7),
	.w1(32'h3b8a8c6f),
	.w2(32'h3bc531f1),
	.w3(32'h3b6d9b13),
	.w4(32'h3c1a26ea),
	.w5(32'h3af33362),
	.w6(32'h3a822ad1),
	.w7(32'h3bb69b45),
	.w8(32'h3a85ad88),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601437),
	.w1(32'hbbb39a80),
	.w2(32'hbb094af5),
	.w3(32'hbb214336),
	.w4(32'hbbc0fbd3),
	.w5(32'h3869a44d),
	.w6(32'hbb191b26),
	.w7(32'hbb5a9b45),
	.w8(32'hb9639e5f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c84f6),
	.w1(32'hbbb41648),
	.w2(32'hbabf1248),
	.w3(32'h3a548b15),
	.w4(32'hba71bbd9),
	.w5(32'h3b1d7e50),
	.w6(32'h370d18f5),
	.w7(32'hbb37c6aa),
	.w8(32'h3a4feed9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e26d),
	.w1(32'h3b9a461b),
	.w2(32'h3a33ae69),
	.w3(32'hbbf17672),
	.w4(32'h3b93716d),
	.w5(32'h3b7155b3),
	.w6(32'hbbeecdc0),
	.w7(32'h3c0a6967),
	.w8(32'h3b8595f5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fee5d),
	.w1(32'hbb955e9d),
	.w2(32'hbbf6b952),
	.w3(32'h3bbc3d03),
	.w4(32'hbc0e8cbe),
	.w5(32'hbc36154f),
	.w6(32'h3bc6c0a8),
	.w7(32'hbbf45dd9),
	.w8(32'hbc0274d2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7d458),
	.w1(32'hbb3637f6),
	.w2(32'hbbc681de),
	.w3(32'hbbb962e0),
	.w4(32'hbaad58a4),
	.w5(32'h3906cdba),
	.w6(32'hbc01cefc),
	.w7(32'hbb8a829a),
	.w8(32'hbb5bc8dd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43f5f0),
	.w1(32'h3acee551),
	.w2(32'hbc19df52),
	.w3(32'hbb9d3313),
	.w4(32'hbad55a54),
	.w5(32'hbc1128c7),
	.w6(32'hbc4140b5),
	.w7(32'hbacbb604),
	.w8(32'hbc3e9c2d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842b6c),
	.w1(32'h3a9c8ed2),
	.w2(32'h3b99830a),
	.w3(32'hbc90ca2e),
	.w4(32'h3b7df2d9),
	.w5(32'h3c64af29),
	.w6(32'hbcbcaf2e),
	.w7(32'hbb3b43c8),
	.w8(32'hbb22a8ee),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab34187),
	.w1(32'h3c0d4941),
	.w2(32'hbb32f376),
	.w3(32'hbb5f8401),
	.w4(32'h3c3f827e),
	.w5(32'hbbcc8221),
	.w6(32'hba794162),
	.w7(32'h3b61aa23),
	.w8(32'hbb27c4ff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7235e),
	.w1(32'hbb6af22c),
	.w2(32'hbc2df857),
	.w3(32'hbb3dffe3),
	.w4(32'hbc006cb9),
	.w5(32'h3b8383ea),
	.w6(32'h3ab7200f),
	.w7(32'h3b1628d8),
	.w8(32'hbb2af948),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0729ca),
	.w1(32'h3ca38b8c),
	.w2(32'h3d081dfc),
	.w3(32'hbb9e8b3d),
	.w4(32'h3c81443e),
	.w5(32'h3d66e0d9),
	.w6(32'hba2fc9cb),
	.w7(32'h3c62967c),
	.w8(32'h3d2b67f9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392d31),
	.w1(32'h3ab2ed91),
	.w2(32'h3af880b7),
	.w3(32'h3ca6ada6),
	.w4(32'hbb9d65de),
	.w5(32'h3b91c048),
	.w6(32'h3ce8ae9c),
	.w7(32'hbaaee9f6),
	.w8(32'h3b2ef23c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b929671),
	.w1(32'hbb6456fd),
	.w2(32'hbc22bbf5),
	.w3(32'h3bc019c8),
	.w4(32'h3bc88e05),
	.w5(32'h3a994e54),
	.w6(32'h3b5faec2),
	.w7(32'hbb61f5fb),
	.w8(32'hbc0f1451),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc243878),
	.w1(32'hbb4aec06),
	.w2(32'hbb79da1a),
	.w3(32'hbc43c69b),
	.w4(32'hbbab2d75),
	.w5(32'hbb086a6d),
	.w6(32'hbae52164),
	.w7(32'hbb8ebcaa),
	.w8(32'hbba81b17),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba391f29),
	.w1(32'h3b2ed99a),
	.w2(32'h3a692704),
	.w3(32'h3a5753a8),
	.w4(32'hba92ba7b),
	.w5(32'hbc305910),
	.w6(32'hba9a4714),
	.w7(32'hba96e4e6),
	.w8(32'hbb2c5690),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b622604),
	.w1(32'h3ab2ee41),
	.w2(32'hbc0337e4),
	.w3(32'h3c1bae6d),
	.w4(32'h3b650d06),
	.w5(32'hbc087d23),
	.w6(32'h3b42e5ea),
	.w7(32'h3a6f88aa),
	.w8(32'hbc18b52c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8680),
	.w1(32'hbbc5ed54),
	.w2(32'hbbc80949),
	.w3(32'hbc07f069),
	.w4(32'hbb46dbde),
	.w5(32'hbc1d1aea),
	.w6(32'hbbe387e3),
	.w7(32'h3a2da29a),
	.w8(32'hbb16715a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04f540),
	.w1(32'hb91f0754),
	.w2(32'hbc3060dd),
	.w3(32'h3ba690ba),
	.w4(32'hbc1cb51c),
	.w5(32'hbc6edfcc),
	.w6(32'h3c1834d4),
	.w7(32'hbc2f5926),
	.w8(32'hbbc69f23),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bbe59),
	.w1(32'hbb6fc3aa),
	.w2(32'hb8ead55f),
	.w3(32'hbc3cd720),
	.w4(32'hbb6a5e2a),
	.w5(32'hbb943dd6),
	.w6(32'hbc31c498),
	.w7(32'h39a76c56),
	.w8(32'h39c0e55b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32ef0a),
	.w1(32'hb9f3e24e),
	.w2(32'h3af452c2),
	.w3(32'h3c63ce62),
	.w4(32'hba116552),
	.w5(32'h3b3e2496),
	.w6(32'h3c26ce40),
	.w7(32'h39e5961d),
	.w8(32'h3b03c81c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b564a53),
	.w1(32'hbb05e800),
	.w2(32'hbb8f1d80),
	.w3(32'h3bbb426f),
	.w4(32'hbb5758a5),
	.w5(32'h3b9f9265),
	.w6(32'h3aeb7c1c),
	.w7(32'hbb6dd40d),
	.w8(32'h3a7eb29e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fbfd),
	.w1(32'hbbce8ed9),
	.w2(32'hbad0dad3),
	.w3(32'h3b8bd03d),
	.w4(32'hbbb05d5a),
	.w5(32'h3ca3fcad),
	.w6(32'h3a06d132),
	.w7(32'hbbe01b1e),
	.w8(32'h3c395776),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5f5b),
	.w1(32'hbb64b7a6),
	.w2(32'h3bd47a6d),
	.w3(32'h3c482e27),
	.w4(32'hba8ed859),
	.w5(32'h3c2f19af),
	.w6(32'h3ba3895a),
	.w7(32'hbb494a0e),
	.w8(32'h3ba58720),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77a81e),
	.w1(32'hbb98ef6d),
	.w2(32'h3a30cdb5),
	.w3(32'h3b8129d9),
	.w4(32'hbb11634a),
	.w5(32'hbbb30c5c),
	.w6(32'h3bf88bd0),
	.w7(32'hbba7aabf),
	.w8(32'hbb5d9dbd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b498345),
	.w1(32'hba5ae509),
	.w2(32'h3b825dde),
	.w3(32'hbb5c27b0),
	.w4(32'hbb482018),
	.w5(32'h3ac21a1d),
	.w6(32'hbad258a0),
	.w7(32'hbb5e8c04),
	.w8(32'hbbf33d20),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc057e15),
	.w1(32'hbb3cbb49),
	.w2(32'hbb9e6ac6),
	.w3(32'hbbea3dc7),
	.w4(32'hbb8b0463),
	.w5(32'h39edf33e),
	.w6(32'hbb96134c),
	.w7(32'hbb71a7be),
	.w8(32'hbb99b7ec),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43caa),
	.w1(32'h3b6573cc),
	.w2(32'hb99a9641),
	.w3(32'hbb36713f),
	.w4(32'h3b60ce14),
	.w5(32'h3a021517),
	.w6(32'hbaa4c87f),
	.w7(32'h3baf0737),
	.w8(32'hbb4166d7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a08a),
	.w1(32'hbbd323bd),
	.w2(32'hbc15da75),
	.w3(32'h3c661d1f),
	.w4(32'hbb2ac21b),
	.w5(32'hbba21331),
	.w6(32'hbb33041b),
	.w7(32'hbb1646c9),
	.w8(32'hbbacecdb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d6dd),
	.w1(32'h3a892e83),
	.w2(32'h3bb27789),
	.w3(32'hbb939c5a),
	.w4(32'hb9b086b0),
	.w5(32'h3ace9452),
	.w6(32'hbbd2780d),
	.w7(32'hbaf398f0),
	.w8(32'h3b27cac1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af52118),
	.w1(32'hbb471fe8),
	.w2(32'h3993f6e6),
	.w3(32'h3bffd037),
	.w4(32'h3c10518f),
	.w5(32'hb93b1dcb),
	.w6(32'hbabef674),
	.w7(32'h3a6ff32c),
	.w8(32'h3add7424),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb42a),
	.w1(32'hbb849cc7),
	.w2(32'hbb19af78),
	.w3(32'hbc12025c),
	.w4(32'hbb3c808a),
	.w5(32'hbaaa290f),
	.w6(32'hbb6cca36),
	.w7(32'hbae7d5fa),
	.w8(32'h3becd9dd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c260628),
	.w1(32'hbab3e539),
	.w2(32'h38aa3d71),
	.w3(32'h3c45128f),
	.w4(32'hb98374a6),
	.w5(32'h3ba21216),
	.w6(32'h3c7cc70d),
	.w7(32'h3b2f09bb),
	.w8(32'h3bed6c49),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0bfdd),
	.w1(32'hba0e87e8),
	.w2(32'hbb71be86),
	.w3(32'h3b6143ec),
	.w4(32'h3b4afeec),
	.w5(32'hba8b7d45),
	.w6(32'h37de8ad2),
	.w7(32'h3b3b61e8),
	.w8(32'h3b1c518c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a0467),
	.w1(32'hbbaa150f),
	.w2(32'hba66c1f2),
	.w3(32'hbbdc6b3c),
	.w4(32'hbb894f60),
	.w5(32'h3bb68d2f),
	.w6(32'hbb272210),
	.w7(32'h3ae7966d),
	.w8(32'hba2ad812),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825d4f),
	.w1(32'hbb6b78d2),
	.w2(32'h3a0a49b2),
	.w3(32'hbbeab84e),
	.w4(32'hbc19ed23),
	.w5(32'h3bcf305e),
	.w6(32'hbba6d6a8),
	.w7(32'hbaf902d4),
	.w8(32'h3898b69f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc080d),
	.w1(32'hbb330f96),
	.w2(32'hbc112c87),
	.w3(32'hbbc55b5e),
	.w4(32'hbb5ea461),
	.w5(32'hbc08c386),
	.w6(32'hbba82556),
	.w7(32'h3ab28ca6),
	.w8(32'hbbbb9c70),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cbde6),
	.w1(32'hbbd65536),
	.w2(32'h3c205723),
	.w3(32'h3c1ccbf3),
	.w4(32'hbc002827),
	.w5(32'h3c76ab3c),
	.w6(32'h3bd132fe),
	.w7(32'h3ba389e5),
	.w8(32'h3c64f1d0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46b46c),
	.w1(32'h37e1c7a1),
	.w2(32'hbbb15c79),
	.w3(32'h3d1e79c6),
	.w4(32'h3b40750f),
	.w5(32'hbb90b615),
	.w6(32'h3ca58251),
	.w7(32'hbb90e650),
	.w8(32'hbba9015c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82a2d1),
	.w1(32'hbad41775),
	.w2(32'h3a6b7241),
	.w3(32'hbbfa7ee8),
	.w4(32'h398f139a),
	.w5(32'h3bc22aa8),
	.w6(32'hbc0eb444),
	.w7(32'h3ba5792f),
	.w8(32'hbaebd9cd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98145b),
	.w1(32'hbb1af2cd),
	.w2(32'hbb4f7b08),
	.w3(32'h3b13f364),
	.w4(32'hbaaeccc3),
	.w5(32'h3a4f0548),
	.w6(32'hbb35baec),
	.w7(32'hbb82eb67),
	.w8(32'h3a854049),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39feb125),
	.w1(32'hbb978754),
	.w2(32'hbb438cdf),
	.w3(32'hba432a85),
	.w4(32'hbbc06e38),
	.w5(32'h3b523686),
	.w6(32'h3afc27f1),
	.w7(32'hbb973bd9),
	.w8(32'hba9a013e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5244cf),
	.w1(32'hbbc2f0cd),
	.w2(32'h3b16ed82),
	.w3(32'h3bbe1e92),
	.w4(32'hbb1cfaab),
	.w5(32'h3b928546),
	.w6(32'hbb002d59),
	.w7(32'h3927b4c9),
	.w8(32'h3ba1007d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45494e),
	.w1(32'hbb4bdc59),
	.w2(32'h3a2af72c),
	.w3(32'hbb82eed3),
	.w4(32'h3b885020),
	.w5(32'h3c52b24f),
	.w6(32'hbae31f45),
	.w7(32'h3c1f181c),
	.w8(32'h3b0b530d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d990),
	.w1(32'hbbcc0e1a),
	.w2(32'h3b704b08),
	.w3(32'hbb76ea04),
	.w4(32'hbb2682ea),
	.w5(32'h3c33655f),
	.w6(32'hbc28e1c7),
	.w7(32'h3b2753a6),
	.w8(32'h3b92ee9e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f472),
	.w1(32'h3c2497a9),
	.w2(32'h3b9249a4),
	.w3(32'h3c03ec90),
	.w4(32'h3c1f97d6),
	.w5(32'hbac2922c),
	.w6(32'h3bb95a0e),
	.w7(32'h3a180701),
	.w8(32'h3add093b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6307cc),
	.w1(32'h3b87b937),
	.w2(32'h3bb844ca),
	.w3(32'hba8afc7b),
	.w4(32'h3bc91dd4),
	.w5(32'h3c46eb86),
	.w6(32'hbb760a4c),
	.w7(32'hbb9003d1),
	.w8(32'h3b32c558),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f55d),
	.w1(32'hbbac22b2),
	.w2(32'h3b1af689),
	.w3(32'h3ba315cf),
	.w4(32'hbb163ddf),
	.w5(32'h3c163a7b),
	.w6(32'h3ab89877),
	.w7(32'h3adc4b09),
	.w8(32'h3abb7e9a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdc4e0),
	.w1(32'hb9f2fe08),
	.w2(32'hbbe31667),
	.w3(32'h3bf8721e),
	.w4(32'h3b2fb0f0),
	.w5(32'hbba26420),
	.w6(32'hba1cd2e1),
	.w7(32'h3b33e20b),
	.w8(32'hbb3e81a3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06fdb3),
	.w1(32'hbad5abcc),
	.w2(32'hbbf2bc2c),
	.w3(32'hbbe4618c),
	.w4(32'hbba39fe8),
	.w5(32'hb9e7c133),
	.w6(32'hbba6b563),
	.w7(32'h3b83d090),
	.w8(32'hbb1a6f76),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b62b1),
	.w1(32'h3b50803b),
	.w2(32'hbbc1fbf7),
	.w3(32'h3a284169),
	.w4(32'hbbebdf36),
	.w5(32'h3a47a36d),
	.w6(32'hbc543012),
	.w7(32'hba84058c),
	.w8(32'hbb67b52b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ade0c),
	.w1(32'h3adb853c),
	.w2(32'h3ab7d25d),
	.w3(32'h38dc8b94),
	.w4(32'hbaf83183),
	.w5(32'h3b9c5515),
	.w6(32'hbbb5f248),
	.w7(32'hb9d4257c),
	.w8(32'h3c0f4f1b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6df72),
	.w1(32'h399b20a8),
	.w2(32'hbbf8ff11),
	.w3(32'hb96429b9),
	.w4(32'hbb69eb43),
	.w5(32'hbc5e4767),
	.w6(32'hbba171af),
	.w7(32'hbb98a336),
	.w8(32'hbba57906),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb524f38),
	.w1(32'h3a92254d),
	.w2(32'hbbea8300),
	.w3(32'hbbc7bab2),
	.w4(32'h3a658ad3),
	.w5(32'hbb65feb5),
	.w6(32'h3bd21f77),
	.w7(32'hba612781),
	.w8(32'h3b32befe),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3f3e2),
	.w1(32'h38ad7f2c),
	.w2(32'hb841c928),
	.w3(32'h38c23a75),
	.w4(32'h3c1ea3b4),
	.w5(32'h3c15336f),
	.w6(32'h3a8914b2),
	.w7(32'h3c15e217),
	.w8(32'hba4557d4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1fa17),
	.w1(32'hbbb318d1),
	.w2(32'hb842dcd4),
	.w3(32'hbaadd3b8),
	.w4(32'hbb982720),
	.w5(32'hba63a490),
	.w6(32'h3a8668d7),
	.w7(32'hbb059ad4),
	.w8(32'h3c0571b5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae00bf),
	.w1(32'hbbd1a583),
	.w2(32'hbb2d8924),
	.w3(32'hbbbec839),
	.w4(32'hbc62337e),
	.w5(32'hbaa9cf97),
	.w6(32'h3bbb42e0),
	.w7(32'hbb310017),
	.w8(32'h3c26c37e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b9144),
	.w1(32'hbb011c94),
	.w2(32'hbb75cff0),
	.w3(32'h3be57cf4),
	.w4(32'hbb913899),
	.w5(32'hbb1ea06a),
	.w6(32'h3b841feb),
	.w7(32'h3ae6f8ef),
	.w8(32'hbc099d5c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f50b6),
	.w1(32'hbb4b1c0a),
	.w2(32'h3b6113a6),
	.w3(32'hbb0c2234),
	.w4(32'hbb40cc28),
	.w5(32'h3b469b36),
	.w6(32'hbbaf3a08),
	.w7(32'hbb7a4b31),
	.w8(32'h3b98a88c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28fdd),
	.w1(32'h3bb5ad3b),
	.w2(32'h3bf11f60),
	.w3(32'h3b432e8d),
	.w4(32'h3b76c8a1),
	.w5(32'h3a827d93),
	.w6(32'hbb175677),
	.w7(32'h3b4dbd9c),
	.w8(32'h3b617945),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd78bf),
	.w1(32'hbbbcfaab),
	.w2(32'hbbdaff5f),
	.w3(32'h3bfe32fb),
	.w4(32'h3b1483a7),
	.w5(32'h3c165368),
	.w6(32'h3acbdd2a),
	.w7(32'h3c2df5ed),
	.w8(32'hbbddaf21),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf560e8),
	.w1(32'hba4fe3e1),
	.w2(32'hb623ef63),
	.w3(32'hbbbc958c),
	.w4(32'h3b261f5b),
	.w5(32'h3ac38f15),
	.w6(32'hbc5ab472),
	.w7(32'h3a29c659),
	.w8(32'hba9aba2d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9615a5),
	.w1(32'hbb09351a),
	.w2(32'hbc04e40f),
	.w3(32'hbc20cb5b),
	.w4(32'h3ab70eb8),
	.w5(32'hbc19f417),
	.w6(32'hbbc89d02),
	.w7(32'hb95c7331),
	.w8(32'hbbf52b59),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3dbab),
	.w1(32'hba24e53a),
	.w2(32'hbb4e1d48),
	.w3(32'hbbc3d837),
	.w4(32'hb6d11ec9),
	.w5(32'hbb5ad7ce),
	.w6(32'hbab62cc9),
	.w7(32'hba05a14e),
	.w8(32'hbb865c68),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9fd2),
	.w1(32'hbbbb7636),
	.w2(32'hbb6aad1c),
	.w3(32'hbbc4865c),
	.w4(32'hbbe5e249),
	.w5(32'h3a9886f6),
	.w6(32'h3a8d6f9b),
	.w7(32'hb8cd59e6),
	.w8(32'h3b23a552),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b34d),
	.w1(32'h39d9ee45),
	.w2(32'hbb829781),
	.w3(32'hbbe155b7),
	.w4(32'hbb83142c),
	.w5(32'hbc95ecba),
	.w6(32'h39809be9),
	.w7(32'hbc0fbc91),
	.w8(32'hbbe3d003),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30236),
	.w1(32'hbc46b3a9),
	.w2(32'h3ba213b5),
	.w3(32'hbc4bbeab),
	.w4(32'hbb927e6f),
	.w5(32'h3c029063),
	.w6(32'hbbddae39),
	.w7(32'hbb2c1312),
	.w8(32'hbbdebbf0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0785fa),
	.w1(32'hbb9483bc),
	.w2(32'hbc0ba1a4),
	.w3(32'hbbb520c2),
	.w4(32'hbb2bc8e1),
	.w5(32'hbb8e6c56),
	.w6(32'hbbe051b3),
	.w7(32'hbb97f26c),
	.w8(32'hbc063cb3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b8ef),
	.w1(32'hbbb42cda),
	.w2(32'hbc1218c1),
	.w3(32'h3ae4fa03),
	.w4(32'hbbff3cb3),
	.w5(32'h394a03de),
	.w6(32'hbad388c8),
	.w7(32'hbbb6a0b9),
	.w8(32'h3b80d93e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ce1b6),
	.w1(32'h3add5d65),
	.w2(32'h3b6f60cf),
	.w3(32'h3b0b77a1),
	.w4(32'hb8cee6f6),
	.w5(32'h3b3f5897),
	.w6(32'h3b1298df),
	.w7(32'h3a868614),
	.w8(32'h3b55eed9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ea013),
	.w1(32'h3b265219),
	.w2(32'h3ba1bb35),
	.w3(32'hbb18e793),
	.w4(32'hbb8ab702),
	.w5(32'h3ba985c4),
	.w6(32'hbbd224d8),
	.w7(32'h3b16a27e),
	.w8(32'hba1426ad),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5843d),
	.w1(32'hbbc1b49a),
	.w2(32'hbc0b3e71),
	.w3(32'hbbde2e8a),
	.w4(32'hbbf4dd4c),
	.w5(32'h3a473f80),
	.w6(32'hbb8ece64),
	.w7(32'hbb8ee1e9),
	.w8(32'hbb18db2a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17881a),
	.w1(32'hbaf52b64),
	.w2(32'hbbb31581),
	.w3(32'hbb9ed903),
	.w4(32'hbb3066f1),
	.w5(32'hbc0062fa),
	.w6(32'hb9c194a5),
	.w7(32'hbbc1c5dc),
	.w8(32'h3a2de5ba),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d833),
	.w1(32'h3af0aad5),
	.w2(32'hbba70982),
	.w3(32'hbb504945),
	.w4(32'hbb794947),
	.w5(32'hbaf73d2b),
	.w6(32'hbb05899f),
	.w7(32'hbb865e88),
	.w8(32'hbc16a24d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea481b),
	.w1(32'hbbbebbcd),
	.w2(32'h3b7d72b1),
	.w3(32'hbb5b4a4b),
	.w4(32'hbc16f783),
	.w5(32'h3b254f6f),
	.w6(32'hbb957a56),
	.w7(32'hbb944aae),
	.w8(32'h3b8b57fe),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1538b4),
	.w1(32'hbb5b918f),
	.w2(32'h3b3588db),
	.w3(32'h3c39466d),
	.w4(32'hbb9af97e),
	.w5(32'h3c16548c),
	.w6(32'h3b951c1c),
	.w7(32'h3b3ad3e2),
	.w8(32'h3c2d9287),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c7026),
	.w1(32'h3aa0c115),
	.w2(32'hbbb3a9d8),
	.w3(32'h3bbf981b),
	.w4(32'hbae395d1),
	.w5(32'h3bf0482f),
	.w6(32'h3ba7fc32),
	.w7(32'h3a2ee7b6),
	.w8(32'h3caa7e03),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8cdb7),
	.w1(32'hbb5a21bf),
	.w2(32'hbba9d9e7),
	.w3(32'h3cdff30c),
	.w4(32'hba8a5e88),
	.w5(32'h398ec463),
	.w6(32'h3c26e9cb),
	.w7(32'hbb2856b1),
	.w8(32'hba36dcd0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b7bf1),
	.w1(32'h3ab6f189),
	.w2(32'h3b73e5e8),
	.w3(32'hb99f9e29),
	.w4(32'h3b4c9346),
	.w5(32'h3c078197),
	.w6(32'h3a4d5d7f),
	.w7(32'h3bbb932b),
	.w8(32'h3bbcf3cc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc37b8e),
	.w1(32'hbae81e44),
	.w2(32'h39aa8117),
	.w3(32'h3c0c27ec),
	.w4(32'h3ba708eb),
	.w5(32'h3c4f7ef9),
	.w6(32'h3beefa0e),
	.w7(32'h3bc5b9c3),
	.w8(32'h3b04e40b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf52942),
	.w1(32'hbb82a225),
	.w2(32'hba79cc75),
	.w3(32'hbb8f664a),
	.w4(32'hbb701fb8),
	.w5(32'h3b5812f9),
	.w6(32'hbb68cc40),
	.w7(32'hba81d048),
	.w8(32'h3b6eca4a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba765b8d),
	.w1(32'h3ac13fae),
	.w2(32'h3bc04206),
	.w3(32'h3ae1ba06),
	.w4(32'hb859481f),
	.w5(32'h3b2ec17b),
	.w6(32'h3b1035a8),
	.w7(32'h3a831575),
	.w8(32'hb9a3c45a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88111a),
	.w1(32'h3b42c0d5),
	.w2(32'h3b8bd68a),
	.w3(32'hbb9ae461),
	.w4(32'h3bf4cea4),
	.w5(32'h3b174679),
	.w6(32'hbbb2f32d),
	.w7(32'h39edd7a8),
	.w8(32'hbba8cfc2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56d2c2),
	.w1(32'h3c095177),
	.w2(32'h383e5b89),
	.w3(32'hbb2f9d9f),
	.w4(32'h3c24d05a),
	.w5(32'h3c1edb17),
	.w6(32'hb98d7077),
	.w7(32'h3bbc0fab),
	.w8(32'h3c1685b9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbea3b8),
	.w1(32'hbaffdcd3),
	.w2(32'hbab552f6),
	.w3(32'hbad93de0),
	.w4(32'hbbb66d0b),
	.w5(32'hbc33c46a),
	.w6(32'hbad189ab),
	.w7(32'hbb7f993a),
	.w8(32'hbb4769e6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e39f8),
	.w1(32'h3a55e2f3),
	.w2(32'h3a8219dd),
	.w3(32'h3b655f76),
	.w4(32'hbb088954),
	.w5(32'h3bb9c900),
	.w6(32'h3bcfd330),
	.w7(32'hba6735b6),
	.w8(32'h3abd2eb1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a637499),
	.w1(32'hbc177239),
	.w2(32'h3a3eed75),
	.w3(32'hbb819b27),
	.w4(32'hb9b09f1e),
	.w5(32'h3c1468cb),
	.w6(32'hbb7ac194),
	.w7(32'hbbbfa0c8),
	.w8(32'h3b3db6a6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d8236),
	.w1(32'h3c337c78),
	.w2(32'hba0b8dc1),
	.w3(32'hbbab6e44),
	.w4(32'h3be82c3b),
	.w5(32'hbb4ebdf5),
	.w6(32'hb9b97216),
	.w7(32'hb91f63c0),
	.w8(32'hb74d0060),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60649),
	.w1(32'hbb54bd0c),
	.w2(32'h3abe1051),
	.w3(32'hbb7d5634),
	.w4(32'h3b15d294),
	.w5(32'hbb2fce5c),
	.w6(32'hba1eacaa),
	.w7(32'hbab93535),
	.w8(32'hbb9be1b6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d62d),
	.w1(32'h3b519df1),
	.w2(32'hbc223946),
	.w3(32'hbc276c6c),
	.w4(32'h3c28b195),
	.w5(32'hbbba12ce),
	.w6(32'hbc1092a3),
	.w7(32'hbb52d75b),
	.w8(32'hbb0fe854),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9195b78),
	.w1(32'hb934117d),
	.w2(32'hbbca029b),
	.w3(32'hbbc53118),
	.w4(32'hbacbf6da),
	.w5(32'hbbb7db90),
	.w6(32'hbbec1168),
	.w7(32'h3a283cbe),
	.w8(32'hbb98d9ca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010060),
	.w1(32'h3badb6b7),
	.w2(32'h3bcc873b),
	.w3(32'hbc1810af),
	.w4(32'hba0b02ec),
	.w5(32'hbab2b1c6),
	.w6(32'hbc023d78),
	.w7(32'hbbc736b5),
	.w8(32'h3afc5709),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f8563),
	.w1(32'h3ae7597a),
	.w2(32'h3b2a8dbf),
	.w3(32'hbbb95e4e),
	.w4(32'h3bed8162),
	.w5(32'hbbef90d9),
	.w6(32'hbabeb4c0),
	.w7(32'h3a9a4d8d),
	.w8(32'hbbc516a2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade7ffe),
	.w1(32'hbb508dae),
	.w2(32'hbc10c4c2),
	.w3(32'h3bc9ea4a),
	.w4(32'h3b66d4db),
	.w5(32'h3a94cfdc),
	.w6(32'h3b8a898b),
	.w7(32'h3c199190),
	.w8(32'hbb8a09b5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6a98d),
	.w1(32'h3b318637),
	.w2(32'h3c6c38b8),
	.w3(32'h3b97e163),
	.w4(32'h3a0603ba),
	.w5(32'h3c41544d),
	.w6(32'h3c00afd7),
	.w7(32'h3b371683),
	.w8(32'h3c860d79),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc992de),
	.w1(32'h399cf96f),
	.w2(32'h3a90503d),
	.w3(32'h3cfe17de),
	.w4(32'hbadaab2d),
	.w5(32'hbba1e8e8),
	.w6(32'h3c95fddf),
	.w7(32'hbb6e94f8),
	.w8(32'hbb720c7c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ed50c),
	.w1(32'h3ab1fe8c),
	.w2(32'hbbb0ac24),
	.w3(32'hbb9c7ad9),
	.w4(32'h3b7337f0),
	.w5(32'hbc210975),
	.w6(32'hbbb577b2),
	.w7(32'h3b0a26f5),
	.w8(32'hbb1542cd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a3ac9),
	.w1(32'h3c354953),
	.w2(32'hbbbe5883),
	.w3(32'h3bf2656d),
	.w4(32'hba40664e),
	.w5(32'hbbec2869),
	.w6(32'h3ba45459),
	.w7(32'h3b050c5b),
	.w8(32'hbbff26e3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fe7d2),
	.w1(32'h3bd23152),
	.w2(32'h3c19cdbc),
	.w3(32'hbc18a149),
	.w4(32'h3bb64e77),
	.w5(32'h3bd67a43),
	.w6(32'hbc3b5892),
	.w7(32'h3b10fd49),
	.w8(32'h3be443b2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908ef77),
	.w1(32'hbbc02ad7),
	.w2(32'hbc2cafe1),
	.w3(32'h3b491112),
	.w4(32'hbb3b026f),
	.w5(32'h3bb162f3),
	.w6(32'h39df4471),
	.w7(32'h3aacc8a9),
	.w8(32'h3699ac45),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379529a3),
	.w1(32'hbb0bd8a3),
	.w2(32'hbb2cc7ea),
	.w3(32'h3c7bf7c7),
	.w4(32'hbbad6f6c),
	.w5(32'h3c802fc0),
	.w6(32'h3c05e4c0),
	.w7(32'h3b88b676),
	.w8(32'h3c296b8a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1127a5),
	.w1(32'hbba414a2),
	.w2(32'hbb07e436),
	.w3(32'h3c7b1a29),
	.w4(32'hbb642c50),
	.w5(32'h3b9820d0),
	.w6(32'hbb11fc91),
	.w7(32'hbba3d6a9),
	.w8(32'h3c73b494),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba279cb9),
	.w1(32'hbb01d978),
	.w2(32'hbb7a88c4),
	.w3(32'h3c597524),
	.w4(32'hbb4a763b),
	.w5(32'hbc55100d),
	.w6(32'h3c0793f7),
	.w7(32'h394ce112),
	.w8(32'hbb83dc40),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcbd4e),
	.w1(32'hbad040eb),
	.w2(32'hbbd8cd0c),
	.w3(32'h3bad84bd),
	.w4(32'hbb3885d9),
	.w5(32'h3a2d9349),
	.w6(32'h3c04ef40),
	.w7(32'hbaa53504),
	.w8(32'hbbdb9ad6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55daaf),
	.w1(32'hbaf18f69),
	.w2(32'h3be935c4),
	.w3(32'hbb88df22),
	.w4(32'hbadd849e),
	.w5(32'h3c78b245),
	.w6(32'hbbb73344),
	.w7(32'hbb16ca00),
	.w8(32'h3c465bb4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab71f3e),
	.w1(32'h3a28ee05),
	.w2(32'h39e97e88),
	.w3(32'hb9ae3c25),
	.w4(32'hbb41bab2),
	.w5(32'h371ca525),
	.w6(32'hbb4f8781),
	.w7(32'h3b33f552),
	.w8(32'h3ae574c8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9bee2),
	.w1(32'h3b525a38),
	.w2(32'h3c15fb81),
	.w3(32'hbbf68e9a),
	.w4(32'h3a5782d1),
	.w5(32'h3c477830),
	.w6(32'hbc090c84),
	.w7(32'hbb41eed5),
	.w8(32'h3bc974ff),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f41a4),
	.w1(32'hbbc1b59d),
	.w2(32'hbc12b318),
	.w3(32'h3c2ddd2a),
	.w4(32'hbb9f5583),
	.w5(32'hbc4ac612),
	.w6(32'h3be2a066),
	.w7(32'hbb965389),
	.w8(32'hbbe1d787),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9070),
	.w1(32'hbb5fbf12),
	.w2(32'hbb4113bc),
	.w3(32'h3b0f4995),
	.w4(32'hbbdc3957),
	.w5(32'h396f45c8),
	.w6(32'h3b32bfa4),
	.w7(32'hbb20e9b6),
	.w8(32'hb9278370),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0131b6),
	.w1(32'h3baa8514),
	.w2(32'h3b36f415),
	.w3(32'h3b5ffc3b),
	.w4(32'h3bca723e),
	.w5(32'h3c2c2ee3),
	.w6(32'h3a75383d),
	.w7(32'h3c16c294),
	.w8(32'h3c2e16af),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe91bb),
	.w1(32'hbaaa584a),
	.w2(32'hba70e79e),
	.w3(32'hbbd7bb58),
	.w4(32'hbb1a3cdb),
	.w5(32'h3b068415),
	.w6(32'hbad9e190),
	.w7(32'h3ad4062f),
	.w8(32'hbb0f551a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe83c27),
	.w1(32'h3c75094e),
	.w2(32'h3c539b60),
	.w3(32'hba95fdff),
	.w4(32'h3c3ce2e3),
	.w5(32'h3c64f3a9),
	.w6(32'hb9ddfe76),
	.w7(32'h3be5b6f6),
	.w8(32'h3c917dc2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06bb83),
	.w1(32'h3ae2a324),
	.w2(32'hbb36577b),
	.w3(32'h3c6476e0),
	.w4(32'h3a4b59b7),
	.w5(32'hbb134ad3),
	.w6(32'h3bb14bd5),
	.w7(32'hbb58df12),
	.w8(32'hbabc68c8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09e1d),
	.w1(32'h3b91c60a),
	.w2(32'hbba18f13),
	.w3(32'hbb77ecd6),
	.w4(32'h3b936115),
	.w5(32'h3b1bfeed),
	.w6(32'h3a28dfda),
	.w7(32'h39c53e60),
	.w8(32'hbb83aa35),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad54b7),
	.w1(32'hbbf8c3e3),
	.w2(32'h398fbebc),
	.w3(32'hbc319d38),
	.w4(32'hbbe0bc48),
	.w5(32'h3bc9dbaa),
	.w6(32'hbbf8db9b),
	.w7(32'hbb953939),
	.w8(32'h3b2c6365),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c41a5a),
	.w1(32'hbc3123ac),
	.w2(32'hbbf80c1a),
	.w3(32'h3a308de7),
	.w4(32'hbc1381f0),
	.w5(32'hbc911644),
	.w6(32'hbc0a3036),
	.w7(32'hbbfefb95),
	.w8(32'hbbd63420),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba441c28),
	.w1(32'hbc194950),
	.w2(32'hbc499ae2),
	.w3(32'hba4def7f),
	.w4(32'hbbf15319),
	.w5(32'hbcf9ca30),
	.w6(32'h3bbf6638),
	.w7(32'hbb50686f),
	.w8(32'hbc498952),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3b413),
	.w1(32'hbb75c6a6),
	.w2(32'hbc16e4ea),
	.w3(32'h3bd23f45),
	.w4(32'hbc2dd65a),
	.w5(32'hbc014b65),
	.w6(32'h3bda3f47),
	.w7(32'hbb1678d2),
	.w8(32'hbc0783e6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf563a3),
	.w1(32'hbbb5d55e),
	.w2(32'hbc7e9ddb),
	.w3(32'hbc2baabb),
	.w4(32'hbbd0ad95),
	.w5(32'hbbf7bd36),
	.w6(32'hbc520fef),
	.w7(32'hbb8790d9),
	.w8(32'hbbd510a3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b509716),
	.w1(32'hba18415a),
	.w2(32'hbb783c82),
	.w3(32'h3a35bb8b),
	.w4(32'hbb86a98f),
	.w5(32'hbc68e3eb),
	.w6(32'hbb8672a3),
	.w7(32'h3a7164be),
	.w8(32'hbbf5811c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917990),
	.w1(32'hbb2cba77),
	.w2(32'h398cbd48),
	.w3(32'h3badbb96),
	.w4(32'hbb278533),
	.w5(32'hba26a53e),
	.w6(32'h3bdda5d9),
	.w7(32'hbb029319),
	.w8(32'h3a95bd82),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063f99),
	.w1(32'h3b6ab994),
	.w2(32'h3c868c07),
	.w3(32'h3bce853c),
	.w4(32'h3a276345),
	.w5(32'h3cd26ef1),
	.w6(32'h3a32d2cd),
	.w7(32'hbb83ff42),
	.w8(32'h3c924cc0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6860f1),
	.w1(32'hbc1cb613),
	.w2(32'hba9b35a4),
	.w3(32'h3cae9275),
	.w4(32'hbc19ec21),
	.w5(32'h3b8b3522),
	.w6(32'h3cbcdca3),
	.w7(32'hbb12f97b),
	.w8(32'h3ba7cec7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9ca3),
	.w1(32'hb6cf5e09),
	.w2(32'hbb88e310),
	.w3(32'hbbf38c75),
	.w4(32'h395f1541),
	.w5(32'h3a7857a6),
	.w6(32'h3b1557b4),
	.w7(32'hbb5de4d1),
	.w8(32'hbbd05a08),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe678dc),
	.w1(32'h3acfc294),
	.w2(32'hba75c440),
	.w3(32'hbc279d0f),
	.w4(32'h3957430c),
	.w5(32'hbb18c6a8),
	.w6(32'hbc19b15e),
	.w7(32'hb99e50e1),
	.w8(32'hbaff0f3e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46d95f),
	.w1(32'hbbbd0916),
	.w2(32'h3b173587),
	.w3(32'hbbbb5280),
	.w4(32'hbb0b4e45),
	.w5(32'h3c839fd7),
	.w6(32'hbbc7a181),
	.w7(32'h3966b9bd),
	.w8(32'hbafd231f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9967a),
	.w1(32'hbbb980db),
	.w2(32'hbb8be974),
	.w3(32'hbbd448c7),
	.w4(32'h3b1176b9),
	.w5(32'hba282e5a),
	.w6(32'h395cb8b2),
	.w7(32'hbb73a78d),
	.w8(32'hbbef7c9f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0829f),
	.w1(32'h3b2343d9),
	.w2(32'h3aab3cd6),
	.w3(32'hbb850f80),
	.w4(32'h3b9496f7),
	.w5(32'h3c28965f),
	.w6(32'h3b6725b5),
	.w7(32'hbaa254fa),
	.w8(32'hbaf37374),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf219a),
	.w1(32'h3a729e5f),
	.w2(32'h3b7978af),
	.w3(32'h3cb9d43d),
	.w4(32'hbb22bbbf),
	.w5(32'h3bd8d573),
	.w6(32'h3c1f8ad7),
	.w7(32'hbb4a0d66),
	.w8(32'h3bb1f132),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c052462),
	.w1(32'h3b28acad),
	.w2(32'h3c122eed),
	.w3(32'h3c39cfef),
	.w4(32'h3b85f89a),
	.w5(32'h3b27677a),
	.w6(32'h3c2abfac),
	.w7(32'hbb352000),
	.w8(32'h378a1c96),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14dc2f),
	.w1(32'hb94b8bc7),
	.w2(32'h3adabeed),
	.w3(32'hbc7399b8),
	.w4(32'h3bda1580),
	.w5(32'h3c6e75dd),
	.w6(32'hbc5c1ada),
	.w7(32'h3c3fc9e3),
	.w8(32'h3bb37095),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb303f04),
	.w1(32'hbbd597c2),
	.w2(32'h3b06baf0),
	.w3(32'hba355646),
	.w4(32'hbb8f625b),
	.w5(32'hbb078c18),
	.w6(32'hbb5d5a5d),
	.w7(32'hbb3a65d9),
	.w8(32'h3a9d6d2e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176961),
	.w1(32'hbb4137c0),
	.w2(32'hbb233747),
	.w3(32'h3b343ae3),
	.w4(32'hba163ecb),
	.w5(32'h39265fbe),
	.w6(32'h3aee5d62),
	.w7(32'hba57354e),
	.w8(32'hb9a41da1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66ace1),
	.w1(32'h3b6beaed),
	.w2(32'h39319e35),
	.w3(32'hbaab36cb),
	.w4(32'h39c82fc4),
	.w5(32'h3b88f729),
	.w6(32'h3b4cf7f7),
	.w7(32'h3b1bd75d),
	.w8(32'h3bb5e8a0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3dd1a),
	.w1(32'hbba41ba7),
	.w2(32'hbbcb02bd),
	.w3(32'h3af4a259),
	.w4(32'hb99f3e1b),
	.w5(32'hbc17c1cf),
	.w6(32'hbae74929),
	.w7(32'hbb74df79),
	.w8(32'hba4a1d72),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab292f),
	.w1(32'h3a4e0bba),
	.w2(32'hbadb57f2),
	.w3(32'h3c9ef6a4),
	.w4(32'hbbe43a02),
	.w5(32'h3bdffee2),
	.w6(32'h3b9a10e9),
	.w7(32'hbbb16f26),
	.w8(32'h3bab1616),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9203bf),
	.w1(32'hb98baa09),
	.w2(32'hbaca78f9),
	.w3(32'h3abdb2af),
	.w4(32'hbb3446b5),
	.w5(32'hbb1413d8),
	.w6(32'hbbaf7aaf),
	.w7(32'hba8b7687),
	.w8(32'h3899b6fe),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58bca0),
	.w1(32'hbb6f1120),
	.w2(32'hbbc5ab88),
	.w3(32'h39a114f7),
	.w4(32'h3ba06fa5),
	.w5(32'h3c0faaf1),
	.w6(32'hb9ae99ef),
	.w7(32'hb9b6965e),
	.w8(32'hbb68c907),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba559c5d),
	.w1(32'h3aa996bb),
	.w2(32'h3a3a32a0),
	.w3(32'h3b0f8f5a),
	.w4(32'hbb3de2ea),
	.w5(32'hbb137d39),
	.w6(32'hbaa86278),
	.w7(32'hba60e350),
	.w8(32'hba903c5b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd9d22),
	.w1(32'hbaa55ba4),
	.w2(32'h3a22589d),
	.w3(32'hbae06be6),
	.w4(32'hbb01de15),
	.w5(32'hbb11ac13),
	.w6(32'h39ae33f3),
	.w7(32'hbc052a75),
	.w8(32'hbbcab8ac),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b602e),
	.w1(32'hbb29e17d),
	.w2(32'h3ad9d59a),
	.w3(32'hbb2a9466),
	.w4(32'h3aeb64c6),
	.w5(32'h3aaf75e4),
	.w6(32'hba56c676),
	.w7(32'hbb2738ee),
	.w8(32'hba8527a4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f326),
	.w1(32'hbc31978e),
	.w2(32'hbbc98759),
	.w3(32'hbb6f94f5),
	.w4(32'h3b8bb010),
	.w5(32'h3bec1f3f),
	.w6(32'hbae5e75a),
	.w7(32'hbb091000),
	.w8(32'hbb1b3ce3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96f592),
	.w1(32'h3b0cacfb),
	.w2(32'h3b80f920),
	.w3(32'h3ae1d454),
	.w4(32'h3b02e764),
	.w5(32'h3b5bf32f),
	.w6(32'hbb2b9e05),
	.w7(32'h3b174d5d),
	.w8(32'h3b9d046a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6c92e),
	.w1(32'hbab33ee2),
	.w2(32'hbb563bc1),
	.w3(32'h3ab86f38),
	.w4(32'h38ecef83),
	.w5(32'hbb28c09b),
	.w6(32'h3b049798),
	.w7(32'h39ad95bf),
	.w8(32'hba274e24),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb385d),
	.w1(32'h3b8ab21d),
	.w2(32'hba738c37),
	.w3(32'hbb487bd9),
	.w4(32'hbad23c5a),
	.w5(32'hbbc7de36),
	.w6(32'hbba3a566),
	.w7(32'h3bf51397),
	.w8(32'h3a80d4ad),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59e0fa),
	.w1(32'h3b76797c),
	.w2(32'hba2c8c58),
	.w3(32'hbbeeea2d),
	.w4(32'h3a7dbb57),
	.w5(32'hba8941e0),
	.w6(32'hbbb1ed4f),
	.w7(32'hb8accb9e),
	.w8(32'hba65376a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b19bc),
	.w1(32'hbbf2b258),
	.w2(32'hbc2c1f19),
	.w3(32'h3b13c4f5),
	.w4(32'hbb9945ce),
	.w5(32'hba281c96),
	.w6(32'hbaf73e5d),
	.w7(32'hbb2f2564),
	.w8(32'h3a347230),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349d35),
	.w1(32'hbaa5e5e0),
	.w2(32'h3b07200d),
	.w3(32'hbb1b961a),
	.w4(32'hbbf647df),
	.w5(32'hbba33c16),
	.w6(32'h3a085129),
	.w7(32'h3b2bdf05),
	.w8(32'h3a5ef337),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab04910),
	.w1(32'h3b2a5f86),
	.w2(32'h3b32855b),
	.w3(32'hb9ba1c67),
	.w4(32'h3ad16469),
	.w5(32'h3aa3c77e),
	.w6(32'h3b1bb0c5),
	.w7(32'h3ae3c66e),
	.w8(32'h3b32ee86),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50ca94),
	.w1(32'h3b6f9fd3),
	.w2(32'hbac8a9f3),
	.w3(32'h3b5c2b91),
	.w4(32'h3b9182e4),
	.w5(32'h3b5b4127),
	.w6(32'h3b8f4855),
	.w7(32'h3b6804c3),
	.w8(32'h3bda9fb0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6ad2e),
	.w1(32'h3bb823d3),
	.w2(32'h3b6b8f89),
	.w3(32'h3917ffaf),
	.w4(32'h3bcb9e03),
	.w5(32'h3ac52e50),
	.w6(32'h3c0a8097),
	.w7(32'h3b07e61b),
	.w8(32'hbbea1aa8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c7dbb),
	.w1(32'hbb6529e9),
	.w2(32'hbb7f5832),
	.w3(32'hbbc41098),
	.w4(32'hbb65d05f),
	.w5(32'hbb7be2df),
	.w6(32'hbb243496),
	.w7(32'hbb309174),
	.w8(32'hbc044829),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba376168),
	.w1(32'hbb5db32a),
	.w2(32'h3b8790bd),
	.w3(32'hbb783c78),
	.w4(32'h3ab425ee),
	.w5(32'hb904abc6),
	.w6(32'hbb9416a1),
	.w7(32'hbae014d1),
	.w8(32'hbb8c1b88),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34604f),
	.w1(32'hba517040),
	.w2(32'hbbd56889),
	.w3(32'hbb8a70d3),
	.w4(32'hb9490f79),
	.w5(32'h3a16377b),
	.w6(32'h3aa86315),
	.w7(32'hba6b68ad),
	.w8(32'hbb711033),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959a1d3),
	.w1(32'h3b67b9b3),
	.w2(32'h3a1334cb),
	.w3(32'h3b32aa45),
	.w4(32'h3c673b19),
	.w5(32'h3cbaac3a),
	.w6(32'hbb2b8da6),
	.w7(32'h3bed28d0),
	.w8(32'hbb296179),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad43819),
	.w1(32'hbb1c5621),
	.w2(32'hbb50aa48),
	.w3(32'h3b98bf00),
	.w4(32'h3be6788a),
	.w5(32'h3c96cb16),
	.w6(32'h3909e333),
	.w7(32'h3bd6f149),
	.w8(32'hbb9f5aaf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0f6f7),
	.w1(32'h3a7d5235),
	.w2(32'h3b44adc0),
	.w3(32'h3bce2fa1),
	.w4(32'hbbce765c),
	.w5(32'h3a905be0),
	.w6(32'hbb93e6fe),
	.w7(32'hbb3a8623),
	.w8(32'h393f38c6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9a485),
	.w1(32'h3994c84d),
	.w2(32'hba447068),
	.w3(32'h3b391bb0),
	.w4(32'hba1573ef),
	.w5(32'hbb9bb63e),
	.w6(32'hbad8e918),
	.w7(32'h3aaf38d0),
	.w8(32'hbb890731),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454ec2),
	.w1(32'hba9f55fa),
	.w2(32'hbad194ef),
	.w3(32'hbb8afbc2),
	.w4(32'h3bc50f49),
	.w5(32'hbba19345),
	.w6(32'hb8da9d99),
	.w7(32'h3a6c6cdb),
	.w8(32'hba9a4a05),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c585cc2),
	.w1(32'hba0758f3),
	.w2(32'hbb16758d),
	.w3(32'hbbc0edb9),
	.w4(32'hbb9f5f45),
	.w5(32'hbb013358),
	.w6(32'h39c66792),
	.w7(32'hbac73e8f),
	.w8(32'hbaa829cc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1ef8f),
	.w1(32'hbb3162c7),
	.w2(32'hb8e58a06),
	.w3(32'hba8b6c05),
	.w4(32'hba911b6a),
	.w5(32'hba8e5dae),
	.w6(32'h3b80edb6),
	.w7(32'h3a941150),
	.w8(32'h3952849e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d809),
	.w1(32'hbbc1124b),
	.w2(32'hbbc7aca4),
	.w3(32'hb9f48a82),
	.w4(32'h3c4e51ae),
	.w5(32'h3c938330),
	.w6(32'hb93ac9e7),
	.w7(32'hbb3c8b0c),
	.w8(32'hbb6c5d16),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc394d4),
	.w1(32'hbaf866cf),
	.w2(32'h3c03d7f5),
	.w3(32'h3c4da9c3),
	.w4(32'h3a85c162),
	.w5(32'h3aedec45),
	.w6(32'h39b69d23),
	.w7(32'hbb0279e0),
	.w8(32'hbbe9532e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b1a0),
	.w1(32'hbbb28fc0),
	.w2(32'hbb6b3d18),
	.w3(32'hbbc3018b),
	.w4(32'h3b703cf1),
	.w5(32'h3c4b3368),
	.w6(32'hbbb57ba5),
	.w7(32'hbb4765d6),
	.w8(32'hbbf3142e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae7e5f),
	.w1(32'hba33458d),
	.w2(32'h3b88422f),
	.w3(32'h3b49757e),
	.w4(32'hbb7e9fbf),
	.w5(32'h3ab63c50),
	.w6(32'hbb13a093),
	.w7(32'hbc0882a2),
	.w8(32'hba80ff09),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80469),
	.w1(32'h3aaa8afd),
	.w2(32'h3a65adab),
	.w3(32'hbb2c2e68),
	.w4(32'hba0ac99a),
	.w5(32'h3b95eb77),
	.w6(32'hbba3185d),
	.w7(32'hbb9f93c8),
	.w8(32'hbb840eb6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ffb17),
	.w1(32'hba5af994),
	.w2(32'hbb966126),
	.w3(32'h3a655993),
	.w4(32'hbb9f4327),
	.w5(32'hbb658608),
	.w6(32'hbba1bc63),
	.w7(32'hbab42aa9),
	.w8(32'h3b884f68),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad13ba4),
	.w1(32'hbb33bcd4),
	.w2(32'hbb542583),
	.w3(32'h3ad67fdf),
	.w4(32'h3b16f684),
	.w5(32'h3c22cb05),
	.w6(32'h3b6af848),
	.w7(32'hbb1d637d),
	.w8(32'h3a950658),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbec1),
	.w1(32'hbad4722a),
	.w2(32'h3b213f54),
	.w3(32'h3b5644da),
	.w4(32'hbadb191f),
	.w5(32'hbb8a3b73),
	.w6(32'hbb59ecf8),
	.w7(32'hba279364),
	.w8(32'hbb96b636),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9050),
	.w1(32'h3b953bfd),
	.w2(32'h38861b04),
	.w3(32'hbbb344e6),
	.w4(32'h3bcacb1f),
	.w5(32'h3ca49f62),
	.w6(32'hbb33d4d1),
	.w7(32'h3bb88504),
	.w8(32'hba26b10e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73946),
	.w1(32'hbb076c26),
	.w2(32'hb96539e8),
	.w3(32'h3b34a5b4),
	.w4(32'hbb241abd),
	.w5(32'hbb274adf),
	.w6(32'h3b93b76f),
	.w7(32'hbbb5f646),
	.w8(32'hbb7af62c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3fc82),
	.w1(32'hbb5a97ac),
	.w2(32'hbb912111),
	.w3(32'h3a236710),
	.w4(32'h3b4ff6d0),
	.w5(32'h3c982f09),
	.w6(32'hbbd79c00),
	.w7(32'hbb353356),
	.w8(32'h3b0c0b82),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854056),
	.w1(32'h3a2a8f4e),
	.w2(32'hbb2e3dd5),
	.w3(32'h3b1b99d2),
	.w4(32'hbb3e4147),
	.w5(32'h3a475db3),
	.w6(32'hb9309bc0),
	.w7(32'h35c61bc5),
	.w8(32'h3b3a4a8c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe240c),
	.w1(32'h3bc836a2),
	.w2(32'h3b74abe1),
	.w3(32'h3b532630),
	.w4(32'h3b2413f0),
	.w5(32'h3a87d0a7),
	.w6(32'h3b99adec),
	.w7(32'h3bbd63bd),
	.w8(32'h3a560631),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9966456),
	.w1(32'h3afabdf0),
	.w2(32'hb8fe7895),
	.w3(32'h39f6c449),
	.w4(32'hbb3bf2b5),
	.w5(32'hbad19413),
	.w6(32'hb98cf035),
	.w7(32'h3b2d1730),
	.w8(32'hb98d2419),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8de1ed),
	.w1(32'h3a48e3f1),
	.w2(32'h3b18321b),
	.w3(32'hb9ddd63e),
	.w4(32'hbb71d2b3),
	.w5(32'h3b122103),
	.w6(32'hbaf0bcdf),
	.w7(32'h37c93f5a),
	.w8(32'h3a1239f4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698f8a),
	.w1(32'hbc01dc0b),
	.w2(32'hbbcdd1f0),
	.w3(32'hbb96c9b5),
	.w4(32'hb9b81f29),
	.w5(32'h3bb3d6a7),
	.w6(32'h3b8b0642),
	.w7(32'hb9e23081),
	.w8(32'h3a102b6a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94bcbe),
	.w1(32'h3c63f6ef),
	.w2(32'h3c8acb8f),
	.w3(32'h383c2158),
	.w4(32'hbbe80d9e),
	.w5(32'hbb69fbf7),
	.w6(32'hbb74bded),
	.w7(32'hbba651ae),
	.w8(32'h3b1bb4c3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22d28f),
	.w1(32'hba837ec9),
	.w2(32'h3b342634),
	.w3(32'hbb7292a0),
	.w4(32'hbbd9a045),
	.w5(32'h3b212164),
	.w6(32'hbac95c2a),
	.w7(32'hbb5a479a),
	.w8(32'h3b8bd0a7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91aa3b),
	.w1(32'hbb79ff65),
	.w2(32'h3b280ed2),
	.w3(32'h3b6ce092),
	.w4(32'h3ac749a9),
	.w5(32'h3bff119a),
	.w6(32'h3b46ab7d),
	.w7(32'h3ad9342f),
	.w8(32'hbac8095b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48c17),
	.w1(32'h3bb499c0),
	.w2(32'h3c02794b),
	.w3(32'hbb437f11),
	.w4(32'hba261975),
	.w5(32'h3acfc195),
	.w6(32'hbadf4e9a),
	.w7(32'h3a875875),
	.w8(32'h3bbed7a9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b1d74),
	.w1(32'hbb4b06ce),
	.w2(32'hbbac3302),
	.w3(32'h39aa1b59),
	.w4(32'hbb248271),
	.w5(32'hbbb44700),
	.w6(32'hbae70a72),
	.w7(32'h3b1bb614),
	.w8(32'hb9d0a6bb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395707f3),
	.w1(32'h3b04bc21),
	.w2(32'hbb617dcd),
	.w3(32'h3b6ee230),
	.w4(32'hbb1a68be),
	.w5(32'hba21a216),
	.w6(32'hb85abe2f),
	.w7(32'hbb2cc781),
	.w8(32'hbb173d5e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37df2b),
	.w1(32'hbaf434cf),
	.w2(32'hb948efa0),
	.w3(32'h3a500e53),
	.w4(32'h3b000015),
	.w5(32'hbbc0d086),
	.w6(32'hbb04701a),
	.w7(32'h3b074cac),
	.w8(32'hbb41b762),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1c808),
	.w1(32'h3b37deee),
	.w2(32'hbabc9d5f),
	.w3(32'h39d3f578),
	.w4(32'hbb9a4793),
	.w5(32'hbafefbeb),
	.w6(32'h3ac535a6),
	.w7(32'hb8a0fe43),
	.w8(32'h3bca6b54),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6ece),
	.w1(32'hbac2df4f),
	.w2(32'h3b26a3f7),
	.w3(32'h39f9fb1b),
	.w4(32'hba27dc80),
	.w5(32'h3c0693c7),
	.w6(32'h3bebc50e),
	.w7(32'hbaac33b8),
	.w8(32'hbb5d21b9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d5390),
	.w1(32'h3aef2283),
	.w2(32'hbb237d05),
	.w3(32'hbbca2f4c),
	.w4(32'h38db5be7),
	.w5(32'hbb05046c),
	.w6(32'hbb86b964),
	.w7(32'hbba1caa3),
	.w8(32'hbb751e39),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2081bb),
	.w1(32'h39a4d767),
	.w2(32'hbb87ec8f),
	.w3(32'h3a58eb3d),
	.w4(32'hb96a0166),
	.w5(32'hba53fe07),
	.w6(32'h3a8369df),
	.w7(32'hba867acf),
	.w8(32'hbb965ffc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27b69d),
	.w1(32'hbba670e0),
	.w2(32'hbbff52ab),
	.w3(32'hba270ef2),
	.w4(32'hbb3e5a1a),
	.w5(32'hbbaa1509),
	.w6(32'hbb1a0464),
	.w7(32'h373c53fc),
	.w8(32'hba57ccfd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb5a4),
	.w1(32'hbb525619),
	.w2(32'hbb64d003),
	.w3(32'hbb0a5dc0),
	.w4(32'h3c147057),
	.w5(32'h3c830427),
	.w6(32'h3b239975),
	.w7(32'h3af26255),
	.w8(32'hbb81c529),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad2eed),
	.w1(32'hbb6c9e27),
	.w2(32'hba08450f),
	.w3(32'h3a21ca7e),
	.w4(32'hb92e8019),
	.w5(32'h3b276a22),
	.w6(32'h3ab8104f),
	.w7(32'h3ae76f8b),
	.w8(32'h3a7628f4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d256d),
	.w1(32'hbb275426),
	.w2(32'hbb0749c1),
	.w3(32'h3b0db555),
	.w4(32'hbc1b9d35),
	.w5(32'hbb472ffe),
	.w6(32'h3b8c893c),
	.w7(32'h3b849b82),
	.w8(32'h3b5dc318),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e05b),
	.w1(32'hbb079137),
	.w2(32'hbb7e08a8),
	.w3(32'hbb6ec7a5),
	.w4(32'hba19beb5),
	.w5(32'h3c0329bf),
	.w6(32'h3b9c1284),
	.w7(32'hbb87aad1),
	.w8(32'h3ab84ac2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44e9ea),
	.w1(32'h3a79ba23),
	.w2(32'hbbc924fd),
	.w3(32'h3a0505d2),
	.w4(32'hb9ff7647),
	.w5(32'h3be35115),
	.w6(32'h39fdf524),
	.w7(32'h3abba0ef),
	.w8(32'hbb67114c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafec111),
	.w1(32'hbb659dfe),
	.w2(32'h3b85913b),
	.w3(32'hbb22733a),
	.w4(32'h3c305595),
	.w5(32'h3bc5d5fb),
	.w6(32'hba66fd78),
	.w7(32'h3b077867),
	.w8(32'hbbb62a7c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule