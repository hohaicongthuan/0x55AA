module layer_8_featuremap_251(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88773),
	.w1(32'h3bbd2845),
	.w2(32'hbcdd011d),
	.w3(32'hbab3593a),
	.w4(32'h3c814178),
	.w5(32'hbd0ddc6e),
	.w6(32'h3ba73e8f),
	.w7(32'hbc6cfb5c),
	.w8(32'h3bb3af38),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8f633),
	.w1(32'h3b1d79a2),
	.w2(32'h3bbbf5e5),
	.w3(32'h3b64cf74),
	.w4(32'h3b6aec2c),
	.w5(32'h3b9e76d5),
	.w6(32'h3ae4c20a),
	.w7(32'h3b465bb0),
	.w8(32'h3b26616a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aedaa),
	.w1(32'h3c101a34),
	.w2(32'hbbd63ad7),
	.w3(32'h3b23c106),
	.w4(32'h3c61560f),
	.w5(32'hbc129eb6),
	.w6(32'h3c242dea),
	.w7(32'h3b8f9847),
	.w8(32'h3bc2a5f1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb32bc3),
	.w1(32'h3bd798fc),
	.w2(32'hbc459dbd),
	.w3(32'h3bfee09c),
	.w4(32'h3b8c6a85),
	.w5(32'hbc682f92),
	.w6(32'hbb539ff9),
	.w7(32'hba4e502c),
	.w8(32'hbbb2e281),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123857),
	.w1(32'hb7d26914),
	.w2(32'h3adfe2fd),
	.w3(32'h3bdd7a02),
	.w4(32'h3aba9add),
	.w5(32'h3bc34438),
	.w6(32'hbacfbb44),
	.w7(32'h3ac7884a),
	.w8(32'hbb11f522),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40c9a),
	.w1(32'h3add0a18),
	.w2(32'hbbc44d62),
	.w3(32'hbbbcf328),
	.w4(32'hbc37affe),
	.w5(32'hbb46a2ab),
	.w6(32'hbb00e2c5),
	.w7(32'h3a78d213),
	.w8(32'h3c3f2f15),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58f122),
	.w1(32'hb9b2b5aa),
	.w2(32'hbb90b1c9),
	.w3(32'h3c427464),
	.w4(32'hb8da0fcd),
	.w5(32'hbacba857),
	.w6(32'hbb6f7069),
	.w7(32'hbb550698),
	.w8(32'hbb99bb43),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e291b8),
	.w1(32'hbc1c8931),
	.w2(32'hbb774b05),
	.w3(32'hbb3c31e6),
	.w4(32'hbc5d3c4b),
	.w5(32'h3b580604),
	.w6(32'hbb83aed7),
	.w7(32'hbb9dce28),
	.w8(32'h3c8170f4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85cbc8),
	.w1(32'h3b4701d0),
	.w2(32'h3b576ac6),
	.w3(32'h3c846df5),
	.w4(32'h3b5c82de),
	.w5(32'h3c317c95),
	.w6(32'hba56446f),
	.w7(32'hba11a93e),
	.w8(32'hbbd25130),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357f20),
	.w1(32'h3bfbbdc8),
	.w2(32'hbb53427b),
	.w3(32'hbb18d9c2),
	.w4(32'h3bcf9681),
	.w5(32'h3a9472e8),
	.w6(32'h3c2a3d96),
	.w7(32'hbb24f1a1),
	.w8(32'h3acb1dfa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d943),
	.w1(32'h3adcc8d1),
	.w2(32'hbba59e05),
	.w3(32'h3b7a96eb),
	.w4(32'hbb32a530),
	.w5(32'hbc820ab9),
	.w6(32'hbb2e7988),
	.w7(32'hbacc4c4e),
	.w8(32'hbb5842f0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd448),
	.w1(32'h3a42e40d),
	.w2(32'h3c252759),
	.w3(32'hb9525daa),
	.w4(32'hbb565183),
	.w5(32'h3c0b7228),
	.w6(32'hbb09a25e),
	.w7(32'h3c272ae4),
	.w8(32'hbb8b56a0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf892),
	.w1(32'h3c09bd7f),
	.w2(32'h3c87ccf2),
	.w3(32'h3ad935b1),
	.w4(32'h3b890238),
	.w5(32'h3c27242d),
	.w6(32'h3a95e1c6),
	.w7(32'h3c5a482c),
	.w8(32'hbb47920e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15078a),
	.w1(32'h3b1d93cd),
	.w2(32'hbccd95fb),
	.w3(32'hbb5a8884),
	.w4(32'h3c8ee161),
	.w5(32'hbc2e94a9),
	.w6(32'h3ae5ba24),
	.w7(32'hbb664617),
	.w8(32'h3c45a26c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac45e70),
	.w1(32'h38a24b34),
	.w2(32'hbb544285),
	.w3(32'h3c16988b),
	.w4(32'hbb8f2745),
	.w5(32'hbb8d0c4b),
	.w6(32'hbadda9d7),
	.w7(32'hbb12f67e),
	.w8(32'h3a6768e6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba76d75),
	.w1(32'h3c9ed65c),
	.w2(32'hbba96edd),
	.w3(32'h3b4a9715),
	.w4(32'h3c4b3c74),
	.w5(32'hbc624050),
	.w6(32'h3c8d7295),
	.w7(32'hba809c68),
	.w8(32'hbc06e40b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf68de7),
	.w1(32'h39d6af8e),
	.w2(32'h3c8960a0),
	.w3(32'hbc9d9cc5),
	.w4(32'h3bd7424c),
	.w5(32'hbc1c4a60),
	.w6(32'hbbfb043b),
	.w7(32'h3c6b016e),
	.w8(32'hbb81e4c5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eb285),
	.w1(32'h3c528cea),
	.w2(32'h3c430343),
	.w3(32'hbb9eeafe),
	.w4(32'h3be0f84d),
	.w5(32'hba3f06e8),
	.w6(32'h3c433f46),
	.w7(32'h3bfc34b5),
	.w8(32'hbc3cd4d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85e6a1),
	.w1(32'hbc789001),
	.w2(32'h3c677cf5),
	.w3(32'hbc9b0b4f),
	.w4(32'hbc4896dd),
	.w5(32'h3bfb1580),
	.w6(32'hbb8a86fe),
	.w7(32'h3c0071f5),
	.w8(32'h3bf84761),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11820b),
	.w1(32'h3afc37f7),
	.w2(32'h3899811b),
	.w3(32'h3c795c68),
	.w4(32'h3a92e2e1),
	.w5(32'hbb0fe819),
	.w6(32'h3ae0144e),
	.w7(32'hbafb4356),
	.w8(32'hbb24bfe9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b242efd),
	.w1(32'hbc810f46),
	.w2(32'hbc0bdfb8),
	.w3(32'h3b3ea17b),
	.w4(32'h3b44710a),
	.w5(32'hba8feff6),
	.w6(32'hbc0a6194),
	.w7(32'hbbf94cdf),
	.w8(32'hbc363fa1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc438c23),
	.w1(32'hbc0d5c11),
	.w2(32'h3b88f550),
	.w3(32'hbc1c64b6),
	.w4(32'hbc6035e4),
	.w5(32'h3adfd17b),
	.w6(32'hba3d50ce),
	.w7(32'h3a4ae8ca),
	.w8(32'h3c706b22),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdaffd),
	.w1(32'hbb98d259),
	.w2(32'h3a62e854),
	.w3(32'h3b683972),
	.w4(32'hbbb6fb94),
	.w5(32'hbbd8b9b0),
	.w6(32'hbb19dde8),
	.w7(32'hbb9c67b3),
	.w8(32'hbc706f9d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bf9b8),
	.w1(32'hbc1c8f28),
	.w2(32'h3c3acb2c),
	.w3(32'hbc8365de),
	.w4(32'hbb3b9fda),
	.w5(32'h3c358690),
	.w6(32'hbc3672c3),
	.w7(32'hba0b931c),
	.w8(32'h3c131df0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33dc45),
	.w1(32'hbbb109dc),
	.w2(32'h3bd46de7),
	.w3(32'h3c093520),
	.w4(32'hbb783d46),
	.w5(32'h3b84e836),
	.w6(32'hb8ffade1),
	.w7(32'h394d057e),
	.w8(32'h3a7d8449),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdb591),
	.w1(32'hba0bb9ea),
	.w2(32'hbcb72fe0),
	.w3(32'h3a802afc),
	.w4(32'hba80b781),
	.w5(32'hbc9c81ab),
	.w6(32'hbab6bf21),
	.w7(32'hbcaeb0d3),
	.w8(32'hbc6d7fce),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932b6d5),
	.w1(32'h3c2eeca3),
	.w2(32'hbbd9e3de),
	.w3(32'hbb689fc4),
	.w4(32'h3bbd86db),
	.w5(32'hbc1235e0),
	.w6(32'hbb884a9d),
	.w7(32'h3b9bf268),
	.w8(32'hba96add8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5874),
	.w1(32'hbafbed09),
	.w2(32'hbcb5b394),
	.w3(32'hbb584257),
	.w4(32'hbb8b9605),
	.w5(32'hbce3c183),
	.w6(32'hbca6f4cb),
	.w7(32'hbd0225fb),
	.w8(32'hbbdea2a5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eed75),
	.w1(32'hb893903a),
	.w2(32'h3c139fd5),
	.w3(32'h3b3f9717),
	.w4(32'hbafebf39),
	.w5(32'h3c17eb42),
	.w6(32'h3a348ba4),
	.w7(32'hba515de9),
	.w8(32'hbb685ebb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98156a),
	.w1(32'h3a1d1ef2),
	.w2(32'hb94e2782),
	.w3(32'h3c0d836d),
	.w4(32'h3c50cd6f),
	.w5(32'h3c4d55f3),
	.w6(32'hbae0f075),
	.w7(32'hbb20d492),
	.w8(32'hbc62d918),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc638136),
	.w1(32'hbbc6544f),
	.w2(32'hbba88a9a),
	.w3(32'hbb38133f),
	.w4(32'hbb42cb2a),
	.w5(32'h39aa2868),
	.w6(32'hbb99a80c),
	.w7(32'hbb139731),
	.w8(32'hbb1a0510),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0b12),
	.w1(32'hbbbe78f7),
	.w2(32'h3c1285c0),
	.w3(32'h3b656362),
	.w4(32'hbbe90fae),
	.w5(32'h3c0ccef6),
	.w6(32'hbc06ed3f),
	.w7(32'h3b871084),
	.w8(32'h3c06df59),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96462),
	.w1(32'h3c0ee572),
	.w2(32'hbbb8f436),
	.w3(32'h3c17861d),
	.w4(32'hbbcbbaa5),
	.w5(32'hbaf1f1f8),
	.w6(32'h3b9da67f),
	.w7(32'hbacf9707),
	.w8(32'hbbc12818),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21488c),
	.w1(32'h3c79e4ba),
	.w2(32'hbc39d030),
	.w3(32'hba63fec7),
	.w4(32'h3bfc66ae),
	.w5(32'hbbcd761b),
	.w6(32'h3ca8640e),
	.w7(32'hbc46373d),
	.w8(32'h3a63e854),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebfedc),
	.w1(32'h3b5ad094),
	.w2(32'hbace10d8),
	.w3(32'hbc8942a0),
	.w4(32'hbaa781b2),
	.w5(32'hb9311e8d),
	.w6(32'h394803e0),
	.w7(32'hbb470c5c),
	.w8(32'hbb581189),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abecd32),
	.w1(32'hbc7eaba3),
	.w2(32'hbc74cc33),
	.w3(32'h3ab8d2b1),
	.w4(32'hbc807308),
	.w5(32'hbc8dd1f1),
	.w6(32'hbb848521),
	.w7(32'hbbb3d8dc),
	.w8(32'hbb66ebe6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b867843),
	.w1(32'hbb1fd142),
	.w2(32'h3ab528a3),
	.w3(32'h3c760ede),
	.w4(32'hba1a24f4),
	.w5(32'h3a0f3822),
	.w6(32'hbb477335),
	.w7(32'hbb5d2ba2),
	.w8(32'hba99a305),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d447b),
	.w1(32'h3ba53cd3),
	.w2(32'h3b97318b),
	.w3(32'h3b912aa9),
	.w4(32'hbaa3d47b),
	.w5(32'h3ae25d7f),
	.w6(32'h3b1ada6f),
	.w7(32'h3bad34e1),
	.w8(32'h3bfc79a3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51d9e),
	.w1(32'hbb269225),
	.w2(32'h3c4d4859),
	.w3(32'h3af03673),
	.w4(32'h3c052a34),
	.w5(32'h3c70d0fa),
	.w6(32'hbc8a6543),
	.w7(32'h3b8f9028),
	.w8(32'hbbf1295d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc284723),
	.w1(32'hbc65fa17),
	.w2(32'h3b15fcb5),
	.w3(32'hbb975b17),
	.w4(32'hbc0bceae),
	.w5(32'h3bf56d71),
	.w6(32'hbc041e81),
	.w7(32'hbac1ff74),
	.w8(32'h3bafe356),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89339f),
	.w1(32'hbae8456f),
	.w2(32'hbc622c05),
	.w3(32'h3c2a32a1),
	.w4(32'hbb4faaa9),
	.w5(32'hbc657898),
	.w6(32'hba61e368),
	.w7(32'hbc325eef),
	.w8(32'hbbaec62d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63604f),
	.w1(32'hbb04858e),
	.w2(32'hbb167816),
	.w3(32'hbb442c60),
	.w4(32'h3bc1bd0f),
	.w5(32'hbc2230c2),
	.w6(32'hbbb6886e),
	.w7(32'hbb5ac3c7),
	.w8(32'h3bf46845),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb911c7),
	.w1(32'h3a69f0dc),
	.w2(32'h3ae29d85),
	.w3(32'h3beb14be),
	.w4(32'h3b9c46a5),
	.w5(32'h3c10446e),
	.w6(32'h3a70cd87),
	.w7(32'hbb836dac),
	.w8(32'hbb3c7e2f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919da40),
	.w1(32'h3a9cd1a7),
	.w2(32'h3ce2a586),
	.w3(32'h3b6a8762),
	.w4(32'h3b5cf3ae),
	.w5(32'h3cb108e7),
	.w6(32'h3bac90a9),
	.w7(32'h3c6305f5),
	.w8(32'hbc6a20f6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55aa1e),
	.w1(32'hbc045d85),
	.w2(32'hbd1e8c27),
	.w3(32'hbc48358e),
	.w4(32'hbc4bde76),
	.w5(32'hbd01a60b),
	.w6(32'h3a94595c),
	.w7(32'hbcc92291),
	.w8(32'h3b8ae884),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c739eb5),
	.w1(32'h3a2ac32f),
	.w2(32'hba957614),
	.w3(32'h3c882009),
	.w4(32'hb923b2e1),
	.w5(32'hbb9d8531),
	.w6(32'h3b29ef6c),
	.w7(32'hba77a385),
	.w8(32'h3b17a98e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c38b),
	.w1(32'h3a7b66db),
	.w2(32'h3b7fc0c0),
	.w3(32'h3b51ffb1),
	.w4(32'h3b97b527),
	.w5(32'h3c00be9e),
	.w6(32'hbb4d984e),
	.w7(32'h3ac2ec2e),
	.w8(32'hbb07d56c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd76b),
	.w1(32'hbc289a88),
	.w2(32'hbb9f4c09),
	.w3(32'hbc03ca5a),
	.w4(32'hbc8ec8d7),
	.w5(32'h3a80718b),
	.w6(32'h3b149f86),
	.w7(32'hbc127ff2),
	.w8(32'h3c063a55),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab19a1),
	.w1(32'hbc1377db),
	.w2(32'hbc061113),
	.w3(32'h3cc32c60),
	.w4(32'hbc76a95d),
	.w5(32'hbbd1b5dc),
	.w6(32'hbb6d3541),
	.w7(32'hbbc7f8bc),
	.w8(32'h3bd86f09),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce88fce),
	.w1(32'h3b2ec26f),
	.w2(32'h3ac6ed4d),
	.w3(32'h3caa7776),
	.w4(32'h3bfd3b5e),
	.w5(32'h3bcf110f),
	.w6(32'h3a1cb566),
	.w7(32'h3bdfc74b),
	.w8(32'hbb282797),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f4d6e),
	.w1(32'h3bd18897),
	.w2(32'hbb36763c),
	.w3(32'hbb0fca77),
	.w4(32'h3b5ff10c),
	.w5(32'hbb666e09),
	.w6(32'h3ad14792),
	.w7(32'hbbddafa7),
	.w8(32'h3b366f87),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389aa73e),
	.w1(32'hbb0279a5),
	.w2(32'hba61561d),
	.w3(32'hba13f5e7),
	.w4(32'hbae29e76),
	.w5(32'hbb9c9f57),
	.w6(32'hbb83a3b3),
	.w7(32'hba09a696),
	.w8(32'h3b9d9a93),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbee41),
	.w1(32'hb976ed16),
	.w2(32'hba9f30f9),
	.w3(32'h3ae32459),
	.w4(32'hbb2c8658),
	.w5(32'hbb4ff521),
	.w6(32'hbb8b1510),
	.w7(32'hbb88e7ed),
	.w8(32'hb9bdc06e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6377a2),
	.w1(32'hbc9e1c9b),
	.w2(32'h3c918d99),
	.w3(32'hb90a89af),
	.w4(32'hbc5ae84d),
	.w5(32'h3cf76bc1),
	.w6(32'hbc127763),
	.w7(32'h3c39ab8d),
	.w8(32'h3c5436dc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96ca03),
	.w1(32'h3a8e8053),
	.w2(32'h3bb233c3),
	.w3(32'h3c87d295),
	.w4(32'h3b9a35e7),
	.w5(32'h3bca381b),
	.w6(32'hbb088885),
	.w7(32'h3b25d84e),
	.w8(32'hbb2ef4fa),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c61c0),
	.w1(32'h3c01ed12),
	.w2(32'h3c00c7d5),
	.w3(32'h3b2424ab),
	.w4(32'h3bb8adc0),
	.w5(32'hbc02f351),
	.w6(32'h3c9b596a),
	.w7(32'hbae22ab1),
	.w8(32'hbc9618de),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54eb30),
	.w1(32'h3c0ae9f8),
	.w2(32'h3b0e6735),
	.w3(32'hbcdb3367),
	.w4(32'h3b8aaf22),
	.w5(32'h38c3c55e),
	.w6(32'h3ab55ef1),
	.w7(32'h3b855886),
	.w8(32'hbc42e624),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c1b33),
	.w1(32'hbb9d6c64),
	.w2(32'hbc10dc9e),
	.w3(32'hbc94efbf),
	.w4(32'hbb3a760b),
	.w5(32'hbb90aec0),
	.w6(32'hba4be7d7),
	.w7(32'hbc263b12),
	.w8(32'hbbae541f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef0fe0),
	.w1(32'h3a85208d),
	.w2(32'h3b03d020),
	.w3(32'h3aae2e50),
	.w4(32'hbac5025a),
	.w5(32'hbb44aacf),
	.w6(32'hbacc9c7b),
	.w7(32'hb921aafe),
	.w8(32'h3a9a6a6c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b029501),
	.w1(32'hbc199cc3),
	.w2(32'h3c808a71),
	.w3(32'h3a2fad6a),
	.w4(32'hbbcbd494),
	.w5(32'h3b203f7d),
	.w6(32'hbbec8729),
	.w7(32'h3b82c167),
	.w8(32'h3c321736),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0184dc),
	.w1(32'h3c0fc885),
	.w2(32'h3c30ff1f),
	.w3(32'h3b51995e),
	.w4(32'h3bdcf93e),
	.w5(32'hbaf18905),
	.w6(32'h3bf641ad),
	.w7(32'h3c9692f4),
	.w8(32'h3b162e7b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99150),
	.w1(32'h3ad4f40d),
	.w2(32'hbbc76cbd),
	.w3(32'hbc20da1c),
	.w4(32'h3ae8474d),
	.w5(32'hbb452fe4),
	.w6(32'hba9eaf59),
	.w7(32'hbb818a92),
	.w8(32'hbb87a05b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05fc5c),
	.w1(32'h398c51e4),
	.w2(32'h3baa705d),
	.w3(32'hb9722534),
	.w4(32'hbbba7d17),
	.w5(32'h3b4e5d2d),
	.w6(32'h3b1ba280),
	.w7(32'h3bdd3aca),
	.w8(32'h3b3a986a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed0bdd),
	.w1(32'hb9e7a6d2),
	.w2(32'hbb5e6a3e),
	.w3(32'h3c3be154),
	.w4(32'h3a406581),
	.w5(32'hbad35ebb),
	.w6(32'hbb0e06b1),
	.w7(32'hbb956ec4),
	.w8(32'hbbb05d17),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecafd9),
	.w1(32'hbb32df75),
	.w2(32'hbaba3f0d),
	.w3(32'hbbea6bfc),
	.w4(32'hbb55d393),
	.w5(32'hbb603c4e),
	.w6(32'hbb92422c),
	.w7(32'hbb8fdc91),
	.w8(32'hbaac4095),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65dc1c),
	.w1(32'hbc52c7e9),
	.w2(32'h3bc680a1),
	.w3(32'h3b5f2613),
	.w4(32'hbc408599),
	.w5(32'h3bee73ce),
	.w6(32'hbb721fa8),
	.w7(32'hbbed82e5),
	.w8(32'h3c2a260e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44f657),
	.w1(32'hbb979ab7),
	.w2(32'h3bc4d78d),
	.w3(32'h3c558b9a),
	.w4(32'h3bd7959b),
	.w5(32'h3c1afbb2),
	.w6(32'hb9445408),
	.w7(32'h3a0f6504),
	.w8(32'hbbf6a8a1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e277),
	.w1(32'h3b33414c),
	.w2(32'h3c12f60f),
	.w3(32'hbcc2f4af),
	.w4(32'h3be4e34d),
	.w5(32'h3b730b07),
	.w6(32'h3b77facd),
	.w7(32'h3ae24f28),
	.w8(32'hbb1aa7e8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc383457),
	.w1(32'h3c95f3f7),
	.w2(32'hbcd50159),
	.w3(32'hbc35025e),
	.w4(32'h3ba24116),
	.w5(32'hbc813f60),
	.w6(32'h3c9e7b99),
	.w7(32'hbc188540),
	.w8(32'hbb88eaad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd84b4d),
	.w1(32'hbb8d9705),
	.w2(32'hbc2f65f0),
	.w3(32'hbcb4a8b4),
	.w4(32'hbc682f35),
	.w5(32'hbc81d85f),
	.w6(32'hba617d3d),
	.w7(32'hbc1f7ff6),
	.w8(32'h3c1501ff),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc98522),
	.w1(32'hb9539908),
	.w2(32'hbba14263),
	.w3(32'h3bbf49fc),
	.w4(32'hbb6095b1),
	.w5(32'hbbcd83bc),
	.w6(32'hbb064ee1),
	.w7(32'hbb797933),
	.w8(32'h3b339fff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fe3e3),
	.w1(32'hbbb87d96),
	.w2(32'hbc9651e2),
	.w3(32'h3bab54ff),
	.w4(32'h39dc8c0c),
	.w5(32'hbc8ea9f5),
	.w6(32'h39fc6966),
	.w7(32'hbb314020),
	.w8(32'h3bb959ae),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97542b),
	.w1(32'hbbdc594a),
	.w2(32'hbc917456),
	.w3(32'h3ba109d7),
	.w4(32'hbbcdf142),
	.w5(32'hbc647010),
	.w6(32'hbb3c0ba4),
	.w7(32'hbb3f7da4),
	.w8(32'hbb9397f5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0da8ee),
	.w1(32'h3b72ef35),
	.w2(32'h39803abc),
	.w3(32'h3ca0fb2e),
	.w4(32'hbb19a12d),
	.w5(32'hbb66884c),
	.w6(32'h3bd4ace6),
	.w7(32'hbb3d2d6d),
	.w8(32'hbb681863),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7f15b),
	.w1(32'h3b0e57ba),
	.w2(32'hbbbd6d32),
	.w3(32'h3a105cbd),
	.w4(32'hbb3d4055),
	.w5(32'hbc295166),
	.w6(32'h3ae23dfc),
	.w7(32'hbb061f12),
	.w8(32'hbb2f186b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6df2e),
	.w1(32'hbb09584a),
	.w2(32'h3bb50323),
	.w3(32'h3b9860ef),
	.w4(32'hbb31ec90),
	.w5(32'h39da35a4),
	.w6(32'hbb935bb5),
	.w7(32'h3b31a3d4),
	.w8(32'hbc0a313c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7d509),
	.w1(32'hbbd6fc67),
	.w2(32'hb96e67d3),
	.w3(32'hbbcd5bac),
	.w4(32'hbb9b8891),
	.w5(32'h3b6d3fb9),
	.w6(32'hba5ea6e2),
	.w7(32'hbb1294ea),
	.w8(32'hbb3b91e9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0adb44),
	.w1(32'hbbd3ee3c),
	.w2(32'hbbd27802),
	.w3(32'h3b0665bc),
	.w4(32'hbb8cdc54),
	.w5(32'hbc0722a8),
	.w6(32'hbc037307),
	.w7(32'hbc4db775),
	.w8(32'hbc5dd83c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4f91a),
	.w1(32'hbb71cd75),
	.w2(32'hbc46adb4),
	.w3(32'hbb841386),
	.w4(32'hbbb5018b),
	.w5(32'hbc58a32a),
	.w6(32'hbba3adeb),
	.w7(32'hbc332d68),
	.w8(32'h3ba88200),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964bed),
	.w1(32'h3c98465d),
	.w2(32'hbc63e958),
	.w3(32'h3b2d4307),
	.w4(32'h3a2fa79d),
	.w5(32'hbc3f1512),
	.w6(32'h3c03ba30),
	.w7(32'hbc297529),
	.w8(32'hbc187caa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185da7),
	.w1(32'h3b5a303a),
	.w2(32'hbc85fae3),
	.w3(32'hbc5f9b46),
	.w4(32'h3bd2fb90),
	.w5(32'hbc26f6e9),
	.w6(32'h3b8b8f9d),
	.w7(32'hbb6ab2ca),
	.w8(32'h3b049039),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e7441),
	.w1(32'h3c6e4c76),
	.w2(32'hbccf2daf),
	.w3(32'h3b9711df),
	.w4(32'h3c0b1839),
	.w5(32'hbc81848e),
	.w6(32'h3b0d6492),
	.w7(32'hbc3ba151),
	.w8(32'h3b806936),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb10982),
	.w1(32'hbc60d40a),
	.w2(32'hbbb33609),
	.w3(32'hbb5dd0a2),
	.w4(32'hbc025060),
	.w5(32'hbc22cf46),
	.w6(32'h3a60e1a6),
	.w7(32'hba92f12c),
	.w8(32'hb9d5b2fa),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb108a0d),
	.w1(32'hbbc074b6),
	.w2(32'hbb3d26b2),
	.w3(32'hbb913ced),
	.w4(32'h39ef4193),
	.w5(32'h3c243357),
	.w6(32'hbbb8305b),
	.w7(32'hbbac61d6),
	.w8(32'h3bf6a47a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a994683),
	.w1(32'h3b9b54bd),
	.w2(32'hbce091c9),
	.w3(32'h3b45d062),
	.w4(32'h3bd8d02d),
	.w5(32'hbce10a64),
	.w6(32'hbb9a4c96),
	.w7(32'hbc6aab81),
	.w8(32'h3b00fcb1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a78e4),
	.w1(32'h3c342b4c),
	.w2(32'hbbd38d7f),
	.w3(32'h3a2e3299),
	.w4(32'h3b84ff57),
	.w5(32'hbc90dc4e),
	.w6(32'h3bd26ca1),
	.w7(32'hbc1772a9),
	.w8(32'hbc24ad62),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901169),
	.w1(32'hbac44167),
	.w2(32'h3ae8e6cb),
	.w3(32'hbb3185aa),
	.w4(32'h3aa1906a),
	.w5(32'h3b740179),
	.w6(32'h3a68e940),
	.w7(32'h3b29e259),
	.w8(32'h3b9e0e19),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b380ba6),
	.w1(32'hbac2013f),
	.w2(32'h39227cf5),
	.w3(32'h3be74660),
	.w4(32'hbacc4c79),
	.w5(32'hbb509c8d),
	.w6(32'h3bbbca19),
	.w7(32'h3ba1b2f0),
	.w8(32'h3bccc79c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74f831),
	.w1(32'h3ac2da7a),
	.w2(32'h3a42efaa),
	.w3(32'h3b1ecd8c),
	.w4(32'hba680ae3),
	.w5(32'hbafcde60),
	.w6(32'h3b2db537),
	.w7(32'h3b1eb87a),
	.w8(32'h3ab04dac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaedec8),
	.w1(32'hbbe9b170),
	.w2(32'hbbc17160),
	.w3(32'h3b5ebbfa),
	.w4(32'hbb934051),
	.w5(32'hbba07b18),
	.w6(32'h3b1dc0df),
	.w7(32'h3b78b22f),
	.w8(32'h3bf0487e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51c76e),
	.w1(32'hbbefb88d),
	.w2(32'hbc3ff7fd),
	.w3(32'h3c75c293),
	.w4(32'hbba95cf6),
	.w5(32'hbc8e9e9c),
	.w6(32'hba320013),
	.w7(32'hbabbc27f),
	.w8(32'hbbd740ce),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6444b),
	.w1(32'h3c5f523b),
	.w2(32'hbc4ac3cc),
	.w3(32'h3c77969d),
	.w4(32'h3bb72874),
	.w5(32'hbb9f0e62),
	.w6(32'h3bc64e92),
	.w7(32'hbc4b08bb),
	.w8(32'hbb913dfc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dc9b6),
	.w1(32'h3b5828e2),
	.w2(32'h3b8b1994),
	.w3(32'hbba9f36b),
	.w4(32'h3b29e4c6),
	.w5(32'h3b7062de),
	.w6(32'hba5aa51c),
	.w7(32'h3b467112),
	.w8(32'h3b3256d9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade2f62),
	.w1(32'h380c4c7c),
	.w2(32'h3ba1f80f),
	.w3(32'hb983344c),
	.w4(32'h3ab1c9b8),
	.w5(32'h3b65e002),
	.w6(32'hba96233b),
	.w7(32'h3b000cd8),
	.w8(32'h3b1c46cf),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaced1b),
	.w1(32'hbc4ce3ee),
	.w2(32'h3c8ab9ac),
	.w3(32'h3b0e438e),
	.w4(32'hbb9e93bd),
	.w5(32'h3c83b134),
	.w6(32'hbbdfc141),
	.w7(32'h3c553be0),
	.w8(32'h3c1ffe37),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09e986),
	.w1(32'hba2f367b),
	.w2(32'hbbe1442f),
	.w3(32'h3bd68f6f),
	.w4(32'hbb64b6e7),
	.w5(32'hbc0ad21b),
	.w6(32'h3ac32644),
	.w7(32'hbb97d7f0),
	.w8(32'hbbc9bea5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf65b1),
	.w1(32'hbb917303),
	.w2(32'h3b245691),
	.w3(32'hbb6e0f66),
	.w4(32'hbb1531fb),
	.w5(32'h3b7c7fcc),
	.w6(32'hbc3f5779),
	.w7(32'hbaf4310b),
	.w8(32'hbbef2a08),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893bf71),
	.w1(32'hbc0a8b02),
	.w2(32'h3c2d684b),
	.w3(32'hbb4a0d13),
	.w4(32'h3bc463ab),
	.w5(32'h3c5421da),
	.w6(32'hbbbfa02b),
	.w7(32'h3bcc7532),
	.w8(32'hbbb3d47f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc180242),
	.w1(32'hba727179),
	.w2(32'h3c78c04b),
	.w3(32'hbafd7949),
	.w4(32'h3c8045b8),
	.w5(32'h3c68bdef),
	.w6(32'hbbd287e8),
	.w7(32'h3c604dea),
	.w8(32'hbc213f7b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc387615),
	.w1(32'hbc30e497),
	.w2(32'hbc482935),
	.w3(32'hbc59a949),
	.w4(32'hbc23f226),
	.w5(32'hbc688f14),
	.w6(32'h399956e5),
	.w7(32'hbc3be420),
	.w8(32'h3b87080d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14e6bd),
	.w1(32'h3bb8b7e6),
	.w2(32'h3c8c7604),
	.w3(32'h3c27a91a),
	.w4(32'h3b2d2b22),
	.w5(32'h3ca3c86c),
	.w6(32'h3bec3ab5),
	.w7(32'h3abb6780),
	.w8(32'hbb5187f9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8376e),
	.w1(32'h39b84a4e),
	.w2(32'hbc8d5d9c),
	.w3(32'hbc6b269d),
	.w4(32'hbbb445c2),
	.w5(32'hbc5c0b03),
	.w6(32'h3a2ff6d4),
	.w7(32'h3b53014e),
	.w8(32'h3b76718a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c172218),
	.w1(32'h3b88e0a1),
	.w2(32'hbc845967),
	.w3(32'h3c2039e8),
	.w4(32'h3c16d54b),
	.w5(32'hbc338d3e),
	.w6(32'h3a89e484),
	.w7(32'hbb02af2d),
	.w8(32'h3b789feb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc72c0),
	.w1(32'hbc3f15db),
	.w2(32'h3c3ff662),
	.w3(32'hbc0290dc),
	.w4(32'hbbbf4896),
	.w5(32'h3c92defb),
	.w6(32'h3aca6cea),
	.w7(32'h3c17a376),
	.w8(32'h3c3e2979),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9104d),
	.w1(32'h3ca943ee),
	.w2(32'hbc58ad28),
	.w3(32'h37cc7429),
	.w4(32'h3cb04dcc),
	.w5(32'hbc55c970),
	.w6(32'h3c84680c),
	.w7(32'h38b47210),
	.w8(32'hbc223e67),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccae8e),
	.w1(32'hbb03dab3),
	.w2(32'hbb3c16e5),
	.w3(32'hbbc04340),
	.w4(32'hbb558b64),
	.w5(32'hbbf18565),
	.w6(32'hbb5ab001),
	.w7(32'hbb796a2d),
	.w8(32'hba3f9da1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b239178),
	.w1(32'hbbc7fbb9),
	.w2(32'hba3a10e6),
	.w3(32'h3b256745),
	.w4(32'hbb28b125),
	.w5(32'hb9ead081),
	.w6(32'hbb6013df),
	.w7(32'hbbe53607),
	.w8(32'hbc0188d5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc9c84),
	.w1(32'hbc0743e8),
	.w2(32'hbc334f0b),
	.w3(32'h3b49fdc8),
	.w4(32'h39e08697),
	.w5(32'hbc0ee937),
	.w6(32'hbc07c0f3),
	.w7(32'hbc50b2f0),
	.w8(32'hbb92656b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb201279),
	.w1(32'hbb60e7bf),
	.w2(32'h3b0a3cbd),
	.w3(32'h3a8298f4),
	.w4(32'hb969aba3),
	.w5(32'h3b87dc7f),
	.w6(32'h392abd5d),
	.w7(32'h3a429063),
	.w8(32'h3aec8b6d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236bba),
	.w1(32'hba07c2f0),
	.w2(32'h3af05002),
	.w3(32'h3b969dba),
	.w4(32'h3ab10d13),
	.w5(32'h3ae5836b),
	.w6(32'hbad6b0f6),
	.w7(32'hba389782),
	.w8(32'h3a8c0c52),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f2309),
	.w1(32'hbb32edc4),
	.w2(32'hbc445708),
	.w3(32'h3b31da7a),
	.w4(32'h3b6d05cf),
	.w5(32'hbc596aa5),
	.w6(32'hbbd6ae2e),
	.w7(32'hb9ef53f6),
	.w8(32'h3b4f3a95),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9070a2),
	.w1(32'hbafd8315),
	.w2(32'hbabc311e),
	.w3(32'hbab7c82e),
	.w4(32'hba9fbcd4),
	.w5(32'hbabd3da2),
	.w6(32'hba31bef3),
	.w7(32'hbb07a6b7),
	.w8(32'hba9f5f9e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6864b),
	.w1(32'hbb70d0c9),
	.w2(32'h3c40486a),
	.w3(32'hbaf64d62),
	.w4(32'h3b040225),
	.w5(32'h3c0e72b6),
	.w6(32'hbb125be4),
	.w7(32'h3b9a577e),
	.w8(32'h3b5ffa30),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19c2a5),
	.w1(32'hbc0c10e2),
	.w2(32'hbc73d8d7),
	.w3(32'h3ae4c68f),
	.w4(32'hbbabfed2),
	.w5(32'h3b2eb7c4),
	.w6(32'hbbd77623),
	.w7(32'hbc87cbf6),
	.w8(32'h3c70aa69),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0677e),
	.w1(32'hbbe83ffe),
	.w2(32'hbbada771),
	.w3(32'h3c144219),
	.w4(32'hbb67abbf),
	.w5(32'hbbd69e28),
	.w6(32'hbb8eab42),
	.w7(32'hbaa9ddcc),
	.w8(32'h3b4d8e0d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6faad9),
	.w1(32'h3ab696da),
	.w2(32'h3b59cc40),
	.w3(32'h3b1b5474),
	.w4(32'h39da5319),
	.w5(32'h3ac6b6a5),
	.w6(32'hba299c1f),
	.w7(32'h3ab12eda),
	.w8(32'h3adbf156),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2a67),
	.w1(32'h3ba96e98),
	.w2(32'hbacad94d),
	.w3(32'h3b18d284),
	.w4(32'h3ba6ab44),
	.w5(32'hbbb80e4a),
	.w6(32'h3be130dc),
	.w7(32'hbb0b884c),
	.w8(32'hbaee4832),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e41b83),
	.w1(32'h3c20f252),
	.w2(32'h3becbfcd),
	.w3(32'h3b387e32),
	.w4(32'h3b5206a1),
	.w5(32'hbb4e8451),
	.w6(32'h3c1573a8),
	.w7(32'h3ae681a1),
	.w8(32'h3a9bb55c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4272e9),
	.w1(32'h3b3f2f0e),
	.w2(32'hbba8bc27),
	.w3(32'hbbb01121),
	.w4(32'h3bcbcbd6),
	.w5(32'hbc2779f0),
	.w6(32'h3c17e18b),
	.w7(32'h3af5c8f8),
	.w8(32'hbac6d0ff),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81b260),
	.w1(32'hba17c566),
	.w2(32'hbacdd2e2),
	.w3(32'hbc9aeb63),
	.w4(32'h3a8a8745),
	.w5(32'hba817182),
	.w6(32'h3b05e9a6),
	.w7(32'hbb50ff05),
	.w8(32'hbacb95f9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdf933),
	.w1(32'h3cb161fd),
	.w2(32'hbc4fd892),
	.w3(32'h3b4722a1),
	.w4(32'h3bdb2a9d),
	.w5(32'hbc8a3efc),
	.w6(32'h3c8f514d),
	.w7(32'hbc8c6a55),
	.w8(32'hbc4cd034),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd61538),
	.w1(32'h3b4e7cd9),
	.w2(32'hbac68d17),
	.w3(32'hbcb07ec5),
	.w4(32'h3b2d94fc),
	.w5(32'hbc1dee62),
	.w6(32'h3bbbeb7a),
	.w7(32'h3b2728ed),
	.w8(32'h3bac4f20),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48cc0f),
	.w1(32'hbabb402f),
	.w2(32'h3a5142a6),
	.w3(32'hbbdc1b1d),
	.w4(32'hbb06e441),
	.w5(32'h3b171cdf),
	.w6(32'hbb1b0c61),
	.w7(32'h3981251c),
	.w8(32'h3b01db92),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd620e),
	.w1(32'hbbcf86f0),
	.w2(32'h3c00e80c),
	.w3(32'hb938a50c),
	.w4(32'hbbe90439),
	.w5(32'h3b8e0fc5),
	.w6(32'hba9d796e),
	.w7(32'h3c0e5268),
	.w8(32'h3c1b6d59),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841096),
	.w1(32'h3c3ba053),
	.w2(32'hbc8fb0ca),
	.w3(32'h3ad85034),
	.w4(32'h3bcf7bd7),
	.w5(32'hbb563311),
	.w6(32'h3bcf1005),
	.w7(32'hbc4d2849),
	.w8(32'hbc82bee5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52b5ae),
	.w1(32'hbc3cc30a),
	.w2(32'h3a676caa),
	.w3(32'hbc0a408b),
	.w4(32'hbc6a96bf),
	.w5(32'h3b765f35),
	.w6(32'hbab1a3bd),
	.w7(32'hbbb331ed),
	.w8(32'h3c230b2a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc41a6),
	.w1(32'hbae95d55),
	.w2(32'hbb59f665),
	.w3(32'h3ce5199c),
	.w4(32'h39df3379),
	.w5(32'hb982bfbb),
	.w6(32'hb7aa63a8),
	.w7(32'hb87b9b3b),
	.w8(32'hba6fb5c8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66316f),
	.w1(32'h3d099c4b),
	.w2(32'h3d71c33f),
	.w3(32'hbab0d809),
	.w4(32'h3cec68cf),
	.w5(32'h3d33fccd),
	.w6(32'h3cbe9f96),
	.w7(32'h3d20673f),
	.w8(32'h3cd54dd3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule