module layer_10_featuremap_267(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae54dc),
	.w1(32'hba4f712f),
	.w2(32'hbbc76e4a),
	.w3(32'hbaa9a94d),
	.w4(32'hbb5c9128),
	.w5(32'h3c0efa4c),
	.w6(32'h3b8c21aa),
	.w7(32'hbb52c921),
	.w8(32'h3b9f7a96),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9802bb),
	.w1(32'h3bffa336),
	.w2(32'h3cbb54aa),
	.w3(32'h3b46d1a9),
	.w4(32'hbacd4516),
	.w5(32'h3bb6b6e2),
	.w6(32'hbaa12e84),
	.w7(32'hbabbf41c),
	.w8(32'h3a7ca2ee),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c389a),
	.w1(32'hba84fa94),
	.w2(32'hbb74beda),
	.w3(32'h3b55950f),
	.w4(32'h3a13ae13),
	.w5(32'h3b01b4aa),
	.w6(32'h39d4cf1d),
	.w7(32'hbb2d449a),
	.w8(32'h3b22f908),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52814),
	.w1(32'h3bba6bf9),
	.w2(32'h3bf8ebf8),
	.w3(32'h3a38dce2),
	.w4(32'h3aec7628),
	.w5(32'h3afd54fc),
	.w6(32'h3b38a0a2),
	.w7(32'h3a8925b9),
	.w8(32'h37c633b4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b543ede),
	.w1(32'h3bb227ae),
	.w2(32'h3b261cf2),
	.w3(32'h39b01c26),
	.w4(32'hba6b5c4f),
	.w5(32'hba806cc4),
	.w6(32'hb92356ae),
	.w7(32'hbb334ae3),
	.w8(32'hba11a195),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae80ac0),
	.w1(32'hb8036ea7),
	.w2(32'hbacf4361),
	.w3(32'h39574cbb),
	.w4(32'hbac9fb9a),
	.w5(32'h3b81c56a),
	.w6(32'h3accdc35),
	.w7(32'hbab2d1e4),
	.w8(32'h3b7ac570),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33ba6f),
	.w1(32'h3c30d28e),
	.w2(32'hbc1a045c),
	.w3(32'h3b95e503),
	.w4(32'h3b0d2cfd),
	.w5(32'hbc9ebc13),
	.w6(32'h3c32ca59),
	.w7(32'hbab6cc60),
	.w8(32'hbc925116),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babc5b9),
	.w1(32'hbc815f2e),
	.w2(32'hbcc20d81),
	.w3(32'hbc621f91),
	.w4(32'h3c6732c7),
	.w5(32'h3bd7e33a),
	.w6(32'h3b4728c8),
	.w7(32'h3a9cfc5c),
	.w8(32'h3bfb3fe4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56df2),
	.w1(32'h3b6467bf),
	.w2(32'h3b122021),
	.w3(32'h3988cd9f),
	.w4(32'h3abf62ec),
	.w5(32'hbb2c26bf),
	.w6(32'h3b209a34),
	.w7(32'h3a2877c0),
	.w8(32'hbab6158f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87576),
	.w1(32'hbc09e17b),
	.w2(32'hbc77c182),
	.w3(32'hb900e353),
	.w4(32'hbb8f2063),
	.w5(32'hbc0ecaae),
	.w6(32'h3bfbb3e6),
	.w7(32'h39e3dd0e),
	.w8(32'hba7f4faf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a6f2e),
	.w1(32'h3ad3098b),
	.w2(32'hbaa758c8),
	.w3(32'hba877971),
	.w4(32'hba87de82),
	.w5(32'h3bc057b7),
	.w6(32'h3a30b98a),
	.w7(32'hba6bafb4),
	.w8(32'h3afe11c4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3abbf4),
	.w1(32'h3bec5e3c),
	.w2(32'hbcbe6d83),
	.w3(32'h3ba930ad),
	.w4(32'h3be52ecf),
	.w5(32'hbc8d8698),
	.w6(32'h3c3c046f),
	.w7(32'h3a6bff65),
	.w8(32'hbb92c3bf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92bd2),
	.w1(32'hbc476a9a),
	.w2(32'hbc9c41ef),
	.w3(32'h3aab0ebc),
	.w4(32'hbb1e116b),
	.w5(32'hbc3109b3),
	.w6(32'h3b07843a),
	.w7(32'hbb23db40),
	.w8(32'hbbac6a04),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886fde),
	.w1(32'hbbb2ffa0),
	.w2(32'hbc06e305),
	.w3(32'hbc11c7ea),
	.w4(32'hbc2b1070),
	.w5(32'h3a2a664e),
	.w6(32'hbb931831),
	.w7(32'hbc38c59b),
	.w8(32'h3aae337e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9229e),
	.w1(32'h3c3f7665),
	.w2(32'h3c49daae),
	.w3(32'h3ba9104d),
	.w4(32'h3bbd611a),
	.w5(32'h3b5a90b4),
	.w6(32'h3ba41659),
	.w7(32'h3bcf4684),
	.w8(32'h3ad7d16e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a078f),
	.w1(32'hbc143b34),
	.w2(32'hbbbda20c),
	.w3(32'h3a0d310a),
	.w4(32'hbbcac1e3),
	.w5(32'hbb8c8925),
	.w6(32'h39a789ea),
	.w7(32'h3b7b6c56),
	.w8(32'h3bfd2c46),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9819421),
	.w1(32'h3a7c7fdf),
	.w2(32'hb75e2794),
	.w3(32'h3b3a4a4b),
	.w4(32'hb9c9a449),
	.w5(32'hba126b11),
	.w6(32'h3b975b02),
	.w7(32'h39169cd0),
	.w8(32'h3972ca5f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe58633),
	.w1(32'hbc567324),
	.w2(32'hbce27d17),
	.w3(32'h3c0832e6),
	.w4(32'hbaee0b54),
	.w5(32'hbc0ed7a2),
	.w6(32'h3c1b367f),
	.w7(32'h3b907dd8),
	.w8(32'hbb53b565),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4652),
	.w1(32'hbc1159e2),
	.w2(32'hbc829f37),
	.w3(32'h3bb61eaf),
	.w4(32'hb9c1e4ab),
	.w5(32'hbc1ff660),
	.w6(32'h3bf5440d),
	.w7(32'h3b9b7a5c),
	.w8(32'hbb8f8bf1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada11d5),
	.w1(32'hbaa5ee98),
	.w2(32'hb906f143),
	.w3(32'hb9430586),
	.w4(32'h3882371f),
	.w5(32'h38bb0b07),
	.w6(32'hbb16b854),
	.w7(32'h3a2e9b0c),
	.w8(32'h3a6efe97),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067ee4),
	.w1(32'h3b2a6f5d),
	.w2(32'h3ae502a1),
	.w3(32'hba396b56),
	.w4(32'hbaec8989),
	.w5(32'h3aa5843b),
	.w6(32'h3b16f73d),
	.w7(32'h3a3983ac),
	.w8(32'h3b3613cc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf2387),
	.w1(32'h3bf7ef96),
	.w2(32'h3c09da2b),
	.w3(32'h3b7bd935),
	.w4(32'h3b3bb65b),
	.w5(32'h3b281cdb),
	.w6(32'h3acf6d77),
	.w7(32'h3ad29287),
	.w8(32'h3a44d2aa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91b09d),
	.w1(32'hbbd2a15d),
	.w2(32'hbc8c369b),
	.w3(32'h3c50a3ce),
	.w4(32'h3bac13d5),
	.w5(32'hbca57163),
	.w6(32'h3c8a0d83),
	.w7(32'h3c729e8e),
	.w8(32'h3b88d91b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245539),
	.w1(32'h3b2d595c),
	.w2(32'h3a36da18),
	.w3(32'h3a3676bc),
	.w4(32'h3b11bef8),
	.w5(32'h3b98a7d6),
	.w6(32'h3c1bded9),
	.w7(32'h3c1348c5),
	.w8(32'h3ba214e8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c4f7a),
	.w1(32'h3c68ad64),
	.w2(32'h3cef01d1),
	.w3(32'h3aaa0aa3),
	.w4(32'h3bb71072),
	.w5(32'h3c454995),
	.w6(32'hbbd27040),
	.w7(32'hbbba6a34),
	.w8(32'h3b88f2c5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a275da8),
	.w1(32'h3b56cb4d),
	.w2(32'hba405b47),
	.w3(32'h3ad517b6),
	.w4(32'hb8f881c8),
	.w5(32'h3b67b7d7),
	.w6(32'h3b9dfe17),
	.w7(32'h3b3f634e),
	.w8(32'h3b96be81),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cf044),
	.w1(32'h3b627456),
	.w2(32'h3b5b4297),
	.w3(32'h3b5f2968),
	.w4(32'h3b9310c4),
	.w5(32'hbb30ad0d),
	.w6(32'h3b60ca87),
	.w7(32'h3b8be594),
	.w8(32'hba9b6ab8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097d9e),
	.w1(32'hbc52a213),
	.w2(32'hbc153066),
	.w3(32'h3b3c2a15),
	.w4(32'hbcaea7d2),
	.w5(32'hbca26131),
	.w6(32'hbc263f74),
	.w7(32'hbc829511),
	.w8(32'hbc207780),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f98a),
	.w1(32'hb72aa440),
	.w2(32'hbabd8cf0),
	.w3(32'hbb6ffe3f),
	.w4(32'h39ea0df1),
	.w5(32'hbab8b051),
	.w6(32'hbb841443),
	.w7(32'hbaa9d822),
	.w8(32'hba5eaacc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb835946),
	.w1(32'h3b067456),
	.w2(32'h3c5b09b7),
	.w3(32'hbbea8a8a),
	.w4(32'hbc8a6148),
	.w5(32'hbb8c16f8),
	.w6(32'hbc170563),
	.w7(32'hbc632029),
	.w8(32'hbc387cb6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42e1af),
	.w1(32'h3abdb70f),
	.w2(32'h3a68783b),
	.w3(32'hbb0b5776),
	.w4(32'hba9ea16e),
	.w5(32'h3b233f03),
	.w6(32'hbb212471),
	.w7(32'h3b1a58f8),
	.w8(32'h3b49a874),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b7f40),
	.w1(32'hbb082fa8),
	.w2(32'hbb789ee5),
	.w3(32'h3b9c295e),
	.w4(32'h3bc0ce32),
	.w5(32'hbaebbbc6),
	.w6(32'hbb0b866c),
	.w7(32'h3ab49825),
	.w8(32'h3a7ff422),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed1c06),
	.w1(32'hbb3b62b6),
	.w2(32'hbc016744),
	.w3(32'h3b6fb2f4),
	.w4(32'h3b6ff45e),
	.w5(32'hbb6df9c1),
	.w6(32'h3bec2d09),
	.w7(32'h3babe18a),
	.w8(32'hba963701),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb771ce3),
	.w1(32'h3ad033bd),
	.w2(32'h3c01123c),
	.w3(32'hbb8673da),
	.w4(32'hbaf6df88),
	.w5(32'h3b36d128),
	.w6(32'hbbb80151),
	.w7(32'hbb89f15a),
	.w8(32'hba8b79ef),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9761c2),
	.w1(32'hbb41f253),
	.w2(32'hbb3bc369),
	.w3(32'hb9dc3c6a),
	.w4(32'hba12e23a),
	.w5(32'hbab74fc1),
	.w6(32'hb9e1e196),
	.w7(32'hbaaec856),
	.w8(32'hbadb8b5a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb302909),
	.w1(32'hbaaf6245),
	.w2(32'hbbfe00b7),
	.w3(32'h3aa18b29),
	.w4(32'hba18d39b),
	.w5(32'hbc03143c),
	.w6(32'h3b6e3dc2),
	.w7(32'hb9bcf950),
	.w8(32'hbbc1ac44),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc184448),
	.w1(32'h3c5dde0a),
	.w2(32'hba671b15),
	.w3(32'h3a218250),
	.w4(32'h3cc32d58),
	.w5(32'h3bd4d2ab),
	.w6(32'h3b1f08c6),
	.w7(32'h3c64a3fb),
	.w8(32'h3bcd3462),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8de281),
	.w1(32'h3c0f0040),
	.w2(32'h3cf5d7ab),
	.w3(32'hbbf71596),
	.w4(32'hbc73b622),
	.w5(32'h3bf8d35b),
	.w6(32'hbc921b72),
	.w7(32'hbc770bb2),
	.w8(32'h3a54c66d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bc441),
	.w1(32'hbc43a2a2),
	.w2(32'h3bf2ac7a),
	.w3(32'hbc0d9d12),
	.w4(32'hbcb3854d),
	.w5(32'hbc1dfb71),
	.w6(32'hbc2fc905),
	.w7(32'hbc9ce7b0),
	.w8(32'hbc35e9b9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d98a2),
	.w1(32'h3b7d71db),
	.w2(32'h3bc05b61),
	.w3(32'hb990ea69),
	.w4(32'hbb308eeb),
	.w5(32'h3b54fe05),
	.w6(32'hba875479),
	.w7(32'hbb038026),
	.w8(32'h3ad1213c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea2758),
	.w1(32'hb85dcb92),
	.w2(32'h3aa980cb),
	.w3(32'hbb60c540),
	.w4(32'hbaf1ef6b),
	.w5(32'hbb22180a),
	.w6(32'h391b1649),
	.w7(32'h39c149ce),
	.w8(32'h399953ce),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba694353),
	.w1(32'h3a67632e),
	.w2(32'hbab2dac8),
	.w3(32'h38fe77e8),
	.w4(32'h39bbef18),
	.w5(32'hba9c7d93),
	.w6(32'h39f829be),
	.w7(32'h3a02c5c6),
	.w8(32'hbb3240fb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2782d8),
	.w1(32'hbb357be9),
	.w2(32'hb9d7b3c7),
	.w3(32'hbb11968d),
	.w4(32'hb90c04bc),
	.w5(32'h3bd18416),
	.w6(32'hbaf4f93b),
	.w7(32'h3a202db0),
	.w8(32'hba92e810),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd27633),
	.w1(32'hbc942d69),
	.w2(32'hbc7e06da),
	.w3(32'h3c411a85),
	.w4(32'hbb9a4868),
	.w5(32'hbc909d22),
	.w6(32'h3b9acab5),
	.w7(32'h3c1e6e3c),
	.w8(32'hbaf5a14f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c812e),
	.w1(32'h39f43322),
	.w2(32'h3bed254e),
	.w3(32'hbb82e2dd),
	.w4(32'hb98bd354),
	.w5(32'hb8f38bb5),
	.w6(32'hbb03b01c),
	.w7(32'h3b5555a1),
	.w8(32'h3b1afa7b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf89cad),
	.w1(32'h3a13c8ce),
	.w2(32'hb8e5fa12),
	.w3(32'hb9628b70),
	.w4(32'hba30726d),
	.w5(32'h3bac2d8d),
	.w6(32'h3c0b151b),
	.w7(32'h3bf5eaf5),
	.w8(32'h3c1e58e9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3068e7),
	.w1(32'hbaee1ef1),
	.w2(32'h3b80dfef),
	.w3(32'h3b125f2c),
	.w4(32'hbabf19eb),
	.w5(32'h3b6f98aa),
	.w6(32'h3b329302),
	.w7(32'h3b8c20c2),
	.w8(32'h3c13a55b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee92a5),
	.w1(32'hbc3c4143),
	.w2(32'hbcfc5fca),
	.w3(32'h3c546a2d),
	.w4(32'h3b9a559e),
	.w5(32'hbc95f12e),
	.w6(32'h3cb2b772),
	.w7(32'h3c1cf331),
	.w8(32'hbb62cab8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d2ad),
	.w1(32'hba3f9a20),
	.w2(32'hbb525753),
	.w3(32'hbb506f23),
	.w4(32'hbac87ed7),
	.w5(32'h3b9cbace),
	.w6(32'hbb0e949b),
	.w7(32'hbb32f5f6),
	.w8(32'h3bdf353c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9cd8),
	.w1(32'h3ba6a631),
	.w2(32'h3b3ba367),
	.w3(32'h3b9356d9),
	.w4(32'h3b5b1d7c),
	.w5(32'h3b3e9ec6),
	.w6(32'h3b87a566),
	.w7(32'h3b1afcee),
	.w8(32'h3a4c6519),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b866e),
	.w1(32'h3912c603),
	.w2(32'h3b1403a9),
	.w3(32'hb99c6957),
	.w4(32'h3a190e30),
	.w5(32'h3a761640),
	.w6(32'h3a52fd99),
	.w7(32'h3b1e3335),
	.w8(32'hbb2d25f7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03086c),
	.w1(32'hbba0eba3),
	.w2(32'h3a8b7a07),
	.w3(32'hb9ee4f99),
	.w4(32'hbb6fc955),
	.w5(32'h3b04a3f6),
	.w6(32'h3b737b4b),
	.w7(32'h3b32a435),
	.w8(32'hbafbcf2f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6460ff),
	.w1(32'h3a559090),
	.w2(32'hbb9269e5),
	.w3(32'hbacdc374),
	.w4(32'h3a085da6),
	.w5(32'hba8a70fd),
	.w6(32'h39f9a521),
	.w7(32'h3a39d2c4),
	.w8(32'h3a416914),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a73c3),
	.w1(32'hbca02a4e),
	.w2(32'hbd064999),
	.w3(32'h3b084abd),
	.w4(32'hba45fba7),
	.w5(32'hbc705561),
	.w6(32'h3c2febef),
	.w7(32'h3bf37f9b),
	.w8(32'hbba78af3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb480eb),
	.w1(32'hbba9046b),
	.w2(32'hbbec6d0b),
	.w3(32'hba8aa85e),
	.w4(32'hbb0a66fd),
	.w5(32'hbb0b5cff),
	.w6(32'hbb79ef08),
	.w7(32'h39a398d3),
	.w8(32'hba8ed21d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a5a4),
	.w1(32'hbb1bbc41),
	.w2(32'h39e01660),
	.w3(32'hbb7f981d),
	.w4(32'hba8d81b4),
	.w5(32'hbae29894),
	.w6(32'hbac22481),
	.w7(32'hbb3195ca),
	.w8(32'hba391911),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a07c7),
	.w1(32'hba1fb7bb),
	.w2(32'h3a334e3b),
	.w3(32'hbb41e21a),
	.w4(32'hb9b7d0b9),
	.w5(32'hb8d90d5d),
	.w6(32'hbaa2aea7),
	.w7(32'h39a2d940),
	.w8(32'hbaf72324),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63bede),
	.w1(32'hbbdd3f1f),
	.w2(32'hbb451b43),
	.w3(32'hbb3828f8),
	.w4(32'hbb9d3a4d),
	.w5(32'h3b7874ad),
	.w6(32'hbb6c6b02),
	.w7(32'hbb82ebdc),
	.w8(32'h3bcdd076),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01da09),
	.w1(32'h3c0b4b33),
	.w2(32'h3b8cf012),
	.w3(32'h3b952739),
	.w4(32'h3bb854c1),
	.w5(32'hba8e87f8),
	.w6(32'h3b966c41),
	.w7(32'h3b9313cb),
	.w8(32'hba804996),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ab3ff),
	.w1(32'hbb694e1c),
	.w2(32'hbb4cf1dd),
	.w3(32'hb8574ebe),
	.w4(32'hba1cf796),
	.w5(32'hba55cfb3),
	.w6(32'hbbc1bbc4),
	.w7(32'hbb71ef54),
	.w8(32'hba3e9e8f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb415008),
	.w1(32'hbb669fde),
	.w2(32'hbbe39b93),
	.w3(32'h3b8acdaf),
	.w4(32'h38aa94f4),
	.w5(32'hbb964a79),
	.w6(32'h3b9579f0),
	.w7(32'h3a903478),
	.w8(32'hbae8f640),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80e5dc),
	.w1(32'hbc44d2b6),
	.w2(32'hb84dc170),
	.w3(32'hba90a483),
	.w4(32'hbc03835b),
	.w5(32'h3b28e87b),
	.w6(32'hbc2e89fd),
	.w7(32'hbbe48793),
	.w8(32'hbb6aec87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78adc4),
	.w1(32'hbab25857),
	.w2(32'hba8ffb56),
	.w3(32'h39d16e17),
	.w4(32'h394aa2fb),
	.w5(32'h395c6685),
	.w6(32'hba7204bc),
	.w7(32'h39904525),
	.w8(32'hb8a20f10),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e8cc),
	.w1(32'hba475212),
	.w2(32'h3ab927f0),
	.w3(32'hbac97ee9),
	.w4(32'hb92d384f),
	.w5(32'hba4a70a8),
	.w6(32'h3a768017),
	.w7(32'h3aab8bf6),
	.w8(32'hba6367cb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3617e8),
	.w1(32'hbb144b8a),
	.w2(32'h3b18bfaf),
	.w3(32'hbaec9cc7),
	.w4(32'hb74f47d7),
	.w5(32'h3adcd19a),
	.w6(32'h3ac6308d),
	.w7(32'h3b29332b),
	.w8(32'hbb9cdc91),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268e7b),
	.w1(32'hbace1ffc),
	.w2(32'hbb21a355),
	.w3(32'h3a946110),
	.w4(32'h3ad17953),
	.w5(32'h3ae173e1),
	.w6(32'hbb127984),
	.w7(32'hba69e8fc),
	.w8(32'hb920b881),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133195),
	.w1(32'hbc9431ac),
	.w2(32'hbd0f04ff),
	.w3(32'h3c82d798),
	.w4(32'hbb902606),
	.w5(32'hbc570a04),
	.w6(32'h3c24e1cd),
	.w7(32'hba0e792e),
	.w8(32'h3bcb7c8f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78052b),
	.w1(32'h3c6ba431),
	.w2(32'hbaeb66cf),
	.w3(32'hb9138bab),
	.w4(32'hbb998d2e),
	.w5(32'hbb41cb2b),
	.w6(32'h3c2e9b71),
	.w7(32'h3bb94101),
	.w8(32'h3bf0e4fc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1100),
	.w1(32'hbc1b50eb),
	.w2(32'hbc0c82d1),
	.w3(32'hbb4b5d50),
	.w4(32'hbbad6b1b),
	.w5(32'h392c0704),
	.w6(32'hba03d2f6),
	.w7(32'h3aa6f7b4),
	.w8(32'hbbe8007f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a749e18),
	.w1(32'h3c476523),
	.w2(32'h3d0dad14),
	.w3(32'hbbba7572),
	.w4(32'hbbf803cd),
	.w5(32'h3c23850c),
	.w6(32'hbc836711),
	.w7(32'hbc2c3dd7),
	.w8(32'h3a99a68e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0912),
	.w1(32'hbacf8073),
	.w2(32'hbb0aa34b),
	.w3(32'hba5e3747),
	.w4(32'h37e1941e),
	.w5(32'hbb85ea65),
	.w6(32'hb9dead00),
	.w7(32'hb85a9987),
	.w8(32'hb9e00c90),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba81b5),
	.w1(32'hb97dbf46),
	.w2(32'hb91caa1c),
	.w3(32'h3a351ecc),
	.w4(32'hba105a0c),
	.w5(32'hbb64c517),
	.w6(32'h3ad86d5c),
	.w7(32'h3ab7c64d),
	.w8(32'h3ab4f9ae),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4959),
	.w1(32'hb8d45ce2),
	.w2(32'hbb1da54a),
	.w3(32'hbb25cf3e),
	.w4(32'hbb9b3f9e),
	.w5(32'h39b25140),
	.w6(32'hb8cfd29f),
	.w7(32'hbbb7cb34),
	.w8(32'hbb0d0d45),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11150f),
	.w1(32'hbbca2dd9),
	.w2(32'hbb45c6b2),
	.w3(32'h3b8495ae),
	.w4(32'hba83a1cc),
	.w5(32'hbaf22115),
	.w6(32'h3a061a9d),
	.w7(32'h3a4fcd22),
	.w8(32'hba45fa4b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05a5a7),
	.w1(32'hbabe0db0),
	.w2(32'hbb815926),
	.w3(32'hb858e08a),
	.w4(32'hbb7d5b0e),
	.w5(32'hbb3c983d),
	.w6(32'h3b2cc4d0),
	.w7(32'hbb8a2f17),
	.w8(32'hbafe8ecb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95f865),
	.w1(32'hbc1a2bc5),
	.w2(32'hbc6689ff),
	.w3(32'h393ce5af),
	.w4(32'h3b207586),
	.w5(32'hbb77e996),
	.w6(32'h3ba3756e),
	.w7(32'hbacd46f9),
	.w8(32'hba102a66),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c466fd1),
	.w1(32'hba93a611),
	.w2(32'hbc84c352),
	.w3(32'h3beedf10),
	.w4(32'h3c16585a),
	.w5(32'hbbe8792e),
	.w6(32'h3c6afa70),
	.w7(32'h3b3539e2),
	.w8(32'hbbf85066),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3c9d2),
	.w1(32'h3baff63d),
	.w2(32'h3c59708f),
	.w3(32'hb86128b5),
	.w4(32'hba1fbb25),
	.w5(32'h3b4870fa),
	.w6(32'h3aeb7f5d),
	.w7(32'h3b3dc562),
	.w8(32'h3b45a7e7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4c56),
	.w1(32'hbbdc8e61),
	.w2(32'hbbb65c35),
	.w3(32'hb8c03d39),
	.w4(32'hbb33fc7c),
	.w5(32'hbb0379c5),
	.w6(32'hb8d09f43),
	.w7(32'hbabadba7),
	.w8(32'hbab50fbf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b725f61),
	.w1(32'hbbaad2b0),
	.w2(32'hbc3cec08),
	.w3(32'h3ae22f45),
	.w4(32'hbb91eb23),
	.w5(32'hbc18eac9),
	.w6(32'h3b9cfa91),
	.w7(32'hb99179a5),
	.w8(32'hbb2eeb14),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb04a0d),
	.w1(32'hbb65ca47),
	.w2(32'h3a143345),
	.w3(32'h39ddbdd3),
	.w4(32'h3a819995),
	.w5(32'hbb2b202d),
	.w6(32'hbb3c6e02),
	.w7(32'h3b0145b2),
	.w8(32'hba66e380),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2d100),
	.w1(32'hbbb9b277),
	.w2(32'hbc52aa42),
	.w3(32'h3b7e2d3e),
	.w4(32'h399f77ee),
	.w5(32'hbbcdb869),
	.w6(32'h3bbe67b1),
	.w7(32'h3a9f4299),
	.w8(32'hbb52c04b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e625),
	.w1(32'hbaf75723),
	.w2(32'h39d78924),
	.w3(32'hba91d803),
	.w4(32'h3a4e773a),
	.w5(32'hba347643),
	.w6(32'hb99bcc16),
	.w7(32'h3a5bc60c),
	.w8(32'h3b1096ef),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf345),
	.w1(32'h3b8b1343),
	.w2(32'h3ad007ab),
	.w3(32'h394a96a5),
	.w4(32'hb9f95c4e),
	.w5(32'hbaadd044),
	.w6(32'h3b80c2d0),
	.w7(32'h3a474a97),
	.w8(32'hba8c408a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac821eb),
	.w1(32'hbb123336),
	.w2(32'hba8fae2c),
	.w3(32'h39aad5d9),
	.w4(32'h385478e2),
	.w5(32'hbb70f87d),
	.w6(32'hba892daa),
	.w7(32'hba5147bd),
	.w8(32'hbb48720d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44134),
	.w1(32'hbb9dcff8),
	.w2(32'hbb534319),
	.w3(32'hbbc94575),
	.w4(32'hbb3f3df7),
	.w5(32'h3acbd5d3),
	.w6(32'hbb3af39e),
	.w7(32'hbb22e251),
	.w8(32'h3b4780cc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87202c),
	.w1(32'h3bd06dbc),
	.w2(32'h3c20836c),
	.w3(32'hbb5622ac),
	.w4(32'hbb347e95),
	.w5(32'h3b3013d5),
	.w6(32'hbb671877),
	.w7(32'hbb348435),
	.w8(32'h3b274740),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a258f5e),
	.w1(32'h3a4faa41),
	.w2(32'h3a2e8012),
	.w3(32'h3ab35be6),
	.w4(32'h3b0cffff),
	.w5(32'h3bab9d67),
	.w6(32'hba1ead19),
	.w7(32'h39dcdb03),
	.w8(32'h3b9249ab),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983f39),
	.w1(32'h3c56ce50),
	.w2(32'h3c53d27b),
	.w3(32'h3baa9a52),
	.w4(32'h3ba7dd72),
	.w5(32'hbae76d34),
	.w6(32'h3bfb33ee),
	.w7(32'h3be8f76f),
	.w8(32'h3b97cd85),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61fb89),
	.w1(32'hbc12d0ce),
	.w2(32'hbcab861c),
	.w3(32'hbb08a825),
	.w4(32'hbbce2d0a),
	.w5(32'hbc01f483),
	.w6(32'h3bf64eca),
	.w7(32'hbb2ad27f),
	.w8(32'hba92b860),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85870f),
	.w1(32'h3a4a9141),
	.w2(32'h3b466f42),
	.w3(32'hbbdd3be8),
	.w4(32'hbbebcab4),
	.w5(32'hbb5a838f),
	.w6(32'hbaad9421),
	.w7(32'hba346e9d),
	.w8(32'hb9a34d10),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2f07),
	.w1(32'hbc2c8ea9),
	.w2(32'hbce8dfa5),
	.w3(32'h3b9a1a3a),
	.w4(32'h3b448ea1),
	.w5(32'hbc3fe5f1),
	.w6(32'h3c039534),
	.w7(32'hba402135),
	.w8(32'h3b055152),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea3c9e),
	.w1(32'h3b2a5247),
	.w2(32'h3bc6a0ba),
	.w3(32'hbb0f52c2),
	.w4(32'hbad32fe7),
	.w5(32'h3b166359),
	.w6(32'hbbb4cea9),
	.w7(32'hbba37645),
	.w8(32'h3b10dcf2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072883),
	.w1(32'hbc948160),
	.w2(32'hbc5355c0),
	.w3(32'h3a8c1bd4),
	.w4(32'hbc1dbdde),
	.w5(32'hbbc33cdd),
	.w6(32'h3bb1c166),
	.w7(32'hbba1415b),
	.w8(32'hbba6391b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f0cd),
	.w1(32'hbb9bbf87),
	.w2(32'hbc2fc6ca),
	.w3(32'hbb81ea80),
	.w4(32'hbc168a36),
	.w5(32'hbb90ade0),
	.w6(32'h3ab99b86),
	.w7(32'hbaafee1f),
	.w8(32'h3abea6a4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b3f94),
	.w1(32'h3ab1323e),
	.w2(32'h3c425b46),
	.w3(32'hbbb9535b),
	.w4(32'hbc093789),
	.w5(32'h3b88d1c7),
	.w6(32'hbb9d75f1),
	.w7(32'hbb837cd2),
	.w8(32'h3b97ae44),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e9603),
	.w1(32'hb8155da7),
	.w2(32'h3b9b3e73),
	.w3(32'hbaee993f),
	.w4(32'hba7e8edd),
	.w5(32'hbba4362d),
	.w6(32'hbb82f821),
	.w7(32'hbada9ccd),
	.w8(32'hbb8e8064),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d6f7),
	.w1(32'hbba40e6c),
	.w2(32'hbc89dffc),
	.w3(32'h3b7da3f2),
	.w4(32'h3a873af9),
	.w5(32'hbbbca0ab),
	.w6(32'h3c1d9e4f),
	.w7(32'h3bc0ba02),
	.w8(32'hbadba547),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3b5a2),
	.w1(32'hbbe566ad),
	.w2(32'hbca2da87),
	.w3(32'h3c1545af),
	.w4(32'h3b6e68ca),
	.w5(32'hbc289f98),
	.w6(32'h3c36f261),
	.w7(32'h3ad90f76),
	.w8(32'h3a13007e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94a5fd),
	.w1(32'h3c769dc8),
	.w2(32'h3c20b111),
	.w3(32'hbbc51780),
	.w4(32'h3a9928c8),
	.w5(32'hbae2892d),
	.w6(32'h3b515b5e),
	.w7(32'h3b8e0ca1),
	.w8(32'h3c1f84cd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620f3d),
	.w1(32'h3c3c7927),
	.w2(32'h3cdc4666),
	.w3(32'hbc61e25c),
	.w4(32'hbb74202e),
	.w5(32'h3c55a2d2),
	.w6(32'hbc359c03),
	.w7(32'hbb3f9ad1),
	.w8(32'h3c40d0dc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a768d),
	.w1(32'h3c2cd7d7),
	.w2(32'h3c843182),
	.w3(32'hb9e84c1d),
	.w4(32'h3b75184c),
	.w5(32'h3c110fc1),
	.w6(32'hbae76651),
	.w7(32'h3a772b36),
	.w8(32'h3bc0f161),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24684e),
	.w1(32'hbbaa5ba6),
	.w2(32'hbc5636d1),
	.w3(32'hbad178f9),
	.w4(32'h3c184cb7),
	.w5(32'hbbbe4fed),
	.w6(32'h3c5194f4),
	.w7(32'h3bac1c33),
	.w8(32'hba816910),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b348b),
	.w1(32'h3ae9f18b),
	.w2(32'h3ab5bc7f),
	.w3(32'h3ae1cdcc),
	.w4(32'h3ac58c19),
	.w5(32'h3aac3791),
	.w6(32'h3aa6e3e5),
	.w7(32'h3ac3a86e),
	.w8(32'h3aea89e5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85522e),
	.w1(32'hbade9b5e),
	.w2(32'h3c51672c),
	.w3(32'hbc08c006),
	.w4(32'h3c251386),
	.w5(32'h37fbea9c),
	.w6(32'h3c821d13),
	.w7(32'h3bbeda2d),
	.w8(32'h3c36d618),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7cfb5),
	.w1(32'hbbbdfce2),
	.w2(32'hbc2c66ee),
	.w3(32'hba59d19b),
	.w4(32'hbb2bb88d),
	.w5(32'hbbe709c9),
	.w6(32'h3aba5121),
	.w7(32'hbb6b9bb7),
	.w8(32'hbc02d746),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d166c6),
	.w1(32'h3943d7d5),
	.w2(32'h39c49d25),
	.w3(32'hb8c1485b),
	.w4(32'hb91bf657),
	.w5(32'h39903266),
	.w6(32'h3807dccb),
	.w7(32'hb87acbb7),
	.w8(32'h394f2e04),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be023),
	.w1(32'h3afbc701),
	.w2(32'h39e4e2e2),
	.w3(32'hbadc56ea),
	.w4(32'hbb0c1ff5),
	.w5(32'hbaf90df2),
	.w6(32'hbb404b58),
	.w7(32'hba069ba2),
	.w8(32'hba8174c8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efc3a),
	.w1(32'hbb79617c),
	.w2(32'hbc0c7611),
	.w3(32'h3be2cdbb),
	.w4(32'h3b044d52),
	.w5(32'hbba4f669),
	.w6(32'h3c0865c7),
	.w7(32'h3b85bc4e),
	.w8(32'hb96a145e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed3f54),
	.w1(32'h3b9524f3),
	.w2(32'h3c2bb5bd),
	.w3(32'hba44749f),
	.w4(32'hb9e0e573),
	.w5(32'h3b70e2e9),
	.w6(32'h389de112),
	.w7(32'h3a134e5b),
	.w8(32'h3b52d19f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f008f),
	.w1(32'hbc6ce54f),
	.w2(32'hbb99ec5b),
	.w3(32'hba02984a),
	.w4(32'hbc42beb8),
	.w5(32'hbc135ac4),
	.w6(32'hbb9ca64f),
	.w7(32'hbc1d563d),
	.w8(32'hbbc65993),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad693af),
	.w1(32'h3b6be4b5),
	.w2(32'h3c2c62a0),
	.w3(32'hbb10f1bf),
	.w4(32'hba8547c7),
	.w5(32'h3b5f9212),
	.w6(32'hbafb6cfd),
	.w7(32'hba075772),
	.w8(32'h3aeacffc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb5ef),
	.w1(32'h3c8217cb),
	.w2(32'h3c3b74f7),
	.w3(32'hbb73b724),
	.w4(32'h3c1ef119),
	.w5(32'h3c0a499f),
	.w6(32'h3a5acdfa),
	.w7(32'h3b9aeac9),
	.w8(32'h3c0ad345),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d9f56),
	.w1(32'hbc34c358),
	.w2(32'hbbd156f9),
	.w3(32'hbb98f2ed),
	.w4(32'hbc31381c),
	.w5(32'hbbc5e2b0),
	.w6(32'hba1e373f),
	.w7(32'h3b44c750),
	.w8(32'h3b803a1d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3ad4),
	.w1(32'h3a8b409f),
	.w2(32'h3b35d786),
	.w3(32'h3a8ad3f5),
	.w4(32'h3a9b8279),
	.w5(32'h3b1c16fb),
	.w6(32'h3b377f9e),
	.w7(32'h3b4318f2),
	.w8(32'h3b4e736c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ee06a),
	.w1(32'hb89627ab),
	.w2(32'h3815abff),
	.w3(32'hb9a4d625),
	.w4(32'hb927bc28),
	.w5(32'hb7ee8e5a),
	.w6(32'hb987aa4a),
	.w7(32'hb7ef88b4),
	.w8(32'h3851b75e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7ad82),
	.w1(32'hb9e39168),
	.w2(32'h398aa706),
	.w3(32'hba16358a),
	.w4(32'hb9400a23),
	.w5(32'hb9ff0f6a),
	.w6(32'hbad0a8d0),
	.w7(32'hba30915b),
	.w8(32'hb9725248),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38949e5d),
	.w1(32'h382e3267),
	.w2(32'h37255e98),
	.w3(32'h38aa67eb),
	.w4(32'h388d8577),
	.w5(32'h38a19fa8),
	.w6(32'hb7fc8de0),
	.w7(32'hb81fe608),
	.w8(32'h37221896),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce1676),
	.w1(32'h3a0b588b),
	.w2(32'h3a1090ec),
	.w3(32'h39c3b2ea),
	.w4(32'h39e076c8),
	.w5(32'h3a030418),
	.w6(32'h359ca2dc),
	.w7(32'hb7b6de7f),
	.w8(32'h37650216),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a7a55),
	.w1(32'h3ad1adfa),
	.w2(32'h3b831e07),
	.w3(32'h3abe9c31),
	.w4(32'h3b26eff6),
	.w5(32'h3b79b08d),
	.w6(32'h3b5d97b5),
	.w7(32'h3b8d6973),
	.w8(32'h3b8d2e22),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa499e8),
	.w1(32'hba94f032),
	.w2(32'hb9d2328d),
	.w3(32'hba92e732),
	.w4(32'hba850127),
	.w5(32'hb9ff323f),
	.w6(32'hba3334e0),
	.w7(32'hb92f762b),
	.w8(32'hb9f38f02),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1176a5),
	.w1(32'hbb1862d0),
	.w2(32'hbc0caabb),
	.w3(32'h3b7c645b),
	.w4(32'h3bc21124),
	.w5(32'hbaf462d2),
	.w6(32'h3bb9f735),
	.w7(32'h3b8190fc),
	.w8(32'h3ae49a9e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9404),
	.w1(32'h3c2a6ff7),
	.w2(32'h3cd5d8a1),
	.w3(32'hba863b58),
	.w4(32'hbb6791d6),
	.w5(32'h3c0c82f9),
	.w6(32'hbc00ad8b),
	.w7(32'hbbf9ec65),
	.w8(32'hb97e3ec4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843f9bd),
	.w1(32'h3910dfe1),
	.w2(32'h3905f633),
	.w3(32'hb821aadb),
	.w4(32'hb743354e),
	.w5(32'hb65b2603),
	.w6(32'hb8073fc7),
	.w7(32'hb8748bf9),
	.w8(32'h37eea39f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d68373),
	.w1(32'h38865d04),
	.w2(32'hb83b4548),
	.w3(32'h3910f9ca),
	.w4(32'h3902e77a),
	.w5(32'hb88cafa5),
	.w6(32'h386d9458),
	.w7(32'hb716ffd5),
	.w8(32'hb906c1ad),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809979f),
	.w1(32'hb34dc714),
	.w2(32'hb6e0925b),
	.w3(32'h37d72005),
	.w4(32'h37b1064d),
	.w5(32'h37e413af),
	.w6(32'hb7d8efe9),
	.w7(32'hb83db10b),
	.w8(32'hb74cf4ac),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b8f6a),
	.w1(32'h3a055346),
	.w2(32'h3a07ff89),
	.w3(32'h3a0ccfc3),
	.w4(32'h3a3e43ec),
	.w5(32'h3a13e5ea),
	.w6(32'h39bd3509),
	.w7(32'h39de1787),
	.w8(32'h39cc2ecb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92251d),
	.w1(32'h3c1f8174),
	.w2(32'hbc692460),
	.w3(32'hba0932ce),
	.w4(32'hbc064c15),
	.w5(32'hbc114d16),
	.w6(32'h3bf64a6d),
	.w7(32'hbba81ddc),
	.w8(32'hbc01aff3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7774),
	.w1(32'hbc1b4fde),
	.w2(32'hbc9c01be),
	.w3(32'h3b5f7090),
	.w4(32'hbb9204f1),
	.w5(32'hbc1ca91b),
	.w6(32'h3bdb179b),
	.w7(32'h3a861f77),
	.w8(32'hbb244b4e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00665d),
	.w1(32'hbb14c1cd),
	.w2(32'hbb4d8ed3),
	.w3(32'h3ae03675),
	.w4(32'h3a178e1a),
	.w5(32'hbb136126),
	.w6(32'h3b130271),
	.w7(32'h37ef1aaa),
	.w8(32'hb9866473),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f716),
	.w1(32'h3a01ea67),
	.w2(32'hbaffc690),
	.w3(32'hbb2d6098),
	.w4(32'hba8f010b),
	.w5(32'hb9babcaa),
	.w6(32'hbb122653),
	.w7(32'hbb1da744),
	.w8(32'hbacb918a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11ec18),
	.w1(32'h3a79455f),
	.w2(32'h3b0b6ff4),
	.w3(32'hba0001ce),
	.w4(32'hb917c0a1),
	.w5(32'h3a9f434b),
	.w6(32'h3a71bb4a),
	.w7(32'h3ae3fe61),
	.w8(32'h3b027fd1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba920244),
	.w1(32'hbb147e19),
	.w2(32'hbad89417),
	.w3(32'h3b4b53b8),
	.w4(32'hba3aeaea),
	.w5(32'hba321441),
	.w6(32'h3b66d4e7),
	.w7(32'h3ad612ab),
	.w8(32'h3a8295c5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c672),
	.w1(32'hbb6c1233),
	.w2(32'h3b7249c0),
	.w3(32'hbb198337),
	.w4(32'hbbb89aac),
	.w5(32'hb9b770e4),
	.w6(32'hb927b7bb),
	.w7(32'h3ab3f54a),
	.w8(32'h3b04745e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5f6f),
	.w1(32'hbc41d971),
	.w2(32'hbcdffe44),
	.w3(32'h3c28f872),
	.w4(32'h3b34b8a4),
	.w5(32'hbc4b99ee),
	.w6(32'h3c00b50a),
	.w7(32'h3b207cae),
	.w8(32'hbb8a46af),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4870b8),
	.w1(32'h3bced47c),
	.w2(32'h3c41fa4d),
	.w3(32'hbac81fd1),
	.w4(32'hbac88db9),
	.w5(32'h3b59fb9f),
	.w6(32'hbb2d89c2),
	.w7(32'hba8af89b),
	.w8(32'h3ac7be74),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab006c8),
	.w1(32'hbafd05ba),
	.w2(32'hbc088cd7),
	.w3(32'h3aedd434),
	.w4(32'h39a46818),
	.w5(32'hbba444a5),
	.w6(32'h3bb390b2),
	.w7(32'h3b8634f4),
	.w8(32'h3a0814a9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0ff8),
	.w1(32'hbbfaab3b),
	.w2(32'hbc81fc03),
	.w3(32'h3be26677),
	.w4(32'h3b96c137),
	.w5(32'hbc277083),
	.w6(32'h3c4303fd),
	.w7(32'h3be17932),
	.w8(32'hb979f3af),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d640c),
	.w1(32'h3c0ef426),
	.w2(32'h3c17f4d1),
	.w3(32'hb50cd620),
	.w4(32'h3b993fb9),
	.w5(32'h3bcd04f9),
	.w6(32'h3a97f20d),
	.w7(32'h3b8d0ba0),
	.w8(32'h3bd1e39c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7823),
	.w1(32'hbbb1c41a),
	.w2(32'hbc082bfd),
	.w3(32'h3b2cd664),
	.w4(32'h3a68d708),
	.w5(32'hbb4e54f4),
	.w6(32'h3b9cc0db),
	.w7(32'h3a732c34),
	.w8(32'hb914f341),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a287a1),
	.w1(32'h39e62898),
	.w2(32'h3a2a6c6c),
	.w3(32'h397311b6),
	.w4(32'h3a027b79),
	.w5(32'h3a13ca9e),
	.w6(32'h3a7744ae),
	.w7(32'h3a85e0d6),
	.w8(32'h3a4e62f5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071bab),
	.w1(32'h3bb6af2f),
	.w2(32'h3cb24693),
	.w3(32'h374d349c),
	.w4(32'hbc2632ca),
	.w5(32'h3bc106b4),
	.w6(32'h3a8504fd),
	.w7(32'hbc09d927),
	.w8(32'h3b6423fa),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9754f),
	.w1(32'hb96a9883),
	.w2(32'h3a254079),
	.w3(32'hba31d70a),
	.w4(32'hba3f87ea),
	.w5(32'h3a8ae161),
	.w6(32'h3a229f8b),
	.w7(32'hba099fd8),
	.w8(32'h3a2c3c54),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985d861),
	.w1(32'h38dce13a),
	.w2(32'hb8b2316c),
	.w3(32'h372b445a),
	.w4(32'hb99fec43),
	.w5(32'hb9a11e39),
	.w6(32'h39b850fc),
	.w7(32'hb8871a8c),
	.w8(32'h38685ec4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a0a51),
	.w1(32'hb87e07eb),
	.w2(32'h37e31d2d),
	.w3(32'h38fea7a5),
	.w4(32'h399bf5d2),
	.w5(32'h390c90fe),
	.w6(32'hb82b9daf),
	.w7(32'hb84426c3),
	.w8(32'h394b6487),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f8c74),
	.w1(32'hba44217b),
	.w2(32'hb9b108c1),
	.w3(32'hba194b59),
	.w4(32'h394006c7),
	.w5(32'h3a042dbf),
	.w6(32'h3b13f2b3),
	.w7(32'h3a7839d7),
	.w8(32'h3afd252d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b66d),
	.w1(32'h3b7e96a2),
	.w2(32'h3c2d0103),
	.w3(32'hba8563c9),
	.w4(32'h39abe772),
	.w5(32'h3b1bbc77),
	.w6(32'hbbca94c4),
	.w7(32'hbb4c4199),
	.w8(32'h3acb61a5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a925f7e),
	.w1(32'hbb2e208b),
	.w2(32'hbb568750),
	.w3(32'h3b5a0850),
	.w4(32'h3a0f2759),
	.w5(32'hbab8ba71),
	.w6(32'h3bea08eb),
	.w7(32'h3b7a32fb),
	.w8(32'h3a95de92),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ff97a),
	.w1(32'hb8dd8086),
	.w2(32'h3890d713),
	.w3(32'hb8f04b1a),
	.w4(32'hb90a8a45),
	.w5(32'h388fe2bd),
	.w6(32'hb9166816),
	.w7(32'hb8b95c75),
	.w8(32'h39190279),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d838),
	.w1(32'hbc0c5a5c),
	.w2(32'hbc1bba3b),
	.w3(32'h3b3c99e3),
	.w4(32'hba06725a),
	.w5(32'hbbb2054c),
	.w6(32'h3b7e37ee),
	.w7(32'h3a01a80e),
	.w8(32'hbaa80fdd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b276b0d),
	.w1(32'h3ad68844),
	.w2(32'h3a995160),
	.w3(32'h3b2f0683),
	.w4(32'h3ab8e919),
	.w5(32'h3aa3d940),
	.w6(32'h3b6d703e),
	.w7(32'h3b19ec00),
	.w8(32'h3ab7c841),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8cc8a),
	.w1(32'hbbf0c21e),
	.w2(32'hbc8b3d83),
	.w3(32'h3c5e7e92),
	.w4(32'h3c0d7de0),
	.w5(32'hbbab16e8),
	.w6(32'h3c650f50),
	.w7(32'h3bd9c199),
	.w8(32'h3b1838a6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338ab8),
	.w1(32'hbc30b9d0),
	.w2(32'h3a82748f),
	.w3(32'h3c0bc675),
	.w4(32'hbc244059),
	.w5(32'hbc27dc0e),
	.w6(32'hbc4b8a43),
	.w7(32'hbc35f0fc),
	.w8(32'hbbf7666b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56dbfa),
	.w1(32'h3afa9014),
	.w2(32'h3b9f8391),
	.w3(32'hbaea167a),
	.w4(32'hbb38c578),
	.w5(32'h3a623e02),
	.w6(32'hbb85a0db),
	.w7(32'hbb903b68),
	.w8(32'hba473744),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f402b),
	.w1(32'h3b2b6e32),
	.w2(32'h3b11b6a9),
	.w3(32'h3b158d2c),
	.w4(32'h3b19249f),
	.w5(32'h3b0f04c7),
	.w6(32'h3b0122b7),
	.w7(32'h3b07c1b5),
	.w8(32'h3af78990),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c8e19),
	.w1(32'h3b655b50),
	.w2(32'h3bbc2644),
	.w3(32'hbad784bc),
	.w4(32'h3a82aada),
	.w5(32'h3b4a845b),
	.w6(32'hba580564),
	.w7(32'h3ade8bf7),
	.w8(32'h3b721908),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9362f0),
	.w1(32'hbaf1a53d),
	.w2(32'h3b895eca),
	.w3(32'hbb99115a),
	.w4(32'hbb4bfc36),
	.w5(32'h3b0c63bb),
	.w6(32'hb9bd2533),
	.w7(32'h3ab19a4b),
	.w8(32'h3b8e05e3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b417a59),
	.w1(32'h3bc96077),
	.w2(32'h3c25aa27),
	.w3(32'h399c7b5d),
	.w4(32'h3ac6e3b4),
	.w5(32'h3b69a5ab),
	.w6(32'hbb154bb1),
	.w7(32'hb803f859),
	.w8(32'h3b13e725),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74e7afc),
	.w1(32'hbb399bd1),
	.w2(32'hbb892ae3),
	.w3(32'h3b13850d),
	.w4(32'h3a45947b),
	.w5(32'hbb58b995),
	.w6(32'h3b38b379),
	.w7(32'hb990e37d),
	.w8(32'hbab2607f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a164d),
	.w1(32'hb91e0c2c),
	.w2(32'h39d6100d),
	.w3(32'h384dc8e1),
	.w4(32'h387c3d57),
	.w5(32'h398a8f13),
	.w6(32'hb9d01290),
	.w7(32'h39891854),
	.w8(32'h38b7064a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a993502),
	.w1(32'hbba640df),
	.w2(32'hbc0c9a95),
	.w3(32'h3b3d6892),
	.w4(32'h3a82bf64),
	.w5(32'hbb986d08),
	.w6(32'h3bf22e18),
	.w7(32'h3ac3c103),
	.w8(32'hbab3252f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cab66),
	.w1(32'hbb4b1f7f),
	.w2(32'hbb7308c2),
	.w3(32'h3aed8c9e),
	.w4(32'hba6569ee),
	.w5(32'hbafb28a2),
	.w6(32'h3b1f6148),
	.w7(32'hba90147f),
	.w8(32'hba7e536a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11a3b9),
	.w1(32'h3b30cabc),
	.w2(32'h3be2bf2a),
	.w3(32'hbb973ec5),
	.w4(32'hbb7cdcf7),
	.w5(32'h3b7fcc6f),
	.w6(32'hbb6ad755),
	.w7(32'hba968f05),
	.w8(32'h3b487148),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39826aba),
	.w1(32'h3939830f),
	.w2(32'h388288a8),
	.w3(32'hb8e1e3af),
	.w4(32'h39338d75),
	.w5(32'hb71f5bb8),
	.w6(32'hb9c070b5),
	.w7(32'hb92a3db5),
	.w8(32'hb9663131),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71a307),
	.w1(32'h3c17273e),
	.w2(32'hb73c6e60),
	.w3(32'h3a8bd737),
	.w4(32'hbaaabfec),
	.w5(32'hbb76226d),
	.w6(32'h3b05e530),
	.w7(32'hbba73756),
	.w8(32'hbb905fce),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb14b3),
	.w1(32'h38ebe5e2),
	.w2(32'h392ebd5c),
	.w3(32'h38fd7ce4),
	.w4(32'h3944d12f),
	.w5(32'h391f0382),
	.w6(32'h385cc20e),
	.w7(32'h3949d936),
	.w8(32'h3932c10c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37850023),
	.w1(32'hb980c7a3),
	.w2(32'hba31c5eb),
	.w3(32'hb8e48d01),
	.w4(32'hb9c1d0d0),
	.w5(32'hba5e03e4),
	.w6(32'hb9a5877f),
	.w7(32'hb9dc5659),
	.w8(32'hba6ceb42),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebe0ee),
	.w1(32'h3a1e2691),
	.w2(32'h3bd11a07),
	.w3(32'hbb4301e5),
	.w4(32'hbaf5d549),
	.w5(32'h3b4bbc7a),
	.w6(32'hbaf121af),
	.w7(32'h39bf856e),
	.w8(32'h3b24598b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29a2d2),
	.w1(32'h3b47d704),
	.w2(32'hbc3c29ac),
	.w3(32'h3b98449c),
	.w4(32'h3b0cb655),
	.w5(32'hbb64108e),
	.w6(32'h3c668a5d),
	.w7(32'h3b19863e),
	.w8(32'h392aa4da),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc74b5),
	.w1(32'h3ae6ef50),
	.w2(32'h39e4b373),
	.w3(32'h3a818606),
	.w4(32'h3a8fecf1),
	.w5(32'h382a3662),
	.w6(32'h3a2897c6),
	.w7(32'h3a7cddbd),
	.w8(32'h39d639d3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a1b5),
	.w1(32'h3b8e9755),
	.w2(32'h3c169c03),
	.w3(32'hbae1b44a),
	.w4(32'hba977bcb),
	.w5(32'h3b232891),
	.w6(32'hba731d16),
	.w7(32'h3992cdcb),
	.w8(32'h3a3a74d7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba318fcf),
	.w1(32'hbba9c836),
	.w2(32'hbbc8497a),
	.w3(32'hbaa4cb6a),
	.w4(32'hbbbc366e),
	.w5(32'hbc1c2616),
	.w6(32'hbb622b05),
	.w7(32'hbb1edbcf),
	.w8(32'hbb404bc6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ab704),
	.w1(32'hbc7a3bd0),
	.w2(32'hbc704d2e),
	.w3(32'h3c01c206),
	.w4(32'hbbac9535),
	.w5(32'hbb951ccc),
	.w6(32'hb9a87244),
	.w7(32'h3b694c68),
	.w8(32'h3a437d19),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb240fe9),
	.w1(32'hbc2bc90d),
	.w2(32'hbc238229),
	.w3(32'h3ae922e9),
	.w4(32'hba88bb33),
	.w5(32'hbb69e9c7),
	.w6(32'h3b859c9d),
	.w7(32'h3ae3eefe),
	.w8(32'hb8934362),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ca44c),
	.w1(32'hbbd21eaa),
	.w2(32'hbc6828aa),
	.w3(32'h3b89f249),
	.w4(32'hb986bf77),
	.w5(32'hbbd7da90),
	.w6(32'h3bebfb87),
	.w7(32'h3b2f31a1),
	.w8(32'hbb38553a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8289838),
	.w1(32'h39b32062),
	.w2(32'h3a05d3e3),
	.w3(32'h3948c359),
	.w4(32'h3a119d0d),
	.w5(32'h3a309a23),
	.w6(32'h39499587),
	.w7(32'h3a836cfc),
	.w8(32'h3a73163e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0801),
	.w1(32'hbbe5585f),
	.w2(32'hbb9b3afa),
	.w3(32'h3a87611d),
	.w4(32'hbb855de6),
	.w5(32'hbb265000),
	.w6(32'h3af84c3a),
	.w7(32'h3a690f41),
	.w8(32'hb7b1c360),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad9f64),
	.w1(32'hb791a1a4),
	.w2(32'hb6a479c6),
	.w3(32'h379eb09d),
	.w4(32'hb7fd6798),
	.w5(32'h36cb1536),
	.w6(32'h38067609),
	.w7(32'hb67749ad),
	.w8(32'hb61b2d11),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8436ace),
	.w1(32'hba4f181c),
	.w2(32'hba3c30dd),
	.w3(32'h39023a78),
	.w4(32'h39c0448d),
	.w5(32'h38abef68),
	.w6(32'h39d7fbee),
	.w7(32'h39603bf7),
	.w8(32'h39df7d39),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1bab9),
	.w1(32'h3af3c714),
	.w2(32'h3b0c6716),
	.w3(32'hb76fc350),
	.w4(32'hb9bcf576),
	.w5(32'hb88ba999),
	.w6(32'hba8aa4a9),
	.w7(32'hbaccfaa0),
	.w8(32'hba8c289e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc380c1),
	.w1(32'hbc1066bf),
	.w2(32'hbc01c6db),
	.w3(32'h3ad11332),
	.w4(32'hbb1c4882),
	.w5(32'hbaf1992a),
	.w6(32'h3ad7d809),
	.w7(32'h3b01dacb),
	.w8(32'h3b561a5a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79425e1),
	.w1(32'h38bdb3af),
	.w2(32'h377bdac5),
	.w3(32'hb7b03e9b),
	.w4(32'hb77f5aa9),
	.w5(32'h381a8662),
	.w6(32'hb4e76b6e),
	.w7(32'hb856834d),
	.w8(32'h37914031),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8484f3c),
	.w1(32'hb82517d3),
	.w2(32'hb7416439),
	.w3(32'h38483cdf),
	.w4(32'h3855229b),
	.w5(32'h38105139),
	.w6(32'hb6f6b17e),
	.w7(32'h3870943e),
	.w8(32'h38248a16),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d71dc),
	.w1(32'h3b694f13),
	.w2(32'h3b83ea89),
	.w3(32'h3a03a605),
	.w4(32'hbb360ca2),
	.w5(32'hb9178c97),
	.w6(32'hba930b5b),
	.w7(32'hba8934e4),
	.w8(32'h3aaf3ea5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c491),
	.w1(32'hbb704def),
	.w2(32'hbc766efd),
	.w3(32'hb85cfa7a),
	.w4(32'hbaed890b),
	.w5(32'hbbd5b357),
	.w6(32'hba2936fa),
	.w7(32'h3a2757bc),
	.w8(32'hbbde54f8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb950e6c),
	.w1(32'h3b4c4fa5),
	.w2(32'h39e9a125),
	.w3(32'hbbee0ef3),
	.w4(32'h3b78fb33),
	.w5(32'hbaa671b0),
	.w6(32'hbb38dd74),
	.w7(32'hba3a0210),
	.w8(32'h3adbcf63),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4e197),
	.w1(32'hba9a20c5),
	.w2(32'hba441c58),
	.w3(32'hba3f423e),
	.w4(32'hba23300e),
	.w5(32'hba94c727),
	.w6(32'hba6ed8c7),
	.w7(32'hba84e125),
	.w8(32'hba8ff1a3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90f95),
	.w1(32'hbbcd1840),
	.w2(32'hbca513ea),
	.w3(32'h3c1b8945),
	.w4(32'hba13b2af),
	.w5(32'hbc2359a9),
	.w6(32'h3c64f8b7),
	.w7(32'h3be6585b),
	.w8(32'hbb8dd437),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9edb45),
	.w1(32'hbc4dc478),
	.w2(32'h3b9ddcf8),
	.w3(32'h3b98a208),
	.w4(32'hbc6d52f9),
	.w5(32'hbc229f39),
	.w6(32'hbab87675),
	.w7(32'h399e57b9),
	.w8(32'h3bf4feef),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8082e),
	.w1(32'hbaba7579),
	.w2(32'hbbf591b2),
	.w3(32'h3b96ba2a),
	.w4(32'h3b272e73),
	.w5(32'hbb70fc1f),
	.w6(32'h3b525ce7),
	.w7(32'hba7a7e68),
	.w8(32'hbb8307e8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3bd7a),
	.w1(32'hb8af6911),
	.w2(32'hb8a54d77),
	.w3(32'hb711f242),
	.w4(32'hb7dcde52),
	.w5(32'hb8570671),
	.w6(32'hb9254ddc),
	.w7(32'hb9265442),
	.w8(32'hb8c85a0e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939c210),
	.w1(32'hb8d0d5d8),
	.w2(32'hb8138ec3),
	.w3(32'hb8eb2544),
	.w4(32'hb8a18400),
	.w5(32'h373d06c3),
	.w6(32'hb90d1702),
	.w7(32'hb8bd41cd),
	.w8(32'hb680d826),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894d85d),
	.w1(32'hb6b10c30),
	.w2(32'hb690fe6e),
	.w3(32'h376d48ff),
	.w4(32'h37cf8fcd),
	.w5(32'hb7079384),
	.w6(32'hb738c68c),
	.w7(32'h3619af75),
	.w8(32'hb7eeb4d9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fde6),
	.w1(32'h3b3c8168),
	.w2(32'hbc06ebe5),
	.w3(32'h3a0e98cd),
	.w4(32'h3b04e9d2),
	.w5(32'hbbc11e0f),
	.w6(32'h3b90711f),
	.w7(32'hbab5d968),
	.w8(32'hbb7d4875),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e50fc),
	.w1(32'hba906a6f),
	.w2(32'hbb762de2),
	.w3(32'h3b23f2d3),
	.w4(32'hba9bc060),
	.w5(32'hbb0f6e07),
	.w6(32'h3ba162e3),
	.w7(32'h3a9a2d8c),
	.w8(32'hb9c63f2a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7db95e),
	.w1(32'h3c2916e6),
	.w2(32'h3c7be4de),
	.w3(32'hbb68a7a7),
	.w4(32'h3b3c9c5f),
	.w5(32'h3bffb37a),
	.w6(32'hbb264032),
	.w7(32'h3a3788bc),
	.w8(32'h3b7aded0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982c41e),
	.w1(32'h3a850f47),
	.w2(32'h3af53181),
	.w3(32'hba278da2),
	.w4(32'hb8a6f1dc),
	.w5(32'h3aaa6099),
	.w6(32'hba29ffce),
	.w7(32'hb8583b77),
	.w8(32'h3a5cfe93),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adec25d),
	.w1(32'hbb74aba9),
	.w2(32'hbc2cc29a),
	.w3(32'h3bd2ef71),
	.w4(32'h3b025fab),
	.w5(32'hbbfeb594),
	.w6(32'h3c1903f1),
	.w7(32'h3b98dbf3),
	.w8(32'hbb105d25),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb05a),
	.w1(32'h3a87b5be),
	.w2(32'hbac681c8),
	.w3(32'hbb47935d),
	.w4(32'h3ab74c7b),
	.w5(32'hb97c0c8b),
	.w6(32'hbb4b0d6f),
	.w7(32'h3927a744),
	.w8(32'h37145887),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37847075),
	.w1(32'h3887e0f7),
	.w2(32'h38c33904),
	.w3(32'hb7ce41e2),
	.w4(32'h3823887d),
	.w5(32'h387addd2),
	.w6(32'hb7cc896e),
	.w7(32'h3800a733),
	.w8(32'h388d351c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f91c),
	.w1(32'hbb93fdd2),
	.w2(32'h39dba497),
	.w3(32'hbbbb9869),
	.w4(32'hbafaca14),
	.w5(32'hbaf20b18),
	.w6(32'hbb2f68d0),
	.w7(32'h3908c499),
	.w8(32'h3b867de3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34e6382d),
	.w1(32'h38484fe0),
	.w2(32'h3909d9ee),
	.w3(32'hb83e33dc),
	.w4(32'hb593f8a2),
	.w5(32'h38977875),
	.w6(32'hb8a0d7f4),
	.w7(32'hb7b9001e),
	.w8(32'h38be0030),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9e81a),
	.w1(32'hbaba73a3),
	.w2(32'hbb9c4a02),
	.w3(32'h3ac5bd9e),
	.w4(32'h39c7431d),
	.w5(32'hbaff544f),
	.w6(32'h3b6353ab),
	.w7(32'h3b298c95),
	.w8(32'h3853281a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db3db2),
	.w1(32'h3b539052),
	.w2(32'h3c48854c),
	.w3(32'hbacf775f),
	.w4(32'hbb51afe5),
	.w5(32'h3b785a97),
	.w6(32'hbbf60abc),
	.w7(32'hbbc95930),
	.w8(32'hbaab2c94),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38d609),
	.w1(32'h3ab8f00a),
	.w2(32'h3b7af10f),
	.w3(32'hba83aba6),
	.w4(32'h3a1df742),
	.w5(32'h3b46145e),
	.w6(32'h3a6f7d1e),
	.w7(32'h3b2393db),
	.w8(32'h3b708353),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0508a),
	.w1(32'h39ae6d03),
	.w2(32'h390d2d5a),
	.w3(32'hb9289383),
	.w4(32'h38ac39bb),
	.w5(32'hb80612a9),
	.w6(32'hba0936d1),
	.w7(32'hb96f23e1),
	.w8(32'hb91465ea),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce502),
	.w1(32'h3b8560f6),
	.w2(32'h3c5862f7),
	.w3(32'hba7caf2f),
	.w4(32'hba90dcc9),
	.w5(32'h3bbc25ab),
	.w6(32'h3ac47af6),
	.w7(32'h3b87eb72),
	.w8(32'h3bed5af1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c9390),
	.w1(32'hbb8fe70f),
	.w2(32'hbbbe91a4),
	.w3(32'h3b06355a),
	.w4(32'h38ee20ea),
	.w5(32'hbac78fb6),
	.w6(32'h3b98065f),
	.w7(32'h3ac00e93),
	.w8(32'h3a39c33b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31db1a),
	.w1(32'hb9d3acf0),
	.w2(32'hbb035899),
	.w3(32'h3b9771f3),
	.w4(32'h3b01f850),
	.w5(32'hba9ac180),
	.w6(32'h3c12b904),
	.w7(32'h3bb8e5d8),
	.w8(32'h3aa2d35d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e39cb7),
	.w1(32'h38bb4475),
	.w2(32'h38424106),
	.w3(32'h378594c2),
	.w4(32'hb8801c37),
	.w5(32'hb9198efb),
	.w6(32'hb77fa4e1),
	.w7(32'hb8846b80),
	.w8(32'hb80074dd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aaa97b),
	.w1(32'hb9a0c7b5),
	.w2(32'hb9cf9998),
	.w3(32'hb9807ebf),
	.w4(32'hba212e7f),
	.w5(32'hb9e54d23),
	.w6(32'h390d81fc),
	.w7(32'hb9451449),
	.w8(32'hb9a0649b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0667bc),
	.w1(32'h3b629e26),
	.w2(32'hbbcd25b7),
	.w3(32'h3b1165fc),
	.w4(32'hbb7ec4ba),
	.w5(32'hbc06f71d),
	.w6(32'h3c2bef82),
	.w7(32'h3ac13f49),
	.w8(32'h3afae725),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dcfba),
	.w1(32'h3a5ac144),
	.w2(32'hbbf7cea3),
	.w3(32'h3b4cac42),
	.w4(32'hbae9c455),
	.w5(32'hba0d0eea),
	.w6(32'h3c170abd),
	.w7(32'h3b7c44cd),
	.w8(32'h3a86460a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc15c),
	.w1(32'h3b4b5839),
	.w2(32'h3bb018e8),
	.w3(32'h3ae05f06),
	.w4(32'h3b8c4f78),
	.w5(32'h3ba48f06),
	.w6(32'h3b91614a),
	.w7(32'h3bc3eeb3),
	.w8(32'h3bbadf4b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8c912),
	.w1(32'h3b8f54ba),
	.w2(32'hbc7da1d2),
	.w3(32'h3c146d2c),
	.w4(32'h3b73a105),
	.w5(32'hbbbca970),
	.w6(32'h3c098e99),
	.w7(32'h3ab3d66b),
	.w8(32'hb8f4b2fb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b4af4),
	.w1(32'hb81f668d),
	.w2(32'hba19b0ed),
	.w3(32'h392c6c56),
	.w4(32'hbaaaecf2),
	.w5(32'hbae75e3c),
	.w6(32'hbaa3c5cb),
	.w7(32'hbb04c8f8),
	.w8(32'hbab85b06),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e486a),
	.w1(32'hbb419be3),
	.w2(32'hbb427814),
	.w3(32'hbabe2b52),
	.w4(32'hbb22b5ec),
	.w5(32'hbb0a19dc),
	.w6(32'h39ae4192),
	.w7(32'hbad2f923),
	.w8(32'hb9681636),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac672d6),
	.w1(32'h3c26435f),
	.w2(32'hbcc320da),
	.w3(32'hbbe7c7ff),
	.w4(32'h3ac6fecd),
	.w5(32'hbca71935),
	.w6(32'h3b19b3b3),
	.w7(32'hbb651bf1),
	.w8(32'hbbb1c11b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ddafb),
	.w1(32'hbbe820a2),
	.w2(32'hbc93a7c3),
	.w3(32'h3c06cc4a),
	.w4(32'hb98c1004),
	.w5(32'hbbe3b4be),
	.w6(32'h3c3ce2cf),
	.w7(32'h3b97e622),
	.w8(32'hbb59c162),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba005c4),
	.w1(32'hbb0ff68e),
	.w2(32'hbbdd8c0a),
	.w3(32'h3be4dce8),
	.w4(32'h3c0de5d0),
	.w5(32'hbb095927),
	.w6(32'h3c318b7e),
	.w7(32'h3be4ad57),
	.w8(32'h3b6c30a1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab9427),
	.w1(32'h3bb102c6),
	.w2(32'h3c6f0ae1),
	.w3(32'hbb118c81),
	.w4(32'hbb3bdb26),
	.w5(32'h3b8ffa94),
	.w6(32'hbbe44875),
	.w7(32'hbb87ac71),
	.w8(32'h3a021dc1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb573004),
	.w1(32'hba3621d4),
	.w2(32'h3c84e2c9),
	.w3(32'hbbe5ce61),
	.w4(32'hbc075f7d),
	.w5(32'h3b06300f),
	.w6(32'hbbf882c9),
	.w7(32'hbbd386b3),
	.w8(32'h3a4d951a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c21e9),
	.w1(32'h387da955),
	.w2(32'h388a1995),
	.w3(32'h36f747ba),
	.w4(32'h37bc24a0),
	.w5(32'h37d56598),
	.w6(32'h375a9291),
	.w7(32'h381aa053),
	.w8(32'h38932152),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36023b74),
	.w1(32'hb79645b0),
	.w2(32'h3698afd0),
	.w3(32'h37b316c6),
	.w4(32'h37050167),
	.w5(32'h378bac43),
	.w6(32'h3844ffc5),
	.w7(32'h38160abe),
	.w8(32'h3689f5a8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae3dea),
	.w1(32'h3a0c9063),
	.w2(32'hbac7373f),
	.w3(32'hba22dd03),
	.w4(32'hbaa4d6b6),
	.w5(32'hba94d8a3),
	.w6(32'h398bc60d),
	.w7(32'hbaf9d4d4),
	.w8(32'h3a9d510b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817cdd7),
	.w1(32'h379708af),
	.w2(32'h38b0f16d),
	.w3(32'hb7cfe9e2),
	.w4(32'h379075f1),
	.w5(32'h3a0a85c6),
	.w6(32'hb8a6c20c),
	.w7(32'hb6638440),
	.w8(32'h3b4f1d64),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b7d1c),
	.w1(32'hbbc5f57f),
	.w2(32'hbb66080c),
	.w3(32'hbab50751),
	.w4(32'hb9c499ba),
	.w5(32'hbc400fe0),
	.w6(32'hbb7e7be1),
	.w7(32'hbb9325bf),
	.w8(32'hbc793688),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd730),
	.w1(32'h39f69937),
	.w2(32'hbb165a5c),
	.w3(32'hbc3fdf64),
	.w4(32'hbc62f17b),
	.w5(32'hbbcffe8a),
	.w6(32'hbbc7abd9),
	.w7(32'hba81a706),
	.w8(32'hbc809007),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957e6a9),
	.w1(32'h3c849f13),
	.w2(32'h3cc03fe0),
	.w3(32'hbc92560f),
	.w4(32'hbb41937b),
	.w5(32'hbbc169d4),
	.w6(32'hbc11bc0d),
	.w7(32'h3c5c82a0),
	.w8(32'hbbcfef7b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18fea9),
	.w1(32'hba031966),
	.w2(32'h3c1f8fa6),
	.w3(32'hbb95e9c3),
	.w4(32'hba9c74bd),
	.w5(32'hbbbdf246),
	.w6(32'hbc463093),
	.w7(32'hbb2272fc),
	.w8(32'hbb70be74),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73a3bb),
	.w1(32'hbb893a37),
	.w2(32'hbcac5853),
	.w3(32'h3bfd8dd3),
	.w4(32'h3b531567),
	.w5(32'h3c6905b8),
	.w6(32'h3cef6c3f),
	.w7(32'h3b9ea2c5),
	.w8(32'h3cbb1125),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02fab3),
	.w1(32'hbcb0d0f7),
	.w2(32'hbcb0ced6),
	.w3(32'h3ce8b86a),
	.w4(32'h3b5d44f2),
	.w5(32'hbc86b90d),
	.w6(32'h3c290480),
	.w7(32'hbcc9611e),
	.w8(32'hbc97549b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3af81b),
	.w1(32'h3ba3852f),
	.w2(32'h3c36ea72),
	.w3(32'hbc9bc8f9),
	.w4(32'hbc334a99),
	.w5(32'hb982467d),
	.w6(32'hbb9cceea),
	.w7(32'h3c9a0921),
	.w8(32'hbb81af23),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa8e4),
	.w1(32'h3b66162f),
	.w2(32'hbc3dc22b),
	.w3(32'h3baa7011),
	.w4(32'h3b87f6bf),
	.w5(32'hbbc3f0f4),
	.w6(32'h3bd452c9),
	.w7(32'h3c0618ba),
	.w8(32'hbc4651db),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c254da3),
	.w1(32'h3c80acd0),
	.w2(32'h3b73d11b),
	.w3(32'h3bea88c9),
	.w4(32'h3c57a935),
	.w5(32'hba145aa4),
	.w6(32'h3cca13d5),
	.w7(32'h3c0ffb7e),
	.w8(32'hbb5a61da),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2abe),
	.w1(32'h3b98c490),
	.w2(32'h3c2a4c2b),
	.w3(32'hbb946d06),
	.w4(32'h3b118e1a),
	.w5(32'hbbdb463a),
	.w6(32'hba879b0e),
	.w7(32'h3bbbe689),
	.w8(32'hbbb21168),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e424a),
	.w1(32'hbbc8770e),
	.w2(32'h3c1f3e41),
	.w3(32'hbba7a1f5),
	.w4(32'h39d6a404),
	.w5(32'hbb149894),
	.w6(32'hbc1eb323),
	.w7(32'h3b283ab6),
	.w8(32'hbadd647b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f5ac4),
	.w1(32'hbb25e559),
	.w2(32'h3a753511),
	.w3(32'hbb110690),
	.w4(32'hbbd681c8),
	.w5(32'hbb40a32a),
	.w6(32'hbb79cb1f),
	.w7(32'hbb5b3557),
	.w8(32'hbbf87506),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a448475),
	.w1(32'h3c8d41c4),
	.w2(32'h3c092e23),
	.w3(32'hbc58e775),
	.w4(32'h3b8d7df3),
	.w5(32'hbc2f270c),
	.w6(32'hb955d7cb),
	.w7(32'h3c6c80d8),
	.w8(32'h3bb6b61a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7a99),
	.w1(32'hbc2da8ab),
	.w2(32'hbc5da0cc),
	.w3(32'h3c8c26fa),
	.w4(32'hbb566f04),
	.w5(32'hbb775065),
	.w6(32'h3d1e983b),
	.w7(32'hbb8632aa),
	.w8(32'h3bc3fc1e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2081bc),
	.w1(32'hbc235e57),
	.w2(32'hbca631e3),
	.w3(32'h3bb61015),
	.w4(32'hbb6f8ba4),
	.w5(32'hbbd750cc),
	.w6(32'h3b21fb5a),
	.w7(32'h3afcf406),
	.w8(32'hbc23d405),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ee5da),
	.w1(32'hbca679b7),
	.w2(32'hbccac12d),
	.w3(32'hbb102aef),
	.w4(32'hbbdfa2a3),
	.w5(32'hbc8e4b1e),
	.w6(32'h3ba413eb),
	.w7(32'hba91ed8f),
	.w8(32'hbb893a84),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7441c),
	.w1(32'h3b37a088),
	.w2(32'h3bd490f1),
	.w3(32'hbc436045),
	.w4(32'hb84caef4),
	.w5(32'hbc41508b),
	.w6(32'hbbe1624b),
	.w7(32'h3c0564b0),
	.w8(32'hbb2e9590),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9cb9),
	.w1(32'hbc272b76),
	.w2(32'hba9817a0),
	.w3(32'hb93ccf29),
	.w4(32'hbb98ffd9),
	.w5(32'hbbe27669),
	.w6(32'h3ca0686d),
	.w7(32'hbbda3501),
	.w8(32'hbb9d2924),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43681),
	.w1(32'hbaaf0385),
	.w2(32'hbb91e3fb),
	.w3(32'hbbd64c99),
	.w4(32'hbbb13ba4),
	.w5(32'hbc825f73),
	.w6(32'hbb4b8965),
	.w7(32'hbb423730),
	.w8(32'hbbf91af9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b076e11),
	.w1(32'h3c62de90),
	.w2(32'h3c66598e),
	.w3(32'hba561585),
	.w4(32'hbb193d57),
	.w5(32'h3b7e45e5),
	.w6(32'hbbfa13f0),
	.w7(32'h3bf406f6),
	.w8(32'hbae2ce53),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3775f),
	.w1(32'hbc74dfce),
	.w2(32'hbc13a396),
	.w3(32'hbb1eea98),
	.w4(32'hbc116288),
	.w5(32'h3c1d7bd1),
	.w6(32'hbbf4519f),
	.w7(32'hbbc4fe84),
	.w8(32'h3bd441f0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63b59e),
	.w1(32'hbbf8cf11),
	.w2(32'hbc2e9655),
	.w3(32'h3c87e718),
	.w4(32'h3ba1a8ad),
	.w5(32'hbc0a298b),
	.w6(32'hbb79cd0c),
	.w7(32'hbbf55365),
	.w8(32'h39ddd235),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337e75),
	.w1(32'h3ca166c9),
	.w2(32'hba5a2dad),
	.w3(32'hbb3c1806),
	.w4(32'h3c1648bf),
	.w5(32'h3b7b910e),
	.w6(32'h3d5a4ee3),
	.w7(32'h3c9eafa5),
	.w8(32'hbb332d7b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038429),
	.w1(32'hbc40ac83),
	.w2(32'hbb8f0573),
	.w3(32'hbbeeea64),
	.w4(32'hbb814903),
	.w5(32'h3c39175b),
	.w6(32'hbc044a42),
	.w7(32'hbbd1cb03),
	.w8(32'h3bb29b7f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a73e),
	.w1(32'h3b641be1),
	.w2(32'hbbbe4661),
	.w3(32'h3c0a296d),
	.w4(32'h3b5e54c7),
	.w5(32'h3bdbf0e5),
	.w6(32'hbb856584),
	.w7(32'h39e19ace),
	.w8(32'h3a8e8c86),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff1bd8),
	.w1(32'hbbae45c6),
	.w2(32'hbbd52321),
	.w3(32'h3be23571),
	.w4(32'h3b6e74d8),
	.w5(32'h3b36d249),
	.w6(32'h3a72ebd6),
	.w7(32'hba32a0cd),
	.w8(32'h3b4db60e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bbece),
	.w1(32'h3ac3b0bb),
	.w2(32'hbb90cb0e),
	.w3(32'h3a03ddcf),
	.w4(32'hbb4b1bba),
	.w5(32'hbb981216),
	.w6(32'hbb400863),
	.w7(32'hbc16a576),
	.w8(32'hbc669968),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd391c9),
	.w1(32'hbcd02c59),
	.w2(32'hbc4f3c4e),
	.w3(32'h3bea849b),
	.w4(32'hbc1bd72a),
	.w5(32'hbc8fe1d6),
	.w6(32'hbbde9a90),
	.w7(32'hba8d385d),
	.w8(32'hbb7fad1f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa25b0),
	.w1(32'hbb1cb894),
	.w2(32'h3c02ef80),
	.w3(32'hbbab96a6),
	.w4(32'h3b264882),
	.w5(32'hbbbeede7),
	.w6(32'hbc112515),
	.w7(32'h3b9858b8),
	.w8(32'hbc154986),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1160a6),
	.w1(32'h3c339498),
	.w2(32'h3b982356),
	.w3(32'hbc620a84),
	.w4(32'hbb80b973),
	.w5(32'h3c70bb2f),
	.w6(32'hbb970241),
	.w7(32'hbc133349),
	.w8(32'h3c8b234d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule