module layer_8_featuremap_160(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc882e85),
	.w1(32'hbc3d6e43),
	.w2(32'hb95bb46d),
	.w3(32'hbc8cdd72),
	.w4(32'hbcaa69eb),
	.w5(32'hbc668b1d),
	.w6(32'hbbe83224),
	.w7(32'hbc77f123),
	.w8(32'hbb3d4c57),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f6c63),
	.w1(32'hbb85e88e),
	.w2(32'hbb557426),
	.w3(32'hbbbe722d),
	.w4(32'hbac31a0c),
	.w5(32'hbb85b447),
	.w6(32'hbbbb7551),
	.w7(32'hbbc66e45),
	.w8(32'hbb9c79c1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c2db1),
	.w1(32'h3bdc6680),
	.w2(32'h3b15c67a),
	.w3(32'hbb4b9bdd),
	.w4(32'hbae2205d),
	.w5(32'hb924c75c),
	.w6(32'hbc0432d4),
	.w7(32'hbb2f0c67),
	.w8(32'h3b711e7a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4cc85),
	.w1(32'hbc40f74f),
	.w2(32'hbbf99f23),
	.w3(32'hbbbff0aa),
	.w4(32'hbc82ead9),
	.w5(32'hbc9ca464),
	.w6(32'hbad3e2c4),
	.w7(32'hbc0d1ac1),
	.w8(32'hbb52f30d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ccf74),
	.w1(32'hbb8dd7be),
	.w2(32'hbbf50980),
	.w3(32'hbc0a14f0),
	.w4(32'h3b5b873c),
	.w5(32'h3ad081cd),
	.w6(32'h3b02bc31),
	.w7(32'h3a7683ac),
	.w8(32'h3b21a742),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5642),
	.w1(32'h3c721e1d),
	.w2(32'h3cf5e7ae),
	.w3(32'h3bea3d89),
	.w4(32'h3c68a5e8),
	.w5(32'h3a5f6911),
	.w6(32'hbc0b6b8c),
	.w7(32'hbc6829b1),
	.w8(32'hbbfb7fb1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d0367),
	.w1(32'hbbd5f943),
	.w2(32'hbb3024dc),
	.w3(32'h3b8b3359),
	.w4(32'h3a988a87),
	.w5(32'h3b9d8814),
	.w6(32'h3a97d5b2),
	.w7(32'h3af85404),
	.w8(32'h3a3a57df),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996a0c),
	.w1(32'hbbc427aa),
	.w2(32'h3ceaeb36),
	.w3(32'hbba2570d),
	.w4(32'h3b5dbb78),
	.w5(32'hb9ae5dda),
	.w6(32'hbcd8dbdc),
	.w7(32'hbd206e9a),
	.w8(32'hbc552d75),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1906d8),
	.w1(32'hbc1d2e82),
	.w2(32'hbbb37180),
	.w3(32'hbc7f3348),
	.w4(32'h3bde1be3),
	.w5(32'h3c1612a6),
	.w6(32'hbae099be),
	.w7(32'hbb2cb069),
	.w8(32'hb945ede0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1446b7),
	.w1(32'hbc55ca28),
	.w2(32'hbd038f1e),
	.w3(32'h3b19c1a8),
	.w4(32'hbb2ea8af),
	.w5(32'h3ccaa6fb),
	.w6(32'h3c39a014),
	.w7(32'h3cd85341),
	.w8(32'h3bcdfc6f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc610ff8),
	.w1(32'hbb8062b0),
	.w2(32'hbb8b602e),
	.w3(32'h3c6a4765),
	.w4(32'hbc6815e0),
	.w5(32'h3b5cce0e),
	.w6(32'hba1ce56d),
	.w7(32'h3b1fc93b),
	.w8(32'h3c387164),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3a0c9),
	.w1(32'hbb01a3bb),
	.w2(32'h3b184343),
	.w3(32'h3a72262b),
	.w4(32'hbab6869f),
	.w5(32'h3baa4ed7),
	.w6(32'h3a5cc29b),
	.w7(32'h3c012eb1),
	.w8(32'h3a48f9d7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae030db),
	.w1(32'h3a930e12),
	.w2(32'hbc814b54),
	.w3(32'h3bb85e65),
	.w4(32'hbc6c3a2c),
	.w5(32'h3a264fcf),
	.w6(32'hbbac3fd6),
	.w7(32'h3c7a4b9c),
	.w8(32'h3b437aa0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f1ff),
	.w1(32'hbc3f1984),
	.w2(32'hbcceca59),
	.w3(32'hbbb44b2b),
	.w4(32'hbb9e9550),
	.w5(32'hbb988660),
	.w6(32'hbc096a7b),
	.w7(32'hbcc18d10),
	.w8(32'hbc2decdb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81131a),
	.w1(32'hbc09bb75),
	.w2(32'hbb138f3a),
	.w3(32'hbc0bc482),
	.w4(32'hbb6d1a95),
	.w5(32'h3b0a9eae),
	.w6(32'hb9e5b746),
	.w7(32'h3af44ca0),
	.w8(32'hb7fa19b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994160),
	.w1(32'h3b3fd122),
	.w2(32'h3bbf2eab),
	.w3(32'h3a6f9272),
	.w4(32'hbc442112),
	.w5(32'hbc1a4026),
	.w6(32'hbc6c8db3),
	.w7(32'h3c030b03),
	.w8(32'h3c27e574),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb650fe8),
	.w1(32'h3be1e1ea),
	.w2(32'hbc74b405),
	.w3(32'h3b9319dd),
	.w4(32'h3c46d49f),
	.w5(32'h3c981268),
	.w6(32'h3c9bc4e0),
	.w7(32'h3c913de8),
	.w8(32'hbc319f42),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ab93e),
	.w1(32'hbcb3eb3a),
	.w2(32'hbcc2c84c),
	.w3(32'hbb1b8ed2),
	.w4(32'hbb3ba4ad),
	.w5(32'h3bd184a9),
	.w6(32'hbad75a3a),
	.w7(32'h3b3fdad6),
	.w8(32'hbc14133e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb9639),
	.w1(32'hbb092208),
	.w2(32'h3c81103e),
	.w3(32'hbcb4e83a),
	.w4(32'hbba380c1),
	.w5(32'h3b9fcfae),
	.w6(32'h3c38f3ad),
	.w7(32'h3b5ec336),
	.w8(32'h3b17825b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f85e6),
	.w1(32'hbc54b7da),
	.w2(32'hbc3b51f9),
	.w3(32'hbb7101c1),
	.w4(32'hbb543563),
	.w5(32'hbb6966dd),
	.w6(32'h3b85ed64),
	.w7(32'h3b8bf6ca),
	.w8(32'hbaab322c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb378b95),
	.w1(32'h3c174df6),
	.w2(32'h39827a7a),
	.w3(32'h3b9db9c7),
	.w4(32'h39746779),
	.w5(32'h3cb62c70),
	.w6(32'h3af73cba),
	.w7(32'h3c2de9af),
	.w8(32'h3c1d4199),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068ff3),
	.w1(32'h3bf0e772),
	.w2(32'h3bfb0aec),
	.w3(32'h3cc0b8f7),
	.w4(32'h3c0abc72),
	.w5(32'hbaf34080),
	.w6(32'hbc1b2b54),
	.w7(32'h3a68cef6),
	.w8(32'hbb23d5da),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e13a),
	.w1(32'h3bdcf27d),
	.w2(32'h394c1f0c),
	.w3(32'hbc9acd35),
	.w4(32'hbd240da0),
	.w5(32'hbcbfc3bf),
	.w6(32'hba26000c),
	.w7(32'h3c3ca9e2),
	.w8(32'h3cc0749e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef7885),
	.w1(32'hba8a771e),
	.w2(32'hbc70827d),
	.w3(32'hbac08075),
	.w4(32'h3b534aba),
	.w5(32'hbbe34a5a),
	.w6(32'hbc7d7962),
	.w7(32'hbc17218b),
	.w8(32'hbc2b0890),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7016cf),
	.w1(32'h3bea2b5f),
	.w2(32'h3c6cd5a9),
	.w3(32'hbb1de2d8),
	.w4(32'hbbdb750f),
	.w5(32'h3b077797),
	.w6(32'hbc33caaa),
	.w7(32'hbc02fa44),
	.w8(32'hb98c3df1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3e201),
	.w1(32'hbba23fd1),
	.w2(32'hb947162b),
	.w3(32'hbb4594a6),
	.w4(32'hbc4ace55),
	.w5(32'hbbb452f0),
	.w6(32'hbc384534),
	.w7(32'hb9d715b6),
	.w8(32'h3b96f21f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941dbb0),
	.w1(32'h3b021abd),
	.w2(32'h3d645185),
	.w3(32'hbaf78a80),
	.w4(32'h3cb8a245),
	.w5(32'h3c254011),
	.w6(32'h3b046d28),
	.w7(32'hbcb1b4d9),
	.w8(32'hbca7e5ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d895864),
	.w1(32'hbc417d1c),
	.w2(32'hbc18bc04),
	.w3(32'hbd5c44b7),
	.w4(32'hbcc4fe55),
	.w5(32'h38ca1618),
	.w6(32'h3c9f572a),
	.w7(32'h3a6baad8),
	.w8(32'h3c873de2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa279),
	.w1(32'hbb5a5e60),
	.w2(32'h3adb09bb),
	.w3(32'hbb3ab7f6),
	.w4(32'hbc4f7ade),
	.w5(32'hbabb1e1f),
	.w6(32'hbb99c8cd),
	.w7(32'h3ab242a8),
	.w8(32'h3abed67e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9466e1),
	.w1(32'h3b301a4d),
	.w2(32'h3b2f385b),
	.w3(32'hbb222b00),
	.w4(32'h3b0efa8e),
	.w5(32'hb878760f),
	.w6(32'hbb28411d),
	.w7(32'hbb7a511c),
	.w8(32'hba927abc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea31c9),
	.w1(32'h3b6e1196),
	.w2(32'h3b26b185),
	.w3(32'h3b1c49fd),
	.w4(32'hbc869005),
	.w5(32'hbab58658),
	.w6(32'hbc281efd),
	.w7(32'hbaf7fda6),
	.w8(32'h3b72c26c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aac69),
	.w1(32'h3bdddbab),
	.w2(32'h3b8a7515),
	.w3(32'h3c0127a2),
	.w4(32'hbb3031a3),
	.w5(32'hba47eaba),
	.w6(32'hbbbb3d25),
	.w7(32'h3bea5b04),
	.w8(32'hb9fa5e1c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70dab3),
	.w1(32'hbc3719ec),
	.w2(32'hbc23aebc),
	.w3(32'hbbd3e11e),
	.w4(32'h3b13fd45),
	.w5(32'h3c7fb294),
	.w6(32'h3c6d60ad),
	.w7(32'h3b6e68a4),
	.w8(32'hbb8f5d05),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2f64f),
	.w1(32'h3bb0209f),
	.w2(32'hb9989130),
	.w3(32'h3c3bda72),
	.w4(32'h3c09c11d),
	.w5(32'h3c5175b9),
	.w6(32'h3c96a7b7),
	.w7(32'h3c9c4221),
	.w8(32'hbb30fada),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a05eb),
	.w1(32'h3b5b8931),
	.w2(32'hbc2873ff),
	.w3(32'h3ca976ec),
	.w4(32'hba3b329c),
	.w5(32'hbb8e262a),
	.w6(32'h3c92686e),
	.w7(32'h3c8e49f7),
	.w8(32'h3c69ac77),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1ab4e),
	.w1(32'h3bc0dad5),
	.w2(32'h3cfa481e),
	.w3(32'hbbcaa857),
	.w4(32'hbb3479b8),
	.w5(32'hbc7ccda5),
	.w6(32'hbcb020ed),
	.w7(32'hbc5de8e1),
	.w8(32'hbc028b73),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbadff7),
	.w1(32'hb9422141),
	.w2(32'h3b92f93e),
	.w3(32'hbc4aa718),
	.w4(32'h3c04fbca),
	.w5(32'h3c112508),
	.w6(32'h39c26ec5),
	.w7(32'h3ac93f42),
	.w8(32'hba24c519),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff6cf4),
	.w1(32'hbbf49aa0),
	.w2(32'hbb6bc57e),
	.w3(32'h3ac4b8d8),
	.w4(32'hbafdc750),
	.w5(32'h3a96933b),
	.w6(32'h3af70416),
	.w7(32'h3ba15a2a),
	.w8(32'h3b067acf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64a7b0),
	.w1(32'hbb099f74),
	.w2(32'hbbb65765),
	.w3(32'h3a1a1240),
	.w4(32'h3c42c17e),
	.w5(32'h3a903dc5),
	.w6(32'hbb14fd0f),
	.w7(32'hbb6d6a0d),
	.w8(32'h39215054),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c586),
	.w1(32'hbaddad1e),
	.w2(32'h3c2497a6),
	.w3(32'h3bcc67d6),
	.w4(32'h3b143382),
	.w5(32'h3c25c6bc),
	.w6(32'hbc1f21a0),
	.w7(32'hbbad9193),
	.w8(32'hbaebc88a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc404d25),
	.w1(32'hbb54b5e5),
	.w2(32'hbbedbbdc),
	.w3(32'hb84d700b),
	.w4(32'hbb9a209d),
	.w5(32'hbbfdefb7),
	.w6(32'h3a12a7e2),
	.w7(32'h3bc7c3e4),
	.w8(32'hbaa45f2b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f6c2d),
	.w1(32'h3a9bda5d),
	.w2(32'hbb88144f),
	.w3(32'hbb9af890),
	.w4(32'h3b8b96a3),
	.w5(32'h3a1b13e6),
	.w6(32'hbb861c52),
	.w7(32'hbc0d6827),
	.w8(32'hbbb2125e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd17cf),
	.w1(32'hbc347819),
	.w2(32'hbb9da150),
	.w3(32'hba20e7f8),
	.w4(32'h3be0aa74),
	.w5(32'h3bb8e315),
	.w6(32'hbb9b324e),
	.w7(32'hbbaea367),
	.w8(32'hbb106e39),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010891),
	.w1(32'hbc0a60a1),
	.w2(32'hbc69ccca),
	.w3(32'hbc2ca139),
	.w4(32'h3bfeadd8),
	.w5(32'h3b01e516),
	.w6(32'h3b4879d8),
	.w7(32'hbb3db499),
	.w8(32'hbb5eb26f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b737a1b),
	.w1(32'h3b9e9611),
	.w2(32'h3c89961c),
	.w3(32'hbc6d83c3),
	.w4(32'hbd0087ef),
	.w5(32'hbca471ae),
	.w6(32'hbc96afcf),
	.w7(32'h3bb9164b),
	.w8(32'h3c00070a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7feac),
	.w1(32'hbb847d07),
	.w2(32'hbb27e0c0),
	.w3(32'hbb1e1bce),
	.w4(32'h3bbe68f3),
	.w5(32'h3bf03e55),
	.w6(32'h395b1171),
	.w7(32'hbad0fab4),
	.w8(32'hb910006f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b621),
	.w1(32'hbbfc6048),
	.w2(32'hbbcbcabf),
	.w3(32'h3b79751a),
	.w4(32'hbb3ff6b8),
	.w5(32'hbb4cd277),
	.w6(32'hba9e8279),
	.w7(32'h3ac3bdb7),
	.w8(32'h3b4e07c6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf3d1),
	.w1(32'h3c0d56d1),
	.w2(32'h3d0a40ca),
	.w3(32'hbbed37d3),
	.w4(32'hbca364a2),
	.w5(32'hbc363245),
	.w6(32'hbcc008e3),
	.w7(32'hbbc38052),
	.w8(32'h3c9a9d5b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bff870),
	.w1(32'h3d246880),
	.w2(32'h3d8566ed),
	.w3(32'hbbb17433),
	.w4(32'hbc240508),
	.w5(32'hba35140a),
	.w6(32'hbb7e4906),
	.w7(32'h3d06f88d),
	.w8(32'h3d143ffe),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e292c),
	.w1(32'hbc0b035b),
	.w2(32'hbbd49bf9),
	.w3(32'hbba5508c),
	.w4(32'hbacb37f4),
	.w5(32'h3c7b8070),
	.w6(32'h3afcb4d9),
	.w7(32'hbb83bd3f),
	.w8(32'hbc5b5aef),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf370bc),
	.w1(32'h3bbd94e7),
	.w2(32'h3c9bad22),
	.w3(32'h3b838fd2),
	.w4(32'h3b72eb1f),
	.w5(32'h3c2e1f53),
	.w6(32'h3ae7c99c),
	.w7(32'h3c6bcb6b),
	.w8(32'h3b328cf9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d3fbd),
	.w1(32'hbb2bdeb5),
	.w2(32'h3a7f1ccd),
	.w3(32'hbcc81375),
	.w4(32'hbc658b58),
	.w5(32'hbbab9f9a),
	.w6(32'hbbdf2560),
	.w7(32'hbc286345),
	.w8(32'hbc4e9005),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18d6b),
	.w1(32'hbbb2dbbc),
	.w2(32'hbb83543c),
	.w3(32'h3b8257bd),
	.w4(32'hbb19b317),
	.w5(32'hbb659383),
	.w6(32'hba2c0bdf),
	.w7(32'h3a4cb51b),
	.w8(32'h39ed8093),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38548c),
	.w1(32'hbc99b7a7),
	.w2(32'hbc8b9032),
	.w3(32'hbbbc0753),
	.w4(32'hbba8e1ba),
	.w5(32'h3c06ffd9),
	.w6(32'hbbde7c48),
	.w7(32'hbc8f0d2a),
	.w8(32'hbba5006e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02805e),
	.w1(32'hbc84049e),
	.w2(32'hbc488b32),
	.w3(32'h3aa22d93),
	.w4(32'hb8a87957),
	.w5(32'h3c25292d),
	.w6(32'h3bd6d813),
	.w7(32'hbb2e881f),
	.w8(32'hbc546f2c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50599),
	.w1(32'hbcbc36a5),
	.w2(32'hbcdb53bb),
	.w3(32'h3a5e1007),
	.w4(32'hbd015eb0),
	.w5(32'hbc81c9c4),
	.w6(32'h3c11bab8),
	.w7(32'h3b98ab5f),
	.w8(32'hbb19eebe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ca9ff),
	.w1(32'h3c1724d4),
	.w2(32'hbbaa909c),
	.w3(32'hbba18f45),
	.w4(32'h3b829e8d),
	.w5(32'h3873fab5),
	.w6(32'hbb1ce8b2),
	.w7(32'h3c11acf0),
	.w8(32'h3be75986),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b3c2),
	.w1(32'h3bd94aa6),
	.w2(32'hbb087037),
	.w3(32'hbc0b8708),
	.w4(32'h3bb773f0),
	.w5(32'hbb0e4911),
	.w6(32'h3aa9b814),
	.w7(32'hbbf789c0),
	.w8(32'h3b4eec85),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a1d47),
	.w1(32'hbbb7d62d),
	.w2(32'h38beb73a),
	.w3(32'hbba5674e),
	.w4(32'hbc19a299),
	.w5(32'hbbb9c13b),
	.w6(32'hbbacb1ef),
	.w7(32'hba6f12ac),
	.w8(32'h3b378570),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66308a),
	.w1(32'hbc2b6696),
	.w2(32'hbc0a4d3f),
	.w3(32'hbba1522a),
	.w4(32'hbc18e07f),
	.w5(32'hbcd20899),
	.w6(32'hbc8bff15),
	.w7(32'hbca7409c),
	.w8(32'hbc88d697),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dbb6f),
	.w1(32'h3b7e5786),
	.w2(32'h3cd25e98),
	.w3(32'hbbdbbc5d),
	.w4(32'h3c568f3e),
	.w5(32'h3c9390c2),
	.w6(32'hbae7aa93),
	.w7(32'hbc39ab7f),
	.w8(32'hbbf5a8a5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17305b),
	.w1(32'hbc852f47),
	.w2(32'hbb333e93),
	.w3(32'hbb8569ce),
	.w4(32'h3b725ba8),
	.w5(32'h3be99ee1),
	.w6(32'h3a1c16d3),
	.w7(32'hbb761316),
	.w8(32'hbb91630e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b2e5c),
	.w1(32'hbc0968bc),
	.w2(32'hbb1e168f),
	.w3(32'hbbacad90),
	.w4(32'hbc446057),
	.w5(32'hbbef9e31),
	.w6(32'hba74bb35),
	.w7(32'h3a41a985),
	.w8(32'hbb3cd8ce),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2185fc),
	.w1(32'hba342bfa),
	.w2(32'h3a1e8a61),
	.w3(32'hbc1b7b6d),
	.w4(32'hbb884c7c),
	.w5(32'hba9defbb),
	.w6(32'hbb1725ed),
	.w7(32'h3a128903),
	.w8(32'h3af81668),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995a95d),
	.w1(32'h3b7de744),
	.w2(32'h3c066cd3),
	.w3(32'hb5de0bd6),
	.w4(32'h390b72a5),
	.w5(32'h3acbd4bb),
	.w6(32'hbb72d40b),
	.w7(32'h3b38db54),
	.w8(32'h3a65ae08),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befd7a4),
	.w1(32'h3b4d7b54),
	.w2(32'hbad97676),
	.w3(32'hbb12d629),
	.w4(32'hbafb4eb5),
	.w5(32'h3b195efd),
	.w6(32'hbbaece35),
	.w7(32'hbc25e2fc),
	.w8(32'hbc22c659),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696fb5),
	.w1(32'h3c219c54),
	.w2(32'hbc53d7c3),
	.w3(32'h3bde856d),
	.w4(32'hbc8fec8e),
	.w5(32'hbc3314a1),
	.w6(32'h3c012c7e),
	.w7(32'h3d01eadd),
	.w8(32'h3ce85d16),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc96a4),
	.w1(32'hbc2be0fd),
	.w2(32'hbc6f80c9),
	.w3(32'h3c470c3a),
	.w4(32'hbc4af059),
	.w5(32'hbba1e0dc),
	.w6(32'h3af9c39e),
	.w7(32'hbb5a25de),
	.w8(32'hbb996314),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8935f1),
	.w1(32'hbc2deac2),
	.w2(32'hbcc8627c),
	.w3(32'hbc6e4453),
	.w4(32'hba013a73),
	.w5(32'h3a0094e4),
	.w6(32'h3c0fe053),
	.w7(32'hbbce857b),
	.w8(32'hbc0dfe4e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61bc60),
	.w1(32'h3c90db12),
	.w2(32'h3cad7863),
	.w3(32'hbcce1485),
	.w4(32'hbca2af45),
	.w5(32'h3a91baf2),
	.w6(32'hbc3492c7),
	.w7(32'h3c204a24),
	.w8(32'h3bc012cf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be17994),
	.w1(32'hbc05317e),
	.w2(32'hbbfb5e8d),
	.w3(32'h3ade3210),
	.w4(32'h3b189c2b),
	.w5(32'h3b054ac4),
	.w6(32'h3bad4e3e),
	.w7(32'hbba54315),
	.w8(32'hbb968839),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b066064),
	.w1(32'h3aac7073),
	.w2(32'hbc10279f),
	.w3(32'h3bc65298),
	.w4(32'hbc84e544),
	.w5(32'hbc447bb8),
	.w6(32'hbbf7e496),
	.w7(32'h3bb631c0),
	.w8(32'h3bcae7f7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79d57e),
	.w1(32'h3ca81d97),
	.w2(32'h3d14b96d),
	.w3(32'h3c16b0b4),
	.w4(32'hbc2977f5),
	.w5(32'hbc63d12d),
	.w6(32'hbc96315e),
	.w7(32'hbbaeebae),
	.w8(32'h3c186930),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad468c6),
	.w1(32'h3b013e55),
	.w2(32'hbc6b7063),
	.w3(32'hbc3c3181),
	.w4(32'hbc03e32f),
	.w5(32'hbc064644),
	.w6(32'hbb3f3f56),
	.w7(32'h3b43e16f),
	.w8(32'h3bd6505f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08aa2f),
	.w1(32'h3bd5dc73),
	.w2(32'h3b78f16c),
	.w3(32'h3b9004b3),
	.w4(32'h398dc295),
	.w5(32'h3ba59219),
	.w6(32'hbb1ecb79),
	.w7(32'hbbed0ab8),
	.w8(32'h3bc4a8b8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f061a),
	.w1(32'hbb85dd22),
	.w2(32'hbc085eb0),
	.w3(32'h3c5204ac),
	.w4(32'h3b8b4ff0),
	.w5(32'h3bef8159),
	.w6(32'hbb20114f),
	.w7(32'hbab02c42),
	.w8(32'hbbae48ce),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398818d5),
	.w1(32'h3c5aa55f),
	.w2(32'h3c0dfc7f),
	.w3(32'h3ba8a3e1),
	.w4(32'h3af29199),
	.w5(32'h3b409ff3),
	.w6(32'h3ae189c2),
	.w7(32'h3b80fe7e),
	.w8(32'h3be01b98),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0ba0),
	.w1(32'hbbf8ef78),
	.w2(32'hbbcdfce8),
	.w3(32'hbc45abce),
	.w4(32'hbc538f62),
	.w5(32'hbc2f8cc1),
	.w6(32'hbb11a9c0),
	.w7(32'hbb1bc43d),
	.w8(32'hba20b0c9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8668),
	.w1(32'hbba1b3a9),
	.w2(32'hbc2826d8),
	.w3(32'hbc558f76),
	.w4(32'hbb975dd0),
	.w5(32'h3bcc3ed8),
	.w6(32'hbb9cbf39),
	.w7(32'hbaf8c8dc),
	.w8(32'h3a8f076d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc553215),
	.w1(32'hbc9dae67),
	.w2(32'hbc1343ad),
	.w3(32'h3c0c096a),
	.w4(32'h3aa240d9),
	.w5(32'h3bc2502c),
	.w6(32'h3c3ea8e3),
	.w7(32'h3a334637),
	.w8(32'hbbf8b44e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24976),
	.w1(32'h3c02dd4e),
	.w2(32'h3cb22a8b),
	.w3(32'hba01e224),
	.w4(32'h3a0f82d6),
	.w5(32'h3c105a69),
	.w6(32'hbbf57c07),
	.w7(32'h3b3fc63c),
	.w8(32'h3ca2c339),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a787),
	.w1(32'hbbdf69b8),
	.w2(32'hbc633643),
	.w3(32'h3bb3b636),
	.w4(32'h3c06b4a2),
	.w5(32'h3c5666c6),
	.w6(32'h39af36fb),
	.w7(32'hbc690b82),
	.w8(32'hbb2134df),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3279fd),
	.w1(32'hbbf969f6),
	.w2(32'h39ec09bb),
	.w3(32'h3b95233c),
	.w4(32'h3c354937),
	.w5(32'h3c1e2229),
	.w6(32'h3baba33f),
	.w7(32'h3c044bd9),
	.w8(32'hbafa12b7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f3ccc),
	.w1(32'hbcb9b60b),
	.w2(32'hbc1e1a17),
	.w3(32'hbc14e3c5),
	.w4(32'h3bb15672),
	.w5(32'hbacd71c2),
	.w6(32'h3b94dc4b),
	.w7(32'h3a49e2ec),
	.w8(32'hbc098602),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cbe36),
	.w1(32'hbb9ab4f5),
	.w2(32'hbc224a92),
	.w3(32'hbc904980),
	.w4(32'hbcd262f4),
	.w5(32'hbc1eba27),
	.w6(32'hbc23613e),
	.w7(32'h3bf75c5d),
	.w8(32'h3cb0abfc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5d473),
	.w1(32'hbb38e673),
	.w2(32'h3c616a39),
	.w3(32'hbc2a4c8b),
	.w4(32'hbc54c94e),
	.w5(32'hbcba0248),
	.w6(32'hbcd65e8d),
	.w7(32'hbc93e4af),
	.w8(32'h3ae3893d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ac486),
	.w1(32'hbc0287ac),
	.w2(32'hbbcfb651),
	.w3(32'hbcb49f6b),
	.w4(32'hbb61697b),
	.w5(32'hba545d92),
	.w6(32'h3b106871),
	.w7(32'h3b1c7758),
	.w8(32'hbaeaaffb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15a963),
	.w1(32'hbbb7bf4d),
	.w2(32'h3b46c894),
	.w3(32'h3bab9c64),
	.w4(32'h3935dfdc),
	.w5(32'hbb324184),
	.w6(32'hbbbcbed9),
	.w7(32'hbc5b0798),
	.w8(32'hbc48d0fe),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becd243),
	.w1(32'hb941d972),
	.w2(32'h3994d762),
	.w3(32'hbb919eed),
	.w4(32'hbb7eaf2d),
	.w5(32'h3b640f91),
	.w6(32'hbc418776),
	.w7(32'hbb40150c),
	.w8(32'hba52442c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf4a52),
	.w1(32'h3c21edaf),
	.w2(32'h3cd7d567),
	.w3(32'h3c3c1689),
	.w4(32'hbb5fbac3),
	.w5(32'h3bd4db9f),
	.w6(32'hbb1316fe),
	.w7(32'h3c6324eb),
	.w8(32'h3c3e76d9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b1df7),
	.w1(32'hb91cd706),
	.w2(32'h3c42a232),
	.w3(32'h3c3fac15),
	.w4(32'hbc9240e9),
	.w5(32'hbc9900d6),
	.w6(32'hbc6399c9),
	.w7(32'hbc8b8653),
	.w8(32'h3a755357),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d480),
	.w1(32'h3bbd94b7),
	.w2(32'hb99ec389),
	.w3(32'hbc1f595e),
	.w4(32'h3bdb3300),
	.w5(32'h3c525dad),
	.w6(32'h3c7cd122),
	.w7(32'h3c2b7c66),
	.w8(32'h3be4cc53),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a63a2),
	.w1(32'h3aee80be),
	.w2(32'hbb1c455f),
	.w3(32'h3c514e34),
	.w4(32'h3ade89df),
	.w5(32'h3a406ede),
	.w6(32'hba8ac45d),
	.w7(32'h3a02fb56),
	.w8(32'hba290f15),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d34ad),
	.w1(32'hbb825581),
	.w2(32'hbbadf627),
	.w3(32'hbba2ae28),
	.w4(32'hbbb48b83),
	.w5(32'hbba7d9c1),
	.w6(32'hbb373692),
	.w7(32'hbb227699),
	.w8(32'hbb5c1b67),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf730c),
	.w1(32'hbb46d0b3),
	.w2(32'hbcab87fc),
	.w3(32'hba87ff56),
	.w4(32'hbbc65efd),
	.w5(32'hbc20a144),
	.w6(32'h3c887e56),
	.w7(32'h3cb0e014),
	.w8(32'h3c138f6f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc403165),
	.w1(32'hbb647c57),
	.w2(32'hbb388f3c),
	.w3(32'hb9821b4d),
	.w4(32'hbbc22d6e),
	.w5(32'hbb0f4fe5),
	.w6(32'h3bc422af),
	.w7(32'h3b472c8f),
	.w8(32'h39949515),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9bdd),
	.w1(32'hbb97b869),
	.w2(32'hbb963682),
	.w3(32'hbbac3043),
	.w4(32'hba49d32b),
	.w5(32'hbbd3c3ad),
	.w6(32'hbbc7efb6),
	.w7(32'h3ade012a),
	.w8(32'hb9e06ee6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cf329),
	.w1(32'hbb23449f),
	.w2(32'h3a72bbd1),
	.w3(32'h3b5e777d),
	.w4(32'h3c47f708),
	.w5(32'h3c427eff),
	.w6(32'h3c199314),
	.w7(32'h3c20c8fd),
	.w8(32'h3addacad),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d1aa1),
	.w1(32'hbb1d70e5),
	.w2(32'hbbb6c55f),
	.w3(32'h3bf0349c),
	.w4(32'h3ca09390),
	.w5(32'h3bc7ff1c),
	.w6(32'h3b8542c6),
	.w7(32'h3bed3210),
	.w8(32'h3b2a088a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc859),
	.w1(32'h3bb463d5),
	.w2(32'hba0a946b),
	.w3(32'h398cc9e3),
	.w4(32'hba4ac906),
	.w5(32'hbafeda9b),
	.w6(32'h3b7047b1),
	.w7(32'h3be6fb65),
	.w8(32'h3bd61828),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64d728),
	.w1(32'hbc201bc9),
	.w2(32'hbb426b27),
	.w3(32'hbb9f88e1),
	.w4(32'hbb34ed83),
	.w5(32'h3b43b428),
	.w6(32'hbb73689a),
	.w7(32'hbb939dde),
	.w8(32'h3b6641f8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6557b1),
	.w1(32'hbc65b0d0),
	.w2(32'hb939f064),
	.w3(32'h3a3fcf3e),
	.w4(32'h3c098980),
	.w5(32'h3c2bc633),
	.w6(32'h3bfbe2ec),
	.w7(32'hbb389ac7),
	.w8(32'hbbfc3a2a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8db36),
	.w1(32'hbb62134e),
	.w2(32'hbce08f30),
	.w3(32'hbb02013f),
	.w4(32'h3c1a9cbe),
	.w5(32'h3c8dd071),
	.w6(32'h3bea9c62),
	.w7(32'h3bdb25f3),
	.w8(32'h3bdb102a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3794),
	.w1(32'hbbca9db3),
	.w2(32'hbcdbd2ea),
	.w3(32'h3c92e821),
	.w4(32'hbb6c5ca2),
	.w5(32'h3bfb8576),
	.w6(32'h3c947d4f),
	.w7(32'h3cbe2a28),
	.w8(32'hbc72bf89),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca49bfd),
	.w1(32'hbc027e1f),
	.w2(32'hbbed6343),
	.w3(32'hbbd39c59),
	.w4(32'h3c7c18dc),
	.w5(32'h3be94fb2),
	.w6(32'hb9ca8ee7),
	.w7(32'hbbc83ba7),
	.w8(32'hbbbff07c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d57cc),
	.w1(32'hbbbf1904),
	.w2(32'hbba2b783),
	.w3(32'hbc86d3dd),
	.w4(32'hbc1ce1c3),
	.w5(32'hbbbde677),
	.w6(32'hbba522f4),
	.w7(32'hbb5a351b),
	.w8(32'h3b92e2e1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d5359),
	.w1(32'h3c9809e5),
	.w2(32'h3c99f6f5),
	.w3(32'hbac6b1b7),
	.w4(32'hbc1e72b2),
	.w5(32'hbb2a6462),
	.w6(32'hbb1a5411),
	.w7(32'h3c83bbee),
	.w8(32'h3c8d5886),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07991a),
	.w1(32'hbbf712bd),
	.w2(32'hba425933),
	.w3(32'h3ad8e365),
	.w4(32'h3c7efc80),
	.w5(32'h3c876417),
	.w6(32'hbc4bb1d5),
	.w7(32'hbb9e1962),
	.w8(32'hbadfc8a2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af79bda),
	.w1(32'h3b95dcfc),
	.w2(32'h3bad06fc),
	.w3(32'h3ba979e1),
	.w4(32'hba769987),
	.w5(32'hbafd3a2e),
	.w6(32'hbb490bad),
	.w7(32'hbb9dbc46),
	.w8(32'h3aa765bf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0a9f7),
	.w1(32'h3a6be6ea),
	.w2(32'h3b3317ff),
	.w3(32'h39fee87b),
	.w4(32'h3b520c4c),
	.w5(32'h3a5f6f08),
	.w6(32'h3a38dc0a),
	.w7(32'h3b4a0da1),
	.w8(32'h3bbcf899),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94f325),
	.w1(32'hbc37727a),
	.w2(32'hbcb75679),
	.w3(32'h3affcc2c),
	.w4(32'h3b1368ab),
	.w5(32'hbc571e58),
	.w6(32'hbaa7694e),
	.w7(32'hbb7468c4),
	.w8(32'hbba20a29),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f77fa),
	.w1(32'hbb3191d3),
	.w2(32'hb996aa6a),
	.w3(32'hbc0be3dc),
	.w4(32'hbaad08b2),
	.w5(32'hb7de8485),
	.w6(32'hbb948bdf),
	.w7(32'hbb62e02a),
	.w8(32'hbb81cc70),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909454),
	.w1(32'h3aca0b8d),
	.w2(32'h3c39c0cf),
	.w3(32'h3b908129),
	.w4(32'h3b43cde0),
	.w5(32'h3c564122),
	.w6(32'hbc2536a4),
	.w7(32'hbabe6fb1),
	.w8(32'hbc1e9054),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c0991),
	.w1(32'h3c00c486),
	.w2(32'hb9923c27),
	.w3(32'hbacd6440),
	.w4(32'hbc958549),
	.w5(32'h3bd22c4b),
	.w6(32'h3c1df5bf),
	.w7(32'h3d0ed346),
	.w8(32'h3cdba3ad),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b6af8),
	.w1(32'hbb3e132c),
	.w2(32'hbb197f9c),
	.w3(32'h3c579de0),
	.w4(32'hbbd85cac),
	.w5(32'h3a832fb4),
	.w6(32'hbbf0d943),
	.w7(32'hbb82b877),
	.w8(32'hbbbd89c0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054f21),
	.w1(32'h3add46c4),
	.w2(32'h3b91da87),
	.w3(32'h3b919862),
	.w4(32'h3a79525a),
	.w5(32'h3a2a00a4),
	.w6(32'hba942444),
	.w7(32'h3b0f0188),
	.w8(32'h3a21ebd2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35689d),
	.w1(32'hba10df22),
	.w2(32'h3c16e18a),
	.w3(32'hbac36849),
	.w4(32'h3b09e3bf),
	.w5(32'h3b4a6b26),
	.w6(32'hbc1829a7),
	.w7(32'hbc1de81c),
	.w8(32'hbc4d4ed2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d1d2a),
	.w1(32'hbbd78163),
	.w2(32'h3b5a1931),
	.w3(32'hbbcba178),
	.w4(32'h3a7f3bf0),
	.w5(32'h3b9fb4ab),
	.w6(32'hbb687491),
	.w7(32'h3b01bd3a),
	.w8(32'hbb4074fe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a586ef),
	.w1(32'hbb30e32b),
	.w2(32'hbbffa2cd),
	.w3(32'h3b7ff1e8),
	.w4(32'h3bba72e6),
	.w5(32'h3c0bbfc0),
	.w6(32'h3bb269ff),
	.w7(32'h3b03f5ca),
	.w8(32'h3a3b7d8b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb539b15),
	.w1(32'hbb71c152),
	.w2(32'hba2f4927),
	.w3(32'h3c240c93),
	.w4(32'hbaede2ec),
	.w5(32'hba074bc8),
	.w6(32'hbbaed30f),
	.w7(32'hbc1c33ca),
	.w8(32'hbbaf7dd8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6964e5),
	.w1(32'hbc5eff39),
	.w2(32'hbc1f11a4),
	.w3(32'h3b90efe5),
	.w4(32'h389d4a29),
	.w5(32'h3c168d85),
	.w6(32'h3ba2a291),
	.w7(32'hbb27d154),
	.w8(32'hbbd32984),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab6c5),
	.w1(32'h383d2238),
	.w2(32'hbc1ebb9a),
	.w3(32'h3b051232),
	.w4(32'hbb1f1ffe),
	.w5(32'h3b0ad1b4),
	.w6(32'h3ba55dec),
	.w7(32'h3bf0afa2),
	.w8(32'hbb250047),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ace81),
	.w1(32'h3aaf34d5),
	.w2(32'hbac5465c),
	.w3(32'h3bad470f),
	.w4(32'h39cb9f07),
	.w5(32'hbb9d6055),
	.w6(32'hbb06e0e3),
	.w7(32'hbbb4eda0),
	.w8(32'hbac94a38),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ab1a4),
	.w1(32'hb97fdece),
	.w2(32'h3c2d79ca),
	.w3(32'hbb3966fe),
	.w4(32'h3b6fddcb),
	.w5(32'h3b6b083c),
	.w6(32'hbbe16d3f),
	.w7(32'hbae538d9),
	.w8(32'hbc260443),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42d61),
	.w1(32'hbce4e1d6),
	.w2(32'hbcced4d1),
	.w3(32'hb9c39576),
	.w4(32'hbb4e5df1),
	.w5(32'hbc753bca),
	.w6(32'hbb85b864),
	.w7(32'hbc895914),
	.w8(32'hbc6283f4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca67124),
	.w1(32'h3d08fd0d),
	.w2(32'h3d16ac0a),
	.w3(32'hbc3769e5),
	.w4(32'hbc269537),
	.w5(32'hbadb41cc),
	.w6(32'hbca3633b),
	.w7(32'h3b50877a),
	.w8(32'h3c4ee859),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ce0d),
	.w1(32'hbb82bf6e),
	.w2(32'hbb593beb),
	.w3(32'h3b9a4d7a),
	.w4(32'h390193ea),
	.w5(32'h3afa76ab),
	.w6(32'hbb0ca32b),
	.w7(32'hba9fe341),
	.w8(32'hbb00fae6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2eade),
	.w1(32'hba2b6b45),
	.w2(32'h3a85dc8f),
	.w3(32'hba386119),
	.w4(32'hbb687578),
	.w5(32'hbb3b8987),
	.w6(32'hbb12f112),
	.w7(32'h3abbf6d4),
	.w8(32'h3c3526ed),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule