module layer_10_featuremap_187(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34655919),
	.w1(32'hb469ccef),
	.w2(32'h353fda66),
	.w3(32'h341dcc4c),
	.w4(32'hb2a22102),
	.w5(32'hb4bdb1f5),
	.w6(32'h35c21632),
	.w7(32'hb5e12464),
	.w8(32'h34b15bd8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79d106a),
	.w1(32'hb70d738e),
	.w2(32'hb5bbdb8b),
	.w3(32'h366d6a64),
	.w4(32'h3708c38d),
	.w5(32'h382b78de),
	.w6(32'h36491930),
	.w7(32'h37f8c30b),
	.w8(32'h37f78dd1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35656713),
	.w1(32'h352326d5),
	.w2(32'hb3832205),
	.w3(32'h3409b7ef),
	.w4(32'hb38a5ea9),
	.w5(32'hb4b8c0fa),
	.w6(32'h350c596f),
	.w7(32'h359c81c5),
	.w8(32'h348db939),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3757037c),
	.w1(32'h380aa16c),
	.w2(32'h3795e543),
	.w3(32'hb790f5f4),
	.w4(32'h359c66e4),
	.w5(32'hb6cbd72f),
	.w6(32'h3702845f),
	.w7(32'h37256035),
	.w8(32'h37b2870c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35992388),
	.w1(32'h34f5aeb1),
	.w2(32'hb46f22b4),
	.w3(32'h361965d4),
	.w4(32'h35bb22e1),
	.w5(32'h3594508a),
	.w6(32'h3600edc8),
	.w7(32'h35ea2f37),
	.w8(32'h35c20f14),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c1c13f),
	.w1(32'h35940f3e),
	.w2(32'h35445211),
	.w3(32'h3304ae92),
	.w4(32'h35218e2b),
	.w5(32'h35747fdc),
	.w6(32'h35533871),
	.w7(32'hb3e54db1),
	.w8(32'h35690d78),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e5fe8c),
	.w1(32'h37e593af),
	.w2(32'h3864b827),
	.w3(32'hb77a3ffc),
	.w4(32'h366c470e),
	.w5(32'h36cda2ec),
	.w6(32'h3761f41f),
	.w7(32'hb5df2b17),
	.w8(32'h37a82e8b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3797576f),
	.w1(32'hb8fe99dc),
	.w2(32'hb8723675),
	.w3(32'hb83a6a91),
	.w4(32'h3856106b),
	.w5(32'h389aa2cd),
	.w6(32'h381175e5),
	.w7(32'hb88533ee),
	.w8(32'hb754bce7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76e4c4e),
	.w1(32'hb7209f7c),
	.w2(32'h37a67c94),
	.w3(32'h378330b4),
	.w4(32'h38147d99),
	.w5(32'h382b3666),
	.w6(32'hb7bee080),
	.w7(32'hb70eca90),
	.w8(32'h38699b1e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874b43a),
	.w1(32'hb840d2bf),
	.w2(32'hb74edef4),
	.w3(32'h3892a7e8),
	.w4(32'hb7b4166c),
	.w5(32'h36e2d3d8),
	.w6(32'hb86ee97d),
	.w7(32'hb928f19b),
	.w8(32'hb89e436a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8117ab9),
	.w1(32'h38531b8d),
	.w2(32'h38841de6),
	.w3(32'hb87df644),
	.w4(32'h354c66a7),
	.w5(32'h37668575),
	.w6(32'hb857376e),
	.w7(32'hb7f0c076),
	.w8(32'h36a6c7cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f9e6ac),
	.w1(32'h37b3fd5e),
	.w2(32'h375b961d),
	.w3(32'hb8060223),
	.w4(32'h377c36da),
	.w5(32'h37f78645),
	.w6(32'hb6856b54),
	.w7(32'h379f8e31),
	.w8(32'h3854a6a4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e91b7),
	.w1(32'h37fe641a),
	.w2(32'hb80785cd),
	.w3(32'hb8669a8f),
	.w4(32'hb883ef76),
	.w5(32'hb84e11d4),
	.w6(32'hb8518d47),
	.w7(32'hb8daa299),
	.w8(32'hb886f3f0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853ece9),
	.w1(32'h37734f70),
	.w2(32'hb6a4d1d5),
	.w3(32'h3834cbca),
	.w4(32'h37932ac2),
	.w5(32'h3731885a),
	.w6(32'h36b625f2),
	.w7(32'h35b51075),
	.w8(32'h378ebb1a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382ff3f4),
	.w1(32'h378cfdf2),
	.w2(32'hb8575ea0),
	.w3(32'h3883cdb8),
	.w4(32'h3842d1b8),
	.w5(32'h388099e0),
	.w6(32'hb7a12094),
	.w7(32'hb8111e4f),
	.w8(32'hb701f0b8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7945f8c),
	.w1(32'h3864a94e),
	.w2(32'h37927be7),
	.w3(32'h372c6016),
	.w4(32'hb50be6a7),
	.w5(32'h3863a296),
	.w6(32'hb87e1d92),
	.w7(32'hb5796f3a),
	.w8(32'h3751e6bc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d12f3f),
	.w1(32'h367054d9),
	.w2(32'hb4b0aa87),
	.w3(32'h388740b3),
	.w4(32'h3565ed9b),
	.w5(32'hb876bbd1),
	.w6(32'h38ae39ae),
	.w7(32'h3596b8b1),
	.w8(32'h3826fb52),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dda652),
	.w1(32'hb7b505f1),
	.w2(32'h37666f0d),
	.w3(32'hb8b024dd),
	.w4(32'hb8d178f1),
	.w5(32'hb91fe1b0),
	.w6(32'h366e1227),
	.w7(32'hb87abf41),
	.w8(32'h37750058),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6933ab8),
	.w1(32'h37ebccd9),
	.w2(32'h35240bcf),
	.w3(32'hb7855f41),
	.w4(32'hb680457e),
	.w5(32'hb83f0254),
	.w6(32'hb79adfaa),
	.w7(32'hb80092c0),
	.w8(32'h371ff923),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f9c8a2),
	.w1(32'h350d5585),
	.w2(32'hb54be8c1),
	.w3(32'hb4f26be4),
	.w4(32'h34bcacac),
	.w5(32'h35241667),
	.w6(32'h359f5e4b),
	.w7(32'h35cc8756),
	.w8(32'h3463b2e7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ee75f2),
	.w1(32'h35dbd9db),
	.w2(32'hb48c617c),
	.w3(32'h361cd9ec),
	.w4(32'h3606276d),
	.w5(32'h36219f67),
	.w6(32'h3650fd58),
	.w7(32'h364c6df3),
	.w8(32'h36546569),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716220f),
	.w1(32'h375fa708),
	.w2(32'hb5ec04ac),
	.w3(32'h3788d46f),
	.w4(32'h374c9f0f),
	.w5(32'h35f0fde8),
	.w6(32'h379c7771),
	.w7(32'h376ab98d),
	.w8(32'h36b3d3e3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b12256),
	.w1(32'h389798f0),
	.w2(32'h383dad37),
	.w3(32'hb912f070),
	.w4(32'h3823ebf5),
	.w5(32'hb7c92615),
	.w6(32'hb94e73f6),
	.w7(32'h398f89fe),
	.w8(32'h39b30299),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ace16a),
	.w1(32'hb7fbabb9),
	.w2(32'hb6102612),
	.w3(32'hb875f7ba),
	.w4(32'h37203697),
	.w5(32'hb76d3ec8),
	.w6(32'hb8fd1e11),
	.w7(32'hb8a21e2b),
	.w8(32'hb89be030),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883c927),
	.w1(32'h3920321a),
	.w2(32'h3683aace),
	.w3(32'h38c3f770),
	.w4(32'h3960665e),
	.w5(32'h38a7783c),
	.w6(32'h378e356e),
	.w7(32'h38b2e3ba),
	.w8(32'hb8bef285),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7342e5c),
	.w1(32'hb775e757),
	.w2(32'h386cdc04),
	.w3(32'h37ea33b3),
	.w4(32'h37529fa5),
	.w5(32'h388d0113),
	.w6(32'hb6a9854f),
	.w7(32'hb69f15e0),
	.w8(32'h380c8b64),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37841c7e),
	.w1(32'h378037aa),
	.w2(32'h36ec1ef9),
	.w3(32'h3707cde5),
	.w4(32'h374f69c2),
	.w5(32'h36d6ae70),
	.w6(32'h371b5500),
	.w7(32'h3731ec6a),
	.w8(32'h364a9e1d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d12b3b),
	.w1(32'h38888f4f),
	.w2(32'h38215fa0),
	.w3(32'hb8494d4a),
	.w4(32'h389abbc1),
	.w5(32'h38377dac),
	.w6(32'hb8bcb6c9),
	.w7(32'h38bd0391),
	.w8(32'hb7f1dac6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a97320),
	.w1(32'h387a8983),
	.w2(32'h3833e0b4),
	.w3(32'h37a1e9df),
	.w4(32'h3830087e),
	.w5(32'h38a92f94),
	.w6(32'h36afc658),
	.w7(32'h3645e88e),
	.w8(32'h383ce87c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993f3dc),
	.w1(32'hb8dbccb7),
	.w2(32'h38889418),
	.w3(32'hb8b5db34),
	.w4(32'hb6da6afc),
	.w5(32'h3907370a),
	.w6(32'hb916e69b),
	.w7(32'hb8a239ce),
	.w8(32'h38c7e5cc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d32381),
	.w1(32'h36b1b8e0),
	.w2(32'h36ada35f),
	.w3(32'h36787d25),
	.w4(32'h361c3b0c),
	.w5(32'h354ac201),
	.w6(32'h3695dadb),
	.w7(32'h36255f85),
	.w8(32'h357ff809),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fcf523),
	.w1(32'h36aabfd2),
	.w2(32'hb6952ae0),
	.w3(32'h37d60ec0),
	.w4(32'h3672a552),
	.w5(32'h3650a869),
	.w6(32'h37e1a924),
	.w7(32'hb7c3a288),
	.w8(32'h352db93a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cdfc9),
	.w1(32'h37ef4140),
	.w2(32'h37c1b55d),
	.w3(32'hb71841dc),
	.w4(32'hb7ec236a),
	.w5(32'hb7c84aff),
	.w6(32'h3727e267),
	.w7(32'hb807a62a),
	.w8(32'hb7e14dd1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83af63b),
	.w1(32'hb7f5ee19),
	.w2(32'hb822b283),
	.w3(32'hb7e4110b),
	.w4(32'h3754bf92),
	.w5(32'hb7287e99),
	.w6(32'hb86998d9),
	.w7(32'h36fbc05c),
	.w8(32'hb6ba60e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4893259),
	.w1(32'h36dbc8e2),
	.w2(32'h378f0877),
	.w3(32'h36bab9f8),
	.w4(32'h352e864d),
	.w5(32'hb6866446),
	.w6(32'h36c036d9),
	.w7(32'h3756efc5),
	.w8(32'h37852113),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b85d19),
	.w1(32'h37de3385),
	.w2(32'h379d0c6b),
	.w3(32'hb7ea610c),
	.w4(32'hb503e809),
	.w5(32'hb756117a),
	.w6(32'h38206ba4),
	.w7(32'hb72fa2da),
	.w8(32'hb5b16cfa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bc445),
	.w1(32'hb918703d),
	.w2(32'hb859f9e9),
	.w3(32'hb8c119eb),
	.w4(32'hb4c62c13),
	.w5(32'h3802c2b2),
	.w6(32'hb8d005f8),
	.w7(32'hb964cd66),
	.w8(32'h38939586),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78cd13d),
	.w1(32'hb76c111a),
	.w2(32'hb9a4e67b),
	.w3(32'h37df448f),
	.w4(32'h389e7d36),
	.w5(32'h38c21827),
	.w6(32'h38fa3ae9),
	.w7(32'h3897bf44),
	.w8(32'h390906ab),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e51f9f),
	.w1(32'h39311924),
	.w2(32'h38c7bea8),
	.w3(32'h38e237ea),
	.w4(32'h39873ad2),
	.w5(32'h38e754c7),
	.w6(32'hb797423f),
	.w7(32'hb87d377e),
	.w8(32'hb9210eed),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee144a),
	.w1(32'h37bc429f),
	.w2(32'hb864bec8),
	.w3(32'h382df20a),
	.w4(32'h382ec914),
	.w5(32'hb7d80b88),
	.w6(32'h37dff101),
	.w7(32'h37043490),
	.w8(32'hb801fe09),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36168ceb),
	.w1(32'hb7ef0990),
	.w2(32'h378f1541),
	.w3(32'hb7b7a78e),
	.w4(32'h3442378c),
	.w5(32'h381031b3),
	.w6(32'hb672c48d),
	.w7(32'h37482dca),
	.w8(32'h37e72b6d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904f55a),
	.w1(32'hb92de535),
	.w2(32'hb91fd557),
	.w3(32'hb6004013),
	.w4(32'hb84e566f),
	.w5(32'hb8b474bb),
	.w6(32'h34d6f091),
	.w7(32'h3705b890),
	.w8(32'h37c95ad5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e190b5),
	.w1(32'hb832c6a3),
	.w2(32'hb8562d79),
	.w3(32'h3502190d),
	.w4(32'hb6a0b097),
	.w5(32'hb74865d6),
	.w6(32'h37d9f220),
	.w7(32'hb73ce358),
	.w8(32'h37404062),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9744d9c),
	.w1(32'hb923b195),
	.w2(32'h36e84b14),
	.w3(32'hb9875f24),
	.w4(32'hb8ef69f0),
	.w5(32'hb7449b9b),
	.w6(32'hb95d55c1),
	.w7(32'hb88e3cfe),
	.w8(32'hb7ed3f65),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9500f70),
	.w1(32'hb8878364),
	.w2(32'h376a2573),
	.w3(32'hb85aa3e0),
	.w4(32'hb68848fd),
	.w5(32'h380295be),
	.w6(32'hb8a4f0e6),
	.w7(32'hb875c666),
	.w8(32'hb679a2d2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9849775),
	.w1(32'hb90ca466),
	.w2(32'hb81c19cf),
	.w3(32'hb8a304d3),
	.w4(32'h37e2b42b),
	.w5(32'h3724977f),
	.w6(32'hb8f789b9),
	.w7(32'hb8ed7e7c),
	.w8(32'hb6ead930),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ecc03),
	.w1(32'hb98a7d8b),
	.w2(32'hb8e79617),
	.w3(32'h347313e9),
	.w4(32'hb788da76),
	.w5(32'hb7d0594d),
	.w6(32'hb7d1a8e1),
	.w7(32'h37c0c184),
	.w8(32'h387ee1a5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8811b0d),
	.w1(32'hb84cbb22),
	.w2(32'h3884e7d8),
	.w3(32'hb95f49e8),
	.w4(32'hb87e1a2b),
	.w5(32'h38640e8f),
	.w6(32'hb8d5584d),
	.w7(32'hb8acb315),
	.w8(32'h390785b9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e82b27),
	.w1(32'hb91402f0),
	.w2(32'hb735c62a),
	.w3(32'hb8dca242),
	.w4(32'hb8a38233),
	.w5(32'h36dc026c),
	.w6(32'hb8ab2383),
	.w7(32'hb7603e9f),
	.w8(32'h38198d2e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9084ce6),
	.w1(32'hb8ac5f26),
	.w2(32'hb71b148a),
	.w3(32'hb738b654),
	.w4(32'h386630d7),
	.w5(32'h384381bf),
	.w6(32'hb8ec1a79),
	.w7(32'h3834d4ab),
	.w8(32'h385a89b5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f682b4),
	.w1(32'h37d84756),
	.w2(32'h377acc84),
	.w3(32'h3793567d),
	.w4(32'h3888ccf5),
	.w5(32'h353f60c2),
	.w6(32'h377ae680),
	.w7(32'h382365d9),
	.w8(32'h389c1692),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7992110),
	.w1(32'hb8696f66),
	.w2(32'hb78393af),
	.w3(32'hb7650f93),
	.w4(32'hb6d46612),
	.w5(32'h36ce06b4),
	.w6(32'h37e46e5d),
	.w7(32'hb7886dfe),
	.w8(32'hb84ebebd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b34b73),
	.w1(32'hb7355c18),
	.w2(32'hb6eff9f3),
	.w3(32'hb555ed69),
	.w4(32'h3713e26c),
	.w5(32'hb6cdaa28),
	.w6(32'h37450c0f),
	.w7(32'h37b0f775),
	.w8(32'h368dba10),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810921c),
	.w1(32'hb8bbb332),
	.w2(32'h37e6f2a8),
	.w3(32'hb85ac017),
	.w4(32'h381a32c7),
	.w5(32'h36d6f72f),
	.w6(32'hb6875b9e),
	.w7(32'h37022484),
	.w8(32'h379b0ff2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ede728),
	.w1(32'h37739c7c),
	.w2(32'h364ea0b3),
	.w3(32'h36ad9fc0),
	.w4(32'h37d1ec0b),
	.w5(32'h37937bc3),
	.w6(32'h3626cff5),
	.w7(32'h36c10568),
	.w8(32'hb73f19d0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e1e3c6),
	.w1(32'hb3e0b2aa),
	.w2(32'hb5fa274f),
	.w3(32'hb5babea8),
	.w4(32'h351368c3),
	.w5(32'hb54c5526),
	.w6(32'hb5f32e99),
	.w7(32'hb48fee5f),
	.w8(32'hb58709ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36062261),
	.w1(32'h35bf261b),
	.w2(32'h35bd47de),
	.w3(32'h346cdffc),
	.w4(32'hb4db9ca2),
	.w5(32'h3521fec4),
	.w6(32'h35c1e5f8),
	.w7(32'h341f91ce),
	.w8(32'hb53af597),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e97c1c),
	.w1(32'h373cb20b),
	.w2(32'h364995d4),
	.w3(32'hb38a2eac),
	.w4(32'h372b49be),
	.w5(32'h36adf98f),
	.w6(32'hb60fdda2),
	.w7(32'h375d687d),
	.w8(32'hb68afb23),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387213f7),
	.w1(32'h38003cc4),
	.w2(32'h37e42cd4),
	.w3(32'h3820e8a8),
	.w4(32'h3788ca19),
	.w5(32'h379480be),
	.w6(32'h37ced3da),
	.w7(32'h375be537),
	.w8(32'h377fc13d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3be8b89),
	.w1(32'h385bee33),
	.w2(32'h38a3f047),
	.w3(32'hb8146db7),
	.w4(32'h3610d56e),
	.w5(32'h382849ff),
	.w6(32'hb844fdb9),
	.w7(32'h37d88dad),
	.w8(32'h36011251),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88932fa),
	.w1(32'h3800821c),
	.w2(32'h368460dc),
	.w3(32'hb80ff0be),
	.w4(32'h3857b7eb),
	.w5(32'hb801a27e),
	.w6(32'hb7656d84),
	.w7(32'h3831da11),
	.w8(32'hb82f07ca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe918b),
	.w1(32'hb844cdde),
	.w2(32'hb66afd1f),
	.w3(32'hb83a7797),
	.w4(32'hb89a8655),
	.w5(32'h37bbef5c),
	.w6(32'hb81c8a90),
	.w7(32'hb796604b),
	.w8(32'h34beb469),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7987dc1),
	.w1(32'hb7938652),
	.w2(32'hb662029b),
	.w3(32'hb74b8ae9),
	.w4(32'hb72b476e),
	.w5(32'h36bf5831),
	.w6(32'hb6b628da),
	.w7(32'h352a92d2),
	.w8(32'h36174f99),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4e7e239),
	.w1(32'hb3aeaeb0),
	.w2(32'h3549ebe1),
	.w3(32'hb44383d1),
	.w4(32'hb3cb6a2f),
	.w5(32'h3554cd80),
	.w6(32'h35374a32),
	.w7(32'h349f1a9e),
	.w8(32'h352dd706),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ef5c48),
	.w1(32'h36828788),
	.w2(32'hb4a48b87),
	.w3(32'h373aa9b7),
	.w4(32'h3693c418),
	.w5(32'hb64f3006),
	.w6(32'h368bffe1),
	.w7(32'hb71fbdfb),
	.w8(32'hb729e355),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364589d7),
	.w1(32'h35e0e096),
	.w2(32'h36669451),
	.w3(32'h360ecdf7),
	.w4(32'h3571fd7e),
	.w5(32'h3682dd54),
	.w6(32'h361c7647),
	.w7(32'h365f979e),
	.w8(32'h3641c03f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860bba4),
	.w1(32'hb87cf7b7),
	.w2(32'h38b0c987),
	.w3(32'h37ba2f84),
	.w4(32'hb886fb66),
	.w5(32'hb9044d93),
	.w6(32'hb788a2f6),
	.w7(32'h380581d3),
	.w8(32'hb6a99256),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb820b2be),
	.w1(32'hb656ebb3),
	.w2(32'hb7822594),
	.w3(32'hb845414e),
	.w4(32'h3792b6cb),
	.w5(32'h38256914),
	.w6(32'hb74084da),
	.w7(32'hb823db97),
	.w8(32'hb808b7c6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d6526),
	.w1(32'h35b73c3a),
	.w2(32'hb88722aa),
	.w3(32'hb8aee02a),
	.w4(32'hb6930f2d),
	.w5(32'hb80895a1),
	.w6(32'hb7cc1214),
	.w7(32'h37891dea),
	.w8(32'hb883abfc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f36a2),
	.w1(32'h37133c30),
	.w2(32'hb90e76d5),
	.w3(32'hb7974383),
	.w4(32'h37b4775c),
	.w5(32'h383a9da2),
	.w6(32'hb691a0c0),
	.w7(32'h38609647),
	.w8(32'h36391ad0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb55358ec),
	.w1(32'h354458f7),
	.w2(32'h35065a99),
	.w3(32'hb51e31a0),
	.w4(32'h3489d22b),
	.w5(32'h35942985),
	.w6(32'h36122001),
	.w7(32'h35e268cd),
	.w8(32'h35f4cb9b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5de76e9),
	.w1(32'hb612350f),
	.w2(32'h33ae51ce),
	.w3(32'hb5897b6b),
	.w4(32'hb5eefd68),
	.w5(32'h328483e7),
	.w6(32'h35944072),
	.w7(32'h3523c4c4),
	.w8(32'h3676982a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb656f8a2),
	.w1(32'hb61f2801),
	.w2(32'hb5d090a2),
	.w3(32'hb5696762),
	.w4(32'hb627ae63),
	.w5(32'hb635155d),
	.w6(32'h36c5cb50),
	.w7(32'h365aac5f),
	.w8(32'h36306801),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f6d3dd),
	.w1(32'h373f3024),
	.w2(32'hb6acd93a),
	.w3(32'h36ef96b8),
	.w4(32'h372195fc),
	.w5(32'h35843c62),
	.w6(32'h37bc3f64),
	.w7(32'h369c6a6d),
	.w8(32'hb7f459cb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8962e95),
	.w1(32'hb8768d38),
	.w2(32'hb81343c4),
	.w3(32'h360f022e),
	.w4(32'hb6c7d319),
	.w5(32'hb795847b),
	.w6(32'hb7611c80),
	.w7(32'h379479d3),
	.w8(32'h373fb63c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7afaa9b),
	.w1(32'hb7ad3e22),
	.w2(32'h382255b4),
	.w3(32'hb8755075),
	.w4(32'hb752984d),
	.w5(32'hb7ca42fd),
	.w6(32'hb7c9f51e),
	.w7(32'hb74657f4),
	.w8(32'h37d35f47),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37562c7a),
	.w1(32'h37ba86a8),
	.w2(32'hb8823791),
	.w3(32'hb9056acd),
	.w4(32'hb87e8e61),
	.w5(32'hb8a60b37),
	.w6(32'hb7fcd2fb),
	.w7(32'hb80c9564),
	.w8(32'hb8a19d1c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4277c),
	.w1(32'h384d14f1),
	.w2(32'h378b7705),
	.w3(32'hb7ee2db2),
	.w4(32'h3788e543),
	.w5(32'h3810578b),
	.w6(32'hb8904f1f),
	.w7(32'hb898922c),
	.w8(32'hb80b3d69),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b306ba),
	.w1(32'hb70a3ebc),
	.w2(32'hb7e946f5),
	.w3(32'hb8156b5f),
	.w4(32'hb80f3df1),
	.w5(32'hb84294a9),
	.w6(32'hb86d5542),
	.w7(32'hb89c5d39),
	.w8(32'hb89d900b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bdac4b),
	.w1(32'hb638ddd7),
	.w2(32'h38114692),
	.w3(32'h36708eca),
	.w4(32'hb73acddf),
	.w5(32'hb8157a66),
	.w6(32'hb7fb4a58),
	.w7(32'h3782e55d),
	.w8(32'h37d169d1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76513be),
	.w1(32'h376d4929),
	.w2(32'h363ec2ff),
	.w3(32'hb724f63e),
	.w4(32'h3607aacf),
	.w5(32'hb55fa718),
	.w6(32'hb845ec0b),
	.w7(32'hb827a1bb),
	.w8(32'hb84fb41a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acde38),
	.w1(32'h37adaf21),
	.w2(32'h376c0c71),
	.w3(32'hb844919d),
	.w4(32'hb7b2a308),
	.w5(32'hb74cf512),
	.w6(32'hb8088271),
	.w7(32'hb82cc2db),
	.w8(32'hb6ee5ae6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4c0f143),
	.w1(32'hb334c547),
	.w2(32'h3485277c),
	.w3(32'hb395b366),
	.w4(32'h34195d84),
	.w5(32'h3503dc7e),
	.w6(32'h349b487a),
	.w7(32'h34f6e967),
	.w8(32'h34f82d15),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354b4bd6),
	.w1(32'h34e5ba61),
	.w2(32'h364c98f5),
	.w3(32'h3486ba5b),
	.w4(32'hb50bce2b),
	.w5(32'h35d7cba7),
	.w6(32'hb561ac2f),
	.w7(32'hb510a7ce),
	.w8(32'h355ea8c8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3570361a),
	.w1(32'h3592f958),
	.w2(32'h359ec3fa),
	.w3(32'h35a205cc),
	.w4(32'h34964991),
	.w5(32'hb29101fb),
	.w6(32'hb4a49a5e),
	.w7(32'h34d0c540),
	.w8(32'h359139a4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fbb029),
	.w1(32'h367a84f2),
	.w2(32'h371006db),
	.w3(32'hb4ce4d39),
	.w4(32'h374fcc65),
	.w5(32'h3776623b),
	.w6(32'hb71f302a),
	.w7(32'h3602d068),
	.w8(32'h36a0444d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ed0c1),
	.w1(32'h370602fa),
	.w2(32'hb7cabaaf),
	.w3(32'h35fa034d),
	.w4(32'h37b2486b),
	.w5(32'h38815088),
	.w6(32'h374b110a),
	.w7(32'h3767d5c6),
	.w8(32'h36e66cb5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb724e935),
	.w1(32'hb6cb0e62),
	.w2(32'h360e47a9),
	.w3(32'hb65666ac),
	.w4(32'h35e0df1e),
	.w5(32'h36a56947),
	.w6(32'hb68b3eca),
	.w7(32'h364120de),
	.w8(32'h36aec53b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80211f5),
	.w1(32'h376c1a11),
	.w2(32'h36928299),
	.w3(32'hb70b95f8),
	.w4(32'h373b82b9),
	.w5(32'h37e5efe5),
	.w6(32'h377df9bd),
	.w7(32'h37c65f27),
	.w8(32'h37cea7dc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9470b96),
	.w1(32'hb91cdda0),
	.w2(32'hb8ac7e2c),
	.w3(32'hb90677d1),
	.w4(32'hb891b1e5),
	.w5(32'hb89c5731),
	.w6(32'hb7c43557),
	.w7(32'h38db8baa),
	.w8(32'h388fce76),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c471c2),
	.w1(32'h383f2ed6),
	.w2(32'h37f15d1f),
	.w3(32'h35c4ccaf),
	.w4(32'h3887814a),
	.w5(32'h38047311),
	.w6(32'hb8020e7b),
	.w7(32'h385815c6),
	.w8(32'h37c072ed),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38044c4f),
	.w1(32'h38d8887c),
	.w2(32'h38e84164),
	.w3(32'h3621949b),
	.w4(32'h386d3cf1),
	.w5(32'h3821d0aa),
	.w6(32'hb80e4286),
	.w7(32'h37e004d1),
	.w8(32'h3844e083),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a402bc),
	.w1(32'h38d92338),
	.w2(32'hb7e83947),
	.w3(32'h389fbf7e),
	.w4(32'h3833cd3d),
	.w5(32'hb82407bc),
	.w6(32'h38aa4260),
	.w7(32'h37483ed6),
	.w8(32'hb8794164),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a89b8a),
	.w1(32'hb8891fea),
	.w2(32'hb84433ad),
	.w3(32'hb8d31617),
	.w4(32'hb810925f),
	.w5(32'hb898769f),
	.w6(32'hb87c828c),
	.w7(32'h36ddc38b),
	.w8(32'hb760256e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e2a67),
	.w1(32'h3828df7c),
	.w2(32'h38139759),
	.w3(32'hb7df3d7b),
	.w4(32'h36276472),
	.w5(32'h37d6fef5),
	.w6(32'hb8978874),
	.w7(32'hb792244c),
	.w8(32'h379a5104),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8ea69),
	.w1(32'hb6e82e14),
	.w2(32'h35affcf8),
	.w3(32'hb73b109f),
	.w4(32'h384a33a1),
	.w5(32'h37615fac),
	.w6(32'h37db8bdc),
	.w7(32'h38b37ebb),
	.w8(32'h38af2596),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8229c2a),
	.w1(32'hb813403d),
	.w2(32'hb8da50b6),
	.w3(32'h375756bb),
	.w4(32'h36e530cb),
	.w5(32'hb7aa55c3),
	.w6(32'hb7ad0b14),
	.w7(32'h3777d973),
	.w8(32'hb7cfcb7b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f45671),
	.w1(32'hb9473311),
	.w2(32'hb931d705),
	.w3(32'hb8b75399),
	.w4(32'hb90a71ed),
	.w5(32'hb8daf883),
	.w6(32'hb854ed33),
	.w7(32'hb873ea87),
	.w8(32'hb8be5d90),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8112b55),
	.w1(32'hb9072ad8),
	.w2(32'hb8333683),
	.w3(32'h39083bab),
	.w4(32'hb8deb2fc),
	.w5(32'hb898da14),
	.w6(32'h3537e779),
	.w7(32'h38313ca5),
	.w8(32'h37f644ae),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df1bbb),
	.w1(32'hb8c746a6),
	.w2(32'hb82594c0),
	.w3(32'hb976b25e),
	.w4(32'h3766f30f),
	.w5(32'hb7d148d2),
	.w6(32'hb7b74220),
	.w7(32'hb7ea8c78),
	.w8(32'h37d0bed2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84e2d3d),
	.w1(32'hb908ac92),
	.w2(32'h372c9ea1),
	.w3(32'h38f91115),
	.w4(32'hb607ee00),
	.w5(32'hb830b9c1),
	.w6(32'hb91c1f2f),
	.w7(32'hb8952f83),
	.w8(32'hb6b4dafb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eeaa05),
	.w1(32'h390a8b8c),
	.w2(32'h391ad56e),
	.w3(32'h36995c54),
	.w4(32'h390265ae),
	.w5(32'h38bb66fa),
	.w6(32'hb7dfe0a6),
	.w7(32'hb8f96fd4),
	.w8(32'hb80c07d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8755db6),
	.w1(32'h38887b8b),
	.w2(32'h397683ec),
	.w3(32'hb94b003a),
	.w4(32'hb783f109),
	.w5(32'h3885cf2d),
	.w6(32'hb82faeba),
	.w7(32'h3852a9f6),
	.w8(32'h393f7a91),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9373dbe),
	.w1(32'hb8985a59),
	.w2(32'hb9064ae0),
	.w3(32'h37f266d3),
	.w4(32'hb752c82c),
	.w5(32'hb8cfc9f5),
	.w6(32'h381b7b5f),
	.w7(32'h3846998d),
	.w8(32'hb88ef624),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a4896a),
	.w1(32'hb8594262),
	.w2(32'hb8798b85),
	.w3(32'hb9829184),
	.w4(32'hb8926f12),
	.w5(32'hb8822cf1),
	.w6(32'hb83c8f97),
	.w7(32'hb835d782),
	.w8(32'hb8701c24),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3745622a),
	.w1(32'h38845e47),
	.w2(32'hb82bba61),
	.w3(32'hb71fab3e),
	.w4(32'h387f89f5),
	.w5(32'h37ad28b6),
	.w6(32'hb829ead8),
	.w7(32'hb676ab81),
	.w8(32'hb88917e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375c0f69),
	.w1(32'h3781b17e),
	.w2(32'hb4babe0e),
	.w3(32'h37e19a0c),
	.w4(32'h37e9c8c1),
	.w5(32'h36b85208),
	.w6(32'h37690fb0),
	.w7(32'h37ad2359),
	.w8(32'hb7217077),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c9e28),
	.w1(32'h37cbbfab),
	.w2(32'h37fb33ba),
	.w3(32'h35960622),
	.w4(32'h36e4a70a),
	.w5(32'h37f3ab3c),
	.w6(32'hb6a022bb),
	.w7(32'h369a8a36),
	.w8(32'h3813d5eb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbc20f),
	.w1(32'hb8a41409),
	.w2(32'hb8fe8704),
	.w3(32'hb7bc2b70),
	.w4(32'hb86f10ab),
	.w5(32'hb8f7b103),
	.w6(32'hb6fe8534),
	.w7(32'hb8db7a28),
	.w8(32'hb893da0d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93242a6),
	.w1(32'hb88824b6),
	.w2(32'hb7a38f1f),
	.w3(32'hb8a2c4ff),
	.w4(32'hb822db63),
	.w5(32'h37c08f46),
	.w6(32'hb9159838),
	.w7(32'hb8d20dd5),
	.w8(32'hb7ae037b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84bbbc8),
	.w1(32'h35aa2c7f),
	.w2(32'h3821d01c),
	.w3(32'hb8937692),
	.w4(32'h3527e6fb),
	.w5(32'h37b0d959),
	.w6(32'hb8ece3a2),
	.w7(32'h3483e7c9),
	.w8(32'hb72b0995),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f84e85),
	.w1(32'hb7981e45),
	.w2(32'h38f3efef),
	.w3(32'hb859bc16),
	.w4(32'h376fb0ad),
	.w5(32'h38b13380),
	.w6(32'hb8cdee41),
	.w7(32'hb81cc540),
	.w8(32'h38c8075e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb38ee93a),
	.w1(32'h388180d2),
	.w2(32'h37914f19),
	.w3(32'hb81a2c06),
	.w4(32'h37853a29),
	.w5(32'h389eb6ac),
	.w6(32'h389fab2c),
	.w7(32'h37ec1533),
	.w8(32'h3876118d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378270b7),
	.w1(32'h3825c805),
	.w2(32'h39017882),
	.w3(32'hb81b0407),
	.w4(32'h377095d7),
	.w5(32'h382d3261),
	.w6(32'hb81304bf),
	.w7(32'hb7862cfc),
	.w8(32'hb86d6fd8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb784f749),
	.w1(32'h3701fbd7),
	.w2(32'h37c2a043),
	.w3(32'h3734c3bc),
	.w4(32'h37dc95a8),
	.w5(32'h37d62b57),
	.w6(32'h36a04fb8),
	.w7(32'h376314ff),
	.w8(32'h36bea6c6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6881031),
	.w1(32'hb6020679),
	.w2(32'hb5a8ee3a),
	.w3(32'hb5c4551a),
	.w4(32'hb56aca9b),
	.w5(32'h35c19a30),
	.w6(32'hb62238e9),
	.w7(32'hb61bf3d1),
	.w8(32'hb4c9d72f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63c7648),
	.w1(32'h365dd545),
	.w2(32'h3660421a),
	.w3(32'hb716ef4d),
	.w4(32'h36374307),
	.w5(32'h36ce20a5),
	.w6(32'hb70bfc40),
	.w7(32'h36acf14c),
	.w8(32'h3706cd08),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb575b5c0),
	.w1(32'hb61ce5ec),
	.w2(32'hb425a74b),
	.w3(32'hb5898db5),
	.w4(32'hb5ec2d14),
	.w5(32'h35a27269),
	.w6(32'hb590b837),
	.w7(32'hb4dacda1),
	.w8(32'h351e3001),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dca2fa),
	.w1(32'hb67f22e1),
	.w2(32'hb6bac252),
	.w3(32'hb6b6a96d),
	.w4(32'h35b16303),
	.w5(32'h3597f944),
	.w6(32'hb64379e8),
	.w7(32'h36885b87),
	.w8(32'hb14980f1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375fc2fa),
	.w1(32'h384624dc),
	.w2(32'hb739bf35),
	.w3(32'h380aec7c),
	.w4(32'h3802b3c7),
	.w5(32'hb751faac),
	.w6(32'hb80f22f5),
	.w7(32'hb8403738),
	.w8(32'hb85d874e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75b53b8),
	.w1(32'hb77b495a),
	.w2(32'hb4bbea77),
	.w3(32'hb730acf5),
	.w4(32'hb720401e),
	.w5(32'h34d02168),
	.w6(32'hb794b7c8),
	.w7(32'hb7ab2701),
	.w8(32'h36d30d8e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804c0ce),
	.w1(32'h383a7d1b),
	.w2(32'h38343910),
	.w3(32'hb855e8ff),
	.w4(32'h378618d6),
	.w5(32'hb650461d),
	.w6(32'hb7f6e1a4),
	.w7(32'hb7f67bc0),
	.w8(32'h378c6770),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9162cda),
	.w1(32'hb80562cb),
	.w2(32'h3896588a),
	.w3(32'hb8e7453e),
	.w4(32'hb71bef3d),
	.w5(32'h38ac1561),
	.w6(32'hb8bd1396),
	.w7(32'hb82048c1),
	.w8(32'hb6e386dd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35acf389),
	.w1(32'hb326690a),
	.w2(32'h35064be9),
	.w3(32'h35968699),
	.w4(32'hb58e2c05),
	.w5(32'h3509384f),
	.w6(32'h355bbeee),
	.w7(32'h338ce228),
	.w8(32'h35999358),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f4165),
	.w1(32'hb772759d),
	.w2(32'hb71783fb),
	.w3(32'hb6fe422c),
	.w4(32'hb71c5675),
	.w5(32'hb7056bfc),
	.w6(32'hb6b71f3c),
	.w7(32'hb70507a7),
	.w8(32'hb5718998),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3698f685),
	.w1(32'h36a55654),
	.w2(32'h369899ca),
	.w3(32'h36ebec5d),
	.w4(32'h37334e4e),
	.w5(32'h372da09d),
	.w6(32'h371569b7),
	.w7(32'h361fb5ec),
	.w8(32'h36af7d83),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62da497),
	.w1(32'hba1017f6),
	.w2(32'hba317237),
	.w3(32'h372a2764),
	.w4(32'h3927090a),
	.w5(32'hb82d29c0),
	.w6(32'hb8cfc129),
	.w7(32'hb9e5dcde),
	.w8(32'hb87dafca),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39894f65),
	.w1(32'h3841263a),
	.w2(32'hb9a9af0a),
	.w3(32'h3a0a511f),
	.w4(32'h3a03e350),
	.w5(32'h39cd3edf),
	.w6(32'h398c23c7),
	.w7(32'hb8d5ea83),
	.w8(32'h3905958d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380113c8),
	.w1(32'h3b0a977d),
	.w2(32'h3a823e82),
	.w3(32'h3a1d78de),
	.w4(32'h3a007f96),
	.w5(32'hbac2529f),
	.w6(32'h3a65af0a),
	.w7(32'h3a2d315c),
	.w8(32'h3a8ae42c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb801),
	.w1(32'h3913676e),
	.w2(32'h398678c2),
	.w3(32'hba3ea617),
	.w4(32'h39ab6fa5),
	.w5(32'h3942d4e9),
	.w6(32'hb8a55524),
	.w7(32'h399e83ce),
	.w8(32'h38ce426d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394650f8),
	.w1(32'hba0a5cc2),
	.w2(32'hba3a28cf),
	.w3(32'h3931a5f9),
	.w4(32'hb9ec8d8a),
	.w5(32'hba43b7d2),
	.w6(32'h39114713),
	.w7(32'h3923cfb6),
	.w8(32'h37835b64),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d5487),
	.w1(32'hbb22539b),
	.w2(32'hbab71202),
	.w3(32'hb98a08f6),
	.w4(32'h39fcaef6),
	.w5(32'h38912e4c),
	.w6(32'h393ef941),
	.w7(32'hbaa0453d),
	.w8(32'hba497047),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9d0ef),
	.w1(32'hb9564ba7),
	.w2(32'hbab7395d),
	.w3(32'hb9439fc2),
	.w4(32'h394ee7f0),
	.w5(32'hba5d6569),
	.w6(32'h375e24cc),
	.w7(32'hba0f4804),
	.w8(32'h39b1ffc4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98751ab),
	.w1(32'hb7bf6675),
	.w2(32'hb954489c),
	.w3(32'hb9fb69c1),
	.w4(32'h39aeeecb),
	.w5(32'h395d835b),
	.w6(32'hb8dde5b0),
	.w7(32'hba24c5ec),
	.w8(32'hb9e0451c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7693d8b),
	.w1(32'h384a2cd8),
	.w2(32'h3a066b23),
	.w3(32'h399c6ad7),
	.w4(32'hb91a044a),
	.w5(32'hb9dda3b8),
	.w6(32'hb9dfd2f1),
	.w7(32'h38a603fc),
	.w8(32'h38db4a24),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb808ac4a),
	.w1(32'hb9354974),
	.w2(32'hb9c81005),
	.w3(32'hb8e1221e),
	.w4(32'h3a0de4df),
	.w5(32'h3a20315e),
	.w6(32'h3990bd2b),
	.w7(32'h398ae784),
	.w8(32'h3a032e3f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39025a4c),
	.w1(32'hb9a574fb),
	.w2(32'hb985b566),
	.w3(32'h3a43f466),
	.w4(32'h37c591c2),
	.w5(32'h38bf8472),
	.w6(32'hb9a3f6b1),
	.w7(32'hb94635ea),
	.w8(32'hb7e6f144),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e70b8),
	.w1(32'h390eed29),
	.w2(32'h39c65669),
	.w3(32'h3727df36),
	.w4(32'h39bad1e3),
	.w5(32'hb8c309d5),
	.w6(32'hb9174b2b),
	.w7(32'hb9477652),
	.w8(32'hb8ac0047),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39562ee8),
	.w1(32'hbafa48e5),
	.w2(32'hba8ff3d0),
	.w3(32'hb91552af),
	.w4(32'hba17c06b),
	.w5(32'h38ec7aeb),
	.w6(32'hb93fe6a3),
	.w7(32'hba0cabad),
	.w8(32'hba330aa2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e8ddd),
	.w1(32'hba003a60),
	.w2(32'h3a9a8f9b),
	.w3(32'h39ce6cce),
	.w4(32'h385afb72),
	.w5(32'h3a8992db),
	.w6(32'h39079eb0),
	.w7(32'h393baaf6),
	.w8(32'hb98de0d2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23f3bb),
	.w1(32'hba345b42),
	.w2(32'hba1874c8),
	.w3(32'h396d1b3e),
	.w4(32'hb910ef6b),
	.w5(32'h38abc03c),
	.w6(32'hba05d250),
	.w7(32'hba34f6a6),
	.w8(32'hb9c17aa8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999d1fc),
	.w1(32'hb95c41c7),
	.w2(32'h390a18d7),
	.w3(32'h3963efdb),
	.w4(32'h3a95a0bc),
	.w5(32'h3aebe6f6),
	.w6(32'h39c5847b),
	.w7(32'h3a3c8ad9),
	.w8(32'h3abefd13),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a246388),
	.w1(32'hba206d1d),
	.w2(32'h39171eb2),
	.w3(32'h3aef6aad),
	.w4(32'h3a82a784),
	.w5(32'h3a8c2615),
	.w6(32'h3886832f),
	.w7(32'hb94a3be6),
	.w8(32'hb9bed880),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960321f),
	.w1(32'h3808a32a),
	.w2(32'hb98f1944),
	.w3(32'h3a09c987),
	.w4(32'hb7f0cfcd),
	.w5(32'h3837969a),
	.w6(32'h37283981),
	.w7(32'hb9610402),
	.w8(32'hb8f43f96),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9905131),
	.w1(32'h3a2df051),
	.w2(32'h39ef200f),
	.w3(32'h38cd2fb8),
	.w4(32'hba5573ae),
	.w5(32'hbab8d939),
	.w6(32'hb7f917ea),
	.w7(32'hb90abdd6),
	.w8(32'hbab99305),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19bbdb),
	.w1(32'hb9eb3962),
	.w2(32'h3912a12f),
	.w3(32'hbb083b8c),
	.w4(32'hb7ec311d),
	.w5(32'h3844fab0),
	.w6(32'hba16f3d4),
	.w7(32'hb9aa9227),
	.w8(32'hb95d39f1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebff44),
	.w1(32'hb96177d7),
	.w2(32'hb99c8146),
	.w3(32'hb5bf4503),
	.w4(32'hb9388e1b),
	.w5(32'hba000c6e),
	.w6(32'hb9bdb79b),
	.w7(32'h35c0783a),
	.w8(32'hb9ae380a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea30c3),
	.w1(32'hb943405b),
	.w2(32'h36862f33),
	.w3(32'hb9e0259f),
	.w4(32'h36e4aef4),
	.w5(32'h3931e963),
	.w6(32'hb90ab244),
	.w7(32'hb8dd3ce2),
	.w8(32'hb9157bf4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9819c16),
	.w1(32'hb851227f),
	.w2(32'hb931f1e9),
	.w3(32'hb7c47cff),
	.w4(32'h39ede006),
	.w5(32'hb894637b),
	.w6(32'h38bf2595),
	.w7(32'hb934c7ea),
	.w8(32'h37d45a09),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7e7d1),
	.w1(32'hbb24b902),
	.w2(32'h3a8d5c86),
	.w3(32'h38f5b00f),
	.w4(32'h39da6744),
	.w5(32'hb8b4a6e1),
	.w6(32'hba5611bb),
	.w7(32'hba988f1e),
	.w8(32'hba126daa),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce1ad),
	.w1(32'h38ff1a72),
	.w2(32'hb938d7a6),
	.w3(32'hb7b48726),
	.w4(32'hb99e2db6),
	.w5(32'hbaa6f44d),
	.w6(32'h39779f18),
	.w7(32'hb98d3b25),
	.w8(32'hba8b036a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ce03),
	.w1(32'hb7de4fbe),
	.w2(32'hb9b264cc),
	.w3(32'hbb08c3c2),
	.w4(32'h39f63133),
	.w5(32'h3a08485d),
	.w6(32'h392a519a),
	.w7(32'h3911cca0),
	.w8(32'h398f462d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937fd2d),
	.w1(32'h39851e0d),
	.w2(32'h37e77cbf),
	.w3(32'h3a2e6525),
	.w4(32'h39282aba),
	.w5(32'hb70f4288),
	.w6(32'hb8be75e0),
	.w7(32'hba06174a),
	.w8(32'hb8bd7dbc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de75df),
	.w1(32'h39b33f3c),
	.w2(32'h3b2bbb7a),
	.w3(32'h393c9256),
	.w4(32'hbafeb17b),
	.w5(32'hbb0e317a),
	.w6(32'hb8efb6a8),
	.w7(32'hba26accd),
	.w8(32'hb9876d22),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018c3d),
	.w1(32'hb96ed384),
	.w2(32'h398801e3),
	.w3(32'hbaead111),
	.w4(32'h38c3d9a7),
	.w5(32'h39e89e69),
	.w6(32'hb9c214ed),
	.w7(32'h38a186c4),
	.w8(32'hb94025b6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f01e09),
	.w1(32'hb9c269b8),
	.w2(32'hba2511d1),
	.w3(32'h37ee3834),
	.w4(32'hb9b6a721),
	.w5(32'h3960ac46),
	.w6(32'hb8c84753),
	.w7(32'hba4d1ead),
	.w8(32'h39dd4f25),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1b1d4),
	.w1(32'hb9edc069),
	.w2(32'h3935bdba),
	.w3(32'h39bdbd65),
	.w4(32'hba18c20f),
	.w5(32'hb985266b),
	.w6(32'h37b0b6d2),
	.w7(32'h378dedf5),
	.w8(32'h38455f66),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9520d6a),
	.w1(32'h39a06897),
	.w2(32'hb9a1a2a4),
	.w3(32'hba142757),
	.w4(32'hb9eb5b98),
	.w5(32'hbac53093),
	.w6(32'h3a0245d8),
	.w7(32'h39dcceb0),
	.w8(32'h398ef2e5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e096b),
	.w1(32'h38808209),
	.w2(32'hb90b619b),
	.w3(32'hbaa4ff86),
	.w4(32'h39f0bf36),
	.w5(32'h39860911),
	.w6(32'hb8de36b8),
	.w7(32'hb9740ae8),
	.w8(32'hb9738ed5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947f90e),
	.w1(32'hba0b69c7),
	.w2(32'hb9ab3815),
	.w3(32'h3987bbc8),
	.w4(32'hb8ac10d0),
	.w5(32'h389b34df),
	.w6(32'hb9e1b8f6),
	.w7(32'hba2641ac),
	.w8(32'hb9c7fb29),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e2523),
	.w1(32'h39c855f1),
	.w2(32'hba739572),
	.w3(32'h3931f169),
	.w4(32'h38d90abd),
	.w5(32'hba2d6212),
	.w6(32'hb56f7ce6),
	.w7(32'hb95fd0b8),
	.w8(32'hb9b76557),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855f16),
	.w1(32'hbacaaf8d),
	.w2(32'hb916062f),
	.w3(32'hba6acbd7),
	.w4(32'hbab6fc90),
	.w5(32'hba0f980d),
	.w6(32'hb997a634),
	.w7(32'h3983f60c),
	.w8(32'h3a502afb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca7439),
	.w1(32'hba5ecdd8),
	.w2(32'h39b3356b),
	.w3(32'hb8b04280),
	.w4(32'hb94f7f8a),
	.w5(32'h39456554),
	.w6(32'hba53138b),
	.w7(32'hba4dab21),
	.w8(32'hb9c43cfa),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39add94e),
	.w1(32'hb9dbffe9),
	.w2(32'hb7ae9b41),
	.w3(32'h3849824a),
	.w4(32'hb90f124b),
	.w5(32'h36e74784),
	.w6(32'hb9cec504),
	.w7(32'hba1fc050),
	.w8(32'hba09b2ff),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904605b),
	.w1(32'hba096d8b),
	.w2(32'hb8a416d8),
	.w3(32'hb876c4f8),
	.w4(32'h388a591a),
	.w5(32'h3a05f0d2),
	.w6(32'hba32d4cf),
	.w7(32'hb96a78a4),
	.w8(32'hb9661ca3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0c529),
	.w1(32'h3915c838),
	.w2(32'h396eee00),
	.w3(32'h3983cdac),
	.w4(32'hb8310faa),
	.w5(32'hba00a73c),
	.w6(32'hb9817b8c),
	.w7(32'h3976d6da),
	.w8(32'h3663f3e1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371fff48),
	.w1(32'hb82e2369),
	.w2(32'hb9b6104b),
	.w3(32'hb9921cb3),
	.w4(32'h39e123f2),
	.w5(32'h39bd6f8f),
	.w6(32'h39259920),
	.w7(32'h37dd6717),
	.w8(32'h39499a06),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9010d46),
	.w1(32'hb9b9826f),
	.w2(32'hb9589d45),
	.w3(32'h39f44b08),
	.w4(32'hb9e936cf),
	.w5(32'hb92ee0c8),
	.w6(32'hba31e99e),
	.w7(32'hb92d5971),
	.w8(32'hb71b2df4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0772a),
	.w1(32'h382d4fec),
	.w2(32'hb98b3d3a),
	.w3(32'h37b59167),
	.w4(32'hba4daafd),
	.w5(32'hba895949),
	.w6(32'h390593a7),
	.w7(32'h399f3039),
	.w8(32'h39fe6d7d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a107a7),
	.w1(32'hba306991),
	.w2(32'hb832a62c),
	.w3(32'hba538d41),
	.w4(32'hba1ac21a),
	.w5(32'hb7a1483a),
	.w6(32'h39062521),
	.w7(32'h381c455e),
	.w8(32'hb8dd9385),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b6e6),
	.w1(32'hba24df59),
	.w2(32'hb9b8641b),
	.w3(32'h38f20d49),
	.w4(32'hb93fc7f0),
	.w5(32'h39403ba0),
	.w6(32'hb9d1d9fd),
	.w7(32'hb9ee277c),
	.w8(32'hb9c88895),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348229),
	.w1(32'h39b6b845),
	.w2(32'h393c6999),
	.w3(32'hb8bd87d1),
	.w4(32'h3a5114f8),
	.w5(32'hb8bcdcd3),
	.w6(32'h38c8182d),
	.w7(32'h392ffc32),
	.w8(32'h3a0632a1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20f9ae),
	.w1(32'h39b5721f),
	.w2(32'hb9486c78),
	.w3(32'h3a26c247),
	.w4(32'h3a7ca439),
	.w5(32'hb9507425),
	.w6(32'h38ad48c0),
	.w7(32'h39568c78),
	.w8(32'hb7aacc94),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dec1e6),
	.w1(32'hba3b1f77),
	.w2(32'h395d319e),
	.w3(32'h392e6066),
	.w4(32'hb9172a75),
	.w5(32'h38d08528),
	.w6(32'hb9b5f439),
	.w7(32'h38861fd5),
	.w8(32'h399b96c3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf22e8),
	.w1(32'hba170e65),
	.w2(32'h3aa90d03),
	.w3(32'h39831590),
	.w4(32'h3a2db3a3),
	.w5(32'h3a5fc6f9),
	.w6(32'h3a095624),
	.w7(32'hb9299c71),
	.w8(32'hb8a879c9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394585c3),
	.w1(32'hb86833c9),
	.w2(32'h392903a1),
	.w3(32'hb8af7394),
	.w4(32'hba17e6c9),
	.w5(32'hba1349ed),
	.w6(32'hb973387f),
	.w7(32'h381f914d),
	.w8(32'h397d00ea),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce9af),
	.w1(32'hba725a72),
	.w2(32'hb89734dc),
	.w3(32'hb9f69318),
	.w4(32'hb9f28dee),
	.w5(32'hb89cc77c),
	.w6(32'hba1d56ab),
	.w7(32'hba14d6ee),
	.w8(32'hba0c9918),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fd4ff),
	.w1(32'hb75ec321),
	.w2(32'hb9c52ddb),
	.w3(32'hb948cdc2),
	.w4(32'h3a12b79c),
	.w5(32'h3a27ef20),
	.w6(32'h39a03a4c),
	.w7(32'h39a7df48),
	.w8(32'h3a0f545e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39148469),
	.w1(32'h3813d384),
	.w2(32'h3991e5bf),
	.w3(32'h3a64d114),
	.w4(32'hb8183fa2),
	.w5(32'h3924e22a),
	.w6(32'hb8687e40),
	.w7(32'h398b8481),
	.w8(32'h39ba3e61),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cc5371),
	.w1(32'h3670a0d9),
	.w2(32'hbb526740),
	.w3(32'h39b7d1fe),
	.w4(32'h3a9e46d8),
	.w5(32'h3a868dec),
	.w6(32'h3aa10fd4),
	.w7(32'hba948b17),
	.w8(32'h3a113c0e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70b3e1),
	.w1(32'h3a8139df),
	.w2(32'h3a20c3c2),
	.w3(32'h3acff20a),
	.w4(32'h3a62e877),
	.w5(32'h3a00fa7e),
	.w6(32'h3a1ba6f2),
	.w7(32'h38fb7ac8),
	.w8(32'h3956fd0a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dacc84),
	.w1(32'hba591cfd),
	.w2(32'hba30a31e),
	.w3(32'h3a46a106),
	.w4(32'hba0b674e),
	.w5(32'hba2d43fe),
	.w6(32'hba41efc4),
	.w7(32'hb9bbf1ac),
	.w8(32'hb935cdd7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f924ec),
	.w1(32'h3a096f65),
	.w2(32'h3a8357e3),
	.w3(32'hba08593f),
	.w4(32'h381714e0),
	.w5(32'hb954e3d7),
	.w6(32'h39db7a16),
	.w7(32'h39e470d1),
	.w8(32'hb9757d0f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ff487),
	.w1(32'h38fdd5a1),
	.w2(32'hb9a1b289),
	.w3(32'hb9f79a7d),
	.w4(32'hba2cc47d),
	.w5(32'hba07f1df),
	.w6(32'h3a5d078f),
	.w7(32'h3a591089),
	.w8(32'h3a64444c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8663831),
	.w1(32'hb94a9b67),
	.w2(32'h39e6f7f5),
	.w3(32'h37078b25),
	.w4(32'hb9ca4dd4),
	.w5(32'h390c0c0c),
	.w6(32'hb9affaf9),
	.w7(32'h3a20d1f2),
	.w8(32'h391843af),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb646a),
	.w1(32'hba35cfc6),
	.w2(32'hbb07bbaf),
	.w3(32'hb97bfc4b),
	.w4(32'hba0cd19a),
	.w5(32'hbaa7dd59),
	.w6(32'hb9caa2c1),
	.w7(32'hba3dd26d),
	.w8(32'h39f35ccf),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd09a5),
	.w1(32'h397bef75),
	.w2(32'hb9105192),
	.w3(32'h398c4e5d),
	.w4(32'h39ae6930),
	.w5(32'hb9e327ec),
	.w6(32'hb8bc8031),
	.w7(32'h39780cb2),
	.w8(32'h3992d467),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924e351),
	.w1(32'hb9a370ba),
	.w2(32'hba241587),
	.w3(32'h38d75ccb),
	.w4(32'h398b49f7),
	.w5(32'h393463de),
	.w6(32'h3796d85c),
	.w7(32'hb8dbed32),
	.w8(32'hb8d05ac2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7acbd),
	.w1(32'hb97228a7),
	.w2(32'hb994389f),
	.w3(32'h39df7d1f),
	.w4(32'hb9ef8945),
	.w5(32'hba2bcc8e),
	.w6(32'hb923fd14),
	.w7(32'h39c464e8),
	.w8(32'h38ab69f0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a497d7),
	.w1(32'hb962c896),
	.w2(32'hba0ca3aa),
	.w3(32'hb9838c82),
	.w4(32'h3a343cb9),
	.w5(32'h3a61a373),
	.w6(32'hb952d2fd),
	.w7(32'hb910fac8),
	.w8(32'hb91f26be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd36b1),
	.w1(32'h393dbda3),
	.w2(32'hbb25052c),
	.w3(32'h3a58b0b4),
	.w4(32'hb92ada61),
	.w5(32'hba7b2ca2),
	.w6(32'hba9accdf),
	.w7(32'hbacab943),
	.w8(32'hba2f68f0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0800b2),
	.w1(32'h39123881),
	.w2(32'h397f895a),
	.w3(32'hba553808),
	.w4(32'h39d34089),
	.w5(32'hb8c8059b),
	.w6(32'hb6e72720),
	.w7(32'h37622f64),
	.w8(32'h3947d44d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc4efe),
	.w1(32'h3869c786),
	.w2(32'hb9d3b010),
	.w3(32'h39ba1533),
	.w4(32'hb7d56095),
	.w5(32'hb9977876),
	.w6(32'hb994de57),
	.w7(32'hb984fba5),
	.w8(32'hba0ebaa0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29e8c3),
	.w1(32'hba7d840e),
	.w2(32'hbacbe265),
	.w3(32'hb999faf7),
	.w4(32'hba255719),
	.w5(32'hba68990d),
	.w6(32'hb9d3316f),
	.w7(32'hba14061b),
	.w8(32'h39381eae),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09774d),
	.w1(32'h39159cee),
	.w2(32'hb9af43ed),
	.w3(32'h3915bd9d),
	.w4(32'hba2bf05b),
	.w5(32'hba671e9d),
	.w6(32'h39d888c7),
	.w7(32'h38c10ab7),
	.w8(32'h39b2beb2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924594d),
	.w1(32'h3897189b),
	.w2(32'hb7a27479),
	.w3(32'hb9eff8b7),
	.w4(32'hba556662),
	.w5(32'hbad9fea0),
	.w6(32'h37c21375),
	.w7(32'hb88504ba),
	.w8(32'hb88fe81d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c4a70),
	.w1(32'h39e78207),
	.w2(32'h391aa670),
	.w3(32'hbad55cf2),
	.w4(32'h39f631a5),
	.w5(32'h3921a181),
	.w6(32'h39aaea99),
	.w7(32'h390d3fcb),
	.w8(32'h39f791d2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924d2fd),
	.w1(32'hb9e39354),
	.w2(32'hba8839b2),
	.w3(32'h3a165142),
	.w4(32'hb9155fd8),
	.w5(32'hb9423119),
	.w6(32'h395f40bc),
	.w7(32'hb9b99274),
	.w8(32'h39cc5ada),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b72917),
	.w1(32'hb9ba454c),
	.w2(32'h38557fbd),
	.w3(32'h397958fd),
	.w4(32'hb781aa1c),
	.w5(32'hb93e0abf),
	.w6(32'hba38cf3e),
	.w7(32'hb9a5b3e3),
	.w8(32'hb9654d37),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939d019),
	.w1(32'hb9abab75),
	.w2(32'hba0775c6),
	.w3(32'hb882e237),
	.w4(32'h39a14a81),
	.w5(32'h39365041),
	.w6(32'hb907b881),
	.w7(32'hb97fe6a0),
	.w8(32'h368a9859),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912e02b),
	.w1(32'hb75d2ee7),
	.w2(32'hb982c848),
	.w3(32'h3a47c094),
	.w4(32'h39d8191b),
	.w5(32'h39a87de4),
	.w6(32'h39013d3e),
	.w7(32'h3839a952),
	.w8(32'h397b8f17),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90440f8),
	.w1(32'hb9bcc245),
	.w2(32'h3803cc8d),
	.w3(32'h39ed2fbc),
	.w4(32'hb88df626),
	.w5(32'h384ad8b8),
	.w6(32'hba100752),
	.w7(32'hba2e2c4a),
	.w8(32'hb9e36323),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d59c9),
	.w1(32'h3940d06f),
	.w2(32'h38e99672),
	.w3(32'hb7de3da6),
	.w4(32'h38c5b9e5),
	.w5(32'h3911036d),
	.w6(32'h374ba831),
	.w7(32'h3933e6e4),
	.w8(32'h3931c6cf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947f02d),
	.w1(32'h39e2c3b2),
	.w2(32'h3adc323d),
	.w3(32'h39905474),
	.w4(32'h399c3113),
	.w5(32'h37c01b4d),
	.w6(32'h3b013929),
	.w7(32'h3a25dd99),
	.w8(32'h3a0ec3ac),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a04a),
	.w1(32'h38a9ed51),
	.w2(32'hb9af940d),
	.w3(32'h397d7568),
	.w4(32'h3a8a81b3),
	.w5(32'h3a5f12c2),
	.w6(32'h39d3b210),
	.w7(32'h390cb347),
	.w8(32'h3a06e40f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390378c3),
	.w1(32'h386a05dc),
	.w2(32'hba90f1a9),
	.w3(32'h3a8c8de1),
	.w4(32'h38b876fd),
	.w5(32'hba6d6228),
	.w6(32'h38ff7ce7),
	.w7(32'hb8bd72e9),
	.w8(32'h388157b6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92fef1a),
	.w1(32'h3962aeec),
	.w2(32'h3ad1dc16),
	.w3(32'hb9ac24ef),
	.w4(32'hb9fdbd58),
	.w5(32'hba6262d1),
	.w6(32'h39fa3bbe),
	.w7(32'h3a125201),
	.w8(32'hbac6f40e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2c4a),
	.w1(32'hb8934ca6),
	.w2(32'hb967fe8b),
	.w3(32'hbb232320),
	.w4(32'h39e824f0),
	.w5(32'h38d6dcb0),
	.w6(32'h38a8884e),
	.w7(32'hb80aa3d1),
	.w8(32'hb9268288),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97faad8),
	.w1(32'h398d0813),
	.w2(32'hb85aa07a),
	.w3(32'h399169da),
	.w4(32'hb9c901e9),
	.w5(32'hba2e93b0),
	.w6(32'h39a083ae),
	.w7(32'h39fc7ffb),
	.w8(32'h39b7364a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d536cf),
	.w1(32'h3a27d053),
	.w2(32'h3a26f37a),
	.w3(32'hba461c13),
	.w4(32'h39c0331c),
	.w5(32'h3a120082),
	.w6(32'h39fda2aa),
	.w7(32'h3a4d45e6),
	.w8(32'h3a1df898),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fed4a),
	.w1(32'h38e6cf26),
	.w2(32'hb8e99045),
	.w3(32'h39d9775f),
	.w4(32'hb9524df2),
	.w5(32'hb985a799),
	.w6(32'h39a33367),
	.w7(32'hb8b20128),
	.w8(32'hb8ff6425),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c845a),
	.w1(32'h39b10a94),
	.w2(32'h38b03cab),
	.w3(32'hb9a8575d),
	.w4(32'h392cc2c1),
	.w5(32'hb919c807),
	.w6(32'hb819035b),
	.w7(32'h39e1dca3),
	.w8(32'h394bda19),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffbcc8),
	.w1(32'h3a4a09b8),
	.w2(32'h39a4f64b),
	.w3(32'hb891ad81),
	.w4(32'h3a50088a),
	.w5(32'h39d920cd),
	.w6(32'hb9d0307b),
	.w7(32'hb98dfdaa),
	.w8(32'h39fe6d0c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8d234),
	.w1(32'h39f61364),
	.w2(32'hb81347b2),
	.w3(32'hb94df932),
	.w4(32'h39973955),
	.w5(32'h38347c53),
	.w6(32'h39cffed7),
	.w7(32'h39f7ac16),
	.w8(32'h3788a849),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb740b525),
	.w1(32'h399c8dc0),
	.w2(32'h396b688e),
	.w3(32'hb8f885f2),
	.w4(32'hba159174),
	.w5(32'hba350041),
	.w6(32'h39a25d46),
	.w7(32'hb783257a),
	.w8(32'h39dcefdc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69ce62),
	.w1(32'h38d4c612),
	.w2(32'hb62e138f),
	.w3(32'hb931d409),
	.w4(32'h398f2590),
	.w5(32'h39202dbc),
	.w6(32'h388b5ccc),
	.w7(32'hb8879621),
	.w8(32'hb783c5bd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdc260),
	.w1(32'h39b454f0),
	.w2(32'h3a0d0878),
	.w3(32'h392ecb87),
	.w4(32'hb85d9a55),
	.w5(32'hb939faf7),
	.w6(32'h38d151c8),
	.w7(32'h390f872c),
	.w8(32'hb999898c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987fea5),
	.w1(32'hb91d8d3b),
	.w2(32'hb93131ec),
	.w3(32'hb949b29b),
	.w4(32'h3a031be3),
	.w5(32'h393f3894),
	.w6(32'hb8d48e58),
	.w7(32'hb945214c),
	.w8(32'hb91fa5eb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9856591),
	.w1(32'hb966549f),
	.w2(32'hb9b739fd),
	.w3(32'h39884a21),
	.w4(32'h397bec6c),
	.w5(32'h3988bb7a),
	.w6(32'hb948e927),
	.w7(32'hb9def5d6),
	.w8(32'hb9a84da0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955762f),
	.w1(32'h38e008e3),
	.w2(32'h3a141c71),
	.w3(32'h397e69c4),
	.w4(32'h39218c28),
	.w5(32'hb9360191),
	.w6(32'hba049f10),
	.w7(32'hb7b94ebc),
	.w8(32'hb9898d98),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4a82c),
	.w1(32'h397554d3),
	.w2(32'h39c377a9),
	.w3(32'hb9cbf4c2),
	.w4(32'h3994d0f3),
	.w5(32'h38e395bb),
	.w6(32'hb816383c),
	.w7(32'h39286aec),
	.w8(32'hb7913838),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f71d6),
	.w1(32'h39b0b5fd),
	.w2(32'h3a0753ca),
	.w3(32'h39606f7b),
	.w4(32'hb98d592b),
	.w5(32'hb98f5fb9),
	.w6(32'h3a2d4474),
	.w7(32'h3a801e23),
	.w8(32'h39e27a2c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e24cd),
	.w1(32'hba709c61),
	.w2(32'hba25ad68),
	.w3(32'hba1ec58d),
	.w4(32'hba2973e4),
	.w5(32'hba1ee343),
	.w6(32'hb91ddfbf),
	.w7(32'hb971ba86),
	.w8(32'h38bcbd15),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c5e4b),
	.w1(32'h38eac628),
	.w2(32'h3a8428d8),
	.w3(32'hb99bd0b6),
	.w4(32'hb94c6202),
	.w5(32'hba1bae5f),
	.w6(32'h37ba5a66),
	.w7(32'hb95f7f76),
	.w8(32'hb99117aa),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e6365),
	.w1(32'hb9f596ba),
	.w2(32'hba4d30e6),
	.w3(32'hb9c94631),
	.w4(32'hba05e40f),
	.w5(32'hbaa7f936),
	.w6(32'hba3061d5),
	.w7(32'hbaa33240),
	.w8(32'hbaf00b18),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadac1d6),
	.w1(32'hb97008de),
	.w2(32'hbb020809),
	.w3(32'hbb1a378a),
	.w4(32'h391f837f),
	.w5(32'hba7343a3),
	.w6(32'h38e61554),
	.w7(32'hbac486e6),
	.w8(32'h38aa47f5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf6e7c),
	.w1(32'hba16e8f7),
	.w2(32'hb98b8e4a),
	.w3(32'hb9837cf5),
	.w4(32'hba0ee2e8),
	.w5(32'hb9168732),
	.w6(32'hba06c03c),
	.w7(32'hb9383e0e),
	.w8(32'hb8ac90d3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97632c5),
	.w1(32'h3a3354bb),
	.w2(32'h38ecd068),
	.w3(32'hb9752e31),
	.w4(32'h3a041ca4),
	.w5(32'h398ce756),
	.w6(32'h39e1efc5),
	.w7(32'hb9321ce5),
	.w8(32'h3982c939),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4c6f4),
	.w1(32'hba7e1879),
	.w2(32'hbb0b2b61),
	.w3(32'h3a128720),
	.w4(32'hba896cc8),
	.w5(32'hbad4bcbc),
	.w6(32'hbaadc124),
	.w7(32'hba4a8976),
	.w8(32'hba8834de),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55e1ac),
	.w1(32'hba9fcabd),
	.w2(32'hb9078b5f),
	.w3(32'hba54462b),
	.w4(32'hba199056),
	.w5(32'hb944cc0b),
	.w6(32'hba7c2f17),
	.w7(32'hba9833b9),
	.w8(32'hbacaee6d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a970a),
	.w1(32'h391c738e),
	.w2(32'hb9e110f9),
	.w3(32'hb98a4704),
	.w4(32'h3ad31061),
	.w5(32'h3aa6d0f9),
	.w6(32'h3a2ee95c),
	.w7(32'h39923e25),
	.w8(32'h3a80b582),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927eb1b),
	.w1(32'h3883f192),
	.w2(32'hb9791a93),
	.w3(32'h3ad11c79),
	.w4(32'h3a19a74a),
	.w5(32'h398fd626),
	.w6(32'h3943736d),
	.w7(32'h390edd0c),
	.w8(32'h39927bb5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d260f3),
	.w1(32'h37b9204e),
	.w2(32'hb98db184),
	.w3(32'h3a3ec35c),
	.w4(32'h3a4c3df6),
	.w5(32'h3a258f77),
	.w6(32'h399d328e),
	.w7(32'h38325723),
	.w8(32'h39b2ca94),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881e10f),
	.w1(32'hb98f41f3),
	.w2(32'h39896295),
	.w3(32'h3a4edb00),
	.w4(32'h37eeb3f8),
	.w5(32'h39caf3b1),
	.w6(32'hb9664034),
	.w7(32'h390b465a),
	.w8(32'hb9bcd85d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01f62a),
	.w1(32'hba81e7fc),
	.w2(32'hba6bcb5f),
	.w3(32'hb8ac3907),
	.w4(32'hb8f0e4a9),
	.w5(32'hb9cd4c2b),
	.w6(32'hb931b504),
	.w7(32'hb7b9ae87),
	.w8(32'h394f17ab),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d09cb),
	.w1(32'h3945dc01),
	.w2(32'h3882407f),
	.w3(32'hb9eea13e),
	.w4(32'h3a1f72f8),
	.w5(32'h39d88c52),
	.w6(32'h37fb2806),
	.w7(32'hb9058b4a),
	.w8(32'hb900aae1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9629f),
	.w1(32'h37ead02e),
	.w2(32'hb98a5160),
	.w3(32'h3986783b),
	.w4(32'h3a527f6a),
	.w5(32'h3a2cec39),
	.w6(32'h39b2fe8d),
	.w7(32'h390b34eb),
	.w8(32'h39f32b83),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909355f),
	.w1(32'h39b3220a),
	.w2(32'hb9a9d384),
	.w3(32'h3a64acd1),
	.w4(32'h3a25e847),
	.w5(32'hb9f8cda2),
	.w6(32'h39986f3f),
	.w7(32'h396ec2c3),
	.w8(32'h39f1198e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a42a7),
	.w1(32'h396aceed),
	.w2(32'hb8b7db86),
	.w3(32'hb91dd739),
	.w4(32'h39d8dfd5),
	.w5(32'h3a0683eb),
	.w6(32'h39957f11),
	.w7(32'h396a5bf8),
	.w8(32'h39ee2dd4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857b9e9),
	.w1(32'h3aa1c250),
	.w2(32'hbadb2d87),
	.w3(32'h39ae8fed),
	.w4(32'h3a8096b9),
	.w5(32'hba7c130b),
	.w6(32'h3a8e414b),
	.w7(32'hb9b8b24d),
	.w8(32'h39c70b93),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866a3b0),
	.w1(32'h39aac12c),
	.w2(32'hb8552dae),
	.w3(32'h39aaf489),
	.w4(32'h39de76ef),
	.w5(32'h3a0c3a68),
	.w6(32'h3a000fc2),
	.w7(32'h398e3f3d),
	.w8(32'h39c77beb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936d053),
	.w1(32'hba37a3f1),
	.w2(32'hb9dc2e11),
	.w3(32'h3a306d16),
	.w4(32'h38da686c),
	.w5(32'hb80efc2a),
	.w6(32'h393fda03),
	.w7(32'h392df95a),
	.w8(32'h38abb4b0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a0b05),
	.w1(32'hba48ccba),
	.w2(32'hb92120e4),
	.w3(32'h3a06fdee),
	.w4(32'hb81d260a),
	.w5(32'h398e90d7),
	.w6(32'hba5afea2),
	.w7(32'hba0b99a6),
	.w8(32'h38729b38),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1be07),
	.w1(32'h388d99f5),
	.w2(32'hb9c69c17),
	.w3(32'h3955bb2e),
	.w4(32'h3a993016),
	.w5(32'h3a7558e7),
	.w6(32'h39f958af),
	.w7(32'h391dff87),
	.w8(32'h3a1aee86),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eaa7a7),
	.w1(32'hb8690eaa),
	.w2(32'hb9d1a561),
	.w3(32'h3a9d1d7e),
	.w4(32'h39e2cb0a),
	.w5(32'h399e6ad1),
	.w6(32'h3881ee1d),
	.w7(32'hb8e99c20),
	.w8(32'h38156f4a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b7fbc),
	.w1(32'hb710b8ce),
	.w2(32'hb9ce9c5e),
	.w3(32'h3a0d2e82),
	.w4(32'h3a1f3be1),
	.w5(32'h3a045281),
	.w6(32'h38f3809f),
	.w7(32'hb930a474),
	.w8(32'hb79f3819),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955e516),
	.w1(32'hba2b92f2),
	.w2(32'h3a18af81),
	.w3(32'h39fed7d2),
	.w4(32'h3a9336c8),
	.w5(32'h3ab567fc),
	.w6(32'h37dc1e77),
	.w7(32'hba41ac12),
	.w8(32'hba81dabe),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9905d50),
	.w1(32'hba33b97c),
	.w2(32'hba9f78c5),
	.w3(32'h3a6c0b5a),
	.w4(32'hba726762),
	.w5(32'hba68d5f9),
	.w6(32'hba55b2a1),
	.w7(32'hb932f74e),
	.w8(32'hba47e9e5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba448c94),
	.w1(32'hba028dc2),
	.w2(32'hba233e51),
	.w3(32'hb97f14e0),
	.w4(32'hb8a264d8),
	.w5(32'h392e8453),
	.w6(32'hba099bd2),
	.w7(32'hb9ed9e8d),
	.w8(32'hba4ee644),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35178e),
	.w1(32'hba0034cb),
	.w2(32'hba612dff),
	.w3(32'h39b4308c),
	.w4(32'hb99f275c),
	.w5(32'hb8e10e69),
	.w6(32'hba2329e4),
	.w7(32'hba3aca91),
	.w8(32'hba28ed77),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba837531),
	.w1(32'hb88f557d),
	.w2(32'hb990d2c2),
	.w3(32'hb9ce3259),
	.w4(32'h3a09c442),
	.w5(32'h3a1c6cf5),
	.w6(32'h390e6cf1),
	.w7(32'h38ed7b01),
	.w8(32'h3991a1ae),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7467991),
	.w1(32'hba2f283e),
	.w2(32'h3ae4a21a),
	.w3(32'h3a3f8e1e),
	.w4(32'hb9c8684c),
	.w5(32'hbaa94e7c),
	.w6(32'hba45fad6),
	.w7(32'hba7c0950),
	.w8(32'hbadc20e8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f533c),
	.w1(32'h3a376184),
	.w2(32'h3a237d43),
	.w3(32'hbab21ef5),
	.w4(32'h3a9c09c7),
	.w5(32'h3a14c58a),
	.w6(32'h3a0927fe),
	.w7(32'hba052475),
	.w8(32'hb80367a9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f8e39),
	.w1(32'hb890fe5d),
	.w2(32'h37556c2c),
	.w3(32'h3a965faa),
	.w4(32'h3985ac4d),
	.w5(32'h39518fa3),
	.w6(32'hb8c0a664),
	.w7(32'hb94aed04),
	.w8(32'hb9846cb5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979f6aa),
	.w1(32'hb840da37),
	.w2(32'hb89045bb),
	.w3(32'h3957471c),
	.w4(32'hb9094b36),
	.w5(32'hb8435567),
	.w6(32'h3822af54),
	.w7(32'hb836ca37),
	.w8(32'hb82d883c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb830c64c),
	.w1(32'h39045643),
	.w2(32'hb7f9f7a3),
	.w3(32'h38473aef),
	.w4(32'h391ff562),
	.w5(32'h37c1b904),
	.w6(32'h397d7110),
	.w7(32'h38b7a261),
	.w8(32'h390b2888),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule