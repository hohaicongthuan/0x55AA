module layer_10_featuremap_250(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc8f6e),
	.w1(32'h392f12c6),
	.w2(32'hb93c9bef),
	.w3(32'h38b305d6),
	.w4(32'h38c22c82),
	.w5(32'h3a895cdf),
	.w6(32'hba8e74e6),
	.w7(32'hba494577),
	.w8(32'hba56d3d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62fa5d),
	.w1(32'hbb2ada87),
	.w2(32'hba5a5f44),
	.w3(32'h3a0f330d),
	.w4(32'hba98a7c7),
	.w5(32'hba9799d9),
	.w6(32'hbad6c82b),
	.w7(32'hbb0d1f18),
	.w8(32'hbaf22b90),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a178f92),
	.w1(32'h3a8770a9),
	.w2(32'h39f27e60),
	.w3(32'hbb17b60d),
	.w4(32'hbaf53fe7),
	.w5(32'hbaa9812d),
	.w6(32'hbb4c630c),
	.w7(32'hba90334b),
	.w8(32'hba867f2b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6dcc4),
	.w1(32'hb9dc05e0),
	.w2(32'hba063b8b),
	.w3(32'h39044c42),
	.w4(32'hb9c40088),
	.w5(32'hbb1f2910),
	.w6(32'h3ada90e3),
	.w7(32'h39236125),
	.w8(32'hbb6946c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad34d2),
	.w1(32'hbaa268a0),
	.w2(32'hbb2bc3ef),
	.w3(32'hbb5e4fed),
	.w4(32'hba7c2fdb),
	.w5(32'hba121fe1),
	.w6(32'hbab05555),
	.w7(32'hbb8a50de),
	.w8(32'h38101e22),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1ef6a),
	.w1(32'hba0ab366),
	.w2(32'h38683113),
	.w3(32'hb8ac4a89),
	.w4(32'hb8dec42f),
	.w5(32'hbaa66ef0),
	.w6(32'h3a1d4097),
	.w7(32'h3a38d5ba),
	.w8(32'hba5b1a5f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8fe18),
	.w1(32'h3973de64),
	.w2(32'hbb807840),
	.w3(32'h3a305208),
	.w4(32'hb99d455b),
	.w5(32'hbb89c4e8),
	.w6(32'h3b3aee6e),
	.w7(32'h3a5eeffe),
	.w8(32'hbae9f3f8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a023a),
	.w1(32'hbba2acc6),
	.w2(32'hbbae0ff5),
	.w3(32'hbb5c4872),
	.w4(32'hbb7d0403),
	.w5(32'hbb4a732c),
	.w6(32'hba60e50f),
	.w7(32'hbb90b179),
	.w8(32'hbb3fa553),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f260b),
	.w1(32'hba4d4ab4),
	.w2(32'hbab222b8),
	.w3(32'h394d6c37),
	.w4(32'hba2700b1),
	.w5(32'h3a637109),
	.w6(32'h390a4092),
	.w7(32'hba1d93b9),
	.w8(32'h3a3ce069),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b3163),
	.w1(32'hb8d14452),
	.w2(32'h3817eb3c),
	.w3(32'hbb1e46bf),
	.w4(32'h3a16270b),
	.w5(32'hb9de83d4),
	.w6(32'hbae6b6e4),
	.w7(32'h3a400753),
	.w8(32'hb9ae0d85),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9386b3),
	.w1(32'hb667f5fe),
	.w2(32'hba1e9aa4),
	.w3(32'h3a6d555b),
	.w4(32'h379bad9f),
	.w5(32'hbaa3af79),
	.w6(32'h3b1df8c6),
	.w7(32'h3a9d1ce1),
	.w8(32'hb9a2c47d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03fa38),
	.w1(32'h3ab24b65),
	.w2(32'hbabbae74),
	.w3(32'hba150968),
	.w4(32'h3a385fdd),
	.w5(32'h3b801865),
	.w6(32'hbad44fe7),
	.w7(32'h39c97e90),
	.w8(32'h3b65540f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3b1cf),
	.w1(32'h3ae85df3),
	.w2(32'h3aa67dcc),
	.w3(32'h38b250e1),
	.w4(32'h3b0ddf45),
	.w5(32'hb94b5af1),
	.w6(32'hba214a29),
	.w7(32'h3b1d8495),
	.w8(32'hba854617),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97664),
	.w1(32'hbaf9a1a2),
	.w2(32'hba16c829),
	.w3(32'h39cd16e5),
	.w4(32'h3a8f2464),
	.w5(32'hbb3a96ec),
	.w6(32'hbaae1c92),
	.w7(32'h3a9bbe8c),
	.w8(32'hbaaff0f5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15e3b2),
	.w1(32'hb87ae67e),
	.w2(32'h3a04f673),
	.w3(32'hba3db775),
	.w4(32'hba4d6bcd),
	.w5(32'h3a376890),
	.w6(32'hb8a9c121),
	.w7(32'hba0a208c),
	.w8(32'hba8c5f5f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947dbde),
	.w1(32'h389f9215),
	.w2(32'hba05bae3),
	.w3(32'hbadb3ee9),
	.w4(32'h3ad0072d),
	.w5(32'hba2bf938),
	.w6(32'hbb7bd87d),
	.w7(32'hbb114898),
	.w8(32'hbb334505),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d36f31),
	.w1(32'hb9e86e8a),
	.w2(32'hba9664ea),
	.w3(32'h3a02f99e),
	.w4(32'hb8f4f63b),
	.w5(32'h3b2935dc),
	.w6(32'hb91ca5ad),
	.w7(32'h398f6a30),
	.w8(32'h3b0d110b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1925ff),
	.w1(32'h3a1f8905),
	.w2(32'hba169904),
	.w3(32'hba8c01b7),
	.w4(32'hbaa976a9),
	.w5(32'hbb8a61df),
	.w6(32'h39f674f3),
	.w7(32'h3a1a65e5),
	.w8(32'hbabb91e2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab46bf1),
	.w1(32'h3b24d9ed),
	.w2(32'h3a2833fc),
	.w3(32'hba2ce281),
	.w4(32'h3a960c6a),
	.w5(32'h3a30cf2f),
	.w6(32'h3a909eb9),
	.w7(32'h3aa1f557),
	.w8(32'hbac94dbd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a4514),
	.w1(32'h3943f3ca),
	.w2(32'h3ac09418),
	.w3(32'h3a8aca95),
	.w4(32'h39b6e308),
	.w5(32'h3ae582a0),
	.w6(32'h3aa72e98),
	.w7(32'h3aa964b1),
	.w8(32'h3a57a2c9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b507a),
	.w1(32'h3a024f40),
	.w2(32'h3af6faf4),
	.w3(32'hb9125baa),
	.w4(32'h3b37e74f),
	.w5(32'h3a264738),
	.w6(32'h3b0e3541),
	.w7(32'h3afdf356),
	.w8(32'h3a8695dc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffee4d),
	.w1(32'h3a402278),
	.w2(32'hb79e5e90),
	.w3(32'h3ab4cfa7),
	.w4(32'h3a872afd),
	.w5(32'hba93a803),
	.w6(32'h3b055ebd),
	.w7(32'h3a9980b2),
	.w8(32'hbabc8b6f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ce5b),
	.w1(32'hb9a74647),
	.w2(32'hbb5ce483),
	.w3(32'hbb0efa8f),
	.w4(32'hbb049e79),
	.w5(32'hbb96a49f),
	.w6(32'hbb811ce6),
	.w7(32'hba837ce6),
	.w8(32'hbbd6435a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccb48a),
	.w1(32'hbabd979a),
	.w2(32'hba78e6fe),
	.w3(32'hbac97677),
	.w4(32'h39df63b0),
	.w5(32'hba2e4d05),
	.w6(32'hbb7e7be4),
	.w7(32'hbabd55c5),
	.w8(32'hbaf2a5a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e26de),
	.w1(32'hba057da2),
	.w2(32'h3a59921e),
	.w3(32'hbb1c473e),
	.w4(32'h3a89b06f),
	.w5(32'h3add6a9f),
	.w6(32'hbb9b803f),
	.w7(32'hbabaa5c8),
	.w8(32'h3a8fcde1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04289e),
	.w1(32'h3a97f3cd),
	.w2(32'h3a7a366a),
	.w3(32'h3a6abeb0),
	.w4(32'h3aa7260c),
	.w5(32'hba27ebb8),
	.w6(32'h3a9c2746),
	.w7(32'h3ab21048),
	.w8(32'h36c4912b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901f846),
	.w1(32'hbaf6934f),
	.w2(32'hba660cb6),
	.w3(32'hb99046bf),
	.w4(32'h39a63c49),
	.w5(32'hb9128843),
	.w6(32'hb93a560e),
	.w7(32'hba35e593),
	.w8(32'hba515159),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5214f7),
	.w1(32'hba2ac5fc),
	.w2(32'h3af85616),
	.w3(32'hbb518fae),
	.w4(32'hbaa1f181),
	.w5(32'h3ac39e5a),
	.w6(32'hbb83e3cb),
	.w7(32'hbb45a891),
	.w8(32'h3b248872),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab18851),
	.w1(32'h3ae5db6d),
	.w2(32'h3b089689),
	.w3(32'h3ac1f203),
	.w4(32'h3b35efd3),
	.w5(32'h3b120ae3),
	.w6(32'h3abc4aa6),
	.w7(32'h3b0b2e6c),
	.w8(32'hba4b6484),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27839c),
	.w1(32'h3aaa9676),
	.w2(32'h3b1fc083),
	.w3(32'h3ab8b92e),
	.w4(32'h3ad40214),
	.w5(32'hbaa8205a),
	.w6(32'hbb0d8393),
	.w7(32'h3abcb3ec),
	.w8(32'hbb4ca07b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ddbe5),
	.w1(32'hbb074de9),
	.w2(32'hbaff66ee),
	.w3(32'hbb0f9e68),
	.w4(32'hbb0f6528),
	.w5(32'h38631794),
	.w6(32'hbb69a461),
	.w7(32'hbb0fa2b3),
	.w8(32'h39dc2e0f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb7f60),
	.w1(32'h3b1df07c),
	.w2(32'h3ae22214),
	.w3(32'hba8b5e45),
	.w4(32'hbaa00f3d),
	.w5(32'hbb815be1),
	.w6(32'h3b4ec890),
	.w7(32'hb8e5884d),
	.w8(32'hbb18fbd0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9bcbe),
	.w1(32'h3a2b0335),
	.w2(32'hb8e4762e),
	.w3(32'hba9edf25),
	.w4(32'h39b65566),
	.w5(32'h3a908c4b),
	.w6(32'hbb13370d),
	.w7(32'hbae63558),
	.w8(32'h3a73cf52),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cc7a6),
	.w1(32'h3af03e62),
	.w2(32'h3b88a3f1),
	.w3(32'h3b5e0394),
	.w4(32'h3aadebfc),
	.w5(32'hba50bf8e),
	.w6(32'hba62fcc4),
	.w7(32'h3b12cbbf),
	.w8(32'hbaceb585),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dfcd5),
	.w1(32'h3a2b8676),
	.w2(32'h3a7c10bb),
	.w3(32'hba45a47f),
	.w4(32'hb9db8ac3),
	.w5(32'h3b43d396),
	.w6(32'hbad15ad7),
	.w7(32'hb9b1a45f),
	.w8(32'h3a244a94),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933d387),
	.w1(32'h3af4232e),
	.w2(32'hba0c1548),
	.w3(32'hba44d8fc),
	.w4(32'h3964cc4d),
	.w5(32'hbaf3e76b),
	.w6(32'h3a1cc381),
	.w7(32'h3b088c14),
	.w8(32'hbb006c9f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba505bc3),
	.w1(32'hba647a16),
	.w2(32'h3ae5ead9),
	.w3(32'hb9ac9e24),
	.w4(32'h3b97a1ec),
	.w5(32'h3b35a8a5),
	.w6(32'hbb034510),
	.w7(32'h3a43548d),
	.w8(32'h3b919ec5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec6a4),
	.w1(32'hba258ce7),
	.w2(32'h3b15c21f),
	.w3(32'hbaf4a6d8),
	.w4(32'h3b20f20c),
	.w5(32'h3b9e60ce),
	.w6(32'hbabc4c0a),
	.w7(32'hb9eabbc8),
	.w8(32'h3a74dca7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35081),
	.w1(32'h392b54cf),
	.w2(32'h3b930490),
	.w3(32'h3b8beb25),
	.w4(32'h3a7c219a),
	.w5(32'h3ad4a254),
	.w6(32'h3baad028),
	.w7(32'h3ab366e4),
	.w8(32'h3ac2797c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63c28),
	.w1(32'hba2a7431),
	.w2(32'hbaeda338),
	.w3(32'hbb181dac),
	.w4(32'hb9ee8ee0),
	.w5(32'h3b0c84aa),
	.w6(32'hbacf6b20),
	.w7(32'hbafad8e2),
	.w8(32'h3b1e0742),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb75e1),
	.w1(32'h3a8538a9),
	.w2(32'hb91a4237),
	.w3(32'h3a871cbc),
	.w4(32'h3acf137b),
	.w5(32'h3a44bd24),
	.w6(32'h3a294824),
	.w7(32'h3aa34b8c),
	.w8(32'h3aa8f177),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae17073),
	.w1(32'h3aa74d10),
	.w2(32'h3a08448d),
	.w3(32'h3b0468d9),
	.w4(32'h3b08563b),
	.w5(32'h3aec725b),
	.w6(32'h3b30a135),
	.w7(32'h3b098a87),
	.w8(32'h3aec455a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a795),
	.w1(32'h3a664a66),
	.w2(32'h3b1b6dba),
	.w3(32'h3a2ef783),
	.w4(32'h3ad31782),
	.w5(32'hb90ede40),
	.w6(32'h3ace18c4),
	.w7(32'h3b2838ef),
	.w8(32'hb9ee0a7d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae397c6),
	.w1(32'hba620163),
	.w2(32'hbb4add4e),
	.w3(32'hbb1c8dd1),
	.w4(32'hbb596589),
	.w5(32'hbb7ace21),
	.w6(32'hba704bd0),
	.w7(32'hba50a498),
	.w8(32'hbb251557),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba256d64),
	.w1(32'h39c57e2f),
	.w2(32'hba9b36a1),
	.w3(32'hbb8f90aa),
	.w4(32'h3a116c00),
	.w5(32'h3b01ce29),
	.w6(32'hbb737ee9),
	.w7(32'hbb4168ad),
	.w8(32'h3a075d95),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad131a0),
	.w1(32'h382da969),
	.w2(32'hb93b7a75),
	.w3(32'hb9e76827),
	.w4(32'h3b72b80f),
	.w5(32'h3aefe5b6),
	.w6(32'hbb49b10b),
	.w7(32'h3a46f39c),
	.w8(32'h39d1eed1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd5d30),
	.w1(32'h3aa481a6),
	.w2(32'h3ab4dd98),
	.w3(32'hbafb7f27),
	.w4(32'h3a52eb8f),
	.w5(32'h3a52a7c7),
	.w6(32'hbb645dfc),
	.w7(32'hba1df59e),
	.w8(32'hbacdecbe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39873439),
	.w1(32'h3a3f9e63),
	.w2(32'hbb1791b1),
	.w3(32'hbaa66755),
	.w4(32'h39fcdca1),
	.w5(32'h3ae825eb),
	.w6(32'hbac43506),
	.w7(32'h39a6c1e9),
	.w8(32'h3b053357),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c35a3),
	.w1(32'h3af8bc46),
	.w2(32'h3a201a5d),
	.w3(32'h3b4bb023),
	.w4(32'hba4eed28),
	.w5(32'h39f4ed80),
	.w6(32'h3b1264e1),
	.w7(32'hb9f0828f),
	.w8(32'h3a1160f0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eaa6a),
	.w1(32'h3ab7c6c1),
	.w2(32'h3aec41a0),
	.w3(32'h3aa6d73a),
	.w4(32'h3acdb069),
	.w5(32'hbb31a4a9),
	.w6(32'h3a8a0988),
	.w7(32'h3ab2423d),
	.w8(32'hbb32baf1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9e0f9),
	.w1(32'h3a18c4fb),
	.w2(32'h390c8dbb),
	.w3(32'hbab1944d),
	.w4(32'h393f01f3),
	.w5(32'h3a1edb6f),
	.w6(32'hbb3373eb),
	.w7(32'hba8a5d9f),
	.w8(32'h3afbdabc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbce80),
	.w1(32'hbb0e87a6),
	.w2(32'hbb6791b1),
	.w3(32'hba1ff4fd),
	.w4(32'hbaac3ea9),
	.w5(32'hba9fc780),
	.w6(32'h39983c03),
	.w7(32'hb9ae75ca),
	.w8(32'hbad80703),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ec9b0),
	.w1(32'hbb2d3c63),
	.w2(32'hbb4030ca),
	.w3(32'hba7f49d3),
	.w4(32'hbb24a42d),
	.w5(32'h37d35204),
	.w6(32'hbb49175b),
	.w7(32'hbb588e0c),
	.w8(32'hb904d888),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe529),
	.w1(32'hbaa0b32b),
	.w2(32'hbb81988f),
	.w3(32'hbb1940dc),
	.w4(32'h3aa70c6d),
	.w5(32'hbb00c73c),
	.w6(32'hba449a6e),
	.w7(32'h391e1d12),
	.w8(32'hbb05e7ea),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a1f27),
	.w1(32'h3a2bdb9a),
	.w2(32'h3aad0f9a),
	.w3(32'h395083b9),
	.w4(32'hba80d072),
	.w5(32'hbb1b040a),
	.w6(32'h3b588154),
	.w7(32'h3984d0e4),
	.w8(32'hbb4c7121),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a845),
	.w1(32'hba04b8c0),
	.w2(32'hbae73856),
	.w3(32'hbab41fbc),
	.w4(32'hb9e897dd),
	.w5(32'hbaa5f664),
	.w6(32'hbb2e37f7),
	.w7(32'hbb0d8219),
	.w8(32'hb9deebda),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda92d),
	.w1(32'hba951189),
	.w2(32'hbab74fa0),
	.w3(32'hbad2084e),
	.w4(32'hb9a0a242),
	.w5(32'hba972894),
	.w6(32'hba11399b),
	.w7(32'hb9e58863),
	.w8(32'hbb07b190),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa61373),
	.w1(32'hb727ee20),
	.w2(32'h3a31d939),
	.w3(32'h39741610),
	.w4(32'hba94a841),
	.w5(32'h39a6f8b5),
	.w6(32'h3a76a6c4),
	.w7(32'hba106641),
	.w8(32'h39f4d542),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4ee6),
	.w1(32'h3a625e38),
	.w2(32'h399cc767),
	.w3(32'h3a6d819d),
	.w4(32'h3a0560dd),
	.w5(32'hbaa02860),
	.w6(32'h3a883614),
	.w7(32'h39fd4ca4),
	.w8(32'hba15595a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89b715),
	.w1(32'hba4b507d),
	.w2(32'hbb683aec),
	.w3(32'hba842e2c),
	.w4(32'hbb6bdde8),
	.w5(32'hb92df5f8),
	.w6(32'hba8ab8e4),
	.w7(32'hbb9bb702),
	.w8(32'hba1ab66d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d839b4),
	.w1(32'hb9b4d384),
	.w2(32'h3a8e1540),
	.w3(32'h3a32a3f1),
	.w4(32'hba802bf3),
	.w5(32'hbb0f0528),
	.w6(32'h3ade2ec7),
	.w7(32'h3aa638c2),
	.w8(32'hbaef994b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d83b),
	.w1(32'hb9d72f4a),
	.w2(32'h37fb11be),
	.w3(32'hbae8cb80),
	.w4(32'hb9f17f5c),
	.w5(32'hbb032b8a),
	.w6(32'h39bfe667),
	.w7(32'hba1feb4a),
	.w8(32'hbb37eb43),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77de6e4),
	.w1(32'h3ac3a7ce),
	.w2(32'h3ad588ef),
	.w3(32'hba9fccd8),
	.w4(32'hb848fad1),
	.w5(32'h399b275a),
	.w6(32'hbaa2b546),
	.w7(32'hba4de1c3),
	.w8(32'h39f2b5c0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9955f1b),
	.w1(32'h39a9c59a),
	.w2(32'h3a212bd9),
	.w3(32'hba808655),
	.w4(32'h3a7613c3),
	.w5(32'h3ab5cffe),
	.w6(32'hba0e2424),
	.w7(32'h3a45395f),
	.w8(32'h3976eef9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3fd3e),
	.w1(32'h3a95023e),
	.w2(32'h3b28fabe),
	.w3(32'h3a8afbec),
	.w4(32'h3ad50650),
	.w5(32'hb6171664),
	.w6(32'h3aa0aef0),
	.w7(32'h3b0ecb6b),
	.w8(32'h3ae06e39),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872c4d4),
	.w1(32'hba93bd3b),
	.w2(32'hba63dff5),
	.w3(32'hbb3cf19d),
	.w4(32'hbb28e6a7),
	.w5(32'hbab96888),
	.w6(32'h375c6da2),
	.w7(32'hba8ae31d),
	.w8(32'h3a0d6d19),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b656d5c),
	.w1(32'h3acad12d),
	.w2(32'hba6a99db),
	.w3(32'h399f9982),
	.w4(32'hbb25b10b),
	.w5(32'hbb97c4cf),
	.w6(32'hbb0d26cd),
	.w7(32'hbbb5bdfa),
	.w8(32'hbbd4f6e8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e903),
	.w1(32'hbb6ba9b1),
	.w2(32'hbc0b07c2),
	.w3(32'h3b153e7e),
	.w4(32'h3a698b12),
	.w5(32'hbb71a41e),
	.w6(32'hba28c625),
	.w7(32'hbb973f47),
	.w8(32'hbbb4ee9a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9b1b),
	.w1(32'hbb02b916),
	.w2(32'hba4e6912),
	.w3(32'hbafec404),
	.w4(32'h3a8364c2),
	.w5(32'h3b033e82),
	.w6(32'h3a6823b5),
	.w7(32'h380d4168),
	.w8(32'h39c20b5d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1706),
	.w1(32'h372f165b),
	.w2(32'hb9d9f5e1),
	.w3(32'h3b3ac3ee),
	.w4(32'h3abfcb94),
	.w5(32'h3ad96fba),
	.w6(32'h3a9af30a),
	.w7(32'hbabbf02e),
	.w8(32'h3a58131b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852fee),
	.w1(32'hba1ae342),
	.w2(32'hba575c5b),
	.w3(32'hb73c76c5),
	.w4(32'h39ee187d),
	.w5(32'h3a7d391e),
	.w6(32'h39f4af74),
	.w7(32'h38f54d61),
	.w8(32'h3a4536ae),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6f0fa),
	.w1(32'h39f2c43f),
	.w2(32'hba647ab0),
	.w3(32'hba7449a3),
	.w4(32'h3a67426c),
	.w5(32'hb9aa19ed),
	.w6(32'hbac844c0),
	.w7(32'hb8b5aa69),
	.w8(32'h3b0619f5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44f5ee),
	.w1(32'h3a609ca1),
	.w2(32'h3aa41094),
	.w3(32'hba6a9fcf),
	.w4(32'h3a214822),
	.w5(32'h3bc5e958),
	.w6(32'h3b3dbcf9),
	.w7(32'h3b2ef95a),
	.w8(32'h3ba631c5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99a02e),
	.w1(32'h3b51dc03),
	.w2(32'h3b84e883),
	.w3(32'h3bbd9c14),
	.w4(32'h3add8a74),
	.w5(32'hba04c021),
	.w6(32'h3bb7a62c),
	.w7(32'h3b89063b),
	.w8(32'hb9e34d69),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d135d),
	.w1(32'hba78a317),
	.w2(32'hba3422e7),
	.w3(32'hb796f14a),
	.w4(32'h3994c9a6),
	.w5(32'h3bac3d02),
	.w6(32'h39697a73),
	.w7(32'hb93e38c0),
	.w8(32'h3b8fd41f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e46b),
	.w1(32'h3b35d24d),
	.w2(32'h3b36128c),
	.w3(32'h3b18b684),
	.w4(32'h3aed4b0a),
	.w5(32'hbb0d8f66),
	.w6(32'h3ad41e98),
	.w7(32'h3b06ba2d),
	.w8(32'hbac0012a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ce374),
	.w1(32'hbb57a186),
	.w2(32'hbb8728cf),
	.w3(32'hbb76ebea),
	.w4(32'hbafab00f),
	.w5(32'hbb0a7e80),
	.w6(32'hbb9762b7),
	.w7(32'hbb0792be),
	.w8(32'hbaf0131c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7084ab),
	.w1(32'hba96732e),
	.w2(32'hba3584e4),
	.w3(32'hbb84e57f),
	.w4(32'h3abec535),
	.w5(32'h3bb56aae),
	.w6(32'hbb9db68f),
	.w7(32'h3a237e6f),
	.w8(32'h3be72df8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b467307),
	.w1(32'h3b24b6b3),
	.w2(32'hba948b79),
	.w3(32'h3a0a01ee),
	.w4(32'hb998995c),
	.w5(32'hbb700c72),
	.w6(32'h3a8b5199),
	.w7(32'hb98c248b),
	.w8(32'hbb7d5a55),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a103d18),
	.w1(32'hba2030f7),
	.w2(32'hbae1eca2),
	.w3(32'hba95d1d2),
	.w4(32'hbad71011),
	.w5(32'h3b688a07),
	.w6(32'hbb136c85),
	.w7(32'hbb2d1b8e),
	.w8(32'h3b923dc2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b049bfb),
	.w1(32'h3b411b42),
	.w2(32'h3abca37b),
	.w3(32'h3ae4e66f),
	.w4(32'hba8bd96b),
	.w5(32'h3bbe5ef2),
	.w6(32'h3b74fd77),
	.w7(32'hba606ded),
	.w8(32'h3bc1c36f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8600b7),
	.w1(32'h3b686000),
	.w2(32'h3ac66a0c),
	.w3(32'h3b42e1d5),
	.w4(32'h3b5e057e),
	.w5(32'hbaea8a31),
	.w6(32'h3b1f9dd9),
	.w7(32'h3b641db5),
	.w8(32'hba9a886e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904c8c4),
	.w1(32'h3a273f92),
	.w2(32'h3a88dd22),
	.w3(32'hbaa86eb5),
	.w4(32'hba41084f),
	.w5(32'hbb383947),
	.w6(32'hbae653de),
	.w7(32'h398d2ebc),
	.w8(32'hbb3e116e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf2d05),
	.w1(32'hba878636),
	.w2(32'hb7a022a8),
	.w3(32'hbb16e11a),
	.w4(32'hba11d190),
	.w5(32'h3a4e3d41),
	.w6(32'hbaa5a877),
	.w7(32'hbac63373),
	.w8(32'hba9aed9e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43cbdc),
	.w1(32'h3998a50d),
	.w2(32'hb95a9ca8),
	.w3(32'hba11685e),
	.w4(32'hb8db19b7),
	.w5(32'hbacaa8a0),
	.w6(32'hbaf5ff16),
	.w7(32'hba33cdab),
	.w8(32'h3a0cd99a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982a98a),
	.w1(32'hba485168),
	.w2(32'hb8ecff19),
	.w3(32'hbab77451),
	.w4(32'hb9f3c8d9),
	.w5(32'hba9535c4),
	.w6(32'hb8bbb479),
	.w7(32'h3a201913),
	.w8(32'hbaef417f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5cc1b),
	.w1(32'hbad4fa99),
	.w2(32'hba61be8b),
	.w3(32'hba5e698c),
	.w4(32'h398c051d),
	.w5(32'h39b714f2),
	.w6(32'hbab1c5a1),
	.w7(32'hbb13f292),
	.w8(32'hba9f4a76),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9711dd),
	.w1(32'hba9e5f97),
	.w2(32'hba266128),
	.w3(32'hb96c8380),
	.w4(32'h39843eb6),
	.w5(32'hba972a35),
	.w6(32'hba917a43),
	.w7(32'hba75e146),
	.w8(32'hb9d3e514),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac74bb3),
	.w1(32'hbb1d87fe),
	.w2(32'hbb329306),
	.w3(32'hba9ab3f7),
	.w4(32'hbabe9e08),
	.w5(32'h3b715ebc),
	.w6(32'hbb12ed1b),
	.w7(32'hbae85862),
	.w8(32'hba3cb3f9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e10b3),
	.w1(32'h3ac35eff),
	.w2(32'hb9c459b3),
	.w3(32'h39ea1a72),
	.w4(32'hbb142a2b),
	.w5(32'hbb1544b9),
	.w6(32'hb98bd122),
	.w7(32'hbac37cde),
	.w8(32'hbafa241f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9ccff),
	.w1(32'h3b4bc4e9),
	.w2(32'h3b98c7de),
	.w3(32'h3b0e0b75),
	.w4(32'h3b40c7e6),
	.w5(32'h3a9286c3),
	.w6(32'h3b0f5108),
	.w7(32'h3b2d078b),
	.w8(32'hbaa3ec78),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990d265),
	.w1(32'h39aa25e9),
	.w2(32'hbab720cf),
	.w3(32'h3af88a1a),
	.w4(32'h3b01d93a),
	.w5(32'hbbdbfb99),
	.w6(32'hba7c87fd),
	.w7(32'h3b19f7f8),
	.w8(32'hbc136126),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb14b),
	.w1(32'hbb553086),
	.w2(32'hba940453),
	.w3(32'hbaa28a80),
	.w4(32'h3b20f255),
	.w5(32'h3a602f61),
	.w6(32'hbafbf918),
	.w7(32'h3a1bb413),
	.w8(32'hba30ef1a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7031e3),
	.w1(32'hbb9330eb),
	.w2(32'hbb98a48d),
	.w3(32'hba259b25),
	.w4(32'hbb648ca2),
	.w5(32'hbb0d5d83),
	.w6(32'hbb2b0613),
	.w7(32'hbba60ff8),
	.w8(32'hbb982758),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44dc2d),
	.w1(32'h3af6e2b3),
	.w2(32'h3b1fed57),
	.w3(32'h3b542433),
	.w4(32'h3b7dd2e7),
	.w5(32'h3b07a72d),
	.w6(32'h3a3ca8e0),
	.w7(32'h3a05d3c7),
	.w8(32'h3948f824),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44667b),
	.w1(32'hbb132be7),
	.w2(32'hbb043eff),
	.w3(32'hb9534eea),
	.w4(32'h39b06085),
	.w5(32'h3bda1854),
	.w6(32'hbacd2ad5),
	.w7(32'hbb2cb780),
	.w8(32'h3bb49461),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b541fb9),
	.w1(32'h3b5e0fc0),
	.w2(32'h385ecd03),
	.w3(32'h3b05ae63),
	.w4(32'h3ade43f2),
	.w5(32'hbb3892d5),
	.w6(32'h3b58cf17),
	.w7(32'hba8ac658),
	.w8(32'hb9b7c622),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998c6c4),
	.w1(32'h3af62cb9),
	.w2(32'hbb00f813),
	.w3(32'hba9dfd56),
	.w4(32'hbabc30d0),
	.w5(32'hbbc09087),
	.w6(32'hbb189a93),
	.w7(32'hbaf75615),
	.w8(32'hbbbad642),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d170d),
	.w1(32'hbb39ce22),
	.w2(32'hb92b75c9),
	.w3(32'hbb84a710),
	.w4(32'hbb62ad9e),
	.w5(32'h3b6c62c8),
	.w6(32'hbb84ab70),
	.w7(32'hbb8dac70),
	.w8(32'hbaf3072e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ac881),
	.w1(32'h3a9fcf4e),
	.w2(32'hba5012dc),
	.w3(32'hbc141096),
	.w4(32'h3b1eba97),
	.w5(32'h3b12d2c8),
	.w6(32'h3b4cf88e),
	.w7(32'h3bba20f2),
	.w8(32'h3bea9e02),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4668b0),
	.w1(32'hbc33b8ba),
	.w2(32'hbb96ffa2),
	.w3(32'h3a3130c1),
	.w4(32'h3bb3bb4f),
	.w5(32'h3c15260a),
	.w6(32'hbbfd810f),
	.w7(32'h3be4c2a8),
	.w8(32'hbb2edef7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00c090),
	.w1(32'hbbfa6687),
	.w2(32'hbbaa881f),
	.w3(32'h38b0733e),
	.w4(32'hbb31e830),
	.w5(32'h3a1d758f),
	.w6(32'hbbbcda11),
	.w7(32'hbbc796de),
	.w8(32'hb9635572),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a49d3),
	.w1(32'hbc03f1df),
	.w2(32'h3b12129a),
	.w3(32'hbbd8796c),
	.w4(32'h392b382d),
	.w5(32'h3c40eb4d),
	.w6(32'hbbfbea05),
	.w7(32'h39988ded),
	.w8(32'h3c2648a4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be64fc0),
	.w1(32'h3b2fb261),
	.w2(32'h3c469d1f),
	.w3(32'h3c04a003),
	.w4(32'h3c39c61d),
	.w5(32'hbb925deb),
	.w6(32'hbc4d7942),
	.w7(32'h3c2b9982),
	.w8(32'h3be364a4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1febed),
	.w1(32'hbc25d785),
	.w2(32'hbc0485dd),
	.w3(32'hbc0ff3f4),
	.w4(32'hbc24dc58),
	.w5(32'h3bb937b2),
	.w6(32'h3c5e0eaf),
	.w7(32'h3a9dbbd0),
	.w8(32'h3aa336c8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407709),
	.w1(32'h3c150724),
	.w2(32'h3b8b2b20),
	.w3(32'hbba62d01),
	.w4(32'h3a2f7382),
	.w5(32'hbc0269cf),
	.w6(32'h3bb34008),
	.w7(32'h3b7ef4f4),
	.w8(32'hbb3e5580),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad504),
	.w1(32'h39000362),
	.w2(32'hbc5151da),
	.w3(32'hbc843dcc),
	.w4(32'hbc38734c),
	.w5(32'h39bbd4fa),
	.w6(32'h3bd75982),
	.w7(32'hbb6b0f21),
	.w8(32'hbafcd019),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc752c6),
	.w1(32'h3b16fa18),
	.w2(32'hbb2bc1db),
	.w3(32'hba93d268),
	.w4(32'hb9e9d6c1),
	.w5(32'hbb7126d5),
	.w6(32'h3b7f542f),
	.w7(32'hba9e73e3),
	.w8(32'hbbfbddd9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059944),
	.w1(32'hbbbc3787),
	.w2(32'h3a1ab2d8),
	.w3(32'hbb23c88f),
	.w4(32'h394d940a),
	.w5(32'hbae6c3da),
	.w6(32'hbbe03877),
	.w7(32'hba11952e),
	.w8(32'hbbcb0764),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a86bd),
	.w1(32'hbb77b909),
	.w2(32'hbb3569d8),
	.w3(32'hbbdd2713),
	.w4(32'hbb1b5ea5),
	.w5(32'hbbb7ba19),
	.w6(32'hbba371e1),
	.w7(32'hbb94b4f5),
	.w8(32'hbbf2a81c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8b8e),
	.w1(32'h3a324f19),
	.w2(32'hbb36ce3a),
	.w3(32'h393a50f1),
	.w4(32'hbc2057f2),
	.w5(32'h3bdccf04),
	.w6(32'h3c1e876e),
	.w7(32'hbbe44749),
	.w8(32'h3b35eaac),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ea25),
	.w1(32'hb9ac199c),
	.w2(32'h39383d21),
	.w3(32'hb8871fad),
	.w4(32'h3a9af466),
	.w5(32'hbbc9125f),
	.w6(32'hbba08de2),
	.w7(32'hbad2857b),
	.w8(32'hbbe6b457),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ac34),
	.w1(32'hbc331a02),
	.w2(32'hbc88e803),
	.w3(32'hbc487177),
	.w4(32'hbc1d12ec),
	.w5(32'hbb28757b),
	.w6(32'hbb35b131),
	.w7(32'hbc00eb9d),
	.w8(32'h3aaf3d7c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7eac9),
	.w1(32'hbc2fc565),
	.w2(32'hbbea7178),
	.w3(32'hbb523f38),
	.w4(32'hbb9a22dc),
	.w5(32'hbc3d1152),
	.w6(32'h3b04d6fd),
	.w7(32'hbb2482d4),
	.w8(32'hbb75bd0e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8829d3),
	.w1(32'hbc3a36cf),
	.w2(32'hbc083896),
	.w3(32'hbc0db421),
	.w4(32'h3ac953b5),
	.w5(32'h3baa009f),
	.w6(32'hbc341c3d),
	.w7(32'hbb8048d9),
	.w8(32'hbb11e221),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa101b3),
	.w1(32'hbbc7e4c4),
	.w2(32'hbb87cf34),
	.w3(32'hbb5ecd3a),
	.w4(32'hbaa5bba6),
	.w5(32'hbc0c572f),
	.w6(32'hbc5ac15a),
	.w7(32'hbbb8bdfd),
	.w8(32'hbc12b6b1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdde9a5),
	.w1(32'hbc068de7),
	.w2(32'hbbaf0d20),
	.w3(32'hbc059ea2),
	.w4(32'hbbab5303),
	.w5(32'hbb1e5244),
	.w6(32'hbc2633fe),
	.w7(32'hbbc06e66),
	.w8(32'hbb979175),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e2f3d),
	.w1(32'hbc2a81e4),
	.w2(32'hbb5361a6),
	.w3(32'hbb0fa75d),
	.w4(32'hba6cf199),
	.w5(32'hbb2ac8b0),
	.w6(32'h3b97e750),
	.w7(32'hbc6f743d),
	.w8(32'hba34b016),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c5229),
	.w1(32'hbb550377),
	.w2(32'h3b1afb81),
	.w3(32'hbbc7b230),
	.w4(32'hbb66b029),
	.w5(32'h3bdb9962),
	.w6(32'hbbb540d4),
	.w7(32'hba8e2a57),
	.w8(32'h3b901c4e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406994),
	.w1(32'hbb07ea6f),
	.w2(32'h39b5b643),
	.w3(32'h3b3fb35b),
	.w4(32'h3c113057),
	.w5(32'h3a0818ec),
	.w6(32'hbc179ae4),
	.w7(32'h3bc78b69),
	.w8(32'h3b187eb4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae21258),
	.w1(32'hbad3a946),
	.w2(32'hb8bf4a2b),
	.w3(32'hbba3a96b),
	.w4(32'h3be126ad),
	.w5(32'hba78bde2),
	.w6(32'hbbbffb7c),
	.w7(32'h3be2d05b),
	.w8(32'hbb6b5f8d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2307c6),
	.w1(32'hba3e675a),
	.w2(32'h3ae06b36),
	.w3(32'hbb033c48),
	.w4(32'h3a7898e1),
	.w5(32'hba21db03),
	.w6(32'hbc060f60),
	.w7(32'h39c82942),
	.w8(32'h3b319a70),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cde5b),
	.w1(32'hbb316512),
	.w2(32'hbbbce5f6),
	.w3(32'hbbf5df97),
	.w4(32'hbc2eead9),
	.w5(32'hbb5a29d6),
	.w6(32'h3b3c34f8),
	.w7(32'hbba3630d),
	.w8(32'hbab55db0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcec5dc),
	.w1(32'h3b35709e),
	.w2(32'hbb3c5fa9),
	.w3(32'hbbbee85d),
	.w4(32'hbbdf6e90),
	.w5(32'h3b7bd85d),
	.w6(32'hb9944de1),
	.w7(32'hbb9aa38d),
	.w8(32'h3bc22484),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba82b6),
	.w1(32'h3b0dcd9e),
	.w2(32'hbb94e111),
	.w3(32'hba5d483a),
	.w4(32'hbb3d212c),
	.w5(32'h3acc4540),
	.w6(32'h3b152d55),
	.w7(32'h3b1cb75f),
	.w8(32'h3b9eb7e7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510e71),
	.w1(32'hbbe9e4bc),
	.w2(32'h3826bcaf),
	.w3(32'h3ba3a442),
	.w4(32'hbb092002),
	.w5(32'h3b0f791a),
	.w6(32'h3b905f7d),
	.w7(32'h3bd9cb1b),
	.w8(32'h39b8c458),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb132a65),
	.w1(32'h3b7d8832),
	.w2(32'h3b231e1d),
	.w3(32'hb4760886),
	.w4(32'h3b2608bf),
	.w5(32'hba16f513),
	.w6(32'hbaeb0471),
	.w7(32'hbaa66bdb),
	.w8(32'h3b6a5709),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b114175),
	.w1(32'hbaa0037c),
	.w2(32'hbb7de940),
	.w3(32'h3ba0d6b3),
	.w4(32'h3b617824),
	.w5(32'h39ece927),
	.w6(32'hbab6a00e),
	.w7(32'h3b45b9e8),
	.w8(32'h388f2598),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8fe5),
	.w1(32'hbae29d04),
	.w2(32'hbc055259),
	.w3(32'hbbcf8a20),
	.w4(32'hbb6747e8),
	.w5(32'hbb9e7b0f),
	.w6(32'hbbe96d6d),
	.w7(32'hbbdf3e3a),
	.w8(32'hbbb32e5a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf17324),
	.w1(32'hbb32e97e),
	.w2(32'hbc29c3f8),
	.w3(32'hbb1befd8),
	.w4(32'hbbb04fde),
	.w5(32'hbb85c05c),
	.w6(32'h3b662837),
	.w7(32'hbbec4347),
	.w8(32'hbad0d1eb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397743),
	.w1(32'h3b9a4eb8),
	.w2(32'h3bf16683),
	.w3(32'hbb97a26d),
	.w4(32'hbada01c1),
	.w5(32'h3ad402a2),
	.w6(32'hbc5b2cc1),
	.w7(32'hbb1cabaa),
	.w8(32'h3b2afd67),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b2429),
	.w1(32'h3b5ee7a6),
	.w2(32'h3ac53c73),
	.w3(32'h3bb089d0),
	.w4(32'h3a27f839),
	.w5(32'h3c2fe7de),
	.w6(32'h3c2b1a61),
	.w7(32'hb929c8f3),
	.w8(32'h3bfd9b91),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39910905),
	.w1(32'hba3b89b1),
	.w2(32'hbc22de51),
	.w3(32'h3c17844d),
	.w4(32'h3b1c7c82),
	.w5(32'hbb9a959f),
	.w6(32'h3a7eb028),
	.w7(32'hbbac9201),
	.w8(32'hbba9f336),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861110),
	.w1(32'hbb7bda49),
	.w2(32'hbaa00b8d),
	.w3(32'hbbd69101),
	.w4(32'hbb4e47c4),
	.w5(32'hbbf62a2a),
	.w6(32'hbb659fde),
	.w7(32'hbb9e06dc),
	.w8(32'hbbaafb15),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd16c),
	.w1(32'hbb6a59e3),
	.w2(32'hbbebd4b8),
	.w3(32'hbbe70b32),
	.w4(32'hbbde8801),
	.w5(32'hbc0f0040),
	.w6(32'hbb3e7b14),
	.w7(32'hbbf54e27),
	.w8(32'hbbaba3c1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9304d0),
	.w1(32'hbbbf81f2),
	.w2(32'hbbcc3f73),
	.w3(32'hbb8ae03f),
	.w4(32'hba7758b8),
	.w5(32'hbbe5bb53),
	.w6(32'hbbc41032),
	.w7(32'hbbfd5b23),
	.w8(32'hbbd8c483),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffde94),
	.w1(32'hbc198b83),
	.w2(32'hbc10010e),
	.w3(32'hbc4839d4),
	.w4(32'hbc07eeb7),
	.w5(32'h3a578393),
	.w6(32'hbc08272d),
	.w7(32'hbbdcbe71),
	.w8(32'hb8c09901),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2f87b),
	.w1(32'hbab2ed8c),
	.w2(32'hbabf0574),
	.w3(32'hbb515389),
	.w4(32'h39f05be3),
	.w5(32'hbb81b715),
	.w6(32'hba65f030),
	.w7(32'hb9ac39fb),
	.w8(32'hba965c92),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153de1),
	.w1(32'h3a2c618d),
	.w2(32'h3ac2a913),
	.w3(32'hb92436b5),
	.w4(32'hbab47702),
	.w5(32'hbb3607f4),
	.w6(32'h3b0dc1ec),
	.w7(32'hbb03f5bb),
	.w8(32'hbb7b30b1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6422),
	.w1(32'hbb8df3f6),
	.w2(32'hbc350885),
	.w3(32'hbbe990e0),
	.w4(32'h3a42e422),
	.w5(32'hbaadeed3),
	.w6(32'hbb03eac7),
	.w7(32'hbbda0584),
	.w8(32'h3bf9c2bd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bdf01),
	.w1(32'h3c363920),
	.w2(32'h3aeeb05b),
	.w3(32'hbb86c50f),
	.w4(32'h3ab76d1f),
	.w5(32'hbb2994ce),
	.w6(32'h3c4bf2f7),
	.w7(32'h3bfbcc09),
	.w8(32'hba3e6255),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc5bd),
	.w1(32'h3a8d173b),
	.w2(32'h3b9fc6b0),
	.w3(32'h3a4ae73a),
	.w4(32'hbbb0929a),
	.w5(32'hbaf1fe6d),
	.w6(32'hba9d2929),
	.w7(32'h3b35dece),
	.w8(32'hbac3afb0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319e50),
	.w1(32'h389e702f),
	.w2(32'h3ae2ace3),
	.w3(32'h3acdb18b),
	.w4(32'h39bfb085),
	.w5(32'hba1abc91),
	.w6(32'h3c42bab6),
	.w7(32'h3b28e95c),
	.w8(32'hbb1a0219),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547a27),
	.w1(32'hba35e05a),
	.w2(32'hbbe27992),
	.w3(32'hb91ab8e2),
	.w4(32'hbb9a86e3),
	.w5(32'hbb23dccc),
	.w6(32'h3bc6cd34),
	.w7(32'hbb60b40c),
	.w8(32'hba7ebf8c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87fe6f),
	.w1(32'hb8c7cde1),
	.w2(32'hbb5eb7ea),
	.w3(32'hbbaab3e0),
	.w4(32'hba28fef5),
	.w5(32'hba84663b),
	.w6(32'h3be29af6),
	.w7(32'h3994d79d),
	.w8(32'h38acd0b3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e5b58),
	.w1(32'h38c46f8d),
	.w2(32'hbabfd295),
	.w3(32'hbbf0d030),
	.w4(32'hbb87c749),
	.w5(32'hba809d46),
	.w6(32'hbb840f73),
	.w7(32'hbb67e839),
	.w8(32'hb9f89ca4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337582),
	.w1(32'hbc1e103a),
	.w2(32'h3ab63b7c),
	.w3(32'hbbf52ee7),
	.w4(32'hbc1aa3dd),
	.w5(32'hbac2fddd),
	.w6(32'hbad7650b),
	.w7(32'hbbe1c96e),
	.w8(32'h3bcd0780),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4843ce),
	.w1(32'hbbb949e5),
	.w2(32'h39b6ae47),
	.w3(32'hbbfdcfcd),
	.w4(32'hbb32cfed),
	.w5(32'h3b84bbb7),
	.w6(32'hbb8ba9ea),
	.w7(32'h3aa1fb57),
	.w8(32'hbab894ec),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4e24),
	.w1(32'h3b0ff3e8),
	.w2(32'hba7ad73d),
	.w3(32'hb7f7051b),
	.w4(32'hbb2104c9),
	.w5(32'hb9051679),
	.w6(32'h3b6bb35f),
	.w7(32'hbaded135),
	.w8(32'hbb40db1f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac48a33),
	.w1(32'hbb4e42e3),
	.w2(32'hb9cdda5d),
	.w3(32'h3a301852),
	.w4(32'h3b8ecc89),
	.w5(32'hbac9f470),
	.w6(32'hbba47b43),
	.w7(32'hba967d2d),
	.w8(32'hba629a8b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f298b),
	.w1(32'hbb865395),
	.w2(32'hbb0e488d),
	.w3(32'hbc0dcaa0),
	.w4(32'hbb5bbf51),
	.w5(32'hb991c5f5),
	.w6(32'hbbb20b69),
	.w7(32'hbb941884),
	.w8(32'h3bd03326),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be46aa8),
	.w1(32'hbac2a6bc),
	.w2(32'hbbb962a8),
	.w3(32'hbad1aac9),
	.w4(32'hbb4c9a66),
	.w5(32'h3b78c399),
	.w6(32'hb92a6278),
	.w7(32'hbb80d130),
	.w8(32'h3ac0a327),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f05ac),
	.w1(32'h395208a3),
	.w2(32'h3b201271),
	.w3(32'h3bd8368f),
	.w4(32'h3b05a672),
	.w5(32'h3a25401a),
	.w6(32'hbb785e3f),
	.w7(32'hbb04c9a6),
	.w8(32'hbb1897e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52603),
	.w1(32'hbb549e37),
	.w2(32'hbab2158e),
	.w3(32'hbaf59f99),
	.w4(32'hbabb87bc),
	.w5(32'hbbbda698),
	.w6(32'h3bf373e1),
	.w7(32'hbaff99e0),
	.w8(32'hbbd52f25),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e537),
	.w1(32'hbbb9d259),
	.w2(32'hbb29328b),
	.w3(32'hbb6d15d7),
	.w4(32'hba76d8be),
	.w5(32'h3af5b05d),
	.w6(32'hbb6c5263),
	.w7(32'h3a40154a),
	.w8(32'hb9916be4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ae31f),
	.w1(32'hbb8c5ef8),
	.w2(32'hbb5306e5),
	.w3(32'hbc002eb8),
	.w4(32'hbb82e888),
	.w5(32'h3b53b1fd),
	.w6(32'hbbc66e55),
	.w7(32'hbbc8b915),
	.w8(32'h3bf3d344),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac210e6),
	.w1(32'h3c34462f),
	.w2(32'h3c1f2eee),
	.w3(32'h3b549868),
	.w4(32'hbb04f07f),
	.w5(32'h3b2535ce),
	.w6(32'h3a9fdc5f),
	.w7(32'h3bbbee0a),
	.w8(32'hba2f2ac4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae84d24),
	.w1(32'h3b762bec),
	.w2(32'h3a04c535),
	.w3(32'h3a5df33d),
	.w4(32'hba97f338),
	.w5(32'h3b50f50d),
	.w6(32'h3aad3769),
	.w7(32'hba8781c2),
	.w8(32'hbc0f7975),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb49b61),
	.w1(32'hbc9b767c),
	.w2(32'hbc1f4698),
	.w3(32'h3bbe822d),
	.w4(32'hb9eb8bba),
	.w5(32'hbbf9bb4f),
	.w6(32'hbb10b344),
	.w7(32'hbc9e02c0),
	.w8(32'hbbafd108),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b719df6),
	.w1(32'hbac7d483),
	.w2(32'h3b4bcbbb),
	.w3(32'hbc28d208),
	.w4(32'hbb713677),
	.w5(32'hbbba8598),
	.w6(32'hbc8d8238),
	.w7(32'hbb8f75ae),
	.w8(32'h3a585192),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d454d2),
	.w1(32'hbc23e7d9),
	.w2(32'hbb6f80d2),
	.w3(32'hbc67abf6),
	.w4(32'hbba51d35),
	.w5(32'h3ba1407b),
	.w6(32'hbbc070d4),
	.w7(32'hbb4ccb86),
	.w8(32'h3955fe98),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d5dc3),
	.w1(32'h3b2535d0),
	.w2(32'hbb3d744e),
	.w3(32'hbbd3bb80),
	.w4(32'hbb75bb29),
	.w5(32'hbb2cce0a),
	.w6(32'hbb0948e9),
	.w7(32'hba7bfc44),
	.w8(32'hbaaadb6e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6ff8),
	.w1(32'hbad455ac),
	.w2(32'hb8bccd9d),
	.w3(32'hbb9550d5),
	.w4(32'hbafc4f3b),
	.w5(32'hba781217),
	.w6(32'hbb895cc0),
	.w7(32'h3946a152),
	.w8(32'hbb780600),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11822e),
	.w1(32'hbbdd21b4),
	.w2(32'hbb66090d),
	.w3(32'hbb863e09),
	.w4(32'h3b18cd61),
	.w5(32'hbbeca4cb),
	.w6(32'hbb385ed0),
	.w7(32'hbb4969f9),
	.w8(32'hbaf6aab0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82dbd66),
	.w1(32'hbbf35612),
	.w2(32'hbbc26289),
	.w3(32'hbb7b741e),
	.w4(32'hbbdb6a87),
	.w5(32'hbb4b1482),
	.w6(32'hbb132f73),
	.w7(32'hbb35e009),
	.w8(32'h3a4c784f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1693d),
	.w1(32'hbb3a907d),
	.w2(32'hbb100def),
	.w3(32'hba12c233),
	.w4(32'hba1c1889),
	.w5(32'hbbe7d63c),
	.w6(32'h3b96ffc2),
	.w7(32'hba359454),
	.w8(32'hb90c1ec4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0b1e),
	.w1(32'hbb875fe3),
	.w2(32'hbb01f3e8),
	.w3(32'hbb9a931c),
	.w4(32'hbbe49d0c),
	.w5(32'hba578274),
	.w6(32'h3a144d94),
	.w7(32'hbc1783e5),
	.w8(32'hbbd9a539),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5788a),
	.w1(32'h39956604),
	.w2(32'h3b91bf25),
	.w3(32'hbb2c333b),
	.w4(32'hbb99a3a2),
	.w5(32'h3ad01375),
	.w6(32'hbc106f77),
	.w7(32'h3bf4f68e),
	.w8(32'hbb2d8fe6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba3645),
	.w1(32'hba7a77ed),
	.w2(32'h3a804547),
	.w3(32'hbb398c35),
	.w4(32'h3a1af3c7),
	.w5(32'h39e722e8),
	.w6(32'hbc823ab4),
	.w7(32'h3b214a6c),
	.w8(32'hbb571125),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57ac55),
	.w1(32'h397f893d),
	.w2(32'hba1750de),
	.w3(32'h3a688512),
	.w4(32'h3b0131f5),
	.w5(32'hbc3afc5d),
	.w6(32'h3b349d96),
	.w7(32'h37f97d86),
	.w8(32'hbc74368e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3951),
	.w1(32'hbc89478b),
	.w2(32'hbcb16ab8),
	.w3(32'hbc8f1b7c),
	.w4(32'hbcd3068a),
	.w5(32'hbc1cc48d),
	.w6(32'hbc4a9bee),
	.w7(32'hbccecd17),
	.w8(32'hbbc2de47),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc040327),
	.w1(32'hbc4afad1),
	.w2(32'hbbe08947),
	.w3(32'hbc54e4b1),
	.w4(32'hbc00a302),
	.w5(32'hbb0dfa47),
	.w6(32'h3c53aaca),
	.w7(32'hbc083a06),
	.w8(32'h3bd7690d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3e4ba),
	.w1(32'hbbf54428),
	.w2(32'hbb169952),
	.w3(32'hbb859bfd),
	.w4(32'hba04a181),
	.w5(32'h3cab9e47),
	.w6(32'hbbe51f69),
	.w7(32'h3b2632a0),
	.w8(32'h3c91420d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e7f78),
	.w1(32'h3c8fea02),
	.w2(32'h3c583358),
	.w3(32'h3cbfe23a),
	.w4(32'h3c9a7d1e),
	.w5(32'h3b15d997),
	.w6(32'h3ca7bcf6),
	.w7(32'h3ca42c0b),
	.w8(32'h3c0c0e30),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbe02e),
	.w1(32'h3c3113cd),
	.w2(32'h3ae0c274),
	.w3(32'h3bb2b7ad),
	.w4(32'h3b2b3be2),
	.w5(32'hbbd1a245),
	.w6(32'h3b668c15),
	.w7(32'h3c308957),
	.w8(32'hbc177656),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaa558),
	.w1(32'hbbd870b8),
	.w2(32'hbc197caa),
	.w3(32'hba997829),
	.w4(32'hbb64446a),
	.w5(32'hbae71b0b),
	.w6(32'hbb53be3a),
	.w7(32'hbc0e80b4),
	.w8(32'h3bb704f6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba4014),
	.w1(32'hbbb42f6e),
	.w2(32'hbbd75608),
	.w3(32'hbbe9eda3),
	.w4(32'hbbae1de7),
	.w5(32'hbb1f04e4),
	.w6(32'hba9373af),
	.w7(32'hbbbd1fef),
	.w8(32'hbb8b980d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65c09c),
	.w1(32'hbb79faad),
	.w2(32'hba5b07fc),
	.w3(32'hbabaf8d1),
	.w4(32'h3b5adcca),
	.w5(32'h3bde2477),
	.w6(32'hbbf7332b),
	.w7(32'h3a45aef8),
	.w8(32'hbba2cd9c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12228),
	.w1(32'hbc26906e),
	.w2(32'hbac5d4ab),
	.w3(32'hbc2e005f),
	.w4(32'h3b954903),
	.w5(32'hbaec880a),
	.w6(32'hbca3eb5d),
	.w7(32'hbbe51750),
	.w8(32'hbaa3fa13),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3dcaa),
	.w1(32'hbb8b6e8c),
	.w2(32'hbaa2d31d),
	.w3(32'hbace3dc0),
	.w4(32'h3b46b8eb),
	.w5(32'h38c52b10),
	.w6(32'h3bd4014d),
	.w7(32'hbb643531),
	.w8(32'hbb790139),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5e387),
	.w1(32'hbae532eb),
	.w2(32'hb965d874),
	.w3(32'hba168be2),
	.w4(32'h3b6466e0),
	.w5(32'hbc1011d6),
	.w6(32'hba06f9b8),
	.w7(32'hb985ebc0),
	.w8(32'hbc7288a7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18cb07),
	.w1(32'hbbe65cf4),
	.w2(32'hba8288b5),
	.w3(32'hbbe36c17),
	.w4(32'hba5dfff6),
	.w5(32'hbb9df784),
	.w6(32'hbc7f28ad),
	.w7(32'h3c2e7214),
	.w8(32'h3a003fc1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3298),
	.w1(32'hbbafb436),
	.w2(32'hbb54209c),
	.w3(32'hbbd673d1),
	.w4(32'hbb8f6bd5),
	.w5(32'h3b3b54c3),
	.w6(32'hbb6d337d),
	.w7(32'hbbb33c89),
	.w8(32'h3b4d5c77),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7197c9),
	.w1(32'h3b0e7556),
	.w2(32'hbb3023e7),
	.w3(32'hba45988a),
	.w4(32'h3a86e3e4),
	.w5(32'hbae7a0b1),
	.w6(32'hbbd34691),
	.w7(32'hbaefb5ad),
	.w8(32'hbb82f960),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025e54),
	.w1(32'hba0e2b55),
	.w2(32'h3ab39906),
	.w3(32'hba246954),
	.w4(32'hba85cf5c),
	.w5(32'hbb0e44b5),
	.w6(32'hbc28da40),
	.w7(32'h3bb4c9ec),
	.w8(32'hbb5556f4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90df259),
	.w1(32'hbb746095),
	.w2(32'hbc0545f8),
	.w3(32'h3b0abf7c),
	.w4(32'hbb8fcbd5),
	.w5(32'hbb9ed469),
	.w6(32'h3c21f062),
	.w7(32'hbb88001f),
	.w8(32'hbbec454e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef1b4c),
	.w1(32'hbbcc01ef),
	.w2(32'hbbadde72),
	.w3(32'hbbc0f00e),
	.w4(32'hbab95f6f),
	.w5(32'h3c78540e),
	.w6(32'hbc1c62b6),
	.w7(32'hbb91f6ee),
	.w8(32'h3c756942),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4d60),
	.w1(32'h3a82a8c1),
	.w2(32'h3b9efc82),
	.w3(32'h3bca8a53),
	.w4(32'h3c90e037),
	.w5(32'hbb2dcfaa),
	.w6(32'hbb885f97),
	.w7(32'h3c023e34),
	.w8(32'hbb176e1d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae32057),
	.w1(32'h3a4f3e5d),
	.w2(32'h3b3ca3ad),
	.w3(32'h3ae43ef5),
	.w4(32'hba6fce70),
	.w5(32'h3bf825e0),
	.w6(32'h3b8e07b6),
	.w7(32'hbbd9f301),
	.w8(32'h3bdb680c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2c9c),
	.w1(32'h3c327d24),
	.w2(32'h3bbe8656),
	.w3(32'h3bd7b082),
	.w4(32'h3bb88e28),
	.w5(32'h3a970bae),
	.w6(32'h3c6ff0c5),
	.w7(32'h3c21802b),
	.w8(32'h3bbc5692),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf39ba),
	.w1(32'hba8b3c3e),
	.w2(32'hbb947693),
	.w3(32'h3b67beab),
	.w4(32'h3991aab9),
	.w5(32'h3b016849),
	.w6(32'h3bd94b46),
	.w7(32'hbacfa2cd),
	.w8(32'hbad7fb53),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb291cc4),
	.w1(32'hbb081213),
	.w2(32'h3b0a3501),
	.w3(32'hba1f2027),
	.w4(32'hba2710dc),
	.w5(32'h39ea7d34),
	.w6(32'hbbe835a8),
	.w7(32'h3b8ff63c),
	.w8(32'hba9f8aaa),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000a89),
	.w1(32'hbb957cc5),
	.w2(32'hbabcef47),
	.w3(32'hbb4b6f25),
	.w4(32'h39f62f88),
	.w5(32'hbb3f2f79),
	.w6(32'hbbec8c2b),
	.w7(32'hbbc1b22e),
	.w8(32'h3a6b7325),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c458),
	.w1(32'h399d167c),
	.w2(32'hba88f191),
	.w3(32'h39e11ab2),
	.w4(32'h3a9f095f),
	.w5(32'hbaea78da),
	.w6(32'h3be88037),
	.w7(32'hbb0745a6),
	.w8(32'hbac99e7b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eca69),
	.w1(32'hbb613d45),
	.w2(32'hbb96ccb5),
	.w3(32'h3bb09312),
	.w4(32'hbb0b2095),
	.w5(32'hbae28a62),
	.w6(32'h3af8f468),
	.w7(32'hbba702cb),
	.w8(32'hbbcd799a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009371),
	.w1(32'hbbd2922e),
	.w2(32'hbbb1a28c),
	.w3(32'hbb3c9cca),
	.w4(32'hbb7509d3),
	.w5(32'h3b139a7f),
	.w6(32'h3baff6bf),
	.w7(32'hbadec0ed),
	.w8(32'h3b9ff47f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0a099),
	.w1(32'hbb136142),
	.w2(32'hb98d1738),
	.w3(32'hbbbfd6bb),
	.w4(32'hb9bc4b8c),
	.w5(32'hba35a3f3),
	.w6(32'hbc40fd75),
	.w7(32'hbbe7f5bd),
	.w8(32'h3a5fbc72),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051d2e),
	.w1(32'h3b235f03),
	.w2(32'hbbfe9a49),
	.w3(32'hbbebd8f6),
	.w4(32'hbbde1bfe),
	.w5(32'hbc3bb9c2),
	.w6(32'h3c4e6fd6),
	.w7(32'hbc0170cb),
	.w8(32'hbc14f043),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ed9b),
	.w1(32'hbbe7ed27),
	.w2(32'hbbee0de3),
	.w3(32'hbc2e2c67),
	.w4(32'hbc49b6de),
	.w5(32'hbb869662),
	.w6(32'hb98ec8be),
	.w7(32'hbc071e21),
	.w8(32'hba342221),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc85a2),
	.w1(32'h3beb1f91),
	.w2(32'hbbcecef0),
	.w3(32'h3ba1827e),
	.w4(32'h3aa24d3a),
	.w5(32'hbb10c37a),
	.w6(32'h3c4d3f76),
	.w7(32'hbc0667fd),
	.w8(32'h3955cc6b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3938e),
	.w1(32'h3a0787f2),
	.w2(32'hbb6cc416),
	.w3(32'h3a8fb070),
	.w4(32'h3b197073),
	.w5(32'h3b477238),
	.w6(32'h3bca31d8),
	.w7(32'hbbacb9ff),
	.w8(32'hbba93ba9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7dd19),
	.w1(32'h3b0ddeea),
	.w2(32'h3bbfbb82),
	.w3(32'h3a982a59),
	.w4(32'h3ab22b7c),
	.w5(32'hbacc1cb5),
	.w6(32'h3b5f6833),
	.w7(32'hb9a12c66),
	.w8(32'h3b083ac5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f93281),
	.w1(32'hbb692788),
	.w2(32'hbb9e8679),
	.w3(32'hbbed0ae0),
	.w4(32'hbc0e5d90),
	.w5(32'h3bf6ae1c),
	.w6(32'h3ae78837),
	.w7(32'hb99d266e),
	.w8(32'h3bd9af52),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92fa33),
	.w1(32'h3bff1a30),
	.w2(32'h3bd62b6d),
	.w3(32'h3b1edaf6),
	.w4(32'h3b9e10fa),
	.w5(32'h3b27a8b7),
	.w6(32'h3bd01cfa),
	.w7(32'h3b8af352),
	.w8(32'h38eeee11),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43817a),
	.w1(32'hbc66681c),
	.w2(32'hbab55afa),
	.w3(32'hbbad620a),
	.w4(32'hbb28dffa),
	.w5(32'h39a9eee4),
	.w6(32'hbbc10417),
	.w7(32'hbbd9ea72),
	.w8(32'h3b58f750),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90aa37),
	.w1(32'hbb2efdcb),
	.w2(32'hbbc38b57),
	.w3(32'h3a8973fd),
	.w4(32'hbab116b1),
	.w5(32'h3c69653a),
	.w6(32'h3c48c8e6),
	.w7(32'h39287543),
	.w8(32'h3b91735a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba06515),
	.w1(32'h3bbcd5e6),
	.w2(32'h3bb8b158),
	.w3(32'h3bc3deb6),
	.w4(32'h3c195104),
	.w5(32'hbb8e4179),
	.w6(32'hbad4be4d),
	.w7(32'h3aa8af38),
	.w8(32'hbbf1f67d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083ed4),
	.w1(32'hbbb6ef0e),
	.w2(32'hbb7d30d1),
	.w3(32'hbbe625af),
	.w4(32'hbad059c5),
	.w5(32'hbad902e1),
	.w6(32'hbb361620),
	.w7(32'hbb66e76a),
	.w8(32'hbc00f382),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c165),
	.w1(32'h3ae429f7),
	.w2(32'hbbf2e396),
	.w3(32'h3aa3fb77),
	.w4(32'hbacc8be9),
	.w5(32'hb97b945d),
	.w6(32'hbc6deee4),
	.w7(32'hbc09131c),
	.w8(32'hbb152a92),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacddd88),
	.w1(32'hbb72e8f5),
	.w2(32'hbbbe768d),
	.w3(32'hbb19efce),
	.w4(32'hbb90dfaa),
	.w5(32'hbae8356e),
	.w6(32'h39063613),
	.w7(32'hbbc4a2a0),
	.w8(32'h3a887936),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3cd8c),
	.w1(32'hbbf7bc33),
	.w2(32'hbad39653),
	.w3(32'hbb72b6ba),
	.w4(32'h3a2209a7),
	.w5(32'h3b3d76f4),
	.w6(32'hbb8e4a0e),
	.w7(32'hbb98babb),
	.w8(32'hbace759a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49809c),
	.w1(32'hb9153605),
	.w2(32'h3c248ecf),
	.w3(32'h3c067fcb),
	.w4(32'h3bb9d21f),
	.w5(32'h3ad9b152),
	.w6(32'h3b6aabf6),
	.w7(32'h3bfef903),
	.w8(32'h3b8306fc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee7d36),
	.w1(32'hbb8adee2),
	.w2(32'hbc027a35),
	.w3(32'hba365f86),
	.w4(32'hbb2362d5),
	.w5(32'h3b491cc6),
	.w6(32'h3b1133ad),
	.w7(32'hbbb66204),
	.w8(32'h3abcfac5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c05db),
	.w1(32'h3b0000c0),
	.w2(32'h3c43b440),
	.w3(32'hbb02ebaf),
	.w4(32'h3bca7765),
	.w5(32'hbc0602d7),
	.w6(32'h39e82b89),
	.w7(32'h3b912355),
	.w8(32'hbbf62934),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520ab5),
	.w1(32'hbb01ab56),
	.w2(32'hbc28c7ad),
	.w3(32'hbba0e292),
	.w4(32'hbb89dffb),
	.w5(32'h3b72304e),
	.w6(32'hbb52347a),
	.w7(32'hbbb73698),
	.w8(32'h3b8eab8d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5da970),
	.w1(32'hbbfc528d),
	.w2(32'hbb336e4d),
	.w3(32'h3b43b69d),
	.w4(32'h3a3ea9b2),
	.w5(32'hbbeb229b),
	.w6(32'hb9810daa),
	.w7(32'hba65e13d),
	.w8(32'hbbec0f52),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046d72),
	.w1(32'hbbfe6f67),
	.w2(32'hbbcdc2fd),
	.w3(32'hbbfac9c8),
	.w4(32'hbb78a72a),
	.w5(32'h3a7197a4),
	.w6(32'hbb2f1f98),
	.w7(32'hbb60fac5),
	.w8(32'hbbd13578),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f81d2),
	.w1(32'h3bda51ac),
	.w2(32'hbabfebd5),
	.w3(32'hbb97b143),
	.w4(32'hbb8b278c),
	.w5(32'h3b521767),
	.w6(32'hbbf93b7b),
	.w7(32'h3b7b3740),
	.w8(32'h3bebece6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dda5e),
	.w1(32'h3aa7cde8),
	.w2(32'hb888aeff),
	.w3(32'hbbecb374),
	.w4(32'h398df97d),
	.w5(32'h3b314033),
	.w6(32'hbc133399),
	.w7(32'h3b86766a),
	.w8(32'h3a8bb220),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd170e3),
	.w1(32'h3b2ba716),
	.w2(32'h3b2d6df2),
	.w3(32'h39561d2c),
	.w4(32'h3b51795f),
	.w5(32'hbc267b7b),
	.w6(32'hbb3cae9e),
	.w7(32'h3b9b860f),
	.w8(32'hbbf5626b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bbe25),
	.w1(32'hbb4ce040),
	.w2(32'hbb83c9cb),
	.w3(32'hba64003a),
	.w4(32'h3b9bf970),
	.w5(32'h3a949646),
	.w6(32'hbc541388),
	.w7(32'hbbd4896e),
	.w8(32'h3b557d1e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277003),
	.w1(32'h3aeb50be),
	.w2(32'h3bbbcd09),
	.w3(32'h3aea771a),
	.w4(32'h397a1f25),
	.w5(32'h3a5d7be7),
	.w6(32'hbaf41971),
	.w7(32'hba970527),
	.w8(32'hbaee6307),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97042c),
	.w1(32'hbb871945),
	.w2(32'hbbd742cd),
	.w3(32'hbafba86e),
	.w4(32'hbb33b52d),
	.w5(32'hbc184329),
	.w6(32'hbb07b584),
	.w7(32'hbbb31610),
	.w8(32'hbb96b59b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a01c30),
	.w1(32'hbbc4060e),
	.w2(32'hbb69b201),
	.w3(32'hbc133836),
	.w4(32'hbc72a9fc),
	.w5(32'h3cbd21b2),
	.w6(32'hbc7a5fa7),
	.w7(32'hbc839b3a),
	.w8(32'h3bff8a42),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c871a71),
	.w1(32'h3c29e6eb),
	.w2(32'h3ca2e00b),
	.w3(32'h3c9d1355),
	.w4(32'h3cbe7575),
	.w5(32'hbc006fa1),
	.w6(32'hbbd0e016),
	.w7(32'h3c6a44ac),
	.w8(32'hbc0a1e96),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2fd3e),
	.w1(32'hbc9e22e0),
	.w2(32'hbb45b5f6),
	.w3(32'hbbfd2b5a),
	.w4(32'hbb60c598),
	.w5(32'hbb9cb4da),
	.w6(32'hbc987d50),
	.w7(32'hbc199f19),
	.w8(32'hbbab39cf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b85bd),
	.w1(32'h3ab5b522),
	.w2(32'hbbb13313),
	.w3(32'h3b989d99),
	.w4(32'hbbbcced7),
	.w5(32'h3b6d68eb),
	.w6(32'h3b277e52),
	.w7(32'hbbdbe56b),
	.w8(32'hbc30edfc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39f4ac),
	.w1(32'h3bbbf063),
	.w2(32'hbb317f7d),
	.w3(32'hbbc6869d),
	.w4(32'hbbcd0c03),
	.w5(32'hbc04d5b1),
	.w6(32'hbb472426),
	.w7(32'hbafb5f7c),
	.w8(32'hbbd03aed),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12a467),
	.w1(32'h3cae244c),
	.w2(32'h3c901b8f),
	.w3(32'h3b7d84c1),
	.w4(32'hba532c4c),
	.w5(32'hbbcfa0cf),
	.w6(32'hbb40729e),
	.w7(32'hba7d4664),
	.w8(32'hba8e3c38),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023231),
	.w1(32'hbb954dc3),
	.w2(32'h3ab737e8),
	.w3(32'h3b1ff44c),
	.w4(32'h3b68e101),
	.w5(32'hbae03c37),
	.w6(32'h3c26ec14),
	.w7(32'h3bdb7c52),
	.w8(32'hbb02281e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47876e),
	.w1(32'h3b12fce2),
	.w2(32'hba9f073c),
	.w3(32'hbaaa1ac1),
	.w4(32'hba7cfabe),
	.w5(32'hbc1fe4fa),
	.w6(32'hba52c1b0),
	.w7(32'h391eeacd),
	.w8(32'h3a287308),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5c63),
	.w1(32'h3afd003b),
	.w2(32'h3c614cf8),
	.w3(32'h3b44690b),
	.w4(32'hbb90ee4c),
	.w5(32'hba80cb89),
	.w6(32'hbca0759b),
	.w7(32'h3c013ed2),
	.w8(32'h3b6464cc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e1b53),
	.w1(32'hbba7cb7b),
	.w2(32'hbaea794c),
	.w3(32'hbc8c7f26),
	.w4(32'h3abb547a),
	.w5(32'hbb3f63f7),
	.w6(32'h3d19cc26),
	.w7(32'h3cb7b193),
	.w8(32'h3c299b5a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859e115),
	.w1(32'h3b9d4a71),
	.w2(32'h3a1a7e77),
	.w3(32'h3b28a6c2),
	.w4(32'h3c15e64f),
	.w5(32'hbb708cce),
	.w6(32'hbb53d2ef),
	.w7(32'h3ba65b67),
	.w8(32'hbb2c9752),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ea3c),
	.w1(32'h3c05ebb3),
	.w2(32'hbc0e628a),
	.w3(32'hbbf691ee),
	.w4(32'hbc4d9c6f),
	.w5(32'hbaaa7400),
	.w6(32'hbbe7cfa8),
	.w7(32'h3baabeae),
	.w8(32'hbb68b9f0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be057),
	.w1(32'hbaada9f3),
	.w2(32'hbb06bc54),
	.w3(32'hbaf3f422),
	.w4(32'hbaf60c99),
	.w5(32'hbbf0fd54),
	.w6(32'h3b8f3144),
	.w7(32'hba893df1),
	.w8(32'hbc1440dc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a5f29),
	.w1(32'h3b88d924),
	.w2(32'h3a22f1bb),
	.w3(32'h3c14ab8a),
	.w4(32'hbbb96173),
	.w5(32'hbb085ec9),
	.w6(32'h3c048c5f),
	.w7(32'hbbf0f159),
	.w8(32'hba1f5ff5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a479344),
	.w1(32'hbb366336),
	.w2(32'hba17bef3),
	.w3(32'hbbd5cf03),
	.w4(32'hbb41e5ee),
	.w5(32'h3bf5433e),
	.w6(32'hbb63f477),
	.w7(32'hba0d9186),
	.w8(32'h3b52a530),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b181),
	.w1(32'h3a9dec0e),
	.w2(32'h3bc48aef),
	.w3(32'h3b5245fd),
	.w4(32'h3aeefff6),
	.w5(32'hbac0c4d8),
	.w6(32'h3c90b58a),
	.w7(32'h3c9219fa),
	.w8(32'h3b058caf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81979),
	.w1(32'hbc0152e4),
	.w2(32'hbba54370),
	.w3(32'hbb8cc843),
	.w4(32'hbba1cc88),
	.w5(32'hbb84b178),
	.w6(32'hbc246a68),
	.w7(32'hbbd85a72),
	.w8(32'hbc1f9047),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016c84),
	.w1(32'hbbbeecc9),
	.w2(32'hbb0b71d0),
	.w3(32'hbbdda8e8),
	.w4(32'hba804287),
	.w5(32'hbb66c702),
	.w6(32'hbc1020a5),
	.w7(32'hbba5bc5e),
	.w8(32'hb9883c03),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b83de),
	.w1(32'h3aea5a3e),
	.w2(32'h3b498677),
	.w3(32'h3adcb307),
	.w4(32'hbb1f200e),
	.w5(32'hbc2b276a),
	.w6(32'hbb0e5552),
	.w7(32'h39a35bbc),
	.w8(32'h3b19a2d5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68d84),
	.w1(32'h3be2a182),
	.w2(32'hbc241bc6),
	.w3(32'hbbed24d2),
	.w4(32'h3b232ec7),
	.w5(32'hbb67120a),
	.w6(32'hba1bfad6),
	.w7(32'h3abc8cde),
	.w8(32'h3ba68ffa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881415),
	.w1(32'hbb1d4172),
	.w2(32'hbb2f58a8),
	.w3(32'h39b858fe),
	.w4(32'hbc2000db),
	.w5(32'hb86c926f),
	.w6(32'h3b2bdeac),
	.w7(32'hbbca4a6f),
	.w8(32'hbb6e9755),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9906),
	.w1(32'hbc02a62d),
	.w2(32'hbba1ba4d),
	.w3(32'h3b783adf),
	.w4(32'h3bc16496),
	.w5(32'hbbd9ef4e),
	.w6(32'hbbd3e0f4),
	.w7(32'hbb3f17e4),
	.w8(32'h3bad3780),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38b3d),
	.w1(32'h3b23285c),
	.w2(32'hbbd476d4),
	.w3(32'hbc4ec20c),
	.w4(32'h3ba6f915),
	.w5(32'hbaf20340),
	.w6(32'h3d044c4a),
	.w7(32'h3bd2e295),
	.w8(32'h3beaeb56),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc892ce),
	.w1(32'hbb87130b),
	.w2(32'hbc1326ca),
	.w3(32'hba9204c7),
	.w4(32'hbbf33e4e),
	.w5(32'hbc44f33a),
	.w6(32'h3bed7712),
	.w7(32'h3b83be68),
	.w8(32'hbba79d91),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe360d),
	.w1(32'h3b9fc919),
	.w2(32'hbb3757e1),
	.w3(32'h3c48f74a),
	.w4(32'hbc4a7de9),
	.w5(32'h3a76ee09),
	.w6(32'h3b8ed63a),
	.w7(32'hbc7ba352),
	.w8(32'h38799000),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16cfd8),
	.w1(32'hbbea81aa),
	.w2(32'hbbba811e),
	.w3(32'h3ba817a6),
	.w4(32'h3a473439),
	.w5(32'h3a973a9c),
	.w6(32'h3b7470a3),
	.w7(32'h3ada3862),
	.w8(32'hbad6dec7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d67f1),
	.w1(32'hbc091c4c),
	.w2(32'hbc0456c9),
	.w3(32'hba461a0f),
	.w4(32'hbbc2eb75),
	.w5(32'hbc265bba),
	.w6(32'hbb1ee509),
	.w7(32'hbc480eb4),
	.w8(32'hbaacc293),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44bf88),
	.w1(32'h3a95a18d),
	.w2(32'hbb957840),
	.w3(32'hba85b02a),
	.w4(32'hb91b82c1),
	.w5(32'hbb888398),
	.w6(32'hbb4e3977),
	.w7(32'hba0d33ca),
	.w8(32'hbbfa228a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e37b),
	.w1(32'hbbc2ee97),
	.w2(32'hbb8f3cd6),
	.w3(32'hbad63cac),
	.w4(32'hbb30e711),
	.w5(32'h3bda9bec),
	.w6(32'h3b06b822),
	.w7(32'hbc656c0f),
	.w8(32'hbbe56f3b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c189080),
	.w1(32'h3c658392),
	.w2(32'h3be9bdb4),
	.w3(32'h3c080f99),
	.w4(32'h3b225484),
	.w5(32'hba5cc5a7),
	.w6(32'hbc0ebe5b),
	.w7(32'hbb75c2d2),
	.w8(32'hbad72d3b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba716c85),
	.w1(32'hbba34805),
	.w2(32'hbc06f3f6),
	.w3(32'hb9c3ee9c),
	.w4(32'hb7d03825),
	.w5(32'hbc3b225b),
	.w6(32'h3ada2d64),
	.w7(32'h3ae9ca9a),
	.w8(32'hbc194dca),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02e59d),
	.w1(32'hbb9639d8),
	.w2(32'hbc0e2ec2),
	.w3(32'hbc346527),
	.w4(32'hbc1f3784),
	.w5(32'hbb9c615d),
	.w6(32'h3ba1fd8f),
	.w7(32'hbbe7fb63),
	.w8(32'hbbc92697),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa84c75),
	.w1(32'hbbc84813),
	.w2(32'h3b7a31aa),
	.w3(32'h3b97c9b0),
	.w4(32'h3a9f5553),
	.w5(32'h3a82845b),
	.w6(32'hbc1dd729),
	.w7(32'h3b344884),
	.w8(32'h3a8b882d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule