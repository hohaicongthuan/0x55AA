module layer_10_featuremap_419(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3904),
	.w1(32'h3b4cc3f7),
	.w2(32'h3a53488a),
	.w3(32'h3bba6a2a),
	.w4(32'h39f38657),
	.w5(32'hbb9bd845),
	.w6(32'hbc00eb04),
	.w7(32'h3b23ac95),
	.w8(32'h3b868fd6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ad46),
	.w1(32'hbc04547a),
	.w2(32'hbb84cb6b),
	.w3(32'h3b3f347a),
	.w4(32'hbbce5264),
	.w5(32'hbb5b04ae),
	.w6(32'h3c01f412),
	.w7(32'hbc055590),
	.w8(32'hbac315b2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a96c),
	.w1(32'h3bc6f648),
	.w2(32'h3b2eee29),
	.w3(32'hbbcb5f90),
	.w4(32'hbb95d2e4),
	.w5(32'hbac2d33a),
	.w6(32'hbc07cb45),
	.w7(32'h3ad230ee),
	.w8(32'h3bdd8e8f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3bb4b),
	.w1(32'h3a1c6407),
	.w2(32'h3b0eb0f4),
	.w3(32'h3b2b5eb2),
	.w4(32'hbb24664f),
	.w5(32'hbc0fd561),
	.w6(32'h39bb75ad),
	.w7(32'hbb8dcf24),
	.w8(32'hb9ab47c6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a930),
	.w1(32'h39a5b302),
	.w2(32'h3afccb8e),
	.w3(32'hbb8cb492),
	.w4(32'h39020420),
	.w5(32'h3aba67c3),
	.w6(32'h3c11e8ca),
	.w7(32'hbaf17cf7),
	.w8(32'h385fefbe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855375),
	.w1(32'hb9b24d02),
	.w2(32'h3b8071d6),
	.w3(32'hbb58aefc),
	.w4(32'h3b29d66b),
	.w5(32'hb9a85a3e),
	.w6(32'hbb17d278),
	.w7(32'h3b007ab4),
	.w8(32'h3c27cbc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1718c),
	.w1(32'hb9099568),
	.w2(32'hbb94e8fa),
	.w3(32'h3b6314b4),
	.w4(32'hbac4c04c),
	.w5(32'h3cd60f10),
	.w6(32'hba8923f1),
	.w7(32'h3bc8aa90),
	.w8(32'hba9a2d55),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b3647),
	.w1(32'h3bb9bb18),
	.w2(32'h3b1d56be),
	.w3(32'h3b66fc20),
	.w4(32'hb976a6fc),
	.w5(32'hbb170002),
	.w6(32'hbaeb23f2),
	.w7(32'h3b81c396),
	.w8(32'h3ba1b390),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a269c95),
	.w1(32'h378752ce),
	.w2(32'hbb139e7e),
	.w3(32'h3af7a204),
	.w4(32'hbb2a3379),
	.w5(32'h3bc8dc4a),
	.w6(32'h3b632fa8),
	.w7(32'hbad780e0),
	.w8(32'h3bb3c101),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5ca3c),
	.w1(32'h3bbd1c04),
	.w2(32'h3c1828e7),
	.w3(32'h3c28c993),
	.w4(32'h3af8f436),
	.w5(32'h38254c4a),
	.w6(32'h3b2ffc9e),
	.w7(32'h3aa9fbaa),
	.w8(32'h3b785ef1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c19f7c),
	.w1(32'hbb8caa87),
	.w2(32'hbae9fa3d),
	.w3(32'hb9a4b054),
	.w4(32'hb9f69b82),
	.w5(32'h3ad9bee3),
	.w6(32'h3b79b81b),
	.w7(32'h39900974),
	.w8(32'hbb884418),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa1f5c),
	.w1(32'hba8a5eaf),
	.w2(32'hbad8572a),
	.w3(32'h3b5431be),
	.w4(32'hbb520289),
	.w5(32'hbc1ce4db),
	.w6(32'hbb496cee),
	.w7(32'hbb13764f),
	.w8(32'hbb858049),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c0e1),
	.w1(32'hbbbcd968),
	.w2(32'h3b9eb7c2),
	.w3(32'h3b5dd87d),
	.w4(32'h3a874ac8),
	.w5(32'h3c19f579),
	.w6(32'h3b5a4d46),
	.w7(32'h381d68fe),
	.w8(32'h3c3901e1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f9a5),
	.w1(32'hbb9e96ce),
	.w2(32'h3b30e633),
	.w3(32'h3badf3d9),
	.w4(32'h3ab071d9),
	.w5(32'h39fc3d75),
	.w6(32'hbac111f5),
	.w7(32'h3b037243),
	.w8(32'h3b0a7825),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b7d0c),
	.w1(32'hbb125a96),
	.w2(32'hbb18e8ec),
	.w3(32'h3b5baeb3),
	.w4(32'hbb6ef0bd),
	.w5(32'hbb9189bb),
	.w6(32'h3b9ed47c),
	.w7(32'hb9a7e86e),
	.w8(32'hbad39bfc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84de98),
	.w1(32'h3b0ea731),
	.w2(32'h3b382dd4),
	.w3(32'hbc24f744),
	.w4(32'hbb0b91b4),
	.w5(32'hba54d345),
	.w6(32'h395ca068),
	.w7(32'hbba487ed),
	.w8(32'hbb96c88c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eec05),
	.w1(32'hb986b8bd),
	.w2(32'hbb561394),
	.w3(32'hbbf1be44),
	.w4(32'hb9cccb0c),
	.w5(32'hb93364df),
	.w6(32'hbbebd900),
	.w7(32'hbb8b1d63),
	.w8(32'hbb892a46),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1cb27),
	.w1(32'h3baac47b),
	.w2(32'h3bff0762),
	.w3(32'hbadf32b2),
	.w4(32'h3ac391b4),
	.w5(32'h3a18f4aa),
	.w6(32'h3926d3c5),
	.w7(32'h3baa4441),
	.w8(32'h3b8ba209),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7750ff),
	.w1(32'hbaca51d2),
	.w2(32'hbb8aad65),
	.w3(32'hbaa3363c),
	.w4(32'hbb80d3dc),
	.w5(32'h3b23f198),
	.w6(32'h3bd98af8),
	.w7(32'hbb30e5fc),
	.w8(32'h3b6dace9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa278bf),
	.w1(32'h3c20dcf1),
	.w2(32'h39025ed5),
	.w3(32'h3b85cdae),
	.w4(32'hbb2d13f1),
	.w5(32'hbb68cad9),
	.w6(32'hbaa9c92b),
	.w7(32'h3b498c09),
	.w8(32'h3b35e60b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17435c),
	.w1(32'h3bb5dc23),
	.w2(32'h3b5efd64),
	.w3(32'h3bae2b32),
	.w4(32'h3bbc6d82),
	.w5(32'hbb93286d),
	.w6(32'h3c1877f3),
	.w7(32'h3b466c2e),
	.w8(32'h3b86c245),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10710),
	.w1(32'h3b72c5f6),
	.w2(32'h3a1b0e71),
	.w3(32'h3ac057b7),
	.w4(32'h3b1bde37),
	.w5(32'hbb75d276),
	.w6(32'hba84491d),
	.w7(32'h3b49deba),
	.w8(32'h3b6a4af1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3dae),
	.w1(32'hbaac44b6),
	.w2(32'h3b346378),
	.w3(32'h3ae9dcda),
	.w4(32'hbb282450),
	.w5(32'h38eb298a),
	.w6(32'hba04f922),
	.w7(32'h3bbfd921),
	.w8(32'h3b89d118),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cc0e8),
	.w1(32'h3bb51a5e),
	.w2(32'h3b246907),
	.w3(32'h3b80c168),
	.w4(32'hbafb93d9),
	.w5(32'hbb40e5d4),
	.w6(32'h3bd549b1),
	.w7(32'h3b02179e),
	.w8(32'hbadc5866),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3f7e),
	.w1(32'hbb13eaed),
	.w2(32'hbc211a5e),
	.w3(32'h3a93a4bf),
	.w4(32'hbbc71614),
	.w5(32'hbbcc4f22),
	.w6(32'h3b04140d),
	.w7(32'hbb11093e),
	.w8(32'hbbeb7d09),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ff703),
	.w1(32'h395a1322),
	.w2(32'h3b084e42),
	.w3(32'hbbadb83f),
	.w4(32'h3b1fe23b),
	.w5(32'h3c346789),
	.w6(32'hbc1190f1),
	.w7(32'h3b74d8a8),
	.w8(32'h3b1c1361),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69c757),
	.w1(32'h373ef1d4),
	.w2(32'hbbf2b396),
	.w3(32'h3b12ddeb),
	.w4(32'h3b318d54),
	.w5(32'h3be324fe),
	.w6(32'hbb035589),
	.w7(32'hbb709658),
	.w8(32'hbac43035),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278e0e),
	.w1(32'h3b1ad37b),
	.w2(32'h39b9f8b9),
	.w3(32'hbac628db),
	.w4(32'h3ac28eed),
	.w5(32'h3b97561a),
	.w6(32'hbb9bf4d2),
	.w7(32'h3b0f09a4),
	.w8(32'h39b0d572),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0919f8),
	.w1(32'h3af2d5ba),
	.w2(32'hbb8e6b20),
	.w3(32'hb89ffea7),
	.w4(32'hbc296214),
	.w5(32'h3bfc7b9f),
	.w6(32'hba00ae9f),
	.w7(32'hbb09da17),
	.w8(32'hba7aaf1e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e83cf),
	.w1(32'h39459b34),
	.w2(32'h3b5d5662),
	.w3(32'h3b108151),
	.w4(32'h3b29cdab),
	.w5(32'hbc25633b),
	.w6(32'hbb0c92ee),
	.w7(32'h3b4067e6),
	.w8(32'hbaad2d58),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2921fe),
	.w1(32'hb955c238),
	.w2(32'hbb25bd0b),
	.w3(32'h3a9d1b45),
	.w4(32'hbbc647ac),
	.w5(32'hbb044abc),
	.w6(32'h3b859348),
	.w7(32'hbabd2fd5),
	.w8(32'hba8db618),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7ddae),
	.w1(32'h3a791995),
	.w2(32'hb93ffbac),
	.w3(32'hbb6a78f5),
	.w4(32'h3b7905ff),
	.w5(32'hbc00aefa),
	.w6(32'h3b8548c4),
	.w7(32'h39848ac6),
	.w8(32'h389260f5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe9a79),
	.w1(32'hb9b0b8c7),
	.w2(32'hbaacf116),
	.w3(32'hb97aba78),
	.w4(32'hbb4cb562),
	.w5(32'h3bd98dc5),
	.w6(32'h3bd97e57),
	.w7(32'hbadfc693),
	.w8(32'hba330cf0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40384),
	.w1(32'hba253d15),
	.w2(32'hba77590f),
	.w3(32'h3be32a72),
	.w4(32'hba90cd47),
	.w5(32'h3c778a61),
	.w6(32'h3ac84dd0),
	.w7(32'h3b38d1ea),
	.w8(32'hbb4e351d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac336b0),
	.w1(32'h3aa7cb8c),
	.w2(32'h3a69134b),
	.w3(32'h3b138101),
	.w4(32'h3bd22138),
	.w5(32'hbc31858f),
	.w6(32'h3ac0ee5c),
	.w7(32'hbb8e6871),
	.w8(32'hbb7bbbac),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1772),
	.w1(32'hba5f0732),
	.w2(32'h3bcf6765),
	.w3(32'hbbc75c05),
	.w4(32'hbb644fa3),
	.w5(32'hba882891),
	.w6(32'h3aa3c12c),
	.w7(32'hbb824774),
	.w8(32'h3b8d984f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a13de),
	.w1(32'hbb022bc4),
	.w2(32'hbb97ecc7),
	.w3(32'h3ba1bdd4),
	.w4(32'h3b36b3bc),
	.w5(32'h3c26e2c0),
	.w6(32'h3bdb9d71),
	.w7(32'h37b3e1a0),
	.w8(32'h3a286ebb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3a28d),
	.w1(32'hbb85920e),
	.w2(32'hbbe26e94),
	.w3(32'h3c2a3edd),
	.w4(32'hbb56fe04),
	.w5(32'hbc5a5823),
	.w6(32'h3ab1fad0),
	.w7(32'hbc031fa0),
	.w8(32'hbbb618c3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44d64f),
	.w1(32'hbb2603b7),
	.w2(32'hbbe7200d),
	.w3(32'h3a87c197),
	.w4(32'hbb94c1b6),
	.w5(32'hbbbbe7aa),
	.w6(32'hba9c811f),
	.w7(32'hbbb51f63),
	.w8(32'hbbc9df4a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef2721),
	.w1(32'hbae699b2),
	.w2(32'hba93a9b2),
	.w3(32'h3ae0d501),
	.w4(32'hbaf37ae8),
	.w5(32'hbb11b3d5),
	.w6(32'h3b3e61f6),
	.w7(32'hbb787ae8),
	.w8(32'hb9f148f0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41660a),
	.w1(32'hbbca8921),
	.w2(32'h3b6ad50f),
	.w3(32'hbad260d5),
	.w4(32'hbb06e701),
	.w5(32'h3a7c5773),
	.w6(32'h3bb41f8b),
	.w7(32'hbbab8fd7),
	.w8(32'hbb747628),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28431c),
	.w1(32'hbb41f0cf),
	.w2(32'hbb42b3a3),
	.w3(32'hbb23825f),
	.w4(32'hba824a00),
	.w5(32'h3c0e19d1),
	.w6(32'h3b0bf90d),
	.w7(32'hb9e6a041),
	.w8(32'hba966597),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb373e1),
	.w1(32'h3b608f84),
	.w2(32'h3bb112f8),
	.w3(32'h3b0c59af),
	.w4(32'h3bd4f30b),
	.w5(32'h3a070fd6),
	.w6(32'hbbc9422c),
	.w7(32'h3abd14fa),
	.w8(32'h3b8d7014),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f6589),
	.w1(32'h3c0cb6e0),
	.w2(32'h3b846098),
	.w3(32'h3ba600c9),
	.w4(32'h3b438aff),
	.w5(32'hbc093366),
	.w6(32'h3c4cec4a),
	.w7(32'h3b5e7b07),
	.w8(32'hbb90f232),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68fb4f),
	.w1(32'hba9da567),
	.w2(32'h3a285bb4),
	.w3(32'h3b16bb78),
	.w4(32'h3b18e496),
	.w5(32'h3cb0aef4),
	.w6(32'h3c045bb7),
	.w7(32'h3b8827d3),
	.w8(32'h3b1079ac),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1012e8),
	.w1(32'hba89f06e),
	.w2(32'h3b0053df),
	.w3(32'h3be80d72),
	.w4(32'hbb227792),
	.w5(32'hbaedd613),
	.w6(32'hbb0c185e),
	.w7(32'hb71445ee),
	.w8(32'hbc0f9885),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f5fab),
	.w1(32'hbb4468ea),
	.w2(32'hba4c7034),
	.w3(32'hbadaf0ee),
	.w4(32'h3b3a6438),
	.w5(32'h3c21ee8f),
	.w6(32'h3a97b14a),
	.w7(32'h392e226a),
	.w8(32'h3b30b43f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9db2df),
	.w1(32'h3b1d7245),
	.w2(32'hbac02d6e),
	.w3(32'h3b4da414),
	.w4(32'hbb37d3f1),
	.w5(32'h3ba05fb4),
	.w6(32'hb9add966),
	.w7(32'h39c440fb),
	.w8(32'h3b0c1d5b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c86d5),
	.w1(32'h3ba03268),
	.w2(32'h3b19dbf6),
	.w3(32'hbadac793),
	.w4(32'h3b9a45ef),
	.w5(32'hbb2898f2),
	.w6(32'h3a504fc9),
	.w7(32'hbb6e9849),
	.w8(32'hbbb978ed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4ab23),
	.w1(32'h3c0e4ca9),
	.w2(32'h3c2daabb),
	.w3(32'h3ab8747f),
	.w4(32'h3bc2feca),
	.w5(32'hbc013195),
	.w6(32'h3a9eaa01),
	.w7(32'hba993715),
	.w8(32'hbb45349a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75fca9),
	.w1(32'hbb931571),
	.w2(32'hb9879cd9),
	.w3(32'h39300479),
	.w4(32'hbbe48474),
	.w5(32'h3b39b030),
	.w6(32'h3acd53b4),
	.w7(32'hbbf64a7b),
	.w8(32'h3b5aeb29),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf078b),
	.w1(32'h3a69dee9),
	.w2(32'hbba40925),
	.w3(32'h3ae8a1f1),
	.w4(32'hbb13ab32),
	.w5(32'hb9b0e698),
	.w6(32'hba9e3cb7),
	.w7(32'h38c44ad0),
	.w8(32'hbaaa18e4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0d08),
	.w1(32'hbb09d439),
	.w2(32'hbb7ee874),
	.w3(32'hbb98028f),
	.w4(32'hbafb6140),
	.w5(32'h3b06b2f8),
	.w6(32'h3a46a44e),
	.w7(32'h3abc8b3e),
	.w8(32'hbabf040b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe031d),
	.w1(32'hbb017a62),
	.w2(32'hbb0be815),
	.w3(32'h3af4b119),
	.w4(32'hbbbc76b9),
	.w5(32'hbbafd737),
	.w6(32'h3ad958af),
	.w7(32'hbaf5ccf9),
	.w8(32'hbb0d14ed),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f385f),
	.w1(32'h3b00028f),
	.w2(32'hbae3b602),
	.w3(32'hbaf14c9f),
	.w4(32'h3ad7d4b6),
	.w5(32'hbb2df621),
	.w6(32'hbab438ee),
	.w7(32'hbb5d6c72),
	.w8(32'h3b0d9fed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ddbb1),
	.w1(32'hba5a2047),
	.w2(32'hbabd0563),
	.w3(32'hba7e8cdc),
	.w4(32'hbb319147),
	.w5(32'hbbd2ed11),
	.w6(32'h3b93f222),
	.w7(32'h3a8f155d),
	.w8(32'h3b20b5e4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf05ccb),
	.w1(32'hb88bb07a),
	.w2(32'hb9885a2d),
	.w3(32'hb9625864),
	.w4(32'hba81b1a0),
	.w5(32'h3b0fac1e),
	.w6(32'hbb2500ce),
	.w7(32'hba6887ad),
	.w8(32'hba888e4d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4fcb6),
	.w1(32'h3b9a9266),
	.w2(32'h3bd2149e),
	.w3(32'h3b524f66),
	.w4(32'h3b116eb0),
	.w5(32'h3b6fa25d),
	.w6(32'hbab0c37b),
	.w7(32'h39a85b52),
	.w8(32'h3b59cc4d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3e11f),
	.w1(32'h3b677538),
	.w2(32'hbb3d657f),
	.w3(32'hbb84694f),
	.w4(32'h3abca107),
	.w5(32'h3b3a00c6),
	.w6(32'hba965055),
	.w7(32'h3b6add88),
	.w8(32'h3c46525d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bc63f),
	.w1(32'h3b3942c6),
	.w2(32'h3ac113aa),
	.w3(32'h3b6e464b),
	.w4(32'h3c5fbdff),
	.w5(32'h3b9677c6),
	.w6(32'h3aec6c82),
	.w7(32'hba3b3f53),
	.w8(32'h3b9ceab0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5920),
	.w1(32'h3aae7383),
	.w2(32'h383a6799),
	.w3(32'hbbb230ff),
	.w4(32'h3c15bb27),
	.w5(32'h3cd90cde),
	.w6(32'hbad145bb),
	.w7(32'h3bcce2db),
	.w8(32'h3bc17d26),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95124a),
	.w1(32'h3b815ac9),
	.w2(32'hba230cac),
	.w3(32'h3c291d4c),
	.w4(32'h37f6e6af),
	.w5(32'hb75f9c86),
	.w6(32'hbb0139bf),
	.w7(32'hba893b98),
	.w8(32'hbb09e497),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb834e8da),
	.w1(32'h3bfe168d),
	.w2(32'h3ba7319c),
	.w3(32'hbb70c31b),
	.w4(32'h3c08d8bb),
	.w5(32'hba7c85be),
	.w6(32'h3acc91d0),
	.w7(32'h3b11fcef),
	.w8(32'h3ac95af9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a460f),
	.w1(32'hb9ce6abf),
	.w2(32'h3b35a4bf),
	.w3(32'hbb17439c),
	.w4(32'h394e5907),
	.w5(32'h3a944964),
	.w6(32'h3b743723),
	.w7(32'hba072ded),
	.w8(32'h3bdf8c02),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6912),
	.w1(32'h3b59e175),
	.w2(32'h3beb0247),
	.w3(32'h3be2ea72),
	.w4(32'h3b5ede6b),
	.w5(32'hbae81b12),
	.w6(32'h3b85df7c),
	.w7(32'h3a0d8f93),
	.w8(32'h3af28363),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2f12f),
	.w1(32'h3b39f312),
	.w2(32'hbc0a1383),
	.w3(32'h3ba18655),
	.w4(32'h3a400b89),
	.w5(32'h3b9c6ba8),
	.w6(32'h3bf81a06),
	.w7(32'h3b0edc66),
	.w8(32'hbb987b95),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118971),
	.w1(32'hbc15aa1a),
	.w2(32'hbb925904),
	.w3(32'h3b22ab84),
	.w4(32'hbbf275ac),
	.w5(32'hbaa911d4),
	.w6(32'hbb846ced),
	.w7(32'h3b50e034),
	.w8(32'h3bdc165a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b802c4c),
	.w1(32'h3a25aee3),
	.w2(32'h3b863ea5),
	.w3(32'h3c1c88ee),
	.w4(32'hbbcca5dd),
	.w5(32'h3a878568),
	.w6(32'h3bbf4a12),
	.w7(32'hba989bb7),
	.w8(32'h3b308d95),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f3c0f),
	.w1(32'hbaff4b46),
	.w2(32'hbb1116ef),
	.w3(32'hbb2dc834),
	.w4(32'hbc3327a4),
	.w5(32'hbadf151b),
	.w6(32'h3b937f47),
	.w7(32'hbc1b00a0),
	.w8(32'hbb83b571),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa26462),
	.w1(32'hbc26b6b6),
	.w2(32'hbc053c62),
	.w3(32'hbb0c1a6e),
	.w4(32'hbba626dc),
	.w5(32'hbb12c996),
	.w6(32'hba8ae34d),
	.w7(32'hbbac3498),
	.w8(32'hbb7aee63),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00fed),
	.w1(32'hbbae35b8),
	.w2(32'hbb1ae16a),
	.w3(32'hbb2183c0),
	.w4(32'hbb78be6a),
	.w5(32'hbac6bd3b),
	.w6(32'hbba7bb66),
	.w7(32'hbab95afa),
	.w8(32'hba7d7e59),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e38cb5),
	.w1(32'h3b00a962),
	.w2(32'h3aee8c51),
	.w3(32'h3a063d18),
	.w4(32'h3b0b81af),
	.w5(32'h39770d7e),
	.w6(32'h3a870b13),
	.w7(32'h3954c97a),
	.w8(32'h3b517a70),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4686c),
	.w1(32'h3b01d3c7),
	.w2(32'hbb2da10f),
	.w3(32'h3aea4390),
	.w4(32'h3b49952f),
	.w5(32'hba5edb69),
	.w6(32'h3bc4b4f0),
	.w7(32'h3a9f8d03),
	.w8(32'hb973d9c3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba239121),
	.w1(32'hb8bfcdf1),
	.w2(32'hb9cf7f54),
	.w3(32'hbbd62b84),
	.w4(32'hbaae0a1e),
	.w5(32'h3b358178),
	.w6(32'hbafffcc8),
	.w7(32'h3b42d531),
	.w8(32'h3a8871e9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e222f),
	.w1(32'hb9d0da6d),
	.w2(32'hb98a06a1),
	.w3(32'h39e70efa),
	.w4(32'hbac2656e),
	.w5(32'hb8be4ac6),
	.w6(32'hbb475a80),
	.w7(32'hba957986),
	.w8(32'hb9421975),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59e49),
	.w1(32'hba8cf0c4),
	.w2(32'h3a6a81a5),
	.w3(32'hbb9bcc29),
	.w4(32'hbb60a6d9),
	.w5(32'h3ae62fd9),
	.w6(32'hba169d92),
	.w7(32'hba843a19),
	.w8(32'hb986a544),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65e16),
	.w1(32'hbabf080e),
	.w2(32'h3aae2fdc),
	.w3(32'h3b4f4958),
	.w4(32'h3b2ef0ff),
	.w5(32'h3bc8f2f0),
	.w6(32'hbac16416),
	.w7(32'h39c21a8e),
	.w8(32'h3b9b81f5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18146b),
	.w1(32'hbb80d888),
	.w2(32'hbacc9eb9),
	.w3(32'hbb16f659),
	.w4(32'hbbf81301),
	.w5(32'hbbb5e022),
	.w6(32'h3b20faf6),
	.w7(32'hbba4afeb),
	.w8(32'hbb8e4510),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0658),
	.w1(32'hb9da56f5),
	.w2(32'h3a772b4a),
	.w3(32'hba90d770),
	.w4(32'h3abb0491),
	.w5(32'h39852a9f),
	.w6(32'hbac71822),
	.w7(32'h3a76471c),
	.w8(32'h3a057082),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb138def),
	.w1(32'h3a3d6fb6),
	.w2(32'h397ffd26),
	.w3(32'h3b54402e),
	.w4(32'hbb324f63),
	.w5(32'hb98aa5db),
	.w6(32'h3ab1b78e),
	.w7(32'hbae042ea),
	.w8(32'hbae843c0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58a51f),
	.w1(32'h3c1bbf86),
	.w2(32'h3ba4ffaf),
	.w3(32'hbb9c3e50),
	.w4(32'h3c094e57),
	.w5(32'h3aed1089),
	.w6(32'hbb53b5c3),
	.w7(32'h3c165cfa),
	.w8(32'h3b9cd621),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844213),
	.w1(32'h3a225a16),
	.w2(32'hbb306519),
	.w3(32'h3bb0f3ce),
	.w4(32'hb657b622),
	.w5(32'hbaccd607),
	.w6(32'h3bdd82a9),
	.w7(32'h3b0033a6),
	.w8(32'hb9c599ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dd0a9),
	.w1(32'h3b2c98ff),
	.w2(32'h3b097321),
	.w3(32'hbb9197d2),
	.w4(32'h3afb92d2),
	.w5(32'h3b0fe920),
	.w6(32'hbb3c25e5),
	.w7(32'hbaa35d03),
	.w8(32'hba4ade30),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945a9f),
	.w1(32'hb96d3fbf),
	.w2(32'hbb04bfb3),
	.w3(32'h39cc1d45),
	.w4(32'h3b1a34dd),
	.w5(32'hbab9fb40),
	.w6(32'h3bd0403d),
	.w7(32'h3a108312),
	.w8(32'h3a90b335),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3a52a),
	.w1(32'h37830bb7),
	.w2(32'hbad7962a),
	.w3(32'hba9cac28),
	.w4(32'h3924c566),
	.w5(32'h3a7c51f9),
	.w6(32'h3a4e43ff),
	.w7(32'h3a3e3afe),
	.w8(32'hb7a92021),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a332768),
	.w1(32'hbb0c95f5),
	.w2(32'hbb5df5f3),
	.w3(32'h3a812b64),
	.w4(32'hbbd83a1d),
	.w5(32'hbae549ad),
	.w6(32'h3b772b11),
	.w7(32'hbb486c2c),
	.w8(32'hba957a10),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a946),
	.w1(32'h39f6f0ca),
	.w2(32'hb9deba73),
	.w3(32'hbab9c4fc),
	.w4(32'hbb869366),
	.w5(32'hbb5c9c82),
	.w6(32'hbac706e5),
	.w7(32'hbb67486d),
	.w8(32'h36eb4847),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78a85c),
	.w1(32'hb98e0025),
	.w2(32'hbb687fe4),
	.w3(32'hb9f6a80d),
	.w4(32'h39ff6238),
	.w5(32'h3b2b42d5),
	.w6(32'h3a0758c6),
	.w7(32'h3a8bed3d),
	.w8(32'h3b32b66b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b957d5e),
	.w1(32'hbb763031),
	.w2(32'hba86fdea),
	.w3(32'h3a93f1c2),
	.w4(32'hbadcc094),
	.w5(32'h3adbe481),
	.w6(32'h3b35fd6f),
	.w7(32'hbb269f0e),
	.w8(32'hbaa1a5c8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d99964),
	.w1(32'hbadc193b),
	.w2(32'h39102437),
	.w3(32'hbb08b269),
	.w4(32'hbb2c147c),
	.w5(32'h3b938d56),
	.w6(32'h3a09d717),
	.w7(32'hbb8e98f0),
	.w8(32'h3a146508),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a28a),
	.w1(32'hbbac47f4),
	.w2(32'hbb9d5d1e),
	.w3(32'hba1949e6),
	.w4(32'hbb175fe7),
	.w5(32'hbb4acc82),
	.w6(32'h3a4a32e2),
	.w7(32'hbb8c70f5),
	.w8(32'hbb866e37),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff6b64),
	.w1(32'hbb4f019e),
	.w2(32'hba7668bc),
	.w3(32'h3a2b29e4),
	.w4(32'hbb621e26),
	.w5(32'hbb8b4b3c),
	.w6(32'h3a98b1d6),
	.w7(32'hbb8d74bd),
	.w8(32'hbb5158c4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb761b61),
	.w1(32'h3bd43fc7),
	.w2(32'h3b7f52b4),
	.w3(32'hbc11077e),
	.w4(32'h3b847a13),
	.w5(32'h393a5f06),
	.w6(32'hbbb81ef4),
	.w7(32'hba26d210),
	.w8(32'h3abaa77f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945b5b),
	.w1(32'hba27cc49),
	.w2(32'h3b8ee47e),
	.w3(32'h3b844474),
	.w4(32'hbb2164e1),
	.w5(32'hbb0d2f62),
	.w6(32'h3c30db32),
	.w7(32'hbb1ac418),
	.w8(32'h3a5a335d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfb3a7),
	.w1(32'h3982cc92),
	.w2(32'h3a2c72d8),
	.w3(32'h3b8dbe98),
	.w4(32'hbbd63a54),
	.w5(32'hbbc0cf26),
	.w6(32'hbab86908),
	.w7(32'hbb906b4a),
	.w8(32'hbb6b449e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b668f),
	.w1(32'hb9051816),
	.w2(32'h397d7143),
	.w3(32'hbba1a6da),
	.w4(32'hba46c90b),
	.w5(32'h3bdfb074),
	.w6(32'hbad03b82),
	.w7(32'h3b38b405),
	.w8(32'h3a8a8594),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86eb3f),
	.w1(32'h3b00ab9b),
	.w2(32'hbb74e980),
	.w3(32'hbb01f00b),
	.w4(32'hbacab7b2),
	.w5(32'h3b0531e2),
	.w6(32'hbb99afa3),
	.w7(32'h3b72c26d),
	.w8(32'h3ba21599),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becb0c8),
	.w1(32'h3a54b583),
	.w2(32'h3b8ced30),
	.w3(32'h3bd0eefb),
	.w4(32'hbb1a3f0e),
	.w5(32'h3c10e5cd),
	.w6(32'h3bb2030f),
	.w7(32'hba2dc8c7),
	.w8(32'h3b3f6b50),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ed2bc),
	.w1(32'hbb1d74f5),
	.w2(32'h38f0d8de),
	.w3(32'h3b9ee14c),
	.w4(32'h3b9de08d),
	.w5(32'h3c40d4dc),
	.w6(32'h3b698424),
	.w7(32'h3a267b19),
	.w8(32'hb99629fc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cf614),
	.w1(32'hbb5bf721),
	.w2(32'hbb23875d),
	.w3(32'hbb28bf3c),
	.w4(32'hbb339bb8),
	.w5(32'hbb5ce2c0),
	.w6(32'hbb62b975),
	.w7(32'hbb8ee92c),
	.w8(32'hbb816d76),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b903626),
	.w1(32'h3c0770f9),
	.w2(32'h3b05d94d),
	.w3(32'h3b1b51bc),
	.w4(32'h3b03c581),
	.w5(32'h3b7ce391),
	.w6(32'h3a1ad5c2),
	.w7(32'h3b91762a),
	.w8(32'h3aa72edb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e30b1),
	.w1(32'h3badd298),
	.w2(32'h3bf50b4d),
	.w3(32'h3bf7ad54),
	.w4(32'h3b4f0edd),
	.w5(32'h3c284d66),
	.w6(32'h3b222462),
	.w7(32'h3b465a95),
	.w8(32'h3b79658a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb5ffc),
	.w1(32'h3aca17a5),
	.w2(32'h3a088d3d),
	.w3(32'h3c1a6bd8),
	.w4(32'h3ae14430),
	.w5(32'h3b278316),
	.w6(32'h3bd90d5d),
	.w7(32'hb9bed986),
	.w8(32'hbaac50d4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9ad56),
	.w1(32'hbaae062e),
	.w2(32'hbaee7971),
	.w3(32'h3ad34d7a),
	.w4(32'h39d30858),
	.w5(32'h3b37be25),
	.w6(32'h3b21910e),
	.w7(32'h3b254f6c),
	.w8(32'h3a4639ee),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2736),
	.w1(32'h3b1a45d0),
	.w2(32'h3c129fa8),
	.w3(32'h3be0fc4c),
	.w4(32'hba84c0c7),
	.w5(32'h3aac70b4),
	.w6(32'h3a8b381f),
	.w7(32'h3abef336),
	.w8(32'h3b698cc2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ce9c),
	.w1(32'h3b4c98f9),
	.w2(32'h3baadf69),
	.w3(32'h3b322d66),
	.w4(32'h3ad6ed90),
	.w5(32'h39dd7213),
	.w6(32'h3bde547d),
	.w7(32'h3ad2a9f4),
	.w8(32'h3ab9633d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51c879),
	.w1(32'hb979389b),
	.w2(32'hbaac57f7),
	.w3(32'h3ac28e9c),
	.w4(32'hb994ff0d),
	.w5(32'hba446fc7),
	.w6(32'h3a5aa929),
	.w7(32'h3b68be45),
	.w8(32'h3b6aa91c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdadd3),
	.w1(32'hbaeb7780),
	.w2(32'hbb533841),
	.w3(32'h3ad12dfe),
	.w4(32'hbada4d02),
	.w5(32'hbb620a87),
	.w6(32'h3b6d39bb),
	.w7(32'hbba81d05),
	.w8(32'hbb9710cd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9766ba7),
	.w1(32'h3bbaf2d6),
	.w2(32'h3bc9567f),
	.w3(32'h3b15812e),
	.w4(32'h3b27c5f9),
	.w5(32'h3b9fbccc),
	.w6(32'h3b7213b9),
	.w7(32'h3a4c1da0),
	.w8(32'hbaa280be),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e137f),
	.w1(32'hbb273c79),
	.w2(32'hb9770449),
	.w3(32'h3b75ba85),
	.w4(32'hbbbaf1a0),
	.w5(32'hbb71b24d),
	.w6(32'h3bde2869),
	.w7(32'hbb7b7c29),
	.w8(32'hbac41391),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2209ff),
	.w1(32'hbb9de766),
	.w2(32'hbb435615),
	.w3(32'hbacb8a98),
	.w4(32'hbb9c5512),
	.w5(32'hbac3674f),
	.w6(32'h3b6625a7),
	.w7(32'hbb8c3e23),
	.w8(32'hbb59dd6b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb374159),
	.w1(32'h388c5475),
	.w2(32'h3b72077e),
	.w3(32'hba88bc17),
	.w4(32'hbb9a563c),
	.w5(32'h3b90c5e0),
	.w6(32'hbbac87a5),
	.w7(32'hbb2d3418),
	.w8(32'hba78a25d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf7ab6),
	.w1(32'h3a9ae3d2),
	.w2(32'hbabb0db2),
	.w3(32'h3b2cb708),
	.w4(32'hbb8a9143),
	.w5(32'h3a8320d2),
	.w6(32'h3ba1afb4),
	.w7(32'h3b8a86cc),
	.w8(32'h3a915b7d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d1bef),
	.w1(32'h39e1f67d),
	.w2(32'hbbcd3cf3),
	.w3(32'hbb26de21),
	.w4(32'h3aa430aa),
	.w5(32'hbba7d39d),
	.w6(32'h39bf77df),
	.w7(32'hba9df3f5),
	.w8(32'h3b8cda02),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba445e7f),
	.w1(32'h3991afb6),
	.w2(32'h3b9a05f1),
	.w3(32'h3ba594e8),
	.w4(32'h3a8f3eec),
	.w5(32'hbb4e4b6a),
	.w6(32'hb9cae307),
	.w7(32'hbad67cf7),
	.w8(32'hbaa15534),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52a2b1),
	.w1(32'hb9714433),
	.w2(32'h36897dee),
	.w3(32'h3b7ce3c3),
	.w4(32'hbabd500f),
	.w5(32'h39e2aeb4),
	.w6(32'h3b92d71b),
	.w7(32'hb8bb0a7f),
	.w8(32'h39fb5fed),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af90719),
	.w1(32'h3a5d0438),
	.w2(32'hba0bd627),
	.w3(32'h3a5b0ee3),
	.w4(32'hb84dce29),
	.w5(32'hba60c38b),
	.w6(32'h3a3c3e7d),
	.w7(32'h3b17a648),
	.w8(32'h3ac9bfe2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73a87d),
	.w1(32'h3b37244c),
	.w2(32'h3ad15a57),
	.w3(32'h3b879b25),
	.w4(32'h3aefa36d),
	.w5(32'h3a2e7249),
	.w6(32'h3b06799b),
	.w7(32'h3a32a125),
	.w8(32'h3a955aac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d6192),
	.w1(32'hb8e45db1),
	.w2(32'hbb1c8b1b),
	.w3(32'h3b9ae0ba),
	.w4(32'hba71122d),
	.w5(32'h3b76a066),
	.w6(32'h3baede33),
	.w7(32'h3aab19cd),
	.w8(32'h3b29226d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d289c),
	.w1(32'h3b70d729),
	.w2(32'h3b93ffbe),
	.w3(32'h3b19b45d),
	.w4(32'h3a8af0df),
	.w5(32'hbadfbd5d),
	.w6(32'h3a77bf79),
	.w7(32'hbb0b3487),
	.w8(32'hbb7943f3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88045e),
	.w1(32'hbbbb5c2f),
	.w2(32'hbbccda10),
	.w3(32'h3b024c88),
	.w4(32'h398331c1),
	.w5(32'hb923a6f4),
	.w6(32'h3b2928a9),
	.w7(32'hba651120),
	.w8(32'hbb025e54),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1206),
	.w1(32'hbbd9f0bb),
	.w2(32'hbb926e46),
	.w3(32'hbbb6f27b),
	.w4(32'h3b130a27),
	.w5(32'hba4ad4d8),
	.w6(32'hbb3a5019),
	.w7(32'h3b7e698a),
	.w8(32'hbabb14f0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40a5b0),
	.w1(32'h3ae02ed9),
	.w2(32'hbb0fe80e),
	.w3(32'h3a61a8d3),
	.w4(32'hbafc6714),
	.w5(32'hb980e7e3),
	.w6(32'hba83ea69),
	.w7(32'h37d2445e),
	.w8(32'h396ee78a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53ae64),
	.w1(32'hba46753b),
	.w2(32'h3b32c56a),
	.w3(32'h3a283748),
	.w4(32'hbaf1be36),
	.w5(32'h3bd5eac4),
	.w6(32'h3adb8145),
	.w7(32'h3ab22e2f),
	.w8(32'hbaf4fd3d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4fd68),
	.w1(32'h3b2cebaf),
	.w2(32'h3b70f6a4),
	.w3(32'h3a8441e4),
	.w4(32'h3a8d589c),
	.w5(32'h3b667c1b),
	.w6(32'hba890b10),
	.w7(32'h3b051294),
	.w8(32'h3ac62cc4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a107b1e),
	.w1(32'hbb927810),
	.w2(32'hbb52ed12),
	.w3(32'h3aa40f37),
	.w4(32'hbaefd46b),
	.w5(32'hbb45d0d3),
	.w6(32'h3b8b6366),
	.w7(32'hbb0601d8),
	.w8(32'h397a4b0b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f510),
	.w1(32'hbb8dcb7f),
	.w2(32'hbb1d8d37),
	.w3(32'hbb6b0a8e),
	.w4(32'hbb909f0f),
	.w5(32'hbbb1a9cc),
	.w6(32'hbb6672ff),
	.w7(32'hbb7674b2),
	.w8(32'hbbd9d288),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d13ba4),
	.w1(32'h3b23fdee),
	.w2(32'h3b6c3b1c),
	.w3(32'hbbbe3b3a),
	.w4(32'hb9312766),
	.w5(32'h3b51268b),
	.w6(32'hbbaddcc4),
	.w7(32'hba1bd3b3),
	.w8(32'h3acfa8e4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7912c1),
	.w1(32'h3acfb45b),
	.w2(32'h3a493bdb),
	.w3(32'h3ac6e146),
	.w4(32'h39811a91),
	.w5(32'hb9ff2ae1),
	.w6(32'h3b8e9b4f),
	.w7(32'hba983738),
	.w8(32'hbac10dfd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967f4f9),
	.w1(32'hbb222887),
	.w2(32'hbab2c447),
	.w3(32'hbbcaff6a),
	.w4(32'hbb8c4824),
	.w5(32'hbac39399),
	.w6(32'hbb55b8a5),
	.w7(32'hbb79f278),
	.w8(32'hba1a0af7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71c6de),
	.w1(32'h3adaccec),
	.w2(32'h3b8051c6),
	.w3(32'h3b214292),
	.w4(32'hbb56172a),
	.w5(32'h3bb25112),
	.w6(32'h3a7ad155),
	.w7(32'hbac0409b),
	.w8(32'h3b775dc0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7931),
	.w1(32'hbaa87433),
	.w2(32'hb963c951),
	.w3(32'h3bcb5e38),
	.w4(32'h3b5449b1),
	.w5(32'hbb110ec3),
	.w6(32'h3a8a4ab2),
	.w7(32'hbb4a7fa2),
	.w8(32'hb862b979),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cee75),
	.w1(32'h3aba64ee),
	.w2(32'h3ac454f3),
	.w3(32'h3b5145ec),
	.w4(32'h39a727f0),
	.w5(32'h3beadda4),
	.w6(32'h3a293c9b),
	.w7(32'h38a276bc),
	.w8(32'hb98d86b0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bbec9),
	.w1(32'h3b69fb09),
	.w2(32'h3bd8e392),
	.w3(32'h3a724234),
	.w4(32'h3ad9c316),
	.w5(32'hba60e4ba),
	.w6(32'h3a9df5cd),
	.w7(32'hba1398f4),
	.w8(32'hb9b7f9ed),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2961),
	.w1(32'h3aa16d97),
	.w2(32'h3a08e103),
	.w3(32'h3bd52261),
	.w4(32'hbb6c6d9c),
	.w5(32'h3b868137),
	.w6(32'h3b8f1df2),
	.w7(32'h3b9e2ded),
	.w8(32'h3b9b0194),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84943a),
	.w1(32'hbb41f50f),
	.w2(32'h3b5071f6),
	.w3(32'h3ae2f6ed),
	.w4(32'hbabb0b99),
	.w5(32'h3a7ede93),
	.w6(32'hbac673ed),
	.w7(32'hbaca3600),
	.w8(32'hba7164ec),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc12267),
	.w1(32'hbb315b50),
	.w2(32'h3aa96038),
	.w3(32'h3b8bd57f),
	.w4(32'hbb7f1754),
	.w5(32'h3b860188),
	.w6(32'hbbbd2e93),
	.w7(32'h38e84d81),
	.w8(32'h3abbf47a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5e6b),
	.w1(32'h3b0613d9),
	.w2(32'h3b66ef88),
	.w3(32'h3c0d7df0),
	.w4(32'h3b591295),
	.w5(32'h3af2fe1f),
	.w6(32'h3aa0520b),
	.w7(32'h3b46b2ce),
	.w8(32'h391a2c9e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cba0e),
	.w1(32'h3a15beb4),
	.w2(32'hbb026e4d),
	.w3(32'h3a108874),
	.w4(32'hbb0e01e2),
	.w5(32'hbaa1d2c8),
	.w6(32'h3b2a9225),
	.w7(32'hb9cff58f),
	.w8(32'hbb062308),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0343),
	.w1(32'h3b80a806),
	.w2(32'h3b151473),
	.w3(32'h3a728151),
	.w4(32'h3b757974),
	.w5(32'h3b51f6a5),
	.w6(32'h39f110e3),
	.w7(32'hb9f030da),
	.w8(32'hb8db2d42),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad107da),
	.w1(32'hbba7c4f0),
	.w2(32'hbb2f9980),
	.w3(32'hbab1b876),
	.w4(32'hbb68ae4b),
	.w5(32'hbb798850),
	.w6(32'h3a9cce00),
	.w7(32'h38a06827),
	.w8(32'hba69a813),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5763),
	.w1(32'h3b29691b),
	.w2(32'h3b0ee21b),
	.w3(32'hbb1173d0),
	.w4(32'h3aa2d502),
	.w5(32'h3baaed99),
	.w6(32'hbad20c74),
	.w7(32'hbb6b3ee0),
	.w8(32'hba7c4a34),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484685),
	.w1(32'hbb588036),
	.w2(32'hbac37a7e),
	.w3(32'h3b741f0b),
	.w4(32'hbb92dfad),
	.w5(32'h399fa63c),
	.w6(32'h3bab478f),
	.w7(32'hbaa84fab),
	.w8(32'hbb0f2589),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3563f8),
	.w1(32'h3a2e81d1),
	.w2(32'hbadd5b3b),
	.w3(32'hbb033b5c),
	.w4(32'h3a53d3a2),
	.w5(32'hbb0bbc5a),
	.w6(32'hbb2ff672),
	.w7(32'hbb0e9246),
	.w8(32'hbb18d314),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa951c3),
	.w1(32'hbaf2a634),
	.w2(32'h3a20c7b2),
	.w3(32'hbb037b8f),
	.w4(32'h3ab129d1),
	.w5(32'h3b995067),
	.w6(32'hba85249f),
	.w7(32'h3b2802f1),
	.w8(32'h3b48deb2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a260602),
	.w1(32'h3bbbf46e),
	.w2(32'h3b86f9de),
	.w3(32'h3b50ece2),
	.w4(32'h3c0840cf),
	.w5(32'h3b5f7c51),
	.w6(32'h3b82faa2),
	.w7(32'h3b1feb00),
	.w8(32'h3b854769),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c6d9),
	.w1(32'h3b1dee60),
	.w2(32'h3a72a39d),
	.w3(32'h3b72cbbd),
	.w4(32'h3a54f938),
	.w5(32'h3b8ac38b),
	.w6(32'h3b6d5189),
	.w7(32'h3b621f42),
	.w8(32'h3b534f52),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbadc4b),
	.w1(32'hbbf17f40),
	.w2(32'hbabf8add),
	.w3(32'h3be6990d),
	.w4(32'hbb8908e3),
	.w5(32'hba8674e7),
	.w6(32'h3b9dda0d),
	.w7(32'hbb487a8b),
	.w8(32'hbb07cf51),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2675),
	.w1(32'hbb21418e),
	.w2(32'hbb2e8bf2),
	.w3(32'hbb6705fa),
	.w4(32'hba794f0a),
	.w5(32'hbb760a18),
	.w6(32'hbb7b9fcc),
	.w7(32'hbb5041df),
	.w8(32'hbae61e5d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fd161),
	.w1(32'hbb216b46),
	.w2(32'hbaec1102),
	.w3(32'h3bd1ba21),
	.w4(32'h39c4bf17),
	.w5(32'hbb0f2cf1),
	.w6(32'h3ae85c27),
	.w7(32'hbaa1aca5),
	.w8(32'hba5f783b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe833f5),
	.w1(32'hba9dc9bd),
	.w2(32'h3b4bdac6),
	.w3(32'hbbb353fb),
	.w4(32'h3b05ffbc),
	.w5(32'hbab871f4),
	.w6(32'hbb76bcb0),
	.w7(32'hba78a0a0),
	.w8(32'h3981f3c4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39885e72),
	.w1(32'hbab23ded),
	.w2(32'hb9776b9f),
	.w3(32'hba9b5be3),
	.w4(32'hbb004e0e),
	.w5(32'hbb524aff),
	.w6(32'hbb028362),
	.w7(32'hbb49801d),
	.w8(32'hbb589c01),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef7c63),
	.w1(32'hbbb71f4a),
	.w2(32'hbb4a8a2e),
	.w3(32'hba45cb73),
	.w4(32'hbb51e3a6),
	.w5(32'hbb14ca5a),
	.w6(32'hba469696),
	.w7(32'hbbc7fc8d),
	.w8(32'hbbc2476b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe13df),
	.w1(32'hbb885874),
	.w2(32'hbbaa97e5),
	.w3(32'hbb8e6a18),
	.w4(32'hbaca1e14),
	.w5(32'hbb62f063),
	.w6(32'hbb99cdd2),
	.w7(32'hbaab34ff),
	.w8(32'hbb639e72),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2516f8),
	.w1(32'h3b4a19b5),
	.w2(32'hbbd1d008),
	.w3(32'hbc1afaf7),
	.w4(32'hbb3f8f68),
	.w5(32'hbb998866),
	.w6(32'hbbf36a77),
	.w7(32'h3ac5c80c),
	.w8(32'h3b92b78f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9c360),
	.w1(32'hba94fa16),
	.w2(32'hbac73122),
	.w3(32'h3b4e8a8f),
	.w4(32'h3b2f3ee9),
	.w5(32'h3960d72e),
	.w6(32'h3b880be6),
	.w7(32'h3a4e98f9),
	.w8(32'hbb0439e7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c13b6),
	.w1(32'hbafef7f5),
	.w2(32'hbb0c7b00),
	.w3(32'h3a475e01),
	.w4(32'hbab2cd2f),
	.w5(32'h3b07bf00),
	.w6(32'hbac52db0),
	.w7(32'hbb4f4dc7),
	.w8(32'h3a70f8a2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239108),
	.w1(32'hb98b69a3),
	.w2(32'h384e8fc2),
	.w3(32'hba4a7300),
	.w4(32'h3a59c287),
	.w5(32'hb898c901),
	.w6(32'h3a8ec93c),
	.w7(32'h38d8d351),
	.w8(32'hb922fd97),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3daef),
	.w1(32'hb9fe708a),
	.w2(32'h3a8d88d9),
	.w3(32'h3b026e1a),
	.w4(32'hbb895349),
	.w5(32'hbb824170),
	.w6(32'h3b19923f),
	.w7(32'hbb08bf29),
	.w8(32'hbad229e5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1e4e3),
	.w1(32'h3b62699f),
	.w2(32'h3b8115cf),
	.w3(32'hbb5c00c6),
	.w4(32'h3a8a4b86),
	.w5(32'h3b22d1c2),
	.w6(32'hbaadc12a),
	.w7(32'hba916109),
	.w8(32'hb74509d4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005a4c),
	.w1(32'hba95a4dc),
	.w2(32'hbb0950b5),
	.w3(32'h3b00e356),
	.w4(32'h3a5524c7),
	.w5(32'h3b802ec8),
	.w6(32'h3b7cbaeb),
	.w7(32'hb93081ac),
	.w8(32'hbb56fbe7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296e98),
	.w1(32'h3b90638f),
	.w2(32'h3bbfcdfe),
	.w3(32'h3a6170fc),
	.w4(32'h3b41d02e),
	.w5(32'h3aea3c2e),
	.w6(32'hbac362b4),
	.w7(32'h3b630f3b),
	.w8(32'h3865c919),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc890bb),
	.w1(32'h3bb494c4),
	.w2(32'h3aff823c),
	.w3(32'hbb10f1fe),
	.w4(32'h3bc9f8db),
	.w5(32'hbb193a3c),
	.w6(32'hb91e0762),
	.w7(32'hbadd079b),
	.w8(32'h3ade31a8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4a0aa),
	.w1(32'hbaf54646),
	.w2(32'hbb96b572),
	.w3(32'hba1b19df),
	.w4(32'h3a9073d2),
	.w5(32'hbba6ccb2),
	.w6(32'h3bb64aab),
	.w7(32'hbb608061),
	.w8(32'hbb2434bd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb434a8c),
	.w1(32'hb9d19693),
	.w2(32'hbb1e5f61),
	.w3(32'hb64f301f),
	.w4(32'hbbab6bc1),
	.w5(32'hb9594798),
	.w6(32'hb9edaf4e),
	.w7(32'hbbb1f1d0),
	.w8(32'hbb23c375),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14690d),
	.w1(32'h3a9f3524),
	.w2(32'h3b794920),
	.w3(32'hbabe2cfc),
	.w4(32'hb908e5f8),
	.w5(32'h3aa3abe2),
	.w6(32'hbb459dff),
	.w7(32'h3aa0fe96),
	.w8(32'h3b653b8d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970ac3a),
	.w1(32'h3b21d1fb),
	.w2(32'h3a488f88),
	.w3(32'h3b728285),
	.w4(32'hbae7e231),
	.w5(32'hbb10c127),
	.w6(32'h3b311745),
	.w7(32'hbb0602de),
	.w8(32'hbb7b8ca4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd644a4),
	.w1(32'hbaedb1a6),
	.w2(32'hbb25aae1),
	.w3(32'h374d099c),
	.w4(32'h3ae158eb),
	.w5(32'hbba6006a),
	.w6(32'h3ae463a9),
	.w7(32'hba00ed3a),
	.w8(32'hbb159005),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d4fe2),
	.w1(32'hba2689b6),
	.w2(32'h38a3c8a1),
	.w3(32'h3af36c90),
	.w4(32'hba386366),
	.w5(32'hba8594b3),
	.w6(32'h3a855ac6),
	.w7(32'hbbb9eb12),
	.w8(32'hbba9f613),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51534f),
	.w1(32'hba4a7096),
	.w2(32'hbb654bfc),
	.w3(32'hba6d19bb),
	.w4(32'hba5aef88),
	.w5(32'hba47b2eb),
	.w6(32'hba8905a2),
	.w7(32'hbb58a084),
	.w8(32'hbb709eca),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b17aae),
	.w1(32'h3819927a),
	.w2(32'h3a6a69b3),
	.w3(32'h3afd4fd7),
	.w4(32'h3a2af85e),
	.w5(32'hb99284a7),
	.w6(32'hb8d81786),
	.w7(32'hbb1aac78),
	.w8(32'h37bb4c78),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bcded),
	.w1(32'h3a867fd8),
	.w2(32'h3956632d),
	.w3(32'hbab962ff),
	.w4(32'h3a53dca2),
	.w5(32'hbb69f4c8),
	.w6(32'hba587bda),
	.w7(32'h39ee2bc5),
	.w8(32'hba794e52),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba309),
	.w1(32'h39560e61),
	.w2(32'hb9d1e457),
	.w3(32'hb81113ee),
	.w4(32'hbafae845),
	.w5(32'h38efae76),
	.w6(32'h3a0aad9f),
	.w7(32'h3adb6457),
	.w8(32'hb9b2a5db),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39f438),
	.w1(32'h3aca7e65),
	.w2(32'h3b1a2cf2),
	.w3(32'h39eda825),
	.w4(32'hb9ca7c19),
	.w5(32'hba742e00),
	.w6(32'hba2e0c53),
	.w7(32'hbb8512ec),
	.w8(32'hb8830e1a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01253),
	.w1(32'hba203ac9),
	.w2(32'h3b1a8c7d),
	.w3(32'h3b472345),
	.w4(32'hbb535114),
	.w5(32'hba4b6132),
	.w6(32'h39c19418),
	.w7(32'hbb5917cd),
	.w8(32'h3b43fd27),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0996e),
	.w1(32'hbb3c0897),
	.w2(32'hbb8c28c5),
	.w3(32'hbb2b7870),
	.w4(32'hbb9be24a),
	.w5(32'hbba60c2b),
	.w6(32'h3b7651d9),
	.w7(32'hbb59e4d1),
	.w8(32'hbb970e1f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf282f),
	.w1(32'hbb88c12e),
	.w2(32'h3a4aa3c2),
	.w3(32'hb9847683),
	.w4(32'h3b1c0ecc),
	.w5(32'h3bc213dc),
	.w6(32'hba607619),
	.w7(32'hba45e539),
	.w8(32'hba410787),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2377d),
	.w1(32'hbac9ca38),
	.w2(32'hba295365),
	.w3(32'h3bff0eb7),
	.w4(32'h3ab83bed),
	.w5(32'hbb7aa755),
	.w6(32'h3b097c9f),
	.w7(32'hbb96e186),
	.w8(32'hbbed675b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48dd1d),
	.w1(32'hbac98e7f),
	.w2(32'hb9d31486),
	.w3(32'h3b061157),
	.w4(32'hbaa9dbda),
	.w5(32'h3adc9463),
	.w6(32'h3b90c154),
	.w7(32'hbb29038c),
	.w8(32'hba84cea6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace1078),
	.w1(32'h3ba2c0a2),
	.w2(32'h3a539763),
	.w3(32'h39fc0631),
	.w4(32'hbaa6321d),
	.w5(32'hbb9850fa),
	.w6(32'hbaed9436),
	.w7(32'h3a0c1433),
	.w8(32'h39c15958),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89df8a),
	.w1(32'hbae48f05),
	.w2(32'h39b29640),
	.w3(32'h3b616cdf),
	.w4(32'hba699256),
	.w5(32'hb9a77c7c),
	.w6(32'h3b6c0cbf),
	.w7(32'hbafe3cd2),
	.w8(32'hbb7219aa),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a2d038),
	.w1(32'h3adb1972),
	.w2(32'h3b22782f),
	.w3(32'h3a2579f7),
	.w4(32'h3b0106bb),
	.w5(32'hba9e4ece),
	.w6(32'hbb8f76be),
	.w7(32'h3b48d240),
	.w8(32'h3b7933f9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3d625),
	.w1(32'hb992e0bf),
	.w2(32'h3a1c3ffb),
	.w3(32'h3bd40601),
	.w4(32'hbb2bc377),
	.w5(32'hba8bed61),
	.w6(32'h3ad91697),
	.w7(32'hbb879a0c),
	.w8(32'hb90169cb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6965),
	.w1(32'hbac8249f),
	.w2(32'hba793db7),
	.w3(32'hbb18a3e4),
	.w4(32'hb9ea1eaa),
	.w5(32'h390a98cc),
	.w6(32'hb89f1a42),
	.w7(32'h39a9c1c7),
	.w8(32'h3b8857b0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0239f0),
	.w1(32'h3b69226f),
	.w2(32'h3a4a5c8d),
	.w3(32'h3acb5dcd),
	.w4(32'h3a0cde2a),
	.w5(32'h3a04d82e),
	.w6(32'hba988ae4),
	.w7(32'h3b4d0608),
	.w8(32'hba2c16fc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d9f83),
	.w1(32'hbaf70a26),
	.w2(32'hbb696bc2),
	.w3(32'hbb29962e),
	.w4(32'hbb1a60cf),
	.w5(32'hbb8528d7),
	.w6(32'hba8d8d30),
	.w7(32'hbb97a9f6),
	.w8(32'hbb890e34),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0bc4),
	.w1(32'hbacbf068),
	.w2(32'h3aaecb13),
	.w3(32'hbb9844ff),
	.w4(32'h3a434f4e),
	.w5(32'h3af647b1),
	.w6(32'hbb76ec95),
	.w7(32'hba53729d),
	.w8(32'h3a8f8bd4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26fdcc),
	.w1(32'hbb6dfc1b),
	.w2(32'hbacb4f76),
	.w3(32'hba8ca63e),
	.w4(32'hbbc21b90),
	.w5(32'hbb04cfaf),
	.w6(32'h3ac350d2),
	.w7(32'hbb66bddb),
	.w8(32'hbbc67045),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2751),
	.w1(32'hbbc5d767),
	.w2(32'hbc011108),
	.w3(32'hbb4471c0),
	.w4(32'hbba73176),
	.w5(32'hbad69b50),
	.w6(32'h37ac89cb),
	.w7(32'hbb9ede5f),
	.w8(32'hbb34d1fb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15bf6f),
	.w1(32'h3af3bd98),
	.w2(32'h3a703605),
	.w3(32'hbc059af6),
	.w4(32'h3aa98005),
	.w5(32'h3b95e43b),
	.w6(32'hbbbdc68a),
	.w7(32'h3b781b6d),
	.w8(32'h3ac90b97),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9328e9),
	.w1(32'h3a5032f7),
	.w2(32'h38d217b9),
	.w3(32'h3a23f62b),
	.w4(32'h3b35246f),
	.w5(32'hb79bf4b7),
	.w6(32'h39b612a8),
	.w7(32'hbae4c48c),
	.w8(32'h3881e857),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fd009),
	.w1(32'h3a277d12),
	.w2(32'hb963b688),
	.w3(32'hba999e52),
	.w4(32'hba268f50),
	.w5(32'h39cd09c5),
	.w6(32'h3a970d6f),
	.w7(32'h394c4a27),
	.w8(32'h37ef398f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0f4f1),
	.w1(32'h3bf241e6),
	.w2(32'h3b9cb419),
	.w3(32'hbbbe9473),
	.w4(32'h3bb8ce16),
	.w5(32'h3a37cc32),
	.w6(32'hbb25b659),
	.w7(32'h3bf9f937),
	.w8(32'h3ba2ee7b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08158),
	.w1(32'h3b1135d6),
	.w2(32'h3a1d5f22),
	.w3(32'h3b758eda),
	.w4(32'h3a8fb439),
	.w5(32'h3a948444),
	.w6(32'h3bbddd6d),
	.w7(32'hbab28ba0),
	.w8(32'hbaaea127),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba33663),
	.w1(32'h39bce497),
	.w2(32'hbacd9255),
	.w3(32'h3b37c647),
	.w4(32'h38b65811),
	.w5(32'hbb01598b),
	.w6(32'hba2948a5),
	.w7(32'h3b132df6),
	.w8(32'hbafa966e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbce080),
	.w1(32'hbba0d5d5),
	.w2(32'hb9b4e51a),
	.w3(32'h3b873b8d),
	.w4(32'hbad7eddb),
	.w5(32'h3bcfbadf),
	.w6(32'h3b12726e),
	.w7(32'hbade259d),
	.w8(32'h3a6f00f7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e8bf),
	.w1(32'hbb1aa5bb),
	.w2(32'hbb8bdc05),
	.w3(32'h3b19b321),
	.w4(32'hbb8932da),
	.w5(32'hbb81a1c7),
	.w6(32'hba3f6a87),
	.w7(32'hbb72b89b),
	.w8(32'hbbb59e39),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfe91f),
	.w1(32'h3b6cd4fc),
	.w2(32'hba804d18),
	.w3(32'hbbccce6f),
	.w4(32'hba38def8),
	.w5(32'hbb51c80f),
	.w6(32'hbb825584),
	.w7(32'h3b4d24c0),
	.w8(32'hb8d94f35),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f0d6),
	.w1(32'hbb7b14c5),
	.w2(32'hbb1050a4),
	.w3(32'hbb1c95bf),
	.w4(32'hbaee321d),
	.w5(32'hbb09f6f2),
	.w6(32'hba7a6097),
	.w7(32'hbb00bd91),
	.w8(32'hbaf0ba8b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae82fb1),
	.w1(32'h3b1e2a89),
	.w2(32'h3b823b51),
	.w3(32'hbb00f74d),
	.w4(32'h3bebd9cc),
	.w5(32'h397e7e0b),
	.w6(32'hbb134d8f),
	.w7(32'h3b5d4ebc),
	.w8(32'h3bc678d7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12757),
	.w1(32'h3b3999bb),
	.w2(32'hbaa6f857),
	.w3(32'h3bd07bc3),
	.w4(32'hb98e0a8b),
	.w5(32'hb9e5c427),
	.w6(32'hba7a2901),
	.w7(32'hbb78fb16),
	.w8(32'hbac14c38),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5313),
	.w1(32'h39acbda0),
	.w2(32'h3b247f1a),
	.w3(32'hbb17cdc4),
	.w4(32'h3b30c932),
	.w5(32'h3c0d41f4),
	.w6(32'hbae7d579),
	.w7(32'h3b385e58),
	.w8(32'h3b1622fb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba118cba),
	.w1(32'hbb10c005),
	.w2(32'hbb36b3e6),
	.w3(32'h3af231a0),
	.w4(32'hbbce719b),
	.w5(32'h3ae6180a),
	.w6(32'h39e96287),
	.w7(32'hbad206c4),
	.w8(32'hbbde264b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f0e77),
	.w1(32'hbb79b8e7),
	.w2(32'h3b02bfdf),
	.w3(32'h3a0cc773),
	.w4(32'hba5bdd28),
	.w5(32'hbb389642),
	.w6(32'hbbb0fe84),
	.w7(32'hb985d09a),
	.w8(32'h3ac07848),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545ff3),
	.w1(32'h3b275a5e),
	.w2(32'h39712b7b),
	.w3(32'h3b87b63e),
	.w4(32'hb98c46b0),
	.w5(32'h3b98e67d),
	.w6(32'h3ba92eaa),
	.w7(32'h3b27fca6),
	.w8(32'h3bbf7733),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02fadb),
	.w1(32'h3b8caa33),
	.w2(32'hbb97d3fe),
	.w3(32'hbab2dce3),
	.w4(32'h3aa8b603),
	.w5(32'hbc72364d),
	.w6(32'h3b6df145),
	.w7(32'hbbaadefc),
	.w8(32'hbb1eab15),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8884b1e),
	.w1(32'h3a9f3752),
	.w2(32'h3ae343f7),
	.w3(32'hba33de8a),
	.w4(32'h38619c15),
	.w5(32'hbb8012e2),
	.w6(32'h3b961c91),
	.w7(32'hb9d29bb6),
	.w8(32'h3b84ad6a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeedead),
	.w1(32'h3b11c837),
	.w2(32'h3b959303),
	.w3(32'h395c3a63),
	.w4(32'h3bffc2ad),
	.w5(32'h3b4c3c82),
	.w6(32'h3ba89cc2),
	.w7(32'h3b04f3cf),
	.w8(32'h3a974b67),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e9614),
	.w1(32'h3b8fd55c),
	.w2(32'h3adfe3a1),
	.w3(32'h3b9a15a4),
	.w4(32'hb883300d),
	.w5(32'hbb3e05f8),
	.w6(32'h3b8f2cc7),
	.w7(32'h3b045ac6),
	.w8(32'h38f02512),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9c4d),
	.w1(32'hbae25999),
	.w2(32'hba9947ac),
	.w3(32'h398488c8),
	.w4(32'hbae87684),
	.w5(32'hbb13bb5c),
	.w6(32'h3bb0fb98),
	.w7(32'hbb79b1d5),
	.w8(32'hbbbff0aa),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d479),
	.w1(32'h3a563fc8),
	.w2(32'h39915767),
	.w3(32'hbb3ea071),
	.w4(32'h3b622ea0),
	.w5(32'hbb09889f),
	.w6(32'hbaf3ddef),
	.w7(32'h3adba218),
	.w8(32'hbacfc7b4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba51b0b),
	.w1(32'hba25a2ec),
	.w2(32'hbabb3425),
	.w3(32'h3ba4092f),
	.w4(32'h3a22ed0f),
	.w5(32'hbbb3a43a),
	.w6(32'h3ba95d61),
	.w7(32'hb9fdda70),
	.w8(32'hbb1ecf70),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d2b1d),
	.w1(32'h38c11e8f),
	.w2(32'hbb42b4d8),
	.w3(32'h3bd56b23),
	.w4(32'hbb52052f),
	.w5(32'hbbbd22a6),
	.w6(32'h3ad00818),
	.w7(32'hbb1158db),
	.w8(32'hbb8602ce),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ba3b5),
	.w1(32'hbb986173),
	.w2(32'h3ae3ef8b),
	.w3(32'h3b40b21f),
	.w4(32'hb9bb9353),
	.w5(32'h3bcbadbf),
	.w6(32'h3b69508e),
	.w7(32'h3b75a0bd),
	.w8(32'h3b5e235a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21e682),
	.w1(32'hb98bde25),
	.w2(32'hba826159),
	.w3(32'h387c3c98),
	.w4(32'hbb773c13),
	.w5(32'hbc3c4bb9),
	.w6(32'h3a066ef5),
	.w7(32'hbb870954),
	.w8(32'hbb74bb27),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b65b98),
	.w1(32'h3b68b5ab),
	.w2(32'h3b73fb77),
	.w3(32'h3b09c9fc),
	.w4(32'h3b3d32d5),
	.w5(32'h3cb6d18e),
	.w6(32'h3ba5fb9f),
	.w7(32'h3b3176e6),
	.w8(32'h3bf512a7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841f04),
	.w1(32'hbaf596c3),
	.w2(32'hbb200b14),
	.w3(32'h3b3fc553),
	.w4(32'hbaff32eb),
	.w5(32'h3a1f3ddc),
	.w6(32'h3b129b13),
	.w7(32'hba5d31e4),
	.w8(32'hbac41470),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81d126),
	.w1(32'h3b24c62c),
	.w2(32'h398416cb),
	.w3(32'hbb7b6f9d),
	.w4(32'h3b2e167b),
	.w5(32'hbb3a3527),
	.w6(32'hba6f8f3f),
	.w7(32'hbb7fab72),
	.w8(32'hbb7e26b2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8632250),
	.w1(32'h3aa8507c),
	.w2(32'h3b3bb9e2),
	.w3(32'hbb247c5c),
	.w4(32'hbb6d8e14),
	.w5(32'h3b426369),
	.w6(32'h3b13bb27),
	.w7(32'hba4861d7),
	.w8(32'h3b71a58d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3de595),
	.w1(32'hbafc7819),
	.w2(32'hbb10c8fb),
	.w3(32'hbb766d15),
	.w4(32'hba1bd630),
	.w5(32'hbb5a74b5),
	.w6(32'hbb38080e),
	.w7(32'hba173a15),
	.w8(32'h39987109),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6db14e),
	.w1(32'hba2de66f),
	.w2(32'h394217e8),
	.w3(32'h3b113bdc),
	.w4(32'h3a596cbf),
	.w5(32'hbba19db4),
	.w6(32'h3a4fb37a),
	.w7(32'h3aab477a),
	.w8(32'hbbcbcd9e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37df37),
	.w1(32'h3a2c0317),
	.w2(32'hbb4ab1f7),
	.w3(32'h3be681b8),
	.w4(32'hbb23ad95),
	.w5(32'hbb59c44d),
	.w6(32'h3ad771e4),
	.w7(32'hba30090c),
	.w8(32'hbb407553),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6669),
	.w1(32'hbaa5f898),
	.w2(32'hbb02bfe8),
	.w3(32'hbab12b80),
	.w4(32'hbb23c4b3),
	.w5(32'hbbcae310),
	.w6(32'h3ab36083),
	.w7(32'h3b5b8bc4),
	.w8(32'h3b176f92),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eb7a5),
	.w1(32'hbb1b4cc0),
	.w2(32'h399f2551),
	.w3(32'h3b86e8c3),
	.w4(32'hbb1634a5),
	.w5(32'h3ca5faf7),
	.w6(32'h3b2385ec),
	.w7(32'h3b35b08e),
	.w8(32'h3bc94fd1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8abd59),
	.w1(32'h386ca5ca),
	.w2(32'h3aebefb9),
	.w3(32'hba6d32da),
	.w4(32'h3a6bc3cf),
	.w5(32'h3c80db4e),
	.w6(32'hbbf23765),
	.w7(32'h3b31ccf9),
	.w8(32'h3b81a961),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ccc47),
	.w1(32'hbab61c4a),
	.w2(32'h3b976194),
	.w3(32'h3b8aa418),
	.w4(32'hba383f6e),
	.w5(32'h39433bfd),
	.w6(32'hb8687f4a),
	.w7(32'h39e3b067),
	.w8(32'h39cd9361),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76c17),
	.w1(32'h3abf1ebb),
	.w2(32'hbb063e03),
	.w3(32'hbab08ce8),
	.w4(32'hbb683c5b),
	.w5(32'h3a160b94),
	.w6(32'h3b0124a7),
	.w7(32'hbba799a5),
	.w8(32'h3af59704),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37abfb2a),
	.w1(32'hba066af7),
	.w2(32'h3a537f33),
	.w3(32'hbaf0d911),
	.w4(32'hbb17de66),
	.w5(32'hbb388b69),
	.w6(32'h3b19ba74),
	.w7(32'hbad29cba),
	.w8(32'h3a9be2fe),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23adc2),
	.w1(32'h3acb7256),
	.w2(32'h3a930b87),
	.w3(32'hba828b48),
	.w4(32'hba103097),
	.w5(32'h3b08cfb3),
	.w6(32'h3af2f58e),
	.w7(32'h3ac2bfd9),
	.w8(32'h3b1d26e0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d2e6d),
	.w1(32'hbbca2ecc),
	.w2(32'h3a9e8b08),
	.w3(32'h3b434c45),
	.w4(32'hbbc20f5e),
	.w5(32'h3bc84ddf),
	.w6(32'h3ab035e2),
	.w7(32'hba1708ee),
	.w8(32'hbb0e8b51),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace8c5a),
	.w1(32'hba2cea6b),
	.w2(32'h3a340006),
	.w3(32'hbb24bea4),
	.w4(32'hbb9edaeb),
	.w5(32'h3c58fccb),
	.w6(32'hbb8b9f14),
	.w7(32'h3b2ac4b7),
	.w8(32'h3b4c9169),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58346f),
	.w1(32'hbb20eb91),
	.w2(32'hbabca982),
	.w3(32'hbab2658c),
	.w4(32'hbb89be81),
	.w5(32'hbbe7982b),
	.w6(32'h3991a685),
	.w7(32'hba8e1871),
	.w8(32'hba84196b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01907b),
	.w1(32'h3a663b42),
	.w2(32'h3c10e5f0),
	.w3(32'h3a9031d7),
	.w4(32'h3bd9b062),
	.w5(32'hbbb65b78),
	.w6(32'h3ae7dd6c),
	.w7(32'h3b5f6a39),
	.w8(32'h3af0ebfd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3189),
	.w1(32'hb66aa423),
	.w2(32'hba23952e),
	.w3(32'h3bae6089),
	.w4(32'hbb1e162a),
	.w5(32'hbaa188fc),
	.w6(32'h3b5d42ad),
	.w7(32'hbacaaa58),
	.w8(32'hbb0e380b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6423f6),
	.w1(32'h3b0e54a0),
	.w2(32'h3ac6f971),
	.w3(32'hb918d5ae),
	.w4(32'h3b912365),
	.w5(32'hbb94b3f4),
	.w6(32'h3999bbcb),
	.w7(32'hba1da062),
	.w8(32'hba117445),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6ec87),
	.w1(32'h3a3f9f67),
	.w2(32'hba63f039),
	.w3(32'h39bab8f4),
	.w4(32'hbaf4ef3e),
	.w5(32'hbb9a24ab),
	.w6(32'h3b22785a),
	.w7(32'h381c166b),
	.w8(32'hbb514487),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df45e9),
	.w1(32'hb89f4ada),
	.w2(32'h3b0bbbcb),
	.w3(32'hbae6e23a),
	.w4(32'h399adcb9),
	.w5(32'hbc04b406),
	.w6(32'h3a93e8a2),
	.w7(32'hba5822b4),
	.w8(32'hbb2edf52),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a902667),
	.w1(32'hbb01cc5a),
	.w2(32'h3b7112ec),
	.w3(32'h3b93b5e7),
	.w4(32'hbaec1ed9),
	.w5(32'hbc551247),
	.w6(32'h3b403782),
	.w7(32'h3a27f514),
	.w8(32'hbbac23eb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cb682),
	.w1(32'h3b1bd9d5),
	.w2(32'h3aab4691),
	.w3(32'h3b0d25da),
	.w4(32'h3b124195),
	.w5(32'hbb918178),
	.w6(32'hba365130),
	.w7(32'hba965ecd),
	.w8(32'h3a37b2f5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b787834),
	.w1(32'h38a723ff),
	.w2(32'h3acb78d3),
	.w3(32'hb8be8634),
	.w4(32'hbab942bc),
	.w5(32'hb9dab1f7),
	.w6(32'h3b2b27e6),
	.w7(32'hbabd4922),
	.w8(32'hba055a2a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b940671),
	.w1(32'h3b121982),
	.w2(32'h3aa1926d),
	.w3(32'h3b06ab7e),
	.w4(32'hbb638742),
	.w5(32'h3c77885d),
	.w6(32'hbad89867),
	.w7(32'h3b60589c),
	.w8(32'h3b675230),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0c27c),
	.w1(32'h3a4a8311),
	.w2(32'h3c1a7922),
	.w3(32'h3a5df2ae),
	.w4(32'h3bcb8cf3),
	.w5(32'hbb009715),
	.w6(32'h3b48201f),
	.w7(32'h3ac5ab76),
	.w8(32'h3b084491),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe845d8),
	.w1(32'hba6bc5cc),
	.w2(32'hba9f1748),
	.w3(32'h3a9890d3),
	.w4(32'hbabe1c84),
	.w5(32'hbbc92510),
	.w6(32'h3ba1718d),
	.w7(32'h3a8af4eb),
	.w8(32'hbac590b2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7738c3),
	.w1(32'h3a010dec),
	.w2(32'h3ac069d0),
	.w3(32'hbae80142),
	.w4(32'h3b7d3c09),
	.w5(32'h3ba0f134),
	.w6(32'hbb2cd598),
	.w7(32'h3aa952ea),
	.w8(32'h3a0d650d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c11753),
	.w1(32'hba142271),
	.w2(32'h3bac2266),
	.w3(32'h39e88115),
	.w4(32'hbb3c06a3),
	.w5(32'hba13507c),
	.w6(32'h3ace21fd),
	.w7(32'h3bb67a52),
	.w8(32'h3bb11452),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79523),
	.w1(32'h39b87485),
	.w2(32'h3861de65),
	.w3(32'hb80ebfd4),
	.w4(32'hbb2d7e73),
	.w5(32'hbbbac2a3),
	.w6(32'h39f2d97e),
	.w7(32'hbb3750d8),
	.w8(32'hbb8fe7e5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36ec68),
	.w1(32'hb9c58ff3),
	.w2(32'h3a3429c6),
	.w3(32'h3b0eda9a),
	.w4(32'h3b2ac39e),
	.w5(32'h3cd03c53),
	.w6(32'h3a727c89),
	.w7(32'hba06d268),
	.w8(32'h3b55d67a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c05dc),
	.w1(32'hbb615d8c),
	.w2(32'hb9d0c59d),
	.w3(32'h3b2b759a),
	.w4(32'hba24f434),
	.w5(32'hbad8bd70),
	.w6(32'hbaee5078),
	.w7(32'h3b657bbd),
	.w8(32'hbb1c4b65),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a067a8),
	.w1(32'hb8aec5e8),
	.w2(32'h3a8414da),
	.w3(32'hbae4cfd9),
	.w4(32'hba802e8d),
	.w5(32'h3b6ceff0),
	.w6(32'hba12bfed),
	.w7(32'h3a8609c2),
	.w8(32'hba3a27b7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab25ff1),
	.w1(32'hbb266365),
	.w2(32'hbbe93765),
	.w3(32'h3a8dc2c5),
	.w4(32'hba33f338),
	.w5(32'hbace6967),
	.w6(32'h3b664e47),
	.w7(32'hbb751991),
	.w8(32'hbb843e70),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa32789),
	.w1(32'h3a5b9813),
	.w2(32'h3afdeeac),
	.w3(32'hbbbf17ea),
	.w4(32'hbaec24ee),
	.w5(32'h3c7d95d8),
	.w6(32'h3af65ffa),
	.w7(32'h3aa978f3),
	.w8(32'h3b0e5ccd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec6be8),
	.w1(32'hbb37138a),
	.w2(32'hbb454a04),
	.w3(32'hbaacb736),
	.w4(32'hbbb93858),
	.w5(32'h3b54fc0f),
	.w6(32'h3acd7d5b),
	.w7(32'hba870a1c),
	.w8(32'hbb850c56),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b55f),
	.w1(32'h3aee53bf),
	.w2(32'h39f2694e),
	.w3(32'hbb8abcf0),
	.w4(32'h3b100d36),
	.w5(32'hbc0bbc85),
	.w6(32'hbb31540e),
	.w7(32'h3a9c1329),
	.w8(32'h3a41ea0a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9099a1),
	.w1(32'hba819a92),
	.w2(32'h3bde82fe),
	.w3(32'h3c041851),
	.w4(32'h3b869317),
	.w5(32'h3b468903),
	.w6(32'h3b0b6cbe),
	.w7(32'h3b12b896),
	.w8(32'h3ae6f270),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f6705),
	.w1(32'hb9b5fa1e),
	.w2(32'hbba93762),
	.w3(32'h3bbc8da4),
	.w4(32'hbb00c9b5),
	.w5(32'hbb88b3a7),
	.w6(32'hba21315c),
	.w7(32'hbb3684a9),
	.w8(32'hba1a0659),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2019bf),
	.w1(32'hbb101600),
	.w2(32'hbac43138),
	.w3(32'h3ad1f0c2),
	.w4(32'hb9762345),
	.w5(32'h3bf9b6ba),
	.w6(32'hbaf11bc3),
	.w7(32'h3ba2344c),
	.w8(32'hbae4840f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule