module layer_8_featuremap_109(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c61f4),
	.w1(32'hb9891398),
	.w2(32'h3bdab28d),
	.w3(32'hba85cd48),
	.w4(32'hbbea8377),
	.w5(32'hbbd9cc20),
	.w6(32'hbc069f7a),
	.w7(32'hbbc9cf3c),
	.w8(32'hbb734c02),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48c28),
	.w1(32'h3ab74691),
	.w2(32'hbb96a65f),
	.w3(32'hbb9c6d09),
	.w4(32'h3aa5fe53),
	.w5(32'hbb140e2a),
	.w6(32'hbb95e823),
	.w7(32'hbb60d3e4),
	.w8(32'hbbc39cc4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2be0),
	.w1(32'hba8e3265),
	.w2(32'hbb1aef73),
	.w3(32'h398c5bd4),
	.w4(32'h3b6d179b),
	.w5(32'h3bc18fcb),
	.w6(32'hbb1947a0),
	.w7(32'hbbd0f31c),
	.w8(32'h3b897907),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc19bd),
	.w1(32'hbb70693a),
	.w2(32'hbbcd597d),
	.w3(32'hbbbada21),
	.w4(32'hbad24b0b),
	.w5(32'h3b8c9632),
	.w6(32'hbb3dfdf5),
	.w7(32'hbaf4b08c),
	.w8(32'hba0c3005),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046922),
	.w1(32'h3a3034d1),
	.w2(32'hbc125da2),
	.w3(32'hbba9260b),
	.w4(32'h3b3a07d9),
	.w5(32'h3bf183d7),
	.w6(32'hbb2f6f17),
	.w7(32'hbaece38d),
	.w8(32'h3ac5f8b9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86a51f),
	.w1(32'hbb6f187c),
	.w2(32'hbbb68dd4),
	.w3(32'hba98eeea),
	.w4(32'h3b8c0685),
	.w5(32'h3b1105a3),
	.w6(32'hbb81e9cd),
	.w7(32'h3c0a2559),
	.w8(32'h3c231ac3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756846),
	.w1(32'h3acaa9d7),
	.w2(32'hbab8e5b5),
	.w3(32'hbb2153b0),
	.w4(32'hbb3032a9),
	.w5(32'h39d8f7c7),
	.w6(32'h3a868ab5),
	.w7(32'hbbb66ea7),
	.w8(32'hb94452c7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61dd76),
	.w1(32'h3b44b87c),
	.w2(32'hbb6d6f41),
	.w3(32'hbb9329d5),
	.w4(32'hbb167aa5),
	.w5(32'h3aa9a697),
	.w6(32'hbb562cb1),
	.w7(32'h3b9fc802),
	.w8(32'h39c410e4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb063f66),
	.w1(32'hbb4a1e6f),
	.w2(32'h3b77c42b),
	.w3(32'hbbeb9d15),
	.w4(32'hbb877e92),
	.w5(32'h3976c2eb),
	.w6(32'hbb91d1fd),
	.w7(32'hba5f7c1f),
	.w8(32'h3a1a7203),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e3d3e),
	.w1(32'h3b4523a2),
	.w2(32'hbb914ad9),
	.w3(32'hba96e870),
	.w4(32'hbb4bfab2),
	.w5(32'h3ba8a16d),
	.w6(32'h3967e6e5),
	.w7(32'h3ae8476a),
	.w8(32'h3c09947e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b960),
	.w1(32'hbb861717),
	.w2(32'hbb07dd52),
	.w3(32'hbbfeeb42),
	.w4(32'hbb3d6433),
	.w5(32'hbad0dedc),
	.w6(32'hbc91966c),
	.w7(32'h3b9106a3),
	.w8(32'h3b5e3420),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a0453),
	.w1(32'hbbdcb37c),
	.w2(32'hbbb5a904),
	.w3(32'hbc0de917),
	.w4(32'h3b83333c),
	.w5(32'h39363f38),
	.w6(32'hbbae714d),
	.w7(32'h3b5237f8),
	.w8(32'hba25f9c8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba136a89),
	.w1(32'hbb38f2b5),
	.w2(32'hbb01f4a5),
	.w3(32'hbba68adc),
	.w4(32'hb79322da),
	.w5(32'hba9dfef7),
	.w6(32'hbbd3eede),
	.w7(32'hbb4ced7a),
	.w8(32'hba9d5d18),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa853),
	.w1(32'h3a8fac53),
	.w2(32'hbb5803b2),
	.w3(32'hba71fae1),
	.w4(32'hba8c4c1a),
	.w5(32'hbb20c40f),
	.w6(32'h3ace042e),
	.w7(32'hba1fa40c),
	.w8(32'hba5267a8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad5560),
	.w1(32'hbb00b17f),
	.w2(32'hbb428b2c),
	.w3(32'h395486ca),
	.w4(32'h3a5ce945),
	.w5(32'h38317a8d),
	.w6(32'h3888eefb),
	.w7(32'hbaa0df08),
	.w8(32'hbb0f6622),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381417),
	.w1(32'hbabd94ec),
	.w2(32'hb9f63a79),
	.w3(32'h38f4c0c6),
	.w4(32'hbb3e81e4),
	.w5(32'h3aa4066a),
	.w6(32'hbaa41ef5),
	.w7(32'hb9a6d1a2),
	.w8(32'h3b035b94),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9129d),
	.w1(32'hbb41bbfe),
	.w2(32'h3b57f3c5),
	.w3(32'hba2c3a02),
	.w4(32'hba18aa2f),
	.w5(32'h3a3a5276),
	.w6(32'h3ab32610),
	.w7(32'hbb453893),
	.w8(32'h3b273d9e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ff1a6),
	.w1(32'hba835abf),
	.w2(32'hbc1af9f2),
	.w3(32'hbba9ca82),
	.w4(32'hbc9351ed),
	.w5(32'hbc5a7c64),
	.w6(32'hbc217432),
	.w7(32'hbc9e4b4b),
	.w8(32'hbc4b325a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce2ae93),
	.w1(32'hbcabfc77),
	.w2(32'hbb9a0ce7),
	.w3(32'hbcd3b251),
	.w4(32'hbc929c9c),
	.w5(32'hbb86fcef),
	.w6(32'hbcad39ce),
	.w7(32'hbc5992c5),
	.w8(32'hbba767c1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d9fe9),
	.w1(32'hbc0dd864),
	.w2(32'hbc9c5faa),
	.w3(32'hbc1ec8d8),
	.w4(32'hbc81413a),
	.w5(32'hbc004452),
	.w6(32'hbbb98949),
	.w7(32'hbc7f96ef),
	.w8(32'hbc3cb21d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ee2bb),
	.w1(32'hbbbe3ea3),
	.w2(32'h3b8ed041),
	.w3(32'hbb89e571),
	.w4(32'hbbfc6a7e),
	.w5(32'hbb3635cc),
	.w6(32'hbc009ad9),
	.w7(32'hbbb94623),
	.w8(32'hbc0cb2a3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb028f),
	.w1(32'hbc2e29f3),
	.w2(32'hbb415618),
	.w3(32'hb9a49099),
	.w4(32'h3b1bafe3),
	.w5(32'hbb950deb),
	.w6(32'hbb99a525),
	.w7(32'h3bfde616),
	.w8(32'h3b220f5e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9876),
	.w1(32'h3a14aca2),
	.w2(32'hbb84ba13),
	.w3(32'hbbe7e24c),
	.w4(32'h3aa73c3b),
	.w5(32'h3b08273a),
	.w6(32'hbb8a3fbc),
	.w7(32'hbb112f05),
	.w8(32'hbb92d82d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cd4f6),
	.w1(32'hba8ecb35),
	.w2(32'hbc045b20),
	.w3(32'h3ae5d450),
	.w4(32'hbb9004a2),
	.w5(32'hbad435f6),
	.w6(32'h3b68d5b9),
	.w7(32'hbc0496ef),
	.w8(32'hbc19d949),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512e57),
	.w1(32'h3b4d9339),
	.w2(32'hbbc91c36),
	.w3(32'h3b941032),
	.w4(32'h3bbd41b8),
	.w5(32'h3a206a8d),
	.w6(32'h3b7b7ab7),
	.w7(32'h3aa83249),
	.w8(32'hb91a9dd0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b2e83),
	.w1(32'hbbcaff16),
	.w2(32'hbb3412e9),
	.w3(32'hbbaab0f7),
	.w4(32'hbb1ad72e),
	.w5(32'h3b2a2f6d),
	.w6(32'hbbcdc5c7),
	.w7(32'hba517ad7),
	.w8(32'h3b1ea0fc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadac5fb),
	.w1(32'h3b5c362e),
	.w2(32'h3aed3b52),
	.w3(32'h3c3499d3),
	.w4(32'h3bbbaa17),
	.w5(32'h3b7fcde8),
	.w6(32'hba0d517f),
	.w7(32'h3bf297de),
	.w8(32'h3c3a42db),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b795f),
	.w1(32'hbc297e49),
	.w2(32'hbc09ab99),
	.w3(32'h392ee2f4),
	.w4(32'h3a4ba97a),
	.w5(32'hbc1f76e7),
	.w6(32'hbca7b61f),
	.w7(32'h3cd5da43),
	.w8(32'h3c5d4cc6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b450074),
	.w1(32'h3b9972fe),
	.w2(32'h3be12602),
	.w3(32'h3c82f33c),
	.w4(32'hbaa36ef2),
	.w5(32'hbb95fedf),
	.w6(32'h3c93d0e8),
	.w7(32'h3b56cbd3),
	.w8(32'h396f8372),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b466),
	.w1(32'h3bd2ed1e),
	.w2(32'h3c53ed5a),
	.w3(32'hb9ad985f),
	.w4(32'hbb898ad9),
	.w5(32'hbc2e4124),
	.w6(32'h3b02fdd0),
	.w7(32'h3b8e61e9),
	.w8(32'hbaff2c59),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d3f4c),
	.w1(32'h3b031812),
	.w2(32'h3ac16a5d),
	.w3(32'hbbb3868b),
	.w4(32'h3c21c20b),
	.w5(32'h3c0bf658),
	.w6(32'h3bdbc3de),
	.w7(32'h3bf4dddd),
	.w8(32'h3bae3c6f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63655),
	.w1(32'h3b2626df),
	.w2(32'hbb0c3453),
	.w3(32'h3b98da8b),
	.w4(32'hbb86b501),
	.w5(32'hba802bdd),
	.w6(32'h3aeac143),
	.w7(32'hbb8bd795),
	.w8(32'hbbda29d2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc239a6),
	.w1(32'hbc070390),
	.w2(32'h3b8a8668),
	.w3(32'hbc00ac81),
	.w4(32'hbb0705c4),
	.w5(32'hbb63fc28),
	.w6(32'hba9dd6db),
	.w7(32'hbc1cd4cf),
	.w8(32'hbc00e1ec),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ff22),
	.w1(32'h3a6b758f),
	.w2(32'h3be0d688),
	.w3(32'hbc0ff04c),
	.w4(32'hbbe24f15),
	.w5(32'hbbccb70b),
	.w6(32'hbc52983c),
	.w7(32'hbb698cdc),
	.w8(32'h3b73e77e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca1342),
	.w1(32'hb8b07f58),
	.w2(32'hbb1ce501),
	.w3(32'hb9f65ddb),
	.w4(32'h3a98e22b),
	.w5(32'hbadf53fa),
	.w6(32'hbbc2a1f5),
	.w7(32'hbac53436),
	.w8(32'hbbaba988),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26fc04),
	.w1(32'hbb809fb2),
	.w2(32'hbc06444a),
	.w3(32'h3b26c340),
	.w4(32'h39b2be5d),
	.w5(32'hbc09846c),
	.w6(32'hba448a61),
	.w7(32'hba97a819),
	.w8(32'hbb8180ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aa0ce),
	.w1(32'h3c029a02),
	.w2(32'h3aa048e7),
	.w3(32'hbc360ed4),
	.w4(32'h3b95c394),
	.w5(32'h3b2685a7),
	.w6(32'hbc177340),
	.w7(32'hbc07790d),
	.w8(32'hbbb2ef55),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a24f91),
	.w1(32'h3afdd4ff),
	.w2(32'hbab01e8a),
	.w3(32'h3c100ea3),
	.w4(32'h3b9d0053),
	.w5(32'h3b8d58b1),
	.w6(32'hbbc6c695),
	.w7(32'hba42f341),
	.w8(32'h3b86c0b4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab510b1),
	.w1(32'hba7e401e),
	.w2(32'hbb1a2274),
	.w3(32'hbae51109),
	.w4(32'hba65de1e),
	.w5(32'hbba3be19),
	.w6(32'hbaaacb84),
	.w7(32'hbb6dadf6),
	.w8(32'h3919bfe0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade74f4),
	.w1(32'h3a2a0882),
	.w2(32'hbab7db0f),
	.w3(32'hbb3dec4a),
	.w4(32'h3c72a551),
	.w5(32'h3c68e833),
	.w6(32'h3aa92830),
	.w7(32'h3c78f948),
	.w8(32'h3c9fe9e2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eb4bc),
	.w1(32'hbb5b0f87),
	.w2(32'hbc847ef9),
	.w3(32'hbad8cb93),
	.w4(32'hbbed21af),
	.w5(32'hbc1e6c84),
	.w6(32'h3b7b2858),
	.w7(32'hbb8e8f30),
	.w8(32'hbc318e1f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cff8),
	.w1(32'hbbe033b8),
	.w2(32'h3b12d55a),
	.w3(32'hbb8ad30f),
	.w4(32'h3c7257b6),
	.w5(32'h3c6e9479),
	.w6(32'hbbf4940f),
	.w7(32'h3c1d39b2),
	.w8(32'h3c0cde2a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27d18),
	.w1(32'h3bbf7fa2),
	.w2(32'h3c277633),
	.w3(32'h3c8130b8),
	.w4(32'h3bc2793e),
	.w5(32'hba061804),
	.w6(32'h3c1eacd0),
	.w7(32'hbbb04b6b),
	.w8(32'hbc99f3f9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19bda7),
	.w1(32'h3c135ed8),
	.w2(32'hbba670f6),
	.w3(32'hbbe8ecd2),
	.w4(32'hb9217f07),
	.w5(32'hbb17be45),
	.w6(32'hbb267332),
	.w7(32'hbb6decc9),
	.w8(32'hb990419f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83d69),
	.w1(32'hbb513c4a),
	.w2(32'h3ac4410b),
	.w3(32'hbbeffce6),
	.w4(32'hbbb40676),
	.w5(32'hbbda22ab),
	.w6(32'hbb4bd6c1),
	.w7(32'hbb9b9188),
	.w8(32'h3a5b518b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00a47a),
	.w1(32'hb909a857),
	.w2(32'hbbfb42bf),
	.w3(32'hbb60c910),
	.w4(32'h3c39581e),
	.w5(32'h3b9c047d),
	.w6(32'hbb368ce6),
	.w7(32'h3b9f9895),
	.w8(32'h3b266faf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc16d),
	.w1(32'h3c692ddf),
	.w2(32'hbba21978),
	.w3(32'hbafc452c),
	.w4(32'h3b774f3b),
	.w5(32'hba446459),
	.w6(32'h3bfc97e7),
	.w7(32'hbb859b71),
	.w8(32'hbb9061e3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb732f5e),
	.w1(32'hbb7fe04e),
	.w2(32'h3aa14025),
	.w3(32'hbbb2bd01),
	.w4(32'hbc6801b3),
	.w5(32'hbba0da9f),
	.w6(32'hbbe3bc05),
	.w7(32'hbc0375c2),
	.w8(32'h3abd0e8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319120),
	.w1(32'h3bfbcd7b),
	.w2(32'hbb8a6be6),
	.w3(32'hbb7949f3),
	.w4(32'hbae243c0),
	.w5(32'hb9a13c86),
	.w6(32'h3b03d27f),
	.w7(32'hbb901daa),
	.w8(32'h3bb8c5c9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb631f22),
	.w1(32'hbbbc65db),
	.w2(32'hbae9a2c9),
	.w3(32'h3af9022b),
	.w4(32'hbbdf1c71),
	.w5(32'hbb862664),
	.w6(32'hbb8ed026),
	.w7(32'hbbae22fa),
	.w8(32'h3aaae1f1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e348c),
	.w1(32'h3c29ef9e),
	.w2(32'hbbb3d651),
	.w3(32'h3b71b2cb),
	.w4(32'hba4247dc),
	.w5(32'h3ba3875f),
	.w6(32'h3c027135),
	.w7(32'h3a916514),
	.w8(32'h3c342dd9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc32840),
	.w1(32'hbc92e815),
	.w2(32'hbba64521),
	.w3(32'hbcd5e49c),
	.w4(32'hbca4c76d),
	.w5(32'hbb3abaeb),
	.w6(32'hbca10a30),
	.w7(32'hbc80d1af),
	.w8(32'hbb2eaba9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f6eec),
	.w1(32'hba76f23b),
	.w2(32'h39c98595),
	.w3(32'h3afdd2c8),
	.w4(32'hbbe7eccc),
	.w5(32'h3b12dd37),
	.w6(32'hbba7e78e),
	.w7(32'hbb8fe254),
	.w8(32'h3b6195a7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b995d08),
	.w1(32'h3b5408e8),
	.w2(32'hb9c68df6),
	.w3(32'h3a5f3ab3),
	.w4(32'hbb863d16),
	.w5(32'hbb11cc6e),
	.w6(32'h3b80ea74),
	.w7(32'hbb979a2b),
	.w8(32'hba031502),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ffac),
	.w1(32'h3b29bd83),
	.w2(32'hbc3ea13b),
	.w3(32'h3a7aaa0c),
	.w4(32'hbb37270f),
	.w5(32'hbbcc6a4f),
	.w6(32'h3b59d2fa),
	.w7(32'hbba15ba1),
	.w8(32'hbb02de17),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99402d),
	.w1(32'hba737ea9),
	.w2(32'h3b97f781),
	.w3(32'hbc0626ae),
	.w4(32'hbb8298bf),
	.w5(32'hba4441bf),
	.w6(32'hbb76d42a),
	.w7(32'hbbc0b5b6),
	.w8(32'hbb92db13),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81eabe),
	.w1(32'hbaca5f14),
	.w2(32'h3c128feb),
	.w3(32'hbb92fe6a),
	.w4(32'h3c1496b0),
	.w5(32'h3ca3736f),
	.w6(32'hbbc43e5e),
	.w7(32'h3c939d91),
	.w8(32'h3ce4531c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65659c),
	.w1(32'h3ba04148),
	.w2(32'h3c475653),
	.w3(32'h3ca8b7bf),
	.w4(32'h3c1ac204),
	.w5(32'h3c448bf8),
	.w6(32'h3c3009b4),
	.w7(32'h3c5ea42d),
	.w8(32'h3c2f86f7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aecc5),
	.w1(32'h3c91ee68),
	.w2(32'hba1e523a),
	.w3(32'h3c31a660),
	.w4(32'h399f9d11),
	.w5(32'h399650b3),
	.w6(32'h3c894297),
	.w7(32'hb9c09afb),
	.w8(32'h3b90ccb1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e281),
	.w1(32'h38159ba3),
	.w2(32'hbbe08f3a),
	.w3(32'hbae75792),
	.w4(32'h3b98623d),
	.w5(32'h3c2a6321),
	.w6(32'hb9ad9792),
	.w7(32'h3a9c661c),
	.w8(32'hbbcfcb26),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0241b1),
	.w1(32'hb95936e5),
	.w2(32'hbb520b5d),
	.w3(32'h3c722127),
	.w4(32'h3b8cae9b),
	.w5(32'hbbedaf64),
	.w6(32'hbb807ada),
	.w7(32'h3bc14eb2),
	.w8(32'hbba4bedb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4d77f),
	.w1(32'h3ab0f13f),
	.w2(32'hbb9779f9),
	.w3(32'hbc2a59ba),
	.w4(32'hba625696),
	.w5(32'h39951a42),
	.w6(32'hbc011b5b),
	.w7(32'hbba5a949),
	.w8(32'hbae7d5d9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e9a1a),
	.w1(32'hbbf979b2),
	.w2(32'hbaa2cc6d),
	.w3(32'hbbbb2c09),
	.w4(32'hbb9226fa),
	.w5(32'hbc0f5936),
	.w6(32'hbc18aca2),
	.w7(32'hbb0eb96c),
	.w8(32'hbbf4036c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c3146),
	.w1(32'hbbeb2dac),
	.w2(32'hbb712f06),
	.w3(32'hbbb4cf67),
	.w4(32'hbad0be71),
	.w5(32'hbba3ae1d),
	.w6(32'hbbbd6b49),
	.w7(32'hbb89f00f),
	.w8(32'hbb89c0df),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb301f61),
	.w1(32'hbbb7b991),
	.w2(32'hb9c59cda),
	.w3(32'hbb19ef14),
	.w4(32'h3b6ddea9),
	.w5(32'h3b34904f),
	.w6(32'hba2fe832),
	.w7(32'h3bab1418),
	.w8(32'h3a6ad861),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78ca2a),
	.w1(32'h3a6fed27),
	.w2(32'hbaf9fb48),
	.w3(32'h3bb3e553),
	.w4(32'hbb0d3ca6),
	.w5(32'hbb865824),
	.w6(32'h3bbe79b6),
	.w7(32'hbc01bd45),
	.w8(32'hbc039620),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24a4e),
	.w1(32'hbb332251),
	.w2(32'hbc214bea),
	.w3(32'hbc1ce58d),
	.w4(32'hbc416573),
	.w5(32'hbbb5dc24),
	.w6(32'hbc2a2e77),
	.w7(32'hbc5bf358),
	.w8(32'hbbbcff31),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a64e),
	.w1(32'hbb826193),
	.w2(32'h3bf6990e),
	.w3(32'h3ae19c27),
	.w4(32'h3b8a8244),
	.w5(32'h3ba87b0b),
	.w6(32'h3af699a8),
	.w7(32'hbb9874dc),
	.w8(32'hbc0b53a0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09359f),
	.w1(32'h3b8bce19),
	.w2(32'hbb9e5736),
	.w3(32'h3b06cf1d),
	.w4(32'hbac0ea3d),
	.w5(32'hb931df3b),
	.w6(32'hbae3362d),
	.w7(32'hbba48703),
	.w8(32'hbb876045),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f504),
	.w1(32'hbc388fea),
	.w2(32'h3bd3eb35),
	.w3(32'hbbce86ff),
	.w4(32'hbc901869),
	.w5(32'hbc6c569d),
	.w6(32'hbc260a77),
	.w7(32'hbc329111),
	.w8(32'hbc04fbd3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a363),
	.w1(32'h3b39b020),
	.w2(32'h3b04ff65),
	.w3(32'h3ba9a3c1),
	.w4(32'h3b4c4ddd),
	.w5(32'h3b7d0105),
	.w6(32'hbc0022e0),
	.w7(32'h3a5b1581),
	.w8(32'hbae8fa16),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6acd3c),
	.w1(32'h3b73a69f),
	.w2(32'hbacce771),
	.w3(32'h391a0ec7),
	.w4(32'h3bbbabab),
	.w5(32'hbbb948eb),
	.w6(32'hbb18172c),
	.w7(32'h3afb554d),
	.w8(32'hbb05f1ce),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5242a4),
	.w1(32'h3b01418f),
	.w2(32'h3b70b077),
	.w3(32'hbb23f63c),
	.w4(32'h3be81964),
	.w5(32'h3bd5e2f3),
	.w6(32'hbc0432e8),
	.w7(32'hbbd39ead),
	.w8(32'hbbb50f83),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038374),
	.w1(32'h3c53dd39),
	.w2(32'h3bf32c43),
	.w3(32'h3b947787),
	.w4(32'h3c1d5bb9),
	.w5(32'h3beeb6db),
	.w6(32'hbb63f630),
	.w7(32'hbad5cc88),
	.w8(32'hbbe43f22),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894080),
	.w1(32'hbbaecabc),
	.w2(32'hbbcb7804),
	.w3(32'h3c5897e0),
	.w4(32'hbb161928),
	.w5(32'hbb2770df),
	.w6(32'hbbff9b3f),
	.w7(32'hb80d6930),
	.w8(32'h3b57c0b9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16a7cc),
	.w1(32'h3ba900ec),
	.w2(32'h3b1bcc6a),
	.w3(32'hbb9dbd9a),
	.w4(32'h3bc5ae0b),
	.w5(32'h3b8e69e0),
	.w6(32'h3bf1e3ca),
	.w7(32'h39fe0114),
	.w8(32'hbb69e2f4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ce239),
	.w1(32'h3b44d88f),
	.w2(32'hba7d54b1),
	.w3(32'hb9ef7ca8),
	.w4(32'h3998e66f),
	.w5(32'h3962543e),
	.w6(32'h3a1a4c68),
	.w7(32'hba19de69),
	.w8(32'hba20dacb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc0000),
	.w1(32'hbbc725aa),
	.w2(32'hbc0d8b65),
	.w3(32'hbbe7aed4),
	.w4(32'hbc630f91),
	.w5(32'hbc02f258),
	.w6(32'hbba3c91b),
	.w7(32'hbc042064),
	.w8(32'hbb8ab8d3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9a3fc),
	.w1(32'h3ba2a4b4),
	.w2(32'h3a0cc917),
	.w3(32'hbac70bc7),
	.w4(32'hb9ac1314),
	.w5(32'h3a5a8f6c),
	.w6(32'hb875c993),
	.w7(32'hb9bf7980),
	.w8(32'hbb12a4b1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f27d),
	.w1(32'hbb94329d),
	.w2(32'h3b513f1a),
	.w3(32'hbb942e75),
	.w4(32'h3bdcb101),
	.w5(32'h3acaa50a),
	.w6(32'hbb7e7798),
	.w7(32'h3b6c549d),
	.w8(32'hbaba32c4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dad7de),
	.w1(32'h3c126c5b),
	.w2(32'hba8dc355),
	.w3(32'hbc01297f),
	.w4(32'h3b334860),
	.w5(32'hbbfcc5d5),
	.w6(32'hbc7096db),
	.w7(32'h3bdfbc7e),
	.w8(32'hbc491f0a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82a009),
	.w1(32'hbbddc399),
	.w2(32'hbc0aa463),
	.w3(32'hbba3fea5),
	.w4(32'h3bfc420e),
	.w5(32'hbc46b170),
	.w6(32'hb937059b),
	.w7(32'hbbf5bfb6),
	.w8(32'hbbe61b7c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0056af),
	.w1(32'hbc985265),
	.w2(32'hbc79ef44),
	.w3(32'hbcb15132),
	.w4(32'hbc867dff),
	.w5(32'hbc364f3b),
	.w6(32'hbc64c9ef),
	.w7(32'hbc75935c),
	.w8(32'hbc8326ac),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf685e),
	.w1(32'hbbc653c7),
	.w2(32'hbaa24b55),
	.w3(32'hbbf5227e),
	.w4(32'hbbbd6f96),
	.w5(32'hbc461089),
	.w6(32'hbb964173),
	.w7(32'hbb3b5b20),
	.w8(32'hbcb8b355),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb984d),
	.w1(32'h3c820ee5),
	.w2(32'hbbe3e346),
	.w3(32'hbc867994),
	.w4(32'hbc7451b9),
	.w5(32'hbaf63d73),
	.w6(32'hbc3d0410),
	.w7(32'hbc970d04),
	.w8(32'hbc50795e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a4ddf),
	.w1(32'h3c740664),
	.w2(32'hbca4be28),
	.w3(32'h3b6f62f2),
	.w4(32'hbc524594),
	.w5(32'hbbe41b6a),
	.w6(32'h3c06a8d7),
	.w7(32'hbcd32502),
	.w8(32'hbcf45411),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a4633),
	.w1(32'hbc18bdfc),
	.w2(32'h3a278fa9),
	.w3(32'h3bc8b2f3),
	.w4(32'h3b8a4553),
	.w5(32'hbb2cd980),
	.w6(32'hbc6249e4),
	.w7(32'hb9cf086f),
	.w8(32'hbc2dfb82),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20f98),
	.w1(32'h3b75038f),
	.w2(32'h3bccf682),
	.w3(32'hbb9461fa),
	.w4(32'h3baef59a),
	.w5(32'h3b02a668),
	.w6(32'h3a813e22),
	.w7(32'h3b34f332),
	.w8(32'hbab09eae),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb98fff),
	.w1(32'hb8965135),
	.w2(32'h3b00bc39),
	.w3(32'h3aa62176),
	.w4(32'h3ac83ac2),
	.w5(32'h3afa46fb),
	.w6(32'hb99a01f8),
	.w7(32'hbaa32e56),
	.w8(32'h3aa95257),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f9ff0),
	.w1(32'h39c53bae),
	.w2(32'h3c53e83b),
	.w3(32'h3a4295ca),
	.w4(32'hbba0d404),
	.w5(32'hbc47b0dd),
	.w6(32'hbaf092c7),
	.w7(32'h3b845365),
	.w8(32'hbca04208),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2242),
	.w1(32'h3cb051fb),
	.w2(32'h3bcc13ec),
	.w3(32'hbada2ea8),
	.w4(32'hb9f40ae8),
	.w5(32'h3c070555),
	.w6(32'h3a69025e),
	.w7(32'h3880770a),
	.w8(32'h3c6a80be),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fd4d0),
	.w1(32'h3bdd6388),
	.w2(32'hbbb3045a),
	.w3(32'h39951351),
	.w4(32'hbc22bb0a),
	.w5(32'hbc6e1122),
	.w6(32'h3bdbbc8e),
	.w7(32'hbc4e151c),
	.w8(32'hbc8c1142),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf14bbd),
	.w1(32'hbbeb7ae1),
	.w2(32'h3b4fdf8e),
	.w3(32'hbc8a7691),
	.w4(32'hbac175d4),
	.w5(32'hbc0361f2),
	.w6(32'hbc213d0a),
	.w7(32'h3aa01524),
	.w8(32'hba57ce3d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ce1dc),
	.w1(32'h3ae48ec0),
	.w2(32'hbc2205d1),
	.w3(32'hbb7aed8d),
	.w4(32'hbbd561b5),
	.w5(32'hbc687fad),
	.w6(32'hbc4c58a6),
	.w7(32'hbc9ad0a3),
	.w8(32'h3bfc09f8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30693a),
	.w1(32'hbb06c8af),
	.w2(32'hbbaf361d),
	.w3(32'hbb8d900f),
	.w4(32'hbbb7728c),
	.w5(32'hbb50be35),
	.w6(32'hbb19253b),
	.w7(32'hbb502d5e),
	.w8(32'hbb7cf2ce),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d5e0),
	.w1(32'hba2a2574),
	.w2(32'h3c26e5e3),
	.w3(32'hbaddc96c),
	.w4(32'h3c05c17f),
	.w5(32'h3c597eb8),
	.w6(32'h3a28d7b3),
	.w7(32'hbbd49c78),
	.w8(32'h3c1802a2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5676),
	.w1(32'hbbf6d09d),
	.w2(32'hbb3d4774),
	.w3(32'hbc4291e9),
	.w4(32'hbc16f5f8),
	.w5(32'hbc48cd79),
	.w6(32'hbc1fe2b4),
	.w7(32'hbc1958cf),
	.w8(32'hbc3e98dd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5824d7),
	.w1(32'hbbc69095),
	.w2(32'hbc798b07),
	.w3(32'hbbb62c46),
	.w4(32'hba9df3ec),
	.w5(32'h3a8d2846),
	.w6(32'h3c0f9f7e),
	.w7(32'hbb832f65),
	.w8(32'h3b1e02e2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82db3d),
	.w1(32'hbc83c766),
	.w2(32'h3b18df39),
	.w3(32'hbb001380),
	.w4(32'h39cf130f),
	.w5(32'h3ac4436e),
	.w6(32'hbac6f6a5),
	.w7(32'h3b37c612),
	.w8(32'h3ad7ea0b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fcaab4),
	.w1(32'h3c051114),
	.w2(32'h3b195be4),
	.w3(32'h3c0b945b),
	.w4(32'h3b0da737),
	.w5(32'hbbbe085a),
	.w6(32'h3bf6ba67),
	.w7(32'hbc14e0f1),
	.w8(32'hbca1c9f4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb843e7),
	.w1(32'h3baa2de1),
	.w2(32'h3a322024),
	.w3(32'hbb67bfd1),
	.w4(32'hbc898bd2),
	.w5(32'hba155cc6),
	.w6(32'hbc5a4fc1),
	.w7(32'hbc28f6ac),
	.w8(32'hbc98ba7e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90f181),
	.w1(32'hbbcaa15b),
	.w2(32'hbbeee058),
	.w3(32'hbc62f046),
	.w4(32'hbc1339e5),
	.w5(32'hbc189da2),
	.w6(32'hbc5f5c84),
	.w7(32'hb80dfd58),
	.w8(32'hbc0cd245),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad43b),
	.w1(32'hbba58d1e),
	.w2(32'h3c2b863c),
	.w3(32'h3c55c322),
	.w4(32'h3bd951b6),
	.w5(32'h3b572aae),
	.w6(32'h3b8eb661),
	.w7(32'h3baafb88),
	.w8(32'h3bce67e7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865d46),
	.w1(32'hbb92a5c0),
	.w2(32'hbb500bb3),
	.w3(32'h380a20e3),
	.w4(32'h3bb64019),
	.w5(32'h3afd6276),
	.w6(32'hbba2246d),
	.w7(32'hbba32da8),
	.w8(32'hbbb8cf2f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf90ebf),
	.w1(32'hbbd628dc),
	.w2(32'h39b78b5c),
	.w3(32'hbb00c5bb),
	.w4(32'hbbb431bf),
	.w5(32'hbc61f5fb),
	.w6(32'hbbb4e021),
	.w7(32'hbbcfb9d3),
	.w8(32'hbc2272e6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f156d),
	.w1(32'h3ca22698),
	.w2(32'h3bae139c),
	.w3(32'hbc537cc1),
	.w4(32'hbbb428c7),
	.w5(32'hbc035f07),
	.w6(32'hbc295004),
	.w7(32'hbcf78295),
	.w8(32'hbc8d9d4b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37ca40),
	.w1(32'h3b5d1d86),
	.w2(32'hbc6b0c91),
	.w3(32'hbc967780),
	.w4(32'h3b802812),
	.w5(32'h3b0da500),
	.w6(32'hbc379df5),
	.w7(32'hbbf959d6),
	.w8(32'hbcc94677),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd11a123),
	.w1(32'hbcdc80b3),
	.w2(32'hbab5d7b2),
	.w3(32'hbac544d9),
	.w4(32'hbb750471),
	.w5(32'hbad20102),
	.w6(32'hbca34a29),
	.w7(32'hbae69e51),
	.w8(32'hba26638e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55ef62),
	.w1(32'h3a297e78),
	.w2(32'h3b867b99),
	.w3(32'h3b500bd6),
	.w4(32'h3aedcf52),
	.w5(32'hbc17c93a),
	.w6(32'h3b3aa109),
	.w7(32'h3c89e03d),
	.w8(32'h3a90a18c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8968c1),
	.w1(32'hbc35d1b3),
	.w2(32'h3c74ce10),
	.w3(32'hbc8289df),
	.w4(32'h3b225df5),
	.w5(32'hbc219a08),
	.w6(32'hbc461a99),
	.w7(32'h3b8b54b5),
	.w8(32'hbc681808),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7f263),
	.w1(32'hbc127243),
	.w2(32'hbb15d01e),
	.w3(32'hbc7c6112),
	.w4(32'hbb4894d0),
	.w5(32'hbb3a8e01),
	.w6(32'hbc8bebff),
	.w7(32'hba48f7d5),
	.w8(32'hbc5bb570),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1222d0),
	.w1(32'hbb84d12c),
	.w2(32'hbb863ae4),
	.w3(32'hbb4bacf9),
	.w4(32'hbbc74c81),
	.w5(32'hbc1ac935),
	.w6(32'hbc8629e9),
	.w7(32'h3bda0131),
	.w8(32'hbc597bab),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7953b3),
	.w1(32'hbc5b1ebf),
	.w2(32'h3ba2484d),
	.w3(32'h3bb0761a),
	.w4(32'h3b0ec7c6),
	.w5(32'hbc0143b4),
	.w6(32'hbbb2660a),
	.w7(32'hbb42e9c6),
	.w8(32'h3c321824),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c357038),
	.w1(32'h3c076c73),
	.w2(32'h3bbcf586),
	.w3(32'hbb8baab7),
	.w4(32'h3b3196f4),
	.w5(32'hbbb3c0df),
	.w6(32'hbb50c424),
	.w7(32'h3aa67d72),
	.w8(32'hbab5b5bd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7890a5),
	.w1(32'hbc6283d6),
	.w2(32'h3cb64e66),
	.w3(32'hbc6ba926),
	.w4(32'hbba22436),
	.w5(32'hbc723f18),
	.w6(32'hbc949657),
	.w7(32'h3c8069a6),
	.w8(32'hbaf75a78),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8397d8),
	.w1(32'h3c79d330),
	.w2(32'hba8dfb40),
	.w3(32'hbc86aa8c),
	.w4(32'hbbd1a6af),
	.w5(32'h3b92edb6),
	.w6(32'h3ca88c68),
	.w7(32'hbab01836),
	.w8(32'hbc034674),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa57f95),
	.w1(32'h39c4c02d),
	.w2(32'h3b1d8e1e),
	.w3(32'h3ba2598a),
	.w4(32'h3b53e1a0),
	.w5(32'hbb93e15b),
	.w6(32'hba8fb263),
	.w7(32'h3b04cdd5),
	.w8(32'h3d2551c8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59eb1d),
	.w1(32'h3c67ee1c),
	.w2(32'hbb88ac82),
	.w3(32'h3a8537c8),
	.w4(32'hbb1ead0e),
	.w5(32'hbaf709b5),
	.w6(32'h3cd1df1b),
	.w7(32'hba3d83d5),
	.w8(32'h3aa5a6d5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd28d8),
	.w1(32'h3752f009),
	.w2(32'h3c7972dd),
	.w3(32'hbae4faf2),
	.w4(32'h3a764ddc),
	.w5(32'h3c17ff69),
	.w6(32'hb9070de9),
	.w7(32'h3c000df8),
	.w8(32'hbbefd391),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b2549),
	.w1(32'h3c1d167b),
	.w2(32'h3c291993),
	.w3(32'h3c05e021),
	.w4(32'h3bd76c98),
	.w5(32'hbb96e5b5),
	.w6(32'h3b9eee49),
	.w7(32'h3c9911ee),
	.w8(32'h3aa15b2e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b04f6),
	.w1(32'h3a113807),
	.w2(32'hb9ebb1a4),
	.w3(32'hbc4ed472),
	.w4(32'h3b890efa),
	.w5(32'hbab7ad9e),
	.w6(32'hbc343049),
	.w7(32'hba6abdbb),
	.w8(32'hbb936756),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73325c),
	.w1(32'hbb89452b),
	.w2(32'h3a75b4b6),
	.w3(32'hbae4ea03),
	.w4(32'hbb98af88),
	.w5(32'hbc9d104f),
	.w6(32'hba1aecf7),
	.w7(32'h3c37f3f1),
	.w8(32'hbbbb2b4f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfe0f8),
	.w1(32'h3c3c805e),
	.w2(32'hbb0ec880),
	.w3(32'hbbea20ae),
	.w4(32'h392a1054),
	.w5(32'hb87a4808),
	.w6(32'h3c76887b),
	.w7(32'h3a97c940),
	.w8(32'h3aa21f5c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9ca5a),
	.w1(32'h3b121082),
	.w2(32'h3c912c6a),
	.w3(32'h3ab99979),
	.w4(32'h3c8bfd1b),
	.w5(32'h3b0bf879),
	.w6(32'h395c482f),
	.w7(32'h3c79ac02),
	.w8(32'hbc104b2e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b5cb6),
	.w1(32'h3c5802db),
	.w2(32'hbb903bbe),
	.w3(32'h3ac735b3),
	.w4(32'h3a48a4f4),
	.w5(32'hbb3698e1),
	.w6(32'h3b612b91),
	.w7(32'hbc10fe71),
	.w8(32'hbb2f95cb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc457d51),
	.w1(32'h3bc7e0f5),
	.w2(32'h3b8f262c),
	.w3(32'hbc6ec0c2),
	.w4(32'h3be0cd0f),
	.w5(32'h395b176e),
	.w6(32'hbc446b90),
	.w7(32'h3b585962),
	.w8(32'h3ba17819),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0882),
	.w1(32'h3bc1e2f8),
	.w2(32'hbabb67f0),
	.w3(32'hbbbbb337),
	.w4(32'hbbe3af23),
	.w5(32'h3b8a6ce0),
	.w6(32'hbb43c762),
	.w7(32'h3bd23e77),
	.w8(32'h39bf6d1d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f7bd),
	.w1(32'hbbc1c6c0),
	.w2(32'h3b1b960e),
	.w3(32'h3cc634d2),
	.w4(32'h3baeeb95),
	.w5(32'h3bfd5c7f),
	.w6(32'h3b06ab3d),
	.w7(32'h3c1deef7),
	.w8(32'h3cb046d6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule