module layer_10_featuremap_353(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97bde0),
	.w1(32'hbaf4344c),
	.w2(32'hbaddc79a),
	.w3(32'hbb0d5677),
	.w4(32'hbace2ca9),
	.w5(32'h388db8bc),
	.w6(32'hbab0d341),
	.w7(32'hbaca9ff8),
	.w8(32'h3901aa4a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03069c),
	.w1(32'h39df738e),
	.w2(32'hb86f4501),
	.w3(32'h3a179a5e),
	.w4(32'hb8a0a153),
	.w5(32'hb9d424eb),
	.w6(32'h3abaa70d),
	.w7(32'h37ece4b6),
	.w8(32'hba31fbc6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384773a4),
	.w1(32'hb93c0166),
	.w2(32'hb83cb0b1),
	.w3(32'hba3ebaf8),
	.w4(32'h388bac02),
	.w5(32'hb9860ba8),
	.w6(32'h3a7b4e39),
	.w7(32'h38926c49),
	.w8(32'hb8b40a4b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e1af3),
	.w1(32'hba144f70),
	.w2(32'hba2b753e),
	.w3(32'hba0dae0e),
	.w4(32'hb9ddd2ba),
	.w5(32'hbab6cab6),
	.w6(32'hba9ac2cc),
	.w7(32'hba57b2e2),
	.w8(32'hbb0640d9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79eac4e),
	.w1(32'hb68cacdb),
	.w2(32'h3a4145a7),
	.w3(32'hba61aca8),
	.w4(32'hb947d1d0),
	.w5(32'hb9180ef6),
	.w6(32'hbaf9f5d6),
	.w7(32'hb9e48673),
	.w8(32'hb9bd65da),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aeee5f),
	.w1(32'hb9926a65),
	.w2(32'h38c02451),
	.w3(32'hb951fe21),
	.w4(32'h38b900b7),
	.w5(32'h3ab622d8),
	.w6(32'hba207ee2),
	.w7(32'hb9bf896b),
	.w8(32'h3ab776b9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f9fc),
	.w1(32'h3ab6630e),
	.w2(32'h3a9279ae),
	.w3(32'h3ab95f62),
	.w4(32'h3aae97db),
	.w5(32'hba382a3a),
	.w6(32'h3ac0f795),
	.w7(32'h3ab51375),
	.w8(32'hbab729ba),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa69dd),
	.w1(32'hba9c5d0b),
	.w2(32'hbad17b9c),
	.w3(32'hba72a8c5),
	.w4(32'hba9d1127),
	.w5(32'hba8a22fd),
	.w6(32'hbab7e8d6),
	.w7(32'hbac833c5),
	.w8(32'hbadc6937),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa68071),
	.w1(32'hbaa09d07),
	.w2(32'hba91d437),
	.w3(32'hba46ddf5),
	.w4(32'hba676161),
	.w5(32'hb76006d9),
	.w6(32'hba89fbb3),
	.w7(32'hba5ce75b),
	.w8(32'hb9961898),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb2c9d),
	.w1(32'h3a3a4421),
	.w2(32'hb9324f4e),
	.w3(32'h37cb2cc5),
	.w4(32'h3a97d1a2),
	.w5(32'hb8f4ccb8),
	.w6(32'h37b847a2),
	.w7(32'h3a78db01),
	.w8(32'h398de138),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e05b75),
	.w1(32'hb8d9d7e3),
	.w2(32'h397041b1),
	.w3(32'h38ef67cc),
	.w4(32'hb984b010),
	.w5(32'h3aad4c7c),
	.w6(32'hb9d0274b),
	.w7(32'hba4c2dc3),
	.w8(32'h3a8bd8d6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab70273),
	.w1(32'h3a1cc98b),
	.w2(32'h3880251d),
	.w3(32'h3ab2b2a2),
	.w4(32'h3a65892a),
	.w5(32'h3858186b),
	.w6(32'h3b3c2599),
	.w7(32'h3ab03c7d),
	.w8(32'hb9aa2f4c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb4441),
	.w1(32'h39a9bb4f),
	.w2(32'hba6ef1ce),
	.w3(32'hba26105f),
	.w4(32'h3a52886f),
	.w5(32'hbae3103e),
	.w6(32'hb90d0f51),
	.w7(32'hb93852d5),
	.w8(32'hbace1f4d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fe29e),
	.w1(32'hba9f9c95),
	.w2(32'hb94b2571),
	.w3(32'hbaa30036),
	.w4(32'hba2129a6),
	.w5(32'hb9cfac83),
	.w6(32'hbb0ea60a),
	.w7(32'hba665d38),
	.w8(32'h388f3444),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84fb2b),
	.w1(32'h3a6511bd),
	.w2(32'h381902d6),
	.w3(32'h3a6f9a1a),
	.w4(32'h3a6e2375),
	.w5(32'hba355e80),
	.w6(32'h3a73bea4),
	.w7(32'h3a9554d0),
	.w8(32'hba5e489b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13bcdb),
	.w1(32'h3a8e33cc),
	.w2(32'h3921420f),
	.w3(32'h3a0e2c0c),
	.w4(32'h3a9ba2bf),
	.w5(32'h395a200c),
	.w6(32'hb98633fa),
	.w7(32'h3a85e39d),
	.w8(32'hb9650365),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0cd7e),
	.w1(32'hb84ac3e5),
	.w2(32'h3a00ec65),
	.w3(32'h3861058a),
	.w4(32'hb8c2be9d),
	.w5(32'hb9045c52),
	.w6(32'hba25f467),
	.w7(32'hb9349293),
	.w8(32'h39298a72),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba501ec7),
	.w1(32'hb91941a6),
	.w2(32'hb93a5416),
	.w3(32'hb99100f9),
	.w4(32'hb9f4b165),
	.w5(32'h3ac378a1),
	.w6(32'h3a2d96fc),
	.w7(32'hb8c397e4),
	.w8(32'h3b03ec16),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95b648),
	.w1(32'h3b1e162f),
	.w2(32'h3b0d9ac2),
	.w3(32'h3b211965),
	.w4(32'h3b1ad0be),
	.w5(32'hba6272a3),
	.w6(32'h3b197743),
	.w7(32'h3b3e84a1),
	.w8(32'hb9e293a5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a46fd2),
	.w1(32'hba0d6860),
	.w2(32'hb7e70807),
	.w3(32'hb9e3957b),
	.w4(32'hb939dae2),
	.w5(32'hb960b73e),
	.w6(32'hba99ee09),
	.w7(32'hb9a3e72b),
	.w8(32'hba276aa4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dd304),
	.w1(32'hb9d13945),
	.w2(32'hb89c61dc),
	.w3(32'hb9137212),
	.w4(32'h39b95ba1),
	.w5(32'h3957919f),
	.w6(32'hba626526),
	.w7(32'h38fc56f5),
	.w8(32'h38db57fd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907bcf3),
	.w1(32'hba720a0d),
	.w2(32'hba72fe66),
	.w3(32'h38ab69fc),
	.w4(32'h382e1c46),
	.w5(32'hba07bf64),
	.w6(32'hb905201c),
	.w7(32'h3858ab7c),
	.w8(32'hb9c82b92),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d754a),
	.w1(32'h3a4d941a),
	.w2(32'h390404da),
	.w3(32'hb9e6dd9b),
	.w4(32'h3aeaabaa),
	.w5(32'h39dc6c0a),
	.w6(32'h3a8bf0b8),
	.w7(32'h3a684cf9),
	.w8(32'hba77e2df),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39162b24),
	.w1(32'h3ad41208),
	.w2(32'hb98c1d07),
	.w3(32'hb713aceb),
	.w4(32'h3ab73846),
	.w5(32'hba339e15),
	.w6(32'h3b0987b7),
	.w7(32'h3ae3bb41),
	.w8(32'hb8e1f993),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc60e2),
	.w1(32'hba9ed7e3),
	.w2(32'hbac8ee95),
	.w3(32'h384bf38c),
	.w4(32'hb9c7c1fd),
	.w5(32'hb8705859),
	.w6(32'h3a8217a1),
	.w7(32'hb96d1d5a),
	.w8(32'h3a6c2a7a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985d829),
	.w1(32'h3a2cd4f5),
	.w2(32'h39fb0806),
	.w3(32'hb9e5c403),
	.w4(32'h384b21b0),
	.w5(32'h3a851b77),
	.w6(32'hbab07e36),
	.w7(32'h3984931d),
	.w8(32'hb917a15c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39465835),
	.w1(32'h3a15fb02),
	.w2(32'h3ab1eb3c),
	.w3(32'h3984c5fa),
	.w4(32'h3a336ba5),
	.w5(32'hbafbbb39),
	.w6(32'hba6e43a1),
	.w7(32'h3a40025f),
	.w8(32'hbb11186b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097ba8),
	.w1(32'hbb40360f),
	.w2(32'hbb054a85),
	.w3(32'hbb16075c),
	.w4(32'hbad64620),
	.w5(32'hbacd7636),
	.w6(32'hbb2be821),
	.w7(32'hbb02b05f),
	.w8(32'hbaa69df6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c502e),
	.w1(32'hbaf9189f),
	.w2(32'hba887f83),
	.w3(32'hba7019aa),
	.w4(32'hba36940e),
	.w5(32'hba798759),
	.w6(32'hbaa3e5b4),
	.w7(32'hb8e5654c),
	.w8(32'hb8d23854),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f2a76),
	.w1(32'h3a428f72),
	.w2(32'h393a367a),
	.w3(32'hba667a08),
	.w4(32'h3a0fed6e),
	.w5(32'hba1e5361),
	.w6(32'h394e064e),
	.w7(32'h399b262f),
	.w8(32'h39c29e26),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8a8d1),
	.w1(32'h3a7c018c),
	.w2(32'h3ad9d78f),
	.w3(32'hb9d2dfd8),
	.w4(32'h38a24cf2),
	.w5(32'h38b6fdf8),
	.w6(32'h3a6dd1e2),
	.w7(32'h3a65b422),
	.w8(32'hb9a7d292),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96091a9),
	.w1(32'hba121db2),
	.w2(32'hb9d9f590),
	.w3(32'hb90db171),
	.w4(32'h3a6aacc5),
	.w5(32'h3a966b62),
	.w6(32'hb8f787cd),
	.w7(32'hb992bbef),
	.w8(32'h3ad48003),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8757ea),
	.w1(32'h3ab3c4f7),
	.w2(32'h3a2d847d),
	.w3(32'h3aa33fb0),
	.w4(32'h398ed7b9),
	.w5(32'hba6ce55f),
	.w6(32'h3ac3870e),
	.w7(32'h3a9913e0),
	.w8(32'hba4987f2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5bbb0),
	.w1(32'hba987c3d),
	.w2(32'hbaa1c11a),
	.w3(32'hb9bfa28d),
	.w4(32'hbab7a5b7),
	.w5(32'hba811fa1),
	.w6(32'hb94e1ca6),
	.w7(32'hbaedcbae),
	.w8(32'hba949d45),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a61fc),
	.w1(32'hba7b2756),
	.w2(32'hbac2f09f),
	.w3(32'hbad1afb1),
	.w4(32'hbacc15d9),
	.w5(32'h37ce08b0),
	.w6(32'hbae09a5b),
	.w7(32'hbaf7444d),
	.w8(32'h39e5f390),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169fc4),
	.w1(32'h3ab6bc39),
	.w2(32'h3a1fa20b),
	.w3(32'h3a0cde21),
	.w4(32'hb9862b6d),
	.w5(32'h37bc4355),
	.w6(32'h3aff9a52),
	.w7(32'h3a4848c8),
	.w8(32'hb9a44e64),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8471e4),
	.w1(32'h39d89def),
	.w2(32'h3a958bbd),
	.w3(32'hba9b24ae),
	.w4(32'h3a3a5880),
	.w5(32'h3b0fc265),
	.w6(32'hba956de1),
	.w7(32'h3a06c019),
	.w8(32'h3b1fe598),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f45781),
	.w1(32'hbabcb85d),
	.w2(32'hba958661),
	.w3(32'h37fa9cad),
	.w4(32'hba678bf3),
	.w5(32'hba970f1e),
	.w6(32'h39e36f9d),
	.w7(32'h39a12d50),
	.w8(32'h3a14730f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b75a09),
	.w1(32'hbac18fbe),
	.w2(32'hbacbb934),
	.w3(32'hba646b2d),
	.w4(32'hbadbf0f1),
	.w5(32'hba066711),
	.w6(32'h3b15f7fc),
	.w7(32'h3a1af9fb),
	.w8(32'h3a551295),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19d4ac),
	.w1(32'h386c93fa),
	.w2(32'h394b6689),
	.w3(32'h3a8f120e),
	.w4(32'h3a0cb15d),
	.w5(32'h39e7f116),
	.w6(32'hb96899ef),
	.w7(32'h39be245b),
	.w8(32'h39c0e48c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a0ccc),
	.w1(32'hb9723039),
	.w2(32'hb9b71300),
	.w3(32'hb9a120dd),
	.w4(32'hba19a391),
	.w5(32'h3a26ce9d),
	.w6(32'h3825b8ee),
	.w7(32'hba3bdcfe),
	.w8(32'h3a60ce56),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e0536),
	.w1(32'hb9628b60),
	.w2(32'hb969aac2),
	.w3(32'h388b0aa3),
	.w4(32'h3985e2d5),
	.w5(32'h39fcd431),
	.w6(32'hba81790f),
	.w7(32'hb8fbf0e4),
	.w8(32'h3aa07413),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a9496),
	.w1(32'h3a89943a),
	.w2(32'h3a6f3fac),
	.w3(32'h390c2bd3),
	.w4(32'hbaa2d9b7),
	.w5(32'hb9af16c9),
	.w6(32'h3ab7385e),
	.w7(32'hb924c21c),
	.w8(32'hb9dfeced),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c3427),
	.w1(32'h3a9f9f5a),
	.w2(32'h3aa4492a),
	.w3(32'h3a600728),
	.w4(32'hb84adc4b),
	.w5(32'hbb22478c),
	.w6(32'hba2aa181),
	.w7(32'h3a9ebb57),
	.w8(32'hbad0c4c4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda1b6),
	.w1(32'hbaf98886),
	.w2(32'hbb0cf72c),
	.w3(32'hbb07c3f8),
	.w4(32'hba880fb6),
	.w5(32'h3ad9956f),
	.w6(32'hbb5ea0a3),
	.w7(32'hbabe3c86),
	.w8(32'h3b06af73),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a344f4),
	.w1(32'h393f3b7c),
	.w2(32'h39c6a206),
	.w3(32'h3acedf41),
	.w4(32'h3b2961df),
	.w5(32'h395599e2),
	.w6(32'h3ab0fe8b),
	.w7(32'h3b513dc6),
	.w8(32'h3a04a57a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4e2bb),
	.w1(32'hb9f04b9e),
	.w2(32'h39f07f75),
	.w3(32'h3aa0813c),
	.w4(32'h3add61fd),
	.w5(32'hb9e79c04),
	.w6(32'hb9715433),
	.w7(32'h3aacd77f),
	.w8(32'hba8197d8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba861fec),
	.w1(32'h393a8aff),
	.w2(32'hb9f82b89),
	.w3(32'hba5114b0),
	.w4(32'h3aa5ea33),
	.w5(32'hbac723ac),
	.w6(32'hbabbb03d),
	.w7(32'h3a23030a),
	.w8(32'hba92e7de),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15fd6b),
	.w1(32'hbb2acfd4),
	.w2(32'hbb33b193),
	.w3(32'hbb17cd35),
	.w4(32'hbb0b657e),
	.w5(32'h398ed74c),
	.w6(32'hbacd2bde),
	.w7(32'hbb4d0971),
	.w8(32'h3829d6b6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b1a04),
	.w1(32'hb9049fe1),
	.w2(32'hb9c13abe),
	.w3(32'h3a17d54a),
	.w4(32'h39cd0e9a),
	.w5(32'hbaba453b),
	.w6(32'h3790f6a8),
	.w7(32'hb91cb8ab),
	.w8(32'hbb1f4ce0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7f0fa),
	.w1(32'hba828fd0),
	.w2(32'h3a2a5b04),
	.w3(32'hbac1ead1),
	.w4(32'hba7d6732),
	.w5(32'h3905c77e),
	.w6(32'hbad3c269),
	.w7(32'h3677c256),
	.w8(32'h39c3e19f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4bdec),
	.w1(32'h3aa01d64),
	.w2(32'h3a93bea5),
	.w3(32'hba8659c9),
	.w4(32'h3a64f1dc),
	.w5(32'hba0b0799),
	.w6(32'h39160a94),
	.w7(32'h394cdd4e),
	.w8(32'h38460f6c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840cb68),
	.w1(32'hb9a40420),
	.w2(32'hba1779f1),
	.w3(32'hbaa491a0),
	.w4(32'hba284218),
	.w5(32'hb9b8680b),
	.w6(32'hb970d291),
	.w7(32'hb9b3f298),
	.w8(32'hb85e8b15),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d54662),
	.w1(32'h3a6f073b),
	.w2(32'hb71c8de7),
	.w3(32'h3a5fdfca),
	.w4(32'h3adc07a7),
	.w5(32'h3a9e8486),
	.w6(32'h3b0fd41c),
	.w7(32'h3ab85707),
	.w8(32'h3a946374),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a6f3c),
	.w1(32'h399e0e54),
	.w2(32'h39aa6dbc),
	.w3(32'h390dfdaa),
	.w4(32'hb99ae173),
	.w5(32'hbaa165c2),
	.w6(32'hb848cd27),
	.w7(32'hb9f24aee),
	.w8(32'hba7d23ed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0a218),
	.w1(32'hba21bceb),
	.w2(32'hba5d78af),
	.w3(32'hba9ccf4d),
	.w4(32'hb9ebf34d),
	.w5(32'hba6eaac8),
	.w6(32'hbafe947f),
	.w7(32'hbaa0ab66),
	.w8(32'hba3a86fa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba783808),
	.w1(32'hbab13659),
	.w2(32'hbac7e019),
	.w3(32'hba8f642e),
	.w4(32'hba82d7cf),
	.w5(32'h39a652a3),
	.w6(32'hbabdf136),
	.w7(32'hbae2d3d9),
	.w8(32'h39faeff8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d22f),
	.w1(32'h399f5a0f),
	.w2(32'hb8ece121),
	.w3(32'h3935604c),
	.w4(32'hb7d8a04b),
	.w5(32'h39d84542),
	.w6(32'h398fca86),
	.w7(32'hb8f554c2),
	.w8(32'h39608edf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f89f70),
	.w1(32'h3940dd43),
	.w2(32'hb7d39dea),
	.w3(32'h39d0b45b),
	.w4(32'h39c577c4),
	.w5(32'h3aa3629b),
	.w6(32'h392e5132),
	.w7(32'h39906fb2),
	.w8(32'h39eb28cc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b5ee2),
	.w1(32'hba692748),
	.w2(32'hba49564c),
	.w3(32'h3a6d598a),
	.w4(32'h3a667e0a),
	.w5(32'hb947340e),
	.w6(32'hbb056b5b),
	.w7(32'hba835754),
	.w8(32'hb923d53f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c9d82),
	.w1(32'h37001c1f),
	.w2(32'hb9ebf15c),
	.w3(32'hb8f3520f),
	.w4(32'hba56db75),
	.w5(32'hb940c083),
	.w6(32'hb91a632c),
	.w7(32'h38021cad),
	.w8(32'hb9edd1fb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c1c15),
	.w1(32'hba8fe5dd),
	.w2(32'hb963dff9),
	.w3(32'hba9ebbf4),
	.w4(32'hb9ab2a3f),
	.w5(32'h3915311f),
	.w6(32'hbad9bd9a),
	.w7(32'hba104d32),
	.w8(32'hba7b1204),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7874c7),
	.w1(32'hba496c4b),
	.w2(32'hb92e8741),
	.w3(32'hba8cf5a9),
	.w4(32'hba6b2b49),
	.w5(32'hb89a4e4b),
	.w6(32'hbaecbb95),
	.w7(32'hbadcf575),
	.w8(32'hb9651697),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd06ba),
	.w1(32'hb9ccef8b),
	.w2(32'hba5c4d66),
	.w3(32'hba338dcc),
	.w4(32'hb9ee4e5e),
	.w5(32'hba6663df),
	.w6(32'hba45626a),
	.w7(32'hbaa2a3d6),
	.w8(32'hba6eefe5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8675ae),
	.w1(32'h38846549),
	.w2(32'hb9bc465c),
	.w3(32'hba63e94c),
	.w4(32'hba612c53),
	.w5(32'hb98fde60),
	.w6(32'hba563128),
	.w7(32'hba900ae8),
	.w8(32'hba6e7a26),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0149d9),
	.w1(32'h3a22ff31),
	.w2(32'h3a01ad80),
	.w3(32'hba393405),
	.w4(32'hba17ddc3),
	.w5(32'hb83150a6),
	.w6(32'hb9bf39f2),
	.w7(32'hba4c8f62),
	.w8(32'hba4bcf7d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5bcd),
	.w1(32'hba8f4cd6),
	.w2(32'hbaa5c929),
	.w3(32'hba059ca5),
	.w4(32'hba80d2e8),
	.w5(32'h398f7c14),
	.w6(32'hba7d7eb6),
	.w7(32'hbae339ed),
	.w8(32'hba03ae97),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d2be9),
	.w1(32'hb8647c88),
	.w2(32'h3a1bfa29),
	.w3(32'h3acffe87),
	.w4(32'h3a951bf2),
	.w5(32'h39672289),
	.w6(32'h3a51f75f),
	.w7(32'h3acbd20b),
	.w8(32'h3a67b234),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980f6cb),
	.w1(32'hb9a72667),
	.w2(32'hbaac27ad),
	.w3(32'h38a34471),
	.w4(32'hba537dda),
	.w5(32'h3a4bcad0),
	.w6(32'h3a9d9e59),
	.w7(32'h380fdebc),
	.w8(32'h3ad35de6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393fbf24),
	.w1(32'h38879ccb),
	.w2(32'hba4cc200),
	.w3(32'h3a8aa201),
	.w4(32'h3a25e89b),
	.w5(32'h3a4fdad1),
	.w6(32'h3a92c8f5),
	.w7(32'h39736740),
	.w8(32'h3acbf072),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff2dc8),
	.w1(32'h39b0ce69),
	.w2(32'h39b9454d),
	.w3(32'h39244c96),
	.w4(32'hb944453c),
	.w5(32'h396e488b),
	.w6(32'h386139af),
	.w7(32'h398ba624),
	.w8(32'hba04cc44),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b87c34),
	.w1(32'h3a65c93e),
	.w2(32'h3a923c94),
	.w3(32'hb910f6bc),
	.w4(32'h3a03e17d),
	.w5(32'hb94b2e0c),
	.w6(32'h36f73791),
	.w7(32'h3aef984f),
	.w8(32'hb9c1e190),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c54702),
	.w1(32'h3ab3f83e),
	.w2(32'h399e5a2a),
	.w3(32'hb907eea1),
	.w4(32'hba334cb2),
	.w5(32'hb9c32854),
	.w6(32'h3a211f50),
	.w7(32'hb806faca),
	.w8(32'hba0f64c9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446997),
	.w1(32'hba477c8e),
	.w2(32'hba1d2413),
	.w3(32'hb9323abf),
	.w4(32'hb7baab45),
	.w5(32'hb9acc4ff),
	.w6(32'hba62dbe0),
	.w7(32'hba93feb5),
	.w8(32'hbaab105d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33c4b8),
	.w1(32'hba50e1a2),
	.w2(32'hba58c340),
	.w3(32'hba0b89a3),
	.w4(32'hba93756b),
	.w5(32'h39d30180),
	.w6(32'hba427c41),
	.w7(32'hbaf13c61),
	.w8(32'h3a25b172),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38959e49),
	.w1(32'hb90105da),
	.w2(32'hb90ac0bc),
	.w3(32'h39f11c9b),
	.w4(32'h39e5b067),
	.w5(32'h3a0a55e1),
	.w6(32'h3a34fd43),
	.w7(32'hb92c085a),
	.w8(32'hb922c8c7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab833e4),
	.w1(32'h3a33c501),
	.w2(32'h37b52fad),
	.w3(32'h39b45865),
	.w4(32'hb8b50373),
	.w5(32'hb995c132),
	.w6(32'h398f8084),
	.w7(32'h3999641a),
	.w8(32'h39cea3bb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2817ab),
	.w1(32'h3a3ef24f),
	.w2(32'hb818aaa5),
	.w3(32'hb98b61c5),
	.w4(32'hb99867c5),
	.w5(32'hb84baa11),
	.w6(32'hb9f8d61a),
	.w7(32'hba053f29),
	.w8(32'h3a3af06c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5189b4),
	.w1(32'h3a568d36),
	.w2(32'h39d2b4c9),
	.w3(32'h3a9213d2),
	.w4(32'h3aa8fc6a),
	.w5(32'hba656bee),
	.w6(32'h3a766c4c),
	.w7(32'h3a287a7c),
	.w8(32'hbae2cb12),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29baa),
	.w1(32'hba69647b),
	.w2(32'hb9926d56),
	.w3(32'hba24424c),
	.w4(32'hba13f3e8),
	.w5(32'hbac8f09c),
	.w6(32'hba9d6bd6),
	.w7(32'hba5c4d02),
	.w8(32'hbaea3640),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a06c),
	.w1(32'hbb70c410),
	.w2(32'hbb825bbd),
	.w3(32'hbb15824e),
	.w4(32'hbafa0583),
	.w5(32'hba6ec8ca),
	.w6(32'hbb674c78),
	.w7(32'hbb1fc048),
	.w8(32'hb90e7609),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba640820),
	.w1(32'hb7bdbae2),
	.w2(32'hba2e74e9),
	.w3(32'hba53131b),
	.w4(32'hba6a60d1),
	.w5(32'h38d405ad),
	.w6(32'h379554cb),
	.w7(32'hba91a8d6),
	.w8(32'hb9eac447),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc1c6f),
	.w1(32'h3a4dcfc5),
	.w2(32'hba2c6f0c),
	.w3(32'hb9c1138d),
	.w4(32'hb9f4f7dd),
	.w5(32'h3abbed6b),
	.w6(32'h3a5d1ede),
	.w7(32'hb948ab04),
	.w8(32'h3a3087b7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e52b2),
	.w1(32'h3acc3aee),
	.w2(32'h3ae571d5),
	.w3(32'h3aafa0a1),
	.w4(32'h3ab68104),
	.w5(32'hba66c5cc),
	.w6(32'h3a3228bc),
	.w7(32'h3ad5dbc9),
	.w8(32'hba8c70c4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3804e5e2),
	.w1(32'h3947b45e),
	.w2(32'hba83b71e),
	.w3(32'hba955162),
	.w4(32'hba287a09),
	.w5(32'hb9cff1aa),
	.w6(32'hb8c650c3),
	.w7(32'hba2a64c1),
	.w8(32'hb9811b06),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96600ec),
	.w1(32'hbb04317d),
	.w2(32'hba358f45),
	.w3(32'hb9fcc23c),
	.w4(32'hb9169a03),
	.w5(32'h3a5e9f13),
	.w6(32'hba926fa6),
	.w7(32'hba06b0d5),
	.w8(32'h3a0e065f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f1dd4),
	.w1(32'h38323b63),
	.w2(32'hb9da645d),
	.w3(32'h3981b639),
	.w4(32'hba293c35),
	.w5(32'hb93a7df5),
	.w6(32'h3aac47b4),
	.w7(32'h3a2c9da5),
	.w8(32'hb9cf6d12),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3802da75),
	.w1(32'hb95820a1),
	.w2(32'h38e6243c),
	.w3(32'hb91c2aa4),
	.w4(32'hb9b26dd8),
	.w5(32'h3a243d8c),
	.w6(32'hb9ecda9d),
	.w7(32'hb7d7ab99),
	.w8(32'h38c09807),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53464c),
	.w1(32'h3ac3a54e),
	.w2(32'h3a82d7d9),
	.w3(32'h3a864e1e),
	.w4(32'h3ac07dc2),
	.w5(32'hb998629d),
	.w6(32'h3a4e34f0),
	.w7(32'h3abdca35),
	.w8(32'h39aae7d0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74641f),
	.w1(32'hb9225a04),
	.w2(32'h396a2b13),
	.w3(32'hbb0e17c2),
	.w4(32'hba945050),
	.w5(32'hba1f9149),
	.w6(32'hbad3656c),
	.w7(32'hba9003ec),
	.w8(32'hba7b066f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446127),
	.w1(32'hb9f20d4f),
	.w2(32'hba27a881),
	.w3(32'h3846f6c2),
	.w4(32'hb9b9f7a3),
	.w5(32'h3a3873cb),
	.w6(32'h3a84a9e9),
	.w7(32'hb875503a),
	.w8(32'h3a2d170f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c78173),
	.w1(32'h3918019a),
	.w2(32'h3a03f886),
	.w3(32'hba1bf4f2),
	.w4(32'hb9803d67),
	.w5(32'hba2e77e1),
	.w6(32'hba3a77d6),
	.w7(32'h36e569ea),
	.w8(32'hba87f67d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cfbc3),
	.w1(32'hba5b6ecc),
	.w2(32'hba04aba5),
	.w3(32'hba72e030),
	.w4(32'hba1e5ef9),
	.w5(32'h3a251dfa),
	.w6(32'hbac6f11c),
	.w7(32'hba431e8c),
	.w8(32'h3a364636),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81302f),
	.w1(32'h3b1176e6),
	.w2(32'h3ad57fd3),
	.w3(32'h3b22a55e),
	.w4(32'h3b4da968),
	.w5(32'h3a86f6e4),
	.w6(32'h3ae3cc71),
	.w7(32'h3ad705e4),
	.w8(32'h3947d3d3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50cefa),
	.w1(32'h3a48e671),
	.w2(32'h38c9844d),
	.w3(32'h39bdfa07),
	.w4(32'h390d0d2b),
	.w5(32'h3a9adc2e),
	.w6(32'h372c063a),
	.w7(32'h3a0cc6e4),
	.w8(32'h3a9500a9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b1ee6),
	.w1(32'h3b85c106),
	.w2(32'h3b577294),
	.w3(32'h3acbba3d),
	.w4(32'h3a875b71),
	.w5(32'h3a1d6090),
	.w6(32'h3b14dff9),
	.w7(32'h3b029a18),
	.w8(32'h3a94810a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06eb65),
	.w1(32'hb995ea11),
	.w2(32'h39592010),
	.w3(32'h3a88da80),
	.w4(32'h3a95a904),
	.w5(32'h3a1217d9),
	.w6(32'hb9dec6db),
	.w7(32'h39ddcfb2),
	.w8(32'h3a36649c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8607b),
	.w1(32'h3a1d6631),
	.w2(32'h39b86ea1),
	.w3(32'h3a4bd438),
	.w4(32'h3ad6a84f),
	.w5(32'hba4996dd),
	.w6(32'h3ac88a59),
	.w7(32'h3ae05f72),
	.w8(32'hbaaae10c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e68d3),
	.w1(32'h3b1abc1b),
	.w2(32'h3ba65228),
	.w3(32'hbab57967),
	.w4(32'h3b1c5a4a),
	.w5(32'hbbcbcca4),
	.w6(32'hb9282355),
	.w7(32'h3bc6baba),
	.w8(32'h3b531540),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44a2f6),
	.w1(32'h3b8d693b),
	.w2(32'hbb6a6168),
	.w3(32'h3af1aa77),
	.w4(32'h3ae57456),
	.w5(32'hbbab8d33),
	.w6(32'h3bc6d927),
	.w7(32'hbb08d3ae),
	.w8(32'hbb310d08),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0e14),
	.w1(32'hbbaf2ffe),
	.w2(32'h3acc2acd),
	.w3(32'hbbbda2bc),
	.w4(32'hbb179193),
	.w5(32'h3b636d1b),
	.w6(32'hbb966fe4),
	.w7(32'hbb458caf),
	.w8(32'h3ac73c38),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c0e29),
	.w1(32'h3a849c3a),
	.w2(32'h3a885c15),
	.w3(32'h3b1520a5),
	.w4(32'h38f6e422),
	.w5(32'h38ed06da),
	.w6(32'h3c823e18),
	.w7(32'h3bc46896),
	.w8(32'hba4e1e2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d456f9),
	.w1(32'h3b81a940),
	.w2(32'hbab793e3),
	.w3(32'h3b8fc554),
	.w4(32'h3b7ee43a),
	.w5(32'h3b468fa8),
	.w6(32'h3bc22a7d),
	.w7(32'hba5ad4e1),
	.w8(32'h3bc6c318),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad08ff),
	.w1(32'hbbec1bc9),
	.w2(32'h395a05f6),
	.w3(32'hbb9822ee),
	.w4(32'hbaccbdfd),
	.w5(32'h3b4d67bd),
	.w6(32'hb77af42d),
	.w7(32'hba070c29),
	.w8(32'h3a9d1716),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb280ee),
	.w1(32'hbbeaf33f),
	.w2(32'h3b3505ae),
	.w3(32'hbc4bc096),
	.w4(32'hb9bb596a),
	.w5(32'hbb1bd1a1),
	.w6(32'h3c1b5292),
	.w7(32'h3b00aed9),
	.w8(32'h3b764e68),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab815ae),
	.w1(32'h3be3bd77),
	.w2(32'h3b470feb),
	.w3(32'hbb5af3e2),
	.w4(32'hba1a1731),
	.w5(32'h3b5a6cb7),
	.w6(32'hbbac214b),
	.w7(32'h3b182ca3),
	.w8(32'h3b6998ae),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac46dd9),
	.w1(32'h3a7ddfa0),
	.w2(32'h3c05dce7),
	.w3(32'hbb16e30f),
	.w4(32'hbb183899),
	.w5(32'hbb229bbe),
	.w6(32'hbc0f4b3d),
	.w7(32'hbad4ce6e),
	.w8(32'hbb7a1612),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6499ee),
	.w1(32'h3b98f652),
	.w2(32'h3ae8bbe6),
	.w3(32'h3b2c1589),
	.w4(32'h3b1ccceb),
	.w5(32'hb95fd987),
	.w6(32'h3bfee761),
	.w7(32'h3adf06fe),
	.w8(32'hb9181b72),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de287),
	.w1(32'h3b7ce54f),
	.w2(32'h3bec043c),
	.w3(32'hbad9c9b0),
	.w4(32'h3b6bb906),
	.w5(32'hbb917629),
	.w6(32'hbb81393d),
	.w7(32'h3b9b9a4e),
	.w8(32'hbb2480b2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90b9c),
	.w1(32'hba838c58),
	.w2(32'hbb828b5a),
	.w3(32'hbaf6953f),
	.w4(32'hbba58d72),
	.w5(32'h3b5f32b6),
	.w6(32'h38bee7a2),
	.w7(32'hbb08dc8b),
	.w8(32'hba101d07),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec8c97),
	.w1(32'h3be1569a),
	.w2(32'h3aea8570),
	.w3(32'h3b3d3e7f),
	.w4(32'h3b684be7),
	.w5(32'h3ac9744a),
	.w6(32'h3a5344e5),
	.w7(32'h393d2773),
	.w8(32'hba12ed26),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aeeda),
	.w1(32'hba7fdf5e),
	.w2(32'h3acbaa35),
	.w3(32'h3ba0365f),
	.w4(32'h3bb245d1),
	.w5(32'h3ab792a9),
	.w6(32'h3aa78c36),
	.w7(32'hb98b7112),
	.w8(32'hbadbc8df),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb53c),
	.w1(32'hbadf618b),
	.w2(32'hba8257bc),
	.w3(32'h3996faa2),
	.w4(32'hbb5f8d41),
	.w5(32'hbb59ccbd),
	.w6(32'h3afa9942),
	.w7(32'hbb911905),
	.w8(32'h399f1585),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a287e),
	.w1(32'h3a0827c5),
	.w2(32'h3aa0e1f0),
	.w3(32'hbb9ee1c8),
	.w4(32'hbb000887),
	.w5(32'hbb5b7b0e),
	.w6(32'h3a424b59),
	.w7(32'hbafd13af),
	.w8(32'hba81d891),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92684c),
	.w1(32'h3ba44f20),
	.w2(32'hb938c5f6),
	.w3(32'hbb3b7b7e),
	.w4(32'hbbbf12e3),
	.w5(32'h3b40cfd3),
	.w6(32'hbb9bd7c2),
	.w7(32'h3b80962e),
	.w8(32'h3ab4db91),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342d57),
	.w1(32'h3b4eade6),
	.w2(32'h3a2b187e),
	.w3(32'h3b2c6b88),
	.w4(32'h3b9d7975),
	.w5(32'h3a3712a8),
	.w6(32'h3c13ff30),
	.w7(32'h3afd736a),
	.w8(32'hbb83fc7e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa08849),
	.w1(32'h3b918ba2),
	.w2(32'h39ef93eb),
	.w3(32'hba83c5de),
	.w4(32'h3af0ec14),
	.w5(32'h3b24f742),
	.w6(32'hbaa7282d),
	.w7(32'h3b3dd778),
	.w8(32'h3c027e41),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d4e7),
	.w1(32'h3ac9a322),
	.w2(32'h3b7f2628),
	.w3(32'hbbc82f3b),
	.w4(32'hbb0cb750),
	.w5(32'h3afa1db4),
	.w6(32'h3b32487c),
	.w7(32'h3ad04877),
	.w8(32'h3af80e34),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0633),
	.w1(32'h3b8436ac),
	.w2(32'h388b5c83),
	.w3(32'h39b576f9),
	.w4(32'h39ad067d),
	.w5(32'h3a40ebe1),
	.w6(32'h3b3d7fed),
	.w7(32'h3b888834),
	.w8(32'hb96de29e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba695ef),
	.w1(32'hb8c220b9),
	.w2(32'h3ba96f5a),
	.w3(32'hba7e5995),
	.w4(32'h398d6e40),
	.w5(32'h3a5941aa),
	.w6(32'hbc1d2a2e),
	.w7(32'h3b966599),
	.w8(32'hbac4c4bc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b9de1),
	.w1(32'hbb3b6835),
	.w2(32'hbb350759),
	.w3(32'h386259b2),
	.w4(32'hbb5427b7),
	.w5(32'hbb617ab5),
	.w6(32'hbadd4728),
	.w7(32'hba7b09ec),
	.w8(32'hbae93749),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a747050),
	.w1(32'hbb9fe0cb),
	.w2(32'hbb2b70a0),
	.w3(32'h39a8fd84),
	.w4(32'h39d5e9ea),
	.w5(32'hbb0ff464),
	.w6(32'hbb2b150f),
	.w7(32'hba12d517),
	.w8(32'h3c33b4f8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeca076),
	.w1(32'hbbb0e9bb),
	.w2(32'h3bdbe5aa),
	.w3(32'h3c02c9a3),
	.w4(32'h3bee7daa),
	.w5(32'hbb61e983),
	.w6(32'h3c696a5e),
	.w7(32'h3b0396a1),
	.w8(32'hbbb56792),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce769),
	.w1(32'hbbfc83fc),
	.w2(32'hbb4b004f),
	.w3(32'hba8eb498),
	.w4(32'hbb9ec8a8),
	.w5(32'hbc02c1d5),
	.w6(32'hba1b4009),
	.w7(32'hbbb2762e),
	.w8(32'h3b84daf6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb451b),
	.w1(32'h3b157df3),
	.w2(32'hbb32b0fa),
	.w3(32'hba130816),
	.w4(32'h3b04b5ab),
	.w5(32'hbb5d6b74),
	.w6(32'h3c49c363),
	.w7(32'h39b0818d),
	.w8(32'hbb117599),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b939a),
	.w1(32'hbb9c03e9),
	.w2(32'hbb5f5cdd),
	.w3(32'hbb1b135b),
	.w4(32'hba86e6b9),
	.w5(32'hbb3e22ee),
	.w6(32'h3b5ab2c1),
	.w7(32'h3ab43f6a),
	.w8(32'hbb8f3d7d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518be2),
	.w1(32'h3a676dbe),
	.w2(32'hb9252d55),
	.w3(32'hbb8b2bce),
	.w4(32'hbb407486),
	.w5(32'hbaf5d45e),
	.w6(32'hb9195cad),
	.w7(32'h3aac17d2),
	.w8(32'h3a4202a7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae192de),
	.w1(32'hbbe7688a),
	.w2(32'hb9e4b7e6),
	.w3(32'h39826f8c),
	.w4(32'h3a75ea62),
	.w5(32'hbbe09d51),
	.w6(32'hbb840716),
	.w7(32'h39a183d2),
	.w8(32'h38f35cb7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f5aa1),
	.w1(32'hbb36a0f5),
	.w2(32'hbb0dee08),
	.w3(32'hbc03867e),
	.w4(32'hbb499df5),
	.w5(32'h3a59ac69),
	.w6(32'hbb302c0a),
	.w7(32'hbafc30e8),
	.w8(32'hbb19a9cd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147a1c),
	.w1(32'h38599032),
	.w2(32'h39ceceb8),
	.w3(32'hbb5a7eeb),
	.w4(32'hbb3c0d19),
	.w5(32'h3b251446),
	.w6(32'h39ff8f95),
	.w7(32'hba9ea0ff),
	.w8(32'hbbb10f1d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b255454),
	.w1(32'h3b8a0b62),
	.w2(32'h3ba50467),
	.w3(32'hbb2b9b71),
	.w4(32'hbad2dc2e),
	.w5(32'h3b940958),
	.w6(32'h3b709598),
	.w7(32'hba0fa350),
	.w8(32'h3b89f0f3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e8786),
	.w1(32'h3bef9461),
	.w2(32'h3b5b36ce),
	.w3(32'h3b8a5255),
	.w4(32'h3b6a337f),
	.w5(32'hbb2d32a7),
	.w6(32'h3b3bc462),
	.w7(32'h3b88dbe7),
	.w8(32'hbab1834a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cc8cd),
	.w1(32'h396b6424),
	.w2(32'hbac3f4a1),
	.w3(32'h3b828e0e),
	.w4(32'h3b59f5d2),
	.w5(32'hbb48e221),
	.w6(32'h3bce28c4),
	.w7(32'h3bb2571f),
	.w8(32'hbb57b770),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39876cc1),
	.w1(32'h3b46f00a),
	.w2(32'hbb00cab3),
	.w3(32'hba74925e),
	.w4(32'hbb3caa94),
	.w5(32'hbab8357b),
	.w6(32'h3be33072),
	.w7(32'hb8dcf837),
	.w8(32'hbba3d524),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71477e),
	.w1(32'h3ba9d7cb),
	.w2(32'h3a3f1aaa),
	.w3(32'hbaec572c),
	.w4(32'h3ae98144),
	.w5(32'h3b313bef),
	.w6(32'h3b9c2b39),
	.w7(32'h3b51d2da),
	.w8(32'hbb7773c3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc0691),
	.w1(32'h3c2b6870),
	.w2(32'h3bd27f76),
	.w3(32'h398e6c26),
	.w4(32'h3b44d130),
	.w5(32'hba6a3411),
	.w6(32'h3aa3819f),
	.w7(32'h3c1b7c10),
	.w8(32'hbb8fff05),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bd49c),
	.w1(32'h3b21964d),
	.w2(32'hb9ef72be),
	.w3(32'h39e4c6ab),
	.w4(32'hbab5d9c9),
	.w5(32'hba9da255),
	.w6(32'hba89d6ed),
	.w7(32'hbab1c255),
	.w8(32'hbb51d93a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a7027),
	.w1(32'h3b8449ba),
	.w2(32'h3aac89b2),
	.w3(32'hba82f628),
	.w4(32'hbaa4f992),
	.w5(32'hb9ec96c6),
	.w6(32'h3b86a3da),
	.w7(32'h3a930220),
	.w8(32'hbb6ee2ba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8185bb),
	.w1(32'h3bea8abd),
	.w2(32'hba950ccd),
	.w3(32'hb8f5726f),
	.w4(32'h3b51b7b8),
	.w5(32'hba5f769b),
	.w6(32'h3c6591cf),
	.w7(32'h3b3e6ea2),
	.w8(32'h3ae53ec8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97394c),
	.w1(32'h3babaee5),
	.w2(32'h3b9d009a),
	.w3(32'h3a49589b),
	.w4(32'h3b7bd9bb),
	.w5(32'hbabd981e),
	.w6(32'h3b8e4f43),
	.w7(32'h3b75b63f),
	.w8(32'hbacfe50f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb808),
	.w1(32'hbb16094c),
	.w2(32'h3ab28558),
	.w3(32'hba44e39e),
	.w4(32'h3b04f713),
	.w5(32'hbb9e20da),
	.w6(32'h39fe5f9e),
	.w7(32'hbaebc0ef),
	.w8(32'hbc1a9d66),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf76fd7),
	.w1(32'hbb419355),
	.w2(32'h3bb0dc22),
	.w3(32'hbac0af9f),
	.w4(32'h3b8fb616),
	.w5(32'h3c0e4200),
	.w6(32'h3b095d43),
	.w7(32'h3b9fae2c),
	.w8(32'h3b7276d3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfa861),
	.w1(32'h3bf87829),
	.w2(32'hba5b9651),
	.w3(32'h3bad3614),
	.w4(32'h3b7ec327),
	.w5(32'hb9a81995),
	.w6(32'h3b9150c9),
	.w7(32'h3b49a520),
	.w8(32'hba7da0fd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5be50e),
	.w1(32'hba87c0fb),
	.w2(32'hbb053ba6),
	.w3(32'hbbd7e85f),
	.w4(32'hbabf47f0),
	.w5(32'hbaa2b054),
	.w6(32'h38db0adb),
	.w7(32'hbb48b461),
	.w8(32'hbb9be085),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375539),
	.w1(32'hbb1e825b),
	.w2(32'hbb4f2f48),
	.w3(32'hbb725cd2),
	.w4(32'hba9e72bf),
	.w5(32'hbb8bee77),
	.w6(32'h3b7f91a4),
	.w7(32'hbb0f4122),
	.w8(32'h3abb38e4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd09e13),
	.w1(32'h3bb25544),
	.w2(32'h3b0405ca),
	.w3(32'hba5fd2f2),
	.w4(32'hba108246),
	.w5(32'hbbb416ce),
	.w6(32'h38d3baee),
	.w7(32'h3a12893f),
	.w8(32'h3c33cca6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dcd4e),
	.w1(32'h3b2091c4),
	.w2(32'h3a7ccb1a),
	.w3(32'hbb2e9ed1),
	.w4(32'hb9a5d6eb),
	.w5(32'hbb615421),
	.w6(32'h3bbf1440),
	.w7(32'h3b079e83),
	.w8(32'hbb3aebeb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb263a05),
	.w1(32'hbbb46278),
	.w2(32'hbb1edec6),
	.w3(32'hbbd4423a),
	.w4(32'hbb13038b),
	.w5(32'hba2ebc72),
	.w6(32'hbad52124),
	.w7(32'hbb28eaca),
	.w8(32'hbafc297b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceb017),
	.w1(32'hbaded9cf),
	.w2(32'h3a58a55a),
	.w3(32'hbc0a9aed),
	.w4(32'hbac2e450),
	.w5(32'h3b7c1464),
	.w6(32'hbb796c86),
	.w7(32'hba59507c),
	.w8(32'hbb2a8e6e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa48e48),
	.w1(32'h3b9b3119),
	.w2(32'h3971fd48),
	.w3(32'h385ce94b),
	.w4(32'h3ad91346),
	.w5(32'h3800e64f),
	.w6(32'h3a93333a),
	.w7(32'h3b379a21),
	.w8(32'hbb636c18),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fe69d),
	.w1(32'h3b46a834),
	.w2(32'hbb4b4e86),
	.w3(32'hb9782247),
	.w4(32'h3b76e1c1),
	.w5(32'hbb951114),
	.w6(32'h3b0348be),
	.w7(32'h3a43c3b1),
	.w8(32'hbc41ee2c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7e979),
	.w1(32'h3c689fe9),
	.w2(32'h3b7c510d),
	.w3(32'hbc1e274d),
	.w4(32'h3c112753),
	.w5(32'h39fff98b),
	.w6(32'h3bfe04be),
	.w7(32'h3c414eaf),
	.w8(32'hbb5f38b0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7517f4),
	.w1(32'h3b3104ab),
	.w2(32'h3b05d708),
	.w3(32'hbbb85315),
	.w4(32'hbae9e735),
	.w5(32'h3b1ffe69),
	.w6(32'h3b9ed74d),
	.w7(32'h3b09aebe),
	.w8(32'h3b33fe8c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef0a19),
	.w1(32'h3b02e1bd),
	.w2(32'h3a3c3b3f),
	.w3(32'h3bce4619),
	.w4(32'h3a88124e),
	.w5(32'hba0df182),
	.w6(32'h3b0fe447),
	.w7(32'h3b0510d7),
	.w8(32'hba989135),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918008a),
	.w1(32'h3b11fa6b),
	.w2(32'h3bbdea5a),
	.w3(32'hbb784173),
	.w4(32'h3a424697),
	.w5(32'hbb5293f7),
	.w6(32'h3a4b214e),
	.w7(32'h3b116d4c),
	.w8(32'hbb1138c9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c6f76),
	.w1(32'hbabbfa48),
	.w2(32'hbb3219d6),
	.w3(32'hbb85fde5),
	.w4(32'hbb8bc425),
	.w5(32'hbbb9c0d0),
	.w6(32'hbae46800),
	.w7(32'hba6590c3),
	.w8(32'hbb9ad34d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48fa0e),
	.w1(32'hbb991f55),
	.w2(32'hba62480f),
	.w3(32'hbb993919),
	.w4(32'h39b40c9b),
	.w5(32'h3a630215),
	.w6(32'hbb66541f),
	.w7(32'h3a174cb4),
	.w8(32'h398e480c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba164925),
	.w1(32'hbba69807),
	.w2(32'h3b05d9c2),
	.w3(32'hbb99bd87),
	.w4(32'hbba11b72),
	.w5(32'h3ad9536b),
	.w6(32'hbb42aa56),
	.w7(32'hbb29aaeb),
	.w8(32'h3c4b6b5a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172f44),
	.w1(32'h3c2c6f4b),
	.w2(32'h3a76c95b),
	.w3(32'h3bca0fba),
	.w4(32'h3a501653),
	.w5(32'hbb3e0710),
	.w6(32'h3c496520),
	.w7(32'h3c1f1cdd),
	.w8(32'hbb201ea2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248e99),
	.w1(32'hbbb7fdc7),
	.w2(32'hb663427e),
	.w3(32'hbb28f454),
	.w4(32'hbb6d85db),
	.w5(32'hbb2ab8cc),
	.w6(32'hbba1e560),
	.w7(32'h396c8294),
	.w8(32'h3c615ecc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b9834),
	.w1(32'hbbaa56fa),
	.w2(32'hb99adcee),
	.w3(32'h3c5b86f5),
	.w4(32'hba5aa812),
	.w5(32'hbb93efca),
	.w6(32'h38cecda8),
	.w7(32'h3ab95267),
	.w8(32'h3bb1482c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9d32),
	.w1(32'h3c0552fd),
	.w2(32'h3b3628c1),
	.w3(32'h3b28ec3f),
	.w4(32'h3b0c3ddd),
	.w5(32'hbacbc964),
	.w6(32'h3b7469ca),
	.w7(32'h3b87200c),
	.w8(32'h3a9fa9e6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649ed4),
	.w1(32'hbad63190),
	.w2(32'hb9a1a6c1),
	.w3(32'hbb7c80ee),
	.w4(32'hba73c933),
	.w5(32'hb9a25a54),
	.w6(32'hbb5fd0d7),
	.w7(32'hbb332e06),
	.w8(32'hbb714c1f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42522d),
	.w1(32'h3c1a47f3),
	.w2(32'hba644103),
	.w3(32'hbb4994bf),
	.w4(32'hbafc4f4b),
	.w5(32'h3bad2ca8),
	.w6(32'h3a321960),
	.w7(32'h3bfe0285),
	.w8(32'h3bc7eef5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10129),
	.w1(32'hba8dc876),
	.w2(32'h3a0ebf69),
	.w3(32'h3aa32c62),
	.w4(32'h3b2f0d35),
	.w5(32'hbb2d555a),
	.w6(32'hbb152889),
	.w7(32'hbb445ab1),
	.w8(32'hbb278fd7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb4c4b),
	.w1(32'hb9e60aad),
	.w2(32'hba21daad),
	.w3(32'hbbc271f4),
	.w4(32'hbba72d9a),
	.w5(32'hbbd2d07c),
	.w6(32'h3bc79265),
	.w7(32'hbb50adf6),
	.w8(32'hbbc777ad),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776007),
	.w1(32'hba7dd53b),
	.w2(32'h3a248839),
	.w3(32'hbbeb1edf),
	.w4(32'hbb9194e7),
	.w5(32'h3bfb22d9),
	.w6(32'hbb874823),
	.w7(32'hba9ef2c7),
	.w8(32'hbb818c6c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3368c),
	.w1(32'hbaf70a91),
	.w2(32'h3ac5b058),
	.w3(32'hbb8ec90b),
	.w4(32'hbb029035),
	.w5(32'hbb8a7d7b),
	.w6(32'h3a999cab),
	.w7(32'h3b37f85a),
	.w8(32'hbb8a1a70),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4540d0),
	.w1(32'hbb2de23f),
	.w2(32'h3b910c74),
	.w3(32'h3b4b6683),
	.w4(32'h3b147f8d),
	.w5(32'h3b6dfc0a),
	.w6(32'h3b4fe50f),
	.w7(32'hbb132719),
	.w8(32'hbaf62333),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8949),
	.w1(32'hba8168ef),
	.w2(32'h3900f7fa),
	.w3(32'hbb0976b9),
	.w4(32'hbb1cc69c),
	.w5(32'hbb861ad3),
	.w6(32'h3a93a17e),
	.w7(32'h39eebebf),
	.w8(32'h3bc50244),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fafb),
	.w1(32'h3b889125),
	.w2(32'h3bdbf6f5),
	.w3(32'hba8209d2),
	.w4(32'hba1f6182),
	.w5(32'hbbb622d2),
	.w6(32'h3acbf7b5),
	.w7(32'h3b8e9b34),
	.w8(32'hbbb580c6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a651),
	.w1(32'h3c45c227),
	.w2(32'h3b5d8feb),
	.w3(32'hbb27f120),
	.w4(32'hbb7a153f),
	.w5(32'h3abd48fd),
	.w6(32'h3c90ddf8),
	.w7(32'h3b061f09),
	.w8(32'h3b297639),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374b80),
	.w1(32'h3b24c867),
	.w2(32'h3be2ba4c),
	.w3(32'h3b8421d1),
	.w4(32'h3a2fa681),
	.w5(32'hba313bca),
	.w6(32'h3b0eeee1),
	.w7(32'h3bec53ac),
	.w8(32'hbac98f28),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f3973),
	.w1(32'h3b1182d8),
	.w2(32'h3b506065),
	.w3(32'hbb4464b3),
	.w4(32'h3a637b93),
	.w5(32'h3986347b),
	.w6(32'h374785d4),
	.w7(32'h3b7ffd0c),
	.w8(32'hbac028a1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48b3d4),
	.w1(32'h3b75171f),
	.w2(32'h3b3c2952),
	.w3(32'hbb2dc1ac),
	.w4(32'hbad69e18),
	.w5(32'h3a9e26d6),
	.w6(32'hbad718e4),
	.w7(32'hbaaab992),
	.w8(32'hbb98c0de),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bae7f4),
	.w1(32'hba2edfbc),
	.w2(32'hbb9e87de),
	.w3(32'hb9a0f795),
	.w4(32'hbb1ea87c),
	.w5(32'hbb8adf94),
	.w6(32'hb928026f),
	.w7(32'hbac97777),
	.w8(32'h39212ecd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacfc6c),
	.w1(32'h3b82a48e),
	.w2(32'h3b248da2),
	.w3(32'h39b68720),
	.w4(32'h3b5b4f5e),
	.w5(32'h3bad631a),
	.w6(32'h3baa1009),
	.w7(32'h3bebc409),
	.w8(32'hba4e282a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984cd4d),
	.w1(32'h3b5b1e7f),
	.w2(32'hbabeee21),
	.w3(32'hbad85e51),
	.w4(32'h3ae908d3),
	.w5(32'h3b3882de),
	.w6(32'h3b325ae8),
	.w7(32'h3b2f0525),
	.w8(32'hba210c18),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936edad),
	.w1(32'h3a39bdf2),
	.w2(32'hbb175b74),
	.w3(32'h3acd34b0),
	.w4(32'h3b53e49d),
	.w5(32'hbb8c8742),
	.w6(32'h3bf3ec62),
	.w7(32'h3a83a7a6),
	.w8(32'h3adb239b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75e6c3),
	.w1(32'h3b505bf6),
	.w2(32'h3b101db7),
	.w3(32'hbae6c524),
	.w4(32'hbb981aa2),
	.w5(32'h3b4ddeb4),
	.w6(32'h3a2eb04e),
	.w7(32'h3b0abd36),
	.w8(32'h3b289f5a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf026ba),
	.w1(32'h3bfad288),
	.w2(32'h3b2b4364),
	.w3(32'h3b54c4bc),
	.w4(32'h3bc524fe),
	.w5(32'hbac7c1b6),
	.w6(32'h3c339abc),
	.w7(32'h3bd9268d),
	.w8(32'hba8a1b43),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890346),
	.w1(32'hbb57326b),
	.w2(32'h3b01e36b),
	.w3(32'hba40e8f4),
	.w4(32'hbb27abe3),
	.w5(32'hbbab0b16),
	.w6(32'hbbb0ed46),
	.w7(32'hbabb830f),
	.w8(32'hbacf3341),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e550),
	.w1(32'hbbc587a2),
	.w2(32'hbb62d04f),
	.w3(32'hbbfe8f85),
	.w4(32'hbc0b080c),
	.w5(32'hbb86b015),
	.w6(32'hbbca0303),
	.w7(32'hbbb0681b),
	.w8(32'hbb592add),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ce14e),
	.w1(32'hbb1d994e),
	.w2(32'h38f827c6),
	.w3(32'hbb98399c),
	.w4(32'hbb2ec96e),
	.w5(32'hbaa85259),
	.w6(32'h3a80050b),
	.w7(32'h3ae62714),
	.w8(32'hbb956504),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e66d8),
	.w1(32'hbb028a37),
	.w2(32'h399a5ced),
	.w3(32'h3ad747cd),
	.w4(32'h3b06df18),
	.w5(32'h3b7826a9),
	.w6(32'hbb31a9c5),
	.w7(32'hbb0242cc),
	.w8(32'hbb8de341),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954578),
	.w1(32'hbb5e9ac5),
	.w2(32'h3b015aa6),
	.w3(32'hbbbe18fc),
	.w4(32'hbb8d4b2f),
	.w5(32'h3b0e0338),
	.w6(32'hbb836f26),
	.w7(32'hbb9a210c),
	.w8(32'hbba638c5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09a2b7),
	.w1(32'h3aaf2eb4),
	.w2(32'hbaee4e70),
	.w3(32'hbb150087),
	.w4(32'h3aaaae46),
	.w5(32'h3ba923a2),
	.w6(32'hba2a7e38),
	.w7(32'h3b4c18ba),
	.w8(32'hbb59779f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19858c),
	.w1(32'hbb6a0263),
	.w2(32'hbc57f93b),
	.w3(32'hbb7a65e0),
	.w4(32'h3a4ad876),
	.w5(32'hbbb2aaa7),
	.w6(32'h3ae5f940),
	.w7(32'hbb911f67),
	.w8(32'hbb5baf53),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa29208),
	.w1(32'hba24b253),
	.w2(32'hb9921a4e),
	.w3(32'hbba4c605),
	.w4(32'hbbbfb04c),
	.w5(32'hbab74960),
	.w6(32'hbbf66c12),
	.w7(32'h3ade56de),
	.w8(32'h3b6aba4d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadecf3d),
	.w1(32'hba9ceccd),
	.w2(32'h385a226b),
	.w3(32'h3ba54b4a),
	.w4(32'h3a5f77b8),
	.w5(32'hbbbe1809),
	.w6(32'h3b574c23),
	.w7(32'h3a93c795),
	.w8(32'h3b053dd3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae320),
	.w1(32'h3a5428f1),
	.w2(32'hba2c1348),
	.w3(32'hbbc04879),
	.w4(32'hbb824842),
	.w5(32'hbbc2e3de),
	.w6(32'h3a2d3383),
	.w7(32'hbb077d52),
	.w8(32'hbba51826),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5da1),
	.w1(32'hbbcb3a5a),
	.w2(32'hbb1a1bbb),
	.w3(32'hbb2e53bf),
	.w4(32'hba64c916),
	.w5(32'hbb4fac9c),
	.w6(32'hbb82034a),
	.w7(32'hbb109de6),
	.w8(32'hbabda9c2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97811a),
	.w1(32'hbb618893),
	.w2(32'h3a55edf0),
	.w3(32'hbba95a99),
	.w4(32'hbb7880a3),
	.w5(32'hbad14244),
	.w6(32'hbb2b0a78),
	.w7(32'hb9d91c38),
	.w8(32'h3c0545b5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c0c18),
	.w1(32'h3a109275),
	.w2(32'h3b384529),
	.w3(32'hbb192f7a),
	.w4(32'hbbae82f9),
	.w5(32'h3a880d7f),
	.w6(32'h3bf39d35),
	.w7(32'hbb1abe4b),
	.w8(32'h3b8d05de),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91739),
	.w1(32'h3bbeccc3),
	.w2(32'hb899957b),
	.w3(32'h3b8b9fb5),
	.w4(32'h3ad1ac06),
	.w5(32'h3b11ba3f),
	.w6(32'h3c81a413),
	.w7(32'h3b0230cf),
	.w8(32'h3b4788e4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7bb87),
	.w1(32'hbad47ef0),
	.w2(32'hbb0ba754),
	.w3(32'h3bd48706),
	.w4(32'h377cc6ce),
	.w5(32'hbb0ccff4),
	.w6(32'h3a875b5a),
	.w7(32'hba32fd5f),
	.w8(32'hbb8339e8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd19da2),
	.w1(32'hbba73468),
	.w2(32'h38eafa06),
	.w3(32'hbb5d9df7),
	.w4(32'hbb966c34),
	.w5(32'hbb58d98a),
	.w6(32'hbb338f4f),
	.w7(32'hba5a4a57),
	.w8(32'hba62d75f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48fee2),
	.w1(32'h3c9ada85),
	.w2(32'h3bf678ce),
	.w3(32'hbb2fdf4e),
	.w4(32'h3a39a65e),
	.w5(32'h3ae277fe),
	.w6(32'hb99a8d41),
	.w7(32'h3aa8b2ee),
	.w8(32'h3b989d01),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78af82),
	.w1(32'hbb141829),
	.w2(32'h3aeff099),
	.w3(32'h3b8c4949),
	.w4(32'h3b3a2e48),
	.w5(32'h3baffc74),
	.w6(32'hbb1355c0),
	.w7(32'h3b3073ea),
	.w8(32'hba9168dc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab5a2),
	.w1(32'h3b6d4ed9),
	.w2(32'h3bd72ef3),
	.w3(32'hbbfcc965),
	.w4(32'hba3d9bb8),
	.w5(32'h3b1ec2c0),
	.w6(32'hbc58b532),
	.w7(32'h3c6b0f9b),
	.w8(32'hbc08659c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51a907),
	.w1(32'h3bd31867),
	.w2(32'h3bcaca6d),
	.w3(32'h3ae25751),
	.w4(32'hbbb65ba1),
	.w5(32'hbbdc0a91),
	.w6(32'hbc0225ea),
	.w7(32'h38bb2a60),
	.w8(32'h3984dc31),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d733),
	.w1(32'hbbae0b33),
	.w2(32'h3b22f3dd),
	.w3(32'hbbbc340e),
	.w4(32'hbb89f4d0),
	.w5(32'hbb1f399c),
	.w6(32'hbbca8225),
	.w7(32'hbacbe5a9),
	.w8(32'h3b2bbea9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bd46c),
	.w1(32'hbb3e8faa),
	.w2(32'hbb815128),
	.w3(32'h39fdfb4a),
	.w4(32'h388eb591),
	.w5(32'hbbc46966),
	.w6(32'h3c421820),
	.w7(32'hbbb384a0),
	.w8(32'h3ac9827d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7e9f),
	.w1(32'hba94eed0),
	.w2(32'hbad73bc9),
	.w3(32'hbb82c928),
	.w4(32'hbb03bffb),
	.w5(32'hbb288e9b),
	.w6(32'h3b1fa69e),
	.w7(32'hb94d9154),
	.w8(32'h3b16fed4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b213a),
	.w1(32'h3bc68faf),
	.w2(32'h399bdb81),
	.w3(32'hb9a0789e),
	.w4(32'h3bc35f85),
	.w5(32'hbbdfa98e),
	.w6(32'h3c2e744a),
	.w7(32'h3a827a6d),
	.w8(32'hbaea5fbf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d59fb),
	.w1(32'h3b675a8b),
	.w2(32'h3a63bcd7),
	.w3(32'hba6d65e6),
	.w4(32'hba9e36e8),
	.w5(32'h3b879b9b),
	.w6(32'h3bce9fc0),
	.w7(32'h3a7096e3),
	.w8(32'h3bfa8f4a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a17b),
	.w1(32'h3c0be28e),
	.w2(32'h3bad4951),
	.w3(32'h3bd3b5f5),
	.w4(32'h3bc077f9),
	.w5(32'hb9edebec),
	.w6(32'h3ba9f6ef),
	.w7(32'h3bf9e8d7),
	.w8(32'hba874ecb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f6833),
	.w1(32'h3b92d611),
	.w2(32'hba7d905b),
	.w3(32'h3aa2afbc),
	.w4(32'hba966e93),
	.w5(32'h3b37f1c0),
	.w6(32'h3bf4a354),
	.w7(32'h3b2fdd5c),
	.w8(32'hbbacf072),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc746),
	.w1(32'h3959b0d7),
	.w2(32'h3b5150ee),
	.w3(32'hbba1fc03),
	.w4(32'h3b57af3a),
	.w5(32'hbbac653f),
	.w6(32'hbb3cd312),
	.w7(32'h3bf4d26b),
	.w8(32'h3c15180f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ad36),
	.w1(32'h3bd5d06c),
	.w2(32'h3b225b74),
	.w3(32'hbab87a35),
	.w4(32'h3b287d32),
	.w5(32'h3b82fb5d),
	.w6(32'h3b936921),
	.w7(32'h3be3ba25),
	.w8(32'hbb2e5c2c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3881dd),
	.w1(32'h3b8ebe6b),
	.w2(32'h3a865342),
	.w3(32'h3b063a9e),
	.w4(32'h3a5f4f52),
	.w5(32'hbb26bb03),
	.w6(32'h3c2da2e0),
	.w7(32'h3a54f279),
	.w8(32'hbb235d68),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb501c84),
	.w1(32'hbb351512),
	.w2(32'h3acdbb2c),
	.w3(32'hb98f98d0),
	.w4(32'h3b06ee63),
	.w5(32'h3adf85cd),
	.w6(32'h3c1f02f9),
	.w7(32'h3b14f3da),
	.w8(32'hba9d4a1a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5d53),
	.w1(32'h3a3085e8),
	.w2(32'h3a82e820),
	.w3(32'h3aa7ee3c),
	.w4(32'h3aadcc8f),
	.w5(32'hbb8263b7),
	.w6(32'h3c095427),
	.w7(32'h3b2f623f),
	.w8(32'h3ab6923e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda175a),
	.w1(32'h3bcd5513),
	.w2(32'h3b5e9e6f),
	.w3(32'h3b55532d),
	.w4(32'h3baeec37),
	.w5(32'h3bb1c17b),
	.w6(32'h3c6063b4),
	.w7(32'h3c18838d),
	.w8(32'h3a8d2d91),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81141e),
	.w1(32'h3b9d36c4),
	.w2(32'h3a853df8),
	.w3(32'hbb3930d0),
	.w4(32'hba512be6),
	.w5(32'hbb9d0a89),
	.w6(32'hbc20b6d0),
	.w7(32'hb941e261),
	.w8(32'h3b4f591d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b333),
	.w1(32'hbb3b52bb),
	.w2(32'hbaa411d3),
	.w3(32'hbb8185a2),
	.w4(32'hb82b0275),
	.w5(32'h3a6dc66c),
	.w6(32'h3b5f208b),
	.w7(32'hbb220347),
	.w8(32'hbb9146f8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a358190),
	.w1(32'h3b47a83b),
	.w2(32'hbb336cd4),
	.w3(32'hbaba7507),
	.w4(32'h3937fbf2),
	.w5(32'h3ac0c499),
	.w6(32'h3bbe29c4),
	.w7(32'h3aaac198),
	.w8(32'h3b57e524),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dcc45),
	.w1(32'hbb93cb9f),
	.w2(32'hbb55de77),
	.w3(32'h3c2bbf4f),
	.w4(32'hbb01eaeb),
	.w5(32'hbc15213c),
	.w6(32'hb9b9afab),
	.w7(32'hbb85c130),
	.w8(32'hbc1794ae),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60acf),
	.w1(32'h3b398f0f),
	.w2(32'hbb423dc3),
	.w3(32'hba451de2),
	.w4(32'h39cf7341),
	.w5(32'h3b0441ae),
	.w6(32'h39bfda01),
	.w7(32'h3b523f75),
	.w8(32'h3c62f9ab),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c212853),
	.w1(32'h3ae2c27a),
	.w2(32'h3a669b14),
	.w3(32'h3c8d88aa),
	.w4(32'h3c0729cc),
	.w5(32'hbb82c566),
	.w6(32'h3bd0935d),
	.w7(32'h3b2b5b0a),
	.w8(32'hbb7ec63f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de084),
	.w1(32'hbb524adf),
	.w2(32'h3a99c982),
	.w3(32'h3a76597e),
	.w4(32'h38e33fec),
	.w5(32'h3a6186b3),
	.w6(32'h389a311c),
	.w7(32'hba7fa034),
	.w8(32'h3adc9dd3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27ba4e),
	.w1(32'hb8c122bf),
	.w2(32'hbab6640b),
	.w3(32'h3b5bb788),
	.w4(32'hbbd6fc4f),
	.w5(32'hbba1dbf0),
	.w6(32'h3bea14a1),
	.w7(32'h3ac3ee67),
	.w8(32'hbb0f56fc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbdae9),
	.w1(32'hbb6292a7),
	.w2(32'hb9b0f86c),
	.w3(32'hbb8e7f49),
	.w4(32'hbbafd7cd),
	.w5(32'hbb96ed99),
	.w6(32'hbb91ef44),
	.w7(32'hbb1fee95),
	.w8(32'hb9dc9ce0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913554),
	.w1(32'h39a63c95),
	.w2(32'h3af57637),
	.w3(32'hbab66066),
	.w4(32'hbba53e0e),
	.w5(32'h3b28017f),
	.w6(32'hb9655ded),
	.w7(32'hbb66119e),
	.w8(32'hbb819629),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63ccfa),
	.w1(32'hbaf914f3),
	.w2(32'h3871330a),
	.w3(32'hbb9286e6),
	.w4(32'h3b3455b1),
	.w5(32'hbba1457b),
	.w6(32'h3bc5b4f0),
	.w7(32'h3b891beb),
	.w8(32'h3ae251fe),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf108a),
	.w1(32'hba8183ef),
	.w2(32'h3a65461d),
	.w3(32'h3c4556c1),
	.w4(32'h3bc6a572),
	.w5(32'h3990a884),
	.w6(32'h3c6b9d8b),
	.w7(32'h3ac743ce),
	.w8(32'h39a32a9b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37976456),
	.w1(32'hba733340),
	.w2(32'h39aad88a),
	.w3(32'hb8d15286),
	.w4(32'h39b7ebfe),
	.w5(32'hba205c9d),
	.w6(32'hba521ee4),
	.w7(32'hb8b9b7b2),
	.w8(32'hb9f4b643),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c74112),
	.w1(32'h39d0c390),
	.w2(32'hb90d9f1d),
	.w3(32'h395a74a6),
	.w4(32'h3aafa037),
	.w5(32'h38a64844),
	.w6(32'h38a0d524),
	.w7(32'h3a5dc037),
	.w8(32'h39423675),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0286b3),
	.w1(32'hb9ee5276),
	.w2(32'hba5e5143),
	.w3(32'h398f0f9b),
	.w4(32'hba046a55),
	.w5(32'hb9944869),
	.w6(32'h3b17e337),
	.w7(32'h3a421469),
	.w8(32'h393aa142),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b165107),
	.w1(32'h3b46810d),
	.w2(32'h3ad84a14),
	.w3(32'h38699373),
	.w4(32'hb9789d2e),
	.w5(32'h39cd57d7),
	.w6(32'h3b2f8ca6),
	.w7(32'h3a99d299),
	.w8(32'h3a094153),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a90ea),
	.w1(32'h3a061b43),
	.w2(32'h3ad18e77),
	.w3(32'h3a05e97a),
	.w4(32'h3aba59c2),
	.w5(32'h3b5928ad),
	.w6(32'h3aef6052),
	.w7(32'h3b1796c5),
	.w8(32'h3b2684ef),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afecf97),
	.w1(32'h3a471a26),
	.w2(32'hb9e6d0f9),
	.w3(32'h3a9a05bc),
	.w4(32'h3a916e2a),
	.w5(32'hb8a60fcb),
	.w6(32'h3a429380),
	.w7(32'h3943aafa),
	.w8(32'h3aaefdde),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895baf7),
	.w1(32'hbac44e36),
	.w2(32'hbb05e706),
	.w3(32'hb8610f68),
	.w4(32'hbaca3e64),
	.w5(32'hba0c7eda),
	.w6(32'h39174860),
	.w7(32'h3951f5a3),
	.w8(32'h3a255999),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39739517),
	.w1(32'h3a2dbf2e),
	.w2(32'h3ac47a78),
	.w3(32'h3a93a689),
	.w4(32'h39e3aef5),
	.w5(32'h399200e4),
	.w6(32'h37c8db71),
	.w7(32'hba394fdc),
	.w8(32'h387e10c4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b3d6c),
	.w1(32'h3a5f546e),
	.w2(32'h3a2c31b2),
	.w3(32'h38366e87),
	.w4(32'h3a140a15),
	.w5(32'hb9a76226),
	.w6(32'h388edf32),
	.w7(32'hb9298e8c),
	.w8(32'h3924e48b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8e94),
	.w1(32'hba1f6c7e),
	.w2(32'h3999594a),
	.w3(32'h3745d974),
	.w4(32'h3a533150),
	.w5(32'h39c68e34),
	.w6(32'h3a3810e3),
	.w7(32'h3a37421f),
	.w8(32'h38a962ce),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9546c27),
	.w1(32'hbad20784),
	.w2(32'h39d3a52d),
	.w3(32'hba5708a0),
	.w4(32'h3a2414a0),
	.w5(32'h390cd8fd),
	.w6(32'hbb233d79),
	.w7(32'hba15f0f4),
	.w8(32'hb8a79253),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc8012),
	.w1(32'hb95cde62),
	.w2(32'h3993cb25),
	.w3(32'hba59b624),
	.w4(32'hb93ba9e0),
	.w5(32'h3ab504d0),
	.w6(32'hba3095f3),
	.w7(32'h39d5cecb),
	.w8(32'h3aa18616),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5821eb),
	.w1(32'h3a5aee09),
	.w2(32'h3a99e244),
	.w3(32'h3a080bed),
	.w4(32'h3a9fea1d),
	.w5(32'h3aa4c0fc),
	.w6(32'hba9f3c7d),
	.w7(32'h3a6d3dfa),
	.w8(32'h39ffc21a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d639a4),
	.w1(32'h3b200f60),
	.w2(32'h3a3b3af6),
	.w3(32'h3a6b93b6),
	.w4(32'h3afe038a),
	.w5(32'h394da2a5),
	.w6(32'h3ae715fe),
	.w7(32'h3b217a40),
	.w8(32'h3a67a096),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b3e2c),
	.w1(32'hb8ca2b31),
	.w2(32'h3a6cb024),
	.w3(32'hba33f50a),
	.w4(32'h3a74a7d1),
	.w5(32'h3a5eca9a),
	.w6(32'hba357763),
	.w7(32'h3a71d068),
	.w8(32'h39de8c38),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22df54),
	.w1(32'h3afe2cc0),
	.w2(32'h3979b89c),
	.w3(32'h3aa489db),
	.w4(32'h3a189137),
	.w5(32'hb996ed9f),
	.w6(32'h3a2f8a8f),
	.w7(32'h39978a4c),
	.w8(32'hb9de9275),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf440),
	.w1(32'hbb250cd5),
	.w2(32'hbb2eb938),
	.w3(32'h39717d9e),
	.w4(32'hbaa7a219),
	.w5(32'h3a2fff28),
	.w6(32'hb92b6134),
	.w7(32'hbacd0465),
	.w8(32'h3a28e1af),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db54b1),
	.w1(32'hb9d4da90),
	.w2(32'h39bb460d),
	.w3(32'h3a48361a),
	.w4(32'h3a11b9ba),
	.w5(32'hba0fcd93),
	.w6(32'h3a8f93e3),
	.w7(32'h3a7cfdfe),
	.w8(32'hb97f0933),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811011),
	.w1(32'hb9629877),
	.w2(32'hba77701e),
	.w3(32'hba4593e3),
	.w4(32'hba6f71c2),
	.w5(32'hbafd2f6f),
	.w6(32'hba847b65),
	.w7(32'hba83f1fc),
	.w8(32'hba547431),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0988f8),
	.w1(32'hbadbdc43),
	.w2(32'hbb165951),
	.w3(32'hbadd2bf0),
	.w4(32'hbab1f6b2),
	.w5(32'h3a82eec3),
	.w6(32'hb9f0e964),
	.w7(32'hba97f84a),
	.w8(32'h3ab6bad8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bab0e),
	.w1(32'h3a906839),
	.w2(32'h3a0cf1e1),
	.w3(32'h3abf2aa2),
	.w4(32'h3aafc1d2),
	.w5(32'h3af2891f),
	.w6(32'h3aa7aa09),
	.w7(32'h3a008935),
	.w8(32'h3abee807),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c68fe4),
	.w1(32'hba0e3ec5),
	.w2(32'h39f2b118),
	.w3(32'hbaab0b0c),
	.w4(32'hba3a076b),
	.w5(32'h3b1a0036),
	.w6(32'hbac96292),
	.w7(32'h39c19480),
	.w8(32'h39e61175),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bd0be),
	.w1(32'hb92d4dbb),
	.w2(32'hb9b5b273),
	.w3(32'h3a4475f3),
	.w4(32'h3980f1cf),
	.w5(32'h3a9ecdc2),
	.w6(32'h3a419f18),
	.w7(32'h3a46cf9b),
	.w8(32'h3b188461),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9319cd),
	.w1(32'hbaf6d870),
	.w2(32'hbae39ec3),
	.w3(32'hba4cec50),
	.w4(32'hba035e49),
	.w5(32'h3b4dd54d),
	.w6(32'hb94f2518),
	.w7(32'hba562bd8),
	.w8(32'hbb238d1e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cc94e),
	.w1(32'h3b0fa127),
	.w2(32'h3afd4f39),
	.w3(32'h3b0f65ab),
	.w4(32'hbab6b454),
	.w5(32'hbb10b4fa),
	.w6(32'hbb178ff2),
	.w7(32'hbb725f6b),
	.w8(32'h3a5763da),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394880c2),
	.w1(32'hbb646a2d),
	.w2(32'hba61f8d1),
	.w3(32'hbb4bc191),
	.w4(32'hb9298b3f),
	.w5(32'h3b328f9d),
	.w6(32'hba87d16e),
	.w7(32'h3a9faf85),
	.w8(32'hbaf527a8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac377f1),
	.w1(32'h39280ae0),
	.w2(32'hb88eb6f4),
	.w3(32'h3b485ecc),
	.w4(32'h3a4eacaf),
	.w5(32'hb9ccc7a0),
	.w6(32'hbb119468),
	.w7(32'hbb514b54),
	.w8(32'hba903076),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40eecd),
	.w1(32'h39882d8d),
	.w2(32'h39bba463),
	.w3(32'hb9d4532f),
	.w4(32'h39e7cee4),
	.w5(32'hbac76da7),
	.w6(32'hb9177015),
	.w7(32'hba5268b7),
	.w8(32'hba433188),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ee3a1),
	.w1(32'hba846d66),
	.w2(32'hb9441fc4),
	.w3(32'hba8ce087),
	.w4(32'hba3abfa9),
	.w5(32'h3a45eefc),
	.w6(32'h38f1c713),
	.w7(32'hb98746b0),
	.w8(32'h3a04cb97),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c5ce3f),
	.w1(32'h39ccacec),
	.w2(32'hb9af3f40),
	.w3(32'h395619e5),
	.w4(32'hba36e5dd),
	.w5(32'h3ac2cf1f),
	.w6(32'hb9257965),
	.w7(32'hba68b5bf),
	.w8(32'hb937333d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule