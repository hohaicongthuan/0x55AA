module layer_8_featuremap_172(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82f439),
	.w1(32'h3c08e278),
	.w2(32'hbc8b1dc6),
	.w3(32'h3c5b02af),
	.w4(32'h3aaf2d3f),
	.w5(32'hbc33c29e),
	.w6(32'h3c0d9e06),
	.w7(32'h3bbe3d36),
	.w8(32'hbb2e42c0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8304e8),
	.w1(32'h3830aa31),
	.w2(32'h3bff93eb),
	.w3(32'h3b33d996),
	.w4(32'h3b33d721),
	.w5(32'h3bf60131),
	.w6(32'hbafd4f9f),
	.w7(32'h3b78f0dc),
	.w8(32'h3b31f3b9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43d083),
	.w1(32'h3c4bef9c),
	.w2(32'h3c367eb8),
	.w3(32'hbb2a6c7a),
	.w4(32'h3c2b5b02),
	.w5(32'h3c34ed1a),
	.w6(32'h3bb663db),
	.w7(32'h3c17f41a),
	.w8(32'h3c2787d3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3461),
	.w1(32'hbc1a611e),
	.w2(32'hbc70231b),
	.w3(32'h3c82c5cb),
	.w4(32'h3af9193e),
	.w5(32'hbc38f3c9),
	.w6(32'hbc072e94),
	.w7(32'hbb34e85f),
	.w8(32'h3bde0efd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156146),
	.w1(32'h3bf72bbe),
	.w2(32'h3be89caf),
	.w3(32'hbbb06dc3),
	.w4(32'h3c110f0a),
	.w5(32'h3be4e66c),
	.w6(32'h3b8cc83f),
	.w7(32'h3c09c896),
	.w8(32'h3b159ace),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b8f58),
	.w1(32'h3c2c795e),
	.w2(32'h3c0b4249),
	.w3(32'hbc04e6b2),
	.w4(32'h3b4867eb),
	.w5(32'hbc5f1c32),
	.w6(32'h3c0e9ac8),
	.w7(32'h3c719bba),
	.w8(32'hbbf8a55d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce13b44),
	.w1(32'h3b5b22e9),
	.w2(32'hbaad2f2a),
	.w3(32'hbc898eb5),
	.w4(32'h3aa0aa04),
	.w5(32'hb974935c),
	.w6(32'h3b5f2a8e),
	.w7(32'h3b5b2bf8),
	.w8(32'h3b9d38d0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7b34),
	.w1(32'hbb8a4ba1),
	.w2(32'hbb8b30be),
	.w3(32'h3c444a90),
	.w4(32'h3b1ae7ae),
	.w5(32'hb9eeecc4),
	.w6(32'h3b52b08b),
	.w7(32'h3c3e8ef7),
	.w8(32'h3c88d718),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cada1a6),
	.w1(32'h3c37b354),
	.w2(32'hbb258ef7),
	.w3(32'h3c340bf5),
	.w4(32'h3beea0d8),
	.w5(32'hbb910de8),
	.w6(32'hbb2711b8),
	.w7(32'hbb575f2b),
	.w8(32'hbbdebbea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41d649),
	.w1(32'hbc00d49d),
	.w2(32'hbc9cf0c7),
	.w3(32'hba659455),
	.w4(32'hbb40cd13),
	.w5(32'hbbeb8fe9),
	.w6(32'h3b39c487),
	.w7(32'hbb99b8c3),
	.w8(32'h3baefee2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ab951),
	.w1(32'hbc95bfc5),
	.w2(32'h3d0efd82),
	.w3(32'h3c2373eb),
	.w4(32'hbcae0c3c),
	.w5(32'h3bdc0900),
	.w6(32'hbaf32ecd),
	.w7(32'h3c4c446b),
	.w8(32'h3c11a013),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf5c02e),
	.w1(32'h3b2a594c),
	.w2(32'hbbb64c31),
	.w3(32'h3cd3aea0),
	.w4(32'h3b89816d),
	.w5(32'hbbb7172a),
	.w6(32'h3b961972),
	.w7(32'h3b9a5f49),
	.w8(32'h3b5ee85d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07c09d),
	.w1(32'hb81f41cd),
	.w2(32'h3aec722e),
	.w3(32'hbb8981a3),
	.w4(32'h3c3592c0),
	.w5(32'h3cb678ae),
	.w6(32'hba9167f5),
	.w7(32'hbb50d3f5),
	.w8(32'h3c3a5b88),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae59a),
	.w1(32'h3c0f7ee9),
	.w2(32'h3b560e8b),
	.w3(32'h3bf04945),
	.w4(32'h3b866567),
	.w5(32'hba24d903),
	.w6(32'h3c1f24fc),
	.w7(32'h3c2965d3),
	.w8(32'h3afe5a32),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bb475),
	.w1(32'hbbaf3a8a),
	.w2(32'hbc0f83ce),
	.w3(32'h3b05651b),
	.w4(32'hbb69bf43),
	.w5(32'hbb710a01),
	.w6(32'hbbb4811f),
	.w7(32'hbba6217d),
	.w8(32'hba6990f3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65bb4c),
	.w1(32'hbafc11da),
	.w2(32'hbc4215a4),
	.w3(32'hba158b2a),
	.w4(32'hb8cad223),
	.w5(32'hbc40c41b),
	.w6(32'hbc134dc1),
	.w7(32'hba742a41),
	.w8(32'hbbf42bbc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082df1),
	.w1(32'hbcaa3700),
	.w2(32'hbc381984),
	.w3(32'hbb881395),
	.w4(32'hbc298c71),
	.w5(32'h3b0ef8c1),
	.w6(32'hbc39bac7),
	.w7(32'hbc55aec6),
	.w8(32'hbbb38ef7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55fa59),
	.w1(32'h3b91b351),
	.w2(32'hbc25ec2e),
	.w3(32'hbbd72265),
	.w4(32'h3c00bc05),
	.w5(32'hbb389762),
	.w6(32'hbc000728),
	.w7(32'h3a0f513c),
	.w8(32'h3c409357),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb2dff),
	.w1(32'hbc579f23),
	.w2(32'hbd89883d),
	.w3(32'h3c0f8ba2),
	.w4(32'hbc4f5549),
	.w5(32'hbd486c78),
	.w6(32'h3b87d8f9),
	.w7(32'h3a884aab),
	.w8(32'h3b5433cf),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a792),
	.w1(32'hbbc930d5),
	.w2(32'hbcecdbaa),
	.w3(32'h3bb6ada7),
	.w4(32'hbb1deb05),
	.w5(32'hbc8e3e4e),
	.w6(32'h3c039127),
	.w7(32'hbbe8f837),
	.w8(32'hbbdeece8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67dc8d),
	.w1(32'hbc1eccbe),
	.w2(32'hbaff7b61),
	.w3(32'hbbf2936b),
	.w4(32'h3b05155e),
	.w5(32'h3b2d8cfd),
	.w6(32'h3a16cdeb),
	.w7(32'hbb99a177),
	.w8(32'hbb0af929),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd0b95),
	.w1(32'h3c085cbc),
	.w2(32'h3bb48577),
	.w3(32'h3ac7f010),
	.w4(32'h3c155616),
	.w5(32'h3c8aa7c8),
	.w6(32'h3c535fd5),
	.w7(32'h3c236a34),
	.w8(32'h3c292281),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9dd2f0),
	.w1(32'h3b49a8b1),
	.w2(32'h3822ddbd),
	.w3(32'h3d9397d9),
	.w4(32'h3c7367ba),
	.w5(32'h3ce53030),
	.w6(32'h3cf8a38d),
	.w7(32'h3c27605b),
	.w8(32'h3d1720a0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8b058a),
	.w1(32'hbb407b8e),
	.w2(32'hbc0990d1),
	.w3(32'h3d17901a),
	.w4(32'hbb0ac455),
	.w5(32'hbbd44856),
	.w6(32'h3b8151b4),
	.w7(32'h39a098a8),
	.w8(32'hbc5ef4f2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3093d),
	.w1(32'h3c212516),
	.w2(32'h3ba6d8d7),
	.w3(32'h3c08639e),
	.w4(32'h3ba8f013),
	.w5(32'h3c1a2dbb),
	.w6(32'h3bb00505),
	.w7(32'hbb13cc92),
	.w8(32'h3c10b291),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfe3eb),
	.w1(32'h3ba6d5ef),
	.w2(32'hbc54203e),
	.w3(32'h3ca2bddf),
	.w4(32'h3bd147c5),
	.w5(32'h3b9d36dc),
	.w6(32'hbb32d481),
	.w7(32'hbc3423e7),
	.w8(32'hbb200765),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfbc97),
	.w1(32'hbbddb731),
	.w2(32'hbb2953b0),
	.w3(32'hbb264348),
	.w4(32'hbbc3a32e),
	.w5(32'hbb45d05d),
	.w6(32'h3bbeb468),
	.w7(32'h3b90cca4),
	.w8(32'hbb4f2c50),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bf78b),
	.w1(32'hbc9928d0),
	.w2(32'hbdceab1f),
	.w3(32'h3ca25294),
	.w4(32'hbba1c2bc),
	.w5(32'hbdc15a89),
	.w6(32'hbd8c0dd6),
	.w7(32'hbd5a5873),
	.w8(32'hbc4bc573),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33cadc),
	.w1(32'h3c78cd21),
	.w2(32'hbb25f6e0),
	.w3(32'hbc51d0e8),
	.w4(32'h3c05254e),
	.w5(32'hbc05b92f),
	.w6(32'h3c1b5a8d),
	.w7(32'h3b8cf945),
	.w8(32'hbbefb4c6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99690d),
	.w1(32'h3b4ea7f0),
	.w2(32'h3ac7eb76),
	.w3(32'hbc206f76),
	.w4(32'h3b8f6c44),
	.w5(32'h3b9869e9),
	.w6(32'h3b0b4c30),
	.w7(32'h3a644ceb),
	.w8(32'h3be14af0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5480),
	.w1(32'h3bb3d931),
	.w2(32'h3b1f28a2),
	.w3(32'h3b2e0de3),
	.w4(32'hba99b445),
	.w5(32'hbbc3eb0f),
	.w6(32'h3c225c9c),
	.w7(32'h3be689fe),
	.w8(32'hbb46b445),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886386),
	.w1(32'hbc8bf5cc),
	.w2(32'hbc36d209),
	.w3(32'h3b06d9dd),
	.w4(32'hbc180047),
	.w5(32'h3b36d38b),
	.w6(32'hbc181ccc),
	.w7(32'hbbe3c50f),
	.w8(32'h39fd9232),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c526c0d),
	.w1(32'hb7d96a32),
	.w2(32'h3d08a761),
	.w3(32'h3c7ada29),
	.w4(32'h3a848852),
	.w5(32'h3c39bc64),
	.w6(32'h3c57f99c),
	.w7(32'h3cbc3b1d),
	.w8(32'h3c6f86e0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07feca),
	.w1(32'h3bd89d72),
	.w2(32'h38563171),
	.w3(32'h3cc4f2ef),
	.w4(32'h3c09e0e5),
	.w5(32'h3b9a32ce),
	.w6(32'h3bc34589),
	.w7(32'h3c2d94f3),
	.w8(32'h3bf0841d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9b31),
	.w1(32'h39390580),
	.w2(32'hbbff7f5e),
	.w3(32'h3b5838aa),
	.w4(32'h3baf2179),
	.w5(32'hb93aad73),
	.w6(32'h3bd92598),
	.w7(32'hbb281bd7),
	.w8(32'hbb852355),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8f0b2),
	.w1(32'h3ad2fd23),
	.w2(32'hbc01e9c8),
	.w3(32'hbbc39c98),
	.w4(32'hbc19b3cb),
	.w5(32'hbc03d2e7),
	.w6(32'h3a49be91),
	.w7(32'hbb660b8a),
	.w8(32'hbc0c33d6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f589),
	.w1(32'h3b530866),
	.w2(32'hbba686a3),
	.w3(32'h3bd6d3d0),
	.w4(32'hba689667),
	.w5(32'hbbde802b),
	.w6(32'hbb58f1ca),
	.w7(32'hbb8fae69),
	.w8(32'hbb877e43),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876886),
	.w1(32'h3bd3e249),
	.w2(32'h3c151093),
	.w3(32'hbbf87477),
	.w4(32'h3c19a5ad),
	.w5(32'h3c2c3d28),
	.w6(32'h390ccf52),
	.w7(32'h3bc8f59e),
	.w8(32'h3bfec93f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea0f1e),
	.w1(32'h3b758915),
	.w2(32'h3bdfcc90),
	.w3(32'hb9cdef6b),
	.w4(32'hbadc68d5),
	.w5(32'h3ba8d329),
	.w6(32'h3a694997),
	.w7(32'h3b697a89),
	.w8(32'hbb42a4b9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fc590),
	.w1(32'h3b90a90c),
	.w2(32'h3bc1db3b),
	.w3(32'h3c504466),
	.w4(32'h3b11862d),
	.w5(32'h3bc5b3d2),
	.w6(32'h3b5fb3fa),
	.w7(32'h3b620a44),
	.w8(32'h3bf5c538),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84d12c),
	.w1(32'hbb57cf94),
	.w2(32'hbcef2a96),
	.w3(32'h3b92e248),
	.w4(32'hbc28a752),
	.w5(32'hbcd40960),
	.w6(32'hbc3860b5),
	.w7(32'hbc8252cd),
	.w8(32'hbc00ac56),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd07ea8),
	.w1(32'hbc485dd2),
	.w2(32'hba23c099),
	.w3(32'hbbed8c9f),
	.w4(32'hbc15af9f),
	.w5(32'hbba48240),
	.w6(32'h3b7c71b1),
	.w7(32'h3bad5c8f),
	.w8(32'h3ab69492),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e545),
	.w1(32'h3bbae6e5),
	.w2(32'h3c267066),
	.w3(32'h3b15934a),
	.w4(32'h3c0eb3a6),
	.w5(32'h3c2ffcb4),
	.w6(32'h3b0c1cec),
	.w7(32'h3b1ba30b),
	.w8(32'h3b6653e0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2eda7),
	.w1(32'h3c0e26ab),
	.w2(32'h3a63e4e8),
	.w3(32'hbb2b54bb),
	.w4(32'hbae0cb9b),
	.w5(32'hbb27f4ba),
	.w6(32'h3baf7590),
	.w7(32'h3c160ddb),
	.w8(32'h39f55085),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d083a50),
	.w1(32'h3c0db573),
	.w2(32'hbbaa31a1),
	.w3(32'h3ce46989),
	.w4(32'h3c03f7fb),
	.w5(32'hbc84d2c4),
	.w6(32'h3bf0aef6),
	.w7(32'h3be9b3b8),
	.w8(32'hbb0d88c7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58b944),
	.w1(32'hbbefef1b),
	.w2(32'hbc1007b0),
	.w3(32'hbc0a0f03),
	.w4(32'hbbba9c1c),
	.w5(32'hbbfd5fd6),
	.w6(32'hbb798235),
	.w7(32'h3ab6ee7c),
	.w8(32'hba019ed5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6ab23),
	.w1(32'hbae163e5),
	.w2(32'hbbc34f48),
	.w3(32'hb8d9bf64),
	.w4(32'h3b6b37a8),
	.w5(32'h39ef956c),
	.w6(32'h3ad6b3e1),
	.w7(32'hba44e76b),
	.w8(32'h3c2e50fa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9dab5),
	.w1(32'h3bbaf23f),
	.w2(32'hbcbb46e5),
	.w3(32'h3d0024ed),
	.w4(32'hb9d2a3db),
	.w5(32'hbc028a68),
	.w6(32'h3c8a52b1),
	.w7(32'h3c3c518b),
	.w8(32'h3b8ffa99),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25ffae),
	.w1(32'h3afeec15),
	.w2(32'h3bd4683f),
	.w3(32'h3b832094),
	.w4(32'h3b045847),
	.w5(32'h3c46fb33),
	.w6(32'h3c25ff2a),
	.w7(32'h3c0a181f),
	.w8(32'h3c31e69e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f585b),
	.w1(32'h3bf86972),
	.w2(32'hbcacd74b),
	.w3(32'h3c713c35),
	.w4(32'h3b691a57),
	.w5(32'hbbca78b8),
	.w6(32'hba1385d7),
	.w7(32'hbc2ef1a8),
	.w8(32'hbc79ee13),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf7c60),
	.w1(32'h3c357f3a),
	.w2(32'h3c504004),
	.w3(32'hbcef8c84),
	.w4(32'h3c4844e8),
	.w5(32'h3c96415c),
	.w6(32'h3baab6a2),
	.w7(32'h3bd99b89),
	.w8(32'h3cbf39ea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd98093),
	.w1(32'hbc7c14d5),
	.w2(32'hbcc88595),
	.w3(32'h3c926f78),
	.w4(32'hbcd39204),
	.w5(32'hbd0f06e3),
	.w6(32'h3c7f52ce),
	.w7(32'h3bb24747),
	.w8(32'hbc0d673b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3466),
	.w1(32'hbb859897),
	.w2(32'hbb85f23e),
	.w3(32'h3c309493),
	.w4(32'hbb5448ea),
	.w5(32'hbb8ed2e2),
	.w6(32'h3b987d6c),
	.w7(32'h3b2d3a46),
	.w8(32'h3bb2daae),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2fcd1),
	.w1(32'hbc0dc894),
	.w2(32'h3ad8885c),
	.w3(32'h3c536498),
	.w4(32'hbb8a27ff),
	.w5(32'h3c6e0379),
	.w6(32'h3a99d0d0),
	.w7(32'hbb007af2),
	.w8(32'h3c3281a7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9db703),
	.w1(32'h3b975025),
	.w2(32'h3ca6a30b),
	.w3(32'h3c1612bd),
	.w4(32'h3b4ee97f),
	.w5(32'h3c840fef),
	.w6(32'h3c0d7f9c),
	.w7(32'h3c82804c),
	.w8(32'h3ca10d60),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d52f396),
	.w1(32'h3c818abf),
	.w2(32'hbcc29e23),
	.w3(32'h3d33a526),
	.w4(32'h3cac6bed),
	.w5(32'hbc13bad0),
	.w6(32'h3c66aba0),
	.w7(32'hba301eda),
	.w8(32'h3c2eb651),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951c97),
	.w1(32'hbb5d627a),
	.w2(32'hbd06aed0),
	.w3(32'h3c1111f0),
	.w4(32'hbab02dbc),
	.w5(32'hbc66e13e),
	.w6(32'h3c5065d2),
	.w7(32'hbc92a71e),
	.w8(32'hbc3abea7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d5f81),
	.w1(32'h3aeced27),
	.w2(32'hbc730880),
	.w3(32'hbc099faf),
	.w4(32'hbbd00d73),
	.w5(32'hbcc1cc9c),
	.w6(32'hbac38a61),
	.w7(32'hbbe02447),
	.w8(32'hbc9f9742),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd01cfa),
	.w1(32'hbb655de0),
	.w2(32'hbc1a0324),
	.w3(32'hbcb183f8),
	.w4(32'hbb70be15),
	.w5(32'hbc285291),
	.w6(32'h39c8706d),
	.w7(32'hbb7a0339),
	.w8(32'hbbecdda3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63dd66),
	.w1(32'h3b8b18a5),
	.w2(32'h3bbfe76c),
	.w3(32'hbb294c23),
	.w4(32'hbb63b141),
	.w5(32'h3badf623),
	.w6(32'hbb2029d4),
	.w7(32'h3b7392a8),
	.w8(32'hbb7a16cc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7669b2),
	.w1(32'h3b0a0c1f),
	.w2(32'hbc27024e),
	.w3(32'h3c621c7c),
	.w4(32'hbc51dcd5),
	.w5(32'hbcb8a5fe),
	.w6(32'h3c4b396f),
	.w7(32'h3c088b1e),
	.w8(32'hbc026033),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26415d),
	.w1(32'h3bdef9b6),
	.w2(32'hb7704c98),
	.w3(32'hba8d03d0),
	.w4(32'hbc27a9c4),
	.w5(32'hbbb761a5),
	.w6(32'hbb3189b1),
	.w7(32'hbb945645),
	.w8(32'h3b2f7978),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95cc5d),
	.w1(32'h3c7537fb),
	.w2(32'h3be30f84),
	.w3(32'h3b77b339),
	.w4(32'h3c2c79c4),
	.w5(32'h3a166eb6),
	.w6(32'h3c8078c7),
	.w7(32'h3c854020),
	.w8(32'h3c3baf21),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bc487),
	.w1(32'hbc2b4d3b),
	.w2(32'hbc8b1dad),
	.w3(32'hbc29ffc6),
	.w4(32'hbbea7220),
	.w5(32'hbc83fde3),
	.w6(32'hbb494bfb),
	.w7(32'hbc2ff3dc),
	.w8(32'hbbdea6f0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa9b7c),
	.w1(32'hbc1ab010),
	.w2(32'hbb0dbc70),
	.w3(32'hbb92bc88),
	.w4(32'hbbcd6709),
	.w5(32'hbb68b5e9),
	.w6(32'hbb83442c),
	.w7(32'hbb17f66c),
	.w8(32'h3a92705d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c082e62),
	.w1(32'h3b8f60c3),
	.w2(32'h392152ca),
	.w3(32'h3ba1d37b),
	.w4(32'hbaf17e12),
	.w5(32'h3ad2492a),
	.w6(32'hb9c7f65b),
	.w7(32'h3c0ac93c),
	.w8(32'h3bc2a0db),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89a24b),
	.w1(32'h3cb221d8),
	.w2(32'h3c65f0cf),
	.w3(32'h3c19d3ae),
	.w4(32'h3c52418a),
	.w5(32'h3c238fdb),
	.w6(32'h3c67532f),
	.w7(32'h3c4f3ad6),
	.w8(32'h3b28f13b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1660a),
	.w1(32'h39a754c5),
	.w2(32'hbc36aa34),
	.w3(32'hbbb98d37),
	.w4(32'h3a7ebd71),
	.w5(32'hba291b1d),
	.w6(32'hbc22ed9b),
	.w7(32'h3bb3438d),
	.w8(32'h3c30b658),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c089d66),
	.w1(32'hbc05901a),
	.w2(32'hbc31db2c),
	.w3(32'h3b90237c),
	.w4(32'h3ad077ff),
	.w5(32'hbba0eecf),
	.w6(32'hbaed7f4d),
	.w7(32'h3bb2b06a),
	.w8(32'h3c2f3563),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ddafd),
	.w1(32'h3cc3c5a4),
	.w2(32'hbd1976f8),
	.w3(32'h3cfbf05b),
	.w4(32'hba8d3e96),
	.w5(32'hbd11e924),
	.w6(32'hbb0325a9),
	.w7(32'hbb4cc6fb),
	.w8(32'hbc0891c8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42b9ae),
	.w1(32'h3a89207a),
	.w2(32'hbc44b0ec),
	.w3(32'hba20f16f),
	.w4(32'h3bf667d8),
	.w5(32'hbbf563b8),
	.w6(32'h3bb8e1f6),
	.w7(32'hba9def57),
	.w8(32'hbc0f6ee8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85bd75),
	.w1(32'h3c2e151b),
	.w2(32'h3af4abdb),
	.w3(32'h3b3f60a1),
	.w4(32'h3c33d4d0),
	.w5(32'hba2013a2),
	.w6(32'h3c0c904b),
	.w7(32'hbad3eba3),
	.w8(32'h3ac94516),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd81a8b),
	.w1(32'h3c4ea9d1),
	.w2(32'h3c07c866),
	.w3(32'h3b8895e6),
	.w4(32'h3b2d3fca),
	.w5(32'h3b47bc6d),
	.w6(32'h3c876c4b),
	.w7(32'h3b94f191),
	.w8(32'h3b13b334),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e0695),
	.w1(32'h3c754e59),
	.w2(32'hbc5286d6),
	.w3(32'h3c7be57a),
	.w4(32'h3b9bc457),
	.w5(32'hbc8280cc),
	.w6(32'h3c5b254d),
	.w7(32'h3bb1dcb5),
	.w8(32'hbc14957f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb19612),
	.w1(32'h3b5a3b3f),
	.w2(32'h38d21e39),
	.w3(32'hbcaae4cd),
	.w4(32'hbb6406ef),
	.w5(32'hbb1b1383),
	.w6(32'h3a2de90a),
	.w7(32'hbb5f5e91),
	.w8(32'hbb87ef40),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc9781),
	.w1(32'hbbdf7440),
	.w2(32'hbd2d256d),
	.w3(32'h3c4796c1),
	.w4(32'hbbabcc88),
	.w5(32'hbd0f5d93),
	.w6(32'hb9f575c0),
	.w7(32'hbcea449e),
	.w8(32'hbc73b25f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6578d0),
	.w1(32'h3c65cf88),
	.w2(32'hbbfd613f),
	.w3(32'hbb21e200),
	.w4(32'h3bb3d3c6),
	.w5(32'hbc4e4956),
	.w6(32'h3c38da1f),
	.w7(32'hbaea7cc5),
	.w8(32'hbc41ede5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb653c85),
	.w1(32'h3c86688c),
	.w2(32'hbc8a1288),
	.w3(32'hbb88515a),
	.w4(32'h3c033db3),
	.w5(32'hbc999bd0),
	.w6(32'h399f2572),
	.w7(32'hbbccb025),
	.w8(32'hbaf35223),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c716),
	.w1(32'hbc0e87b2),
	.w2(32'hbceaf27b),
	.w3(32'h3adc6099),
	.w4(32'hbbcd1586),
	.w5(32'hbca97ad1),
	.w6(32'hbba104a6),
	.w7(32'hbb91f3c6),
	.w8(32'hba970d05),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb189ec),
	.w1(32'hbc21e428),
	.w2(32'h3b53979c),
	.w3(32'hbb9d5444),
	.w4(32'hbab342c7),
	.w5(32'hbc250ae7),
	.w6(32'h3b463c46),
	.w7(32'hbb56add5),
	.w8(32'h3c41cbfe),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8db3a0),
	.w1(32'hb9ac2a89),
	.w2(32'hbc00c8ec),
	.w3(32'h3c68139c),
	.w4(32'h3b4dcac4),
	.w5(32'h3b29c27b),
	.w6(32'h3b54bd0c),
	.w7(32'hbbc89829),
	.w8(32'hbb3400a1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08c488),
	.w1(32'h3b90a2f4),
	.w2(32'h3c21882f),
	.w3(32'hbbb7f0b2),
	.w4(32'h3a632ac9),
	.w5(32'h3c290aa6),
	.w6(32'h3b9f4b8c),
	.w7(32'h3bcf98e0),
	.w8(32'hba0ae769),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1ddc6),
	.w1(32'hbb5c4e88),
	.w2(32'hbd2099a9),
	.w3(32'h3cb692e2),
	.w4(32'hbc2331cf),
	.w5(32'hbd19d82c),
	.w6(32'h3b6c11be),
	.w7(32'hbc352fb3),
	.w8(32'hbc09a5a9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc358d95),
	.w1(32'hbc36f3d2),
	.w2(32'h3c392b4d),
	.w3(32'hbcaa6c40),
	.w4(32'hbcb6ed7d),
	.w5(32'h3cb8fe68),
	.w6(32'hbc9b1f37),
	.w7(32'h3c4d6157),
	.w8(32'h3c8c710b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da19083),
	.w1(32'hba794a59),
	.w2(32'hbd110963),
	.w3(32'h3d6d4a0b),
	.w4(32'hbba0d92b),
	.w5(32'hbd234e27),
	.w6(32'h3c8bf43c),
	.w7(32'h3b81af91),
	.w8(32'h3bc4c343),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fa7d6),
	.w1(32'hbba57108),
	.w2(32'hbc4d5de2),
	.w3(32'h3c49d4c0),
	.w4(32'hb8470bfe),
	.w5(32'hbcaa2032),
	.w6(32'h3c2394d2),
	.w7(32'h3c6b2396),
	.w8(32'hbbfc578a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca16ee8),
	.w1(32'hbc13b301),
	.w2(32'hbb30a277),
	.w3(32'hbc40cedd),
	.w4(32'hbb69a7c2),
	.w5(32'h3b3bbffa),
	.w6(32'hbbdf1c52),
	.w7(32'hbbbdfd7c),
	.w8(32'hbc0dcac6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371063),
	.w1(32'h3ad22ad2),
	.w2(32'h3b89f2e3),
	.w3(32'h3b897362),
	.w4(32'hbb74b86f),
	.w5(32'hb838d30a),
	.w6(32'h3b84a2d1),
	.w7(32'h3a212438),
	.w8(32'h3bffe658),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b59fa),
	.w1(32'hbb3eabc2),
	.w2(32'hbbc2b1ab),
	.w3(32'hbc3a3fad),
	.w4(32'hbba42dfe),
	.w5(32'hbaa994a7),
	.w6(32'h3aabbe96),
	.w7(32'h3ab6354b),
	.w8(32'hbc08c01d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22899f),
	.w1(32'h3c93398a),
	.w2(32'h3a146a70),
	.w3(32'h3b9aff06),
	.w4(32'h3c2a0c58),
	.w5(32'h3c16ea83),
	.w6(32'h3c98f5e4),
	.w7(32'h3bea93c6),
	.w8(32'h3c30773d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e9764),
	.w1(32'h3b05925b),
	.w2(32'hbb2dde6e),
	.w3(32'h3c8b0092),
	.w4(32'h3bfb61a6),
	.w5(32'h3bc768f8),
	.w6(32'h3bf0ddea),
	.w7(32'h3af67659),
	.w8(32'h3bf4dbf0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe61264),
	.w1(32'h3b544ef0),
	.w2(32'h3beffe64),
	.w3(32'h3af7bff5),
	.w4(32'h3bdc2677),
	.w5(32'h3b9dc5cb),
	.w6(32'h3a983588),
	.w7(32'hb9f323a8),
	.w8(32'h3c30fda7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb914b),
	.w1(32'hbbc34919),
	.w2(32'h3b4e6781),
	.w3(32'h3c06ce8d),
	.w4(32'hbb784ec9),
	.w5(32'hba5dfe1b),
	.w6(32'hbbc9e2a4),
	.w7(32'hbbe0146a),
	.w8(32'hbb9c43a6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd9ac7),
	.w1(32'h3b27ad22),
	.w2(32'h3bab2cac),
	.w3(32'h3a9b1c2e),
	.w4(32'h3b87ed88),
	.w5(32'h3ba4a13a),
	.w6(32'h3bb53868),
	.w7(32'h3ba4a817),
	.w8(32'h3aef31e1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067dee),
	.w1(32'h3b814c3c),
	.w2(32'hbb1a7a87),
	.w3(32'hbbb834b1),
	.w4(32'h3b617ca6),
	.w5(32'hbabaa7d6),
	.w6(32'h3b6d2a0a),
	.w7(32'h3c1708f2),
	.w8(32'hba9dcd71),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a3bb),
	.w1(32'h3c149714),
	.w2(32'hbc631179),
	.w3(32'hbac0c13f),
	.w4(32'h396de911),
	.w5(32'hbc5c20fe),
	.w6(32'h3c2bfba6),
	.w7(32'h3b0f6941),
	.w8(32'hbc2ffea3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab420),
	.w1(32'h3b5d812b),
	.w2(32'h3c8dfd2d),
	.w3(32'h3a436965),
	.w4(32'h3bd63a32),
	.w5(32'h3cb668f3),
	.w6(32'h3c5649a5),
	.w7(32'h3c7fe7ed),
	.w8(32'h3c000328),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d115efc),
	.w1(32'h3a613caa),
	.w2(32'h3c642827),
	.w3(32'h3cc6c5d9),
	.w4(32'h3c234d19),
	.w5(32'h3c637a60),
	.w6(32'h3bb4af25),
	.w7(32'h3be92bc4),
	.w8(32'h3c22baa7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3808b),
	.w1(32'hbaf23adc),
	.w2(32'hbb593abf),
	.w3(32'h3c6dcaae),
	.w4(32'hbb84c7be),
	.w5(32'h3b7ea79f),
	.w6(32'h3b918479),
	.w7(32'h3a03d784),
	.w8(32'hbafa5463),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade0fac),
	.w1(32'hbc4a983c),
	.w2(32'hbc13a825),
	.w3(32'hbb10af0c),
	.w4(32'hbc2c277f),
	.w5(32'hbbfd1856),
	.w6(32'h3acc9bdd),
	.w7(32'h39dbc447),
	.w8(32'h3c2a9979),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c821982),
	.w1(32'hbc862b61),
	.w2(32'hbba1701d),
	.w3(32'h3c90b894),
	.w4(32'hbbc9842e),
	.w5(32'hbb280380),
	.w6(32'hbbbabf01),
	.w7(32'h3ba2f7bd),
	.w8(32'h3b92a3b9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb761a2),
	.w1(32'h3bbcde2e),
	.w2(32'h3cc3d8b9),
	.w3(32'h3ca76d13),
	.w4(32'h3c42ad64),
	.w5(32'h3c478102),
	.w6(32'hb91891b6),
	.w7(32'h3c100159),
	.w8(32'h3bc74d41),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44160b),
	.w1(32'h3be278bd),
	.w2(32'h3a3f3c3e),
	.w3(32'hbbb044ea),
	.w4(32'h3be7088d),
	.w5(32'h3b70e481),
	.w6(32'hbb685af6),
	.w7(32'hbb7fb25d),
	.w8(32'h3a92e08a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38eee4),
	.w1(32'hbcb73fc4),
	.w2(32'hbd0c6036),
	.w3(32'h3b9ced00),
	.w4(32'hbcaaf440),
	.w5(32'hbc3d4064),
	.w6(32'h3ba85860),
	.w7(32'hbca245d8),
	.w8(32'hbca83891),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca40c2d),
	.w1(32'h3be06221),
	.w2(32'h3d32b286),
	.w3(32'hbababc48),
	.w4(32'h3c197248),
	.w5(32'h3d388af1),
	.w6(32'h3c016ae8),
	.w7(32'h3c894ec0),
	.w8(32'h3d19e7a8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d866942),
	.w1(32'hbc38a820),
	.w2(32'hbce49ca7),
	.w3(32'h3d7b0984),
	.w4(32'hbc6cfd52),
	.w5(32'hbccf1169),
	.w6(32'hbbb8b2d8),
	.w7(32'hbc22f79f),
	.w8(32'hbbbece2c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0d796),
	.w1(32'h3b5010cb),
	.w2(32'hbc9b4172),
	.w3(32'h3b9f6e81),
	.w4(32'hbc00408b),
	.w5(32'hbcb8059f),
	.w6(32'h3b870adb),
	.w7(32'hbabf18ac),
	.w8(32'hbc86b80e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb0a0),
	.w1(32'h3b842357),
	.w2(32'hbc16ed56),
	.w3(32'h3b36c97c),
	.w4(32'h3b92635e),
	.w5(32'h3b0b147c),
	.w6(32'hbbde8254),
	.w7(32'hbc52ba2b),
	.w8(32'hbb607271),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc904549),
	.w1(32'h3c13f1ba),
	.w2(32'h3c186344),
	.w3(32'hbc6f8884),
	.w4(32'h3bc45a72),
	.w5(32'h3bd5ad46),
	.w6(32'h3c77af9d),
	.w7(32'h3c28cb71),
	.w8(32'h3b61135a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba261ccd),
	.w1(32'h3b6cee0e),
	.w2(32'h3c40f162),
	.w3(32'h3b37485a),
	.w4(32'h3c019666),
	.w5(32'h3c5214ad),
	.w6(32'h3b16ebec),
	.w7(32'h3be24a71),
	.w8(32'h3bf71bdd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf05f75),
	.w1(32'h35ed5080),
	.w2(32'hbbfb5665),
	.w3(32'h3a688940),
	.w4(32'hbbaa2e2a),
	.w5(32'hb9d47aa1),
	.w6(32'hb9cfdd60),
	.w7(32'h3b60e9e2),
	.w8(32'h3b77dcfe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2e41),
	.w1(32'hbc2a5274),
	.w2(32'hbc14201a),
	.w3(32'h3baa5ec6),
	.w4(32'hbbe25103),
	.w5(32'hbbc624d1),
	.w6(32'hbba3bde6),
	.w7(32'hbb81e5b5),
	.w8(32'hb9759804),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc3c7d),
	.w1(32'h3bb7705e),
	.w2(32'h3c89a0cc),
	.w3(32'hbba7a492),
	.w4(32'h3b061ea9),
	.w5(32'h3c358383),
	.w6(32'h3acc43dd),
	.w7(32'h3bf69c1c),
	.w8(32'h3c04310b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29f2a7),
	.w1(32'hba8cfc60),
	.w2(32'hbb6c013b),
	.w3(32'h39b418e4),
	.w4(32'h3bd8c55c),
	.w5(32'h3c977d70),
	.w6(32'hba9e6ee6),
	.w7(32'hbc17fdb4),
	.w8(32'h3c6cb424),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86ab77),
	.w1(32'hbb92484a),
	.w2(32'h3af2d514),
	.w3(32'h3c56a15c),
	.w4(32'hbc0d6839),
	.w5(32'hbbd1fdd6),
	.w6(32'h3b54aafe),
	.w7(32'h3c072665),
	.w8(32'h3b81cd5a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50e72f),
	.w1(32'hbb36050f),
	.w2(32'h3bc539ff),
	.w3(32'h3bfae3ff),
	.w4(32'hba4caae6),
	.w5(32'h3bd03017),
	.w6(32'hbbac7621),
	.w7(32'hb99a6560),
	.w8(32'h3baac1b3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c105ed4),
	.w1(32'h391f3c79),
	.w2(32'hbb80e5a3),
	.w3(32'h3b9738d0),
	.w4(32'hbc018548),
	.w5(32'hbc370361),
	.w6(32'h3b2664aa),
	.w7(32'hbc23efc2),
	.w8(32'hbc1283e2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7083),
	.w1(32'h3ba65c9c),
	.w2(32'hb8fb1c9c),
	.w3(32'hb9924326),
	.w4(32'h3b94ab9b),
	.w5(32'hbbdbc562),
	.w6(32'h38e80507),
	.w7(32'h3b51babc),
	.w8(32'h3bb9148f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a22f8),
	.w1(32'h3c67e921),
	.w2(32'hbc02d521),
	.w3(32'h3a6fc33e),
	.w4(32'h3ca29379),
	.w5(32'h3bc3531e),
	.w6(32'h3b9f9128),
	.w7(32'hbb66f926),
	.w8(32'hbb4e5d25),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcee73),
	.w1(32'hbc36b9fd),
	.w2(32'hbc395653),
	.w3(32'hbc1b3356),
	.w4(32'hbb9901e6),
	.w5(32'hbb61547a),
	.w6(32'hbbf018a4),
	.w7(32'hbc1d84dc),
	.w8(32'hbb20c6e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08330),
	.w1(32'h3c2ff764),
	.w2(32'h3afa1ed5),
	.w3(32'h3c4a9851),
	.w4(32'h3bf5804f),
	.w5(32'h3c30af9f),
	.w6(32'h3c08e28b),
	.w7(32'h3b5b0446),
	.w8(32'h3bbf536b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed8b05),
	.w1(32'hbc63af1d),
	.w2(32'hbcc9e441),
	.w3(32'h3b4e27a2),
	.w4(32'hbb983d4a),
	.w5(32'hbc043498),
	.w6(32'h3b5e0f3d),
	.w7(32'h3ba7c305),
	.w8(32'h3c14ebeb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d8a4a),
	.w1(32'hbc15115a),
	.w2(32'hbba809bc),
	.w3(32'h3ba6372b),
	.w4(32'hbbd39170),
	.w5(32'hbb6dd5eb),
	.w6(32'hbbe5bf3b),
	.w7(32'hbc003754),
	.w8(32'hbb5ecb92),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc894),
	.w1(32'h3c235529),
	.w2(32'h3c6a9a56),
	.w3(32'hbbc6d84d),
	.w4(32'h3a8a7eee),
	.w5(32'h3b914214),
	.w6(32'h3bb66a87),
	.w7(32'h3bb4ef68),
	.w8(32'h3a2356a5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba514ee7),
	.w1(32'hbb854ae0),
	.w2(32'hbc811f61),
	.w3(32'h3b81626a),
	.w4(32'h3c0b1cc8),
	.w5(32'hbc4839a4),
	.w6(32'hbbb5a47b),
	.w7(32'hbc44aebe),
	.w8(32'hbb559adf),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc561c29),
	.w1(32'h3c2a55fd),
	.w2(32'h3c8929d2),
	.w3(32'hbba5a88c),
	.w4(32'h3b90036b),
	.w5(32'h3c676c23),
	.w6(32'h3c4ba411),
	.w7(32'h3c4c392b),
	.w8(32'h3cad1fa2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8b9cb),
	.w1(32'h39656872),
	.w2(32'h3a33202d),
	.w3(32'h3c8f2503),
	.w4(32'hba226c8b),
	.w5(32'hbaf534c8),
	.w6(32'hba80a4fa),
	.w7(32'hbaa7dbcf),
	.w8(32'hb9f97a6d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88162a),
	.w1(32'h3a9f9996),
	.w2(32'hba1dc63b),
	.w3(32'h3bac2600),
	.w4(32'hbbae2dc5),
	.w5(32'hbc0bfa46),
	.w6(32'h3b95ae8b),
	.w7(32'h3b35a4b2),
	.w8(32'hbb01da7c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule