module layer_8_featuremap_223(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2a2a0),
	.w1(32'hbadb41ff),
	.w2(32'hbb187c90),
	.w3(32'h3a80bc11),
	.w4(32'h3b9eae8f),
	.w5(32'hbb48340a),
	.w6(32'hba8bf211),
	.w7(32'hbb92c790),
	.w8(32'h3a7a91c2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb132b6d),
	.w1(32'hbaf1c1c6),
	.w2(32'hbb8ee5b5),
	.w3(32'h3b2798f0),
	.w4(32'hba0ba606),
	.w5(32'hbb678842),
	.w6(32'hbb229252),
	.w7(32'hbb90b098),
	.w8(32'hbb6cd6b7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39cb5d),
	.w1(32'h3a9b9ee1),
	.w2(32'h3b1266a5),
	.w3(32'hbb43e392),
	.w4(32'h3b1259f2),
	.w5(32'h3aaeddc1),
	.w6(32'h389359ec),
	.w7(32'h3af219d8),
	.w8(32'h3b4f29c1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4469c1),
	.w1(32'h3b08ad7d),
	.w2(32'h3a2522b2),
	.w3(32'h3a45483e),
	.w4(32'h3aa6bbd1),
	.w5(32'h3b804294),
	.w6(32'h3b91ed83),
	.w7(32'h3b0e3630),
	.w8(32'h3b0618b5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0019d1),
	.w1(32'hbbae923e),
	.w2(32'hbc19e6f3),
	.w3(32'h3adb677d),
	.w4(32'hbb211a48),
	.w5(32'hbbe9ae1a),
	.w6(32'hbb94f154),
	.w7(32'hbbf5bc87),
	.w8(32'hbbba8786),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78e10),
	.w1(32'hbba73b9e),
	.w2(32'hbb2f7833),
	.w3(32'hbba60390),
	.w4(32'hba32a11a),
	.w5(32'hbb72c98f),
	.w6(32'hba3830f0),
	.w7(32'hbb5ff5c1),
	.w8(32'h3b19f934),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc787),
	.w1(32'h3b721c77),
	.w2(32'h3bca6f77),
	.w3(32'hbad7dfa7),
	.w4(32'h3b1ea35b),
	.w5(32'h3bc6d3bc),
	.w6(32'h3b465617),
	.w7(32'h3bb34648),
	.w8(32'h3b56ffc6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8605fe),
	.w1(32'hba8cd92a),
	.w2(32'hb9de3e83),
	.w3(32'h3b8415db),
	.w4(32'h3b379d04),
	.w5(32'h3afd44c5),
	.w6(32'hb9ff537f),
	.w7(32'hbb2b81b2),
	.w8(32'hbabefbd0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f9b7e),
	.w1(32'hbb89a411),
	.w2(32'hbb8b0450),
	.w3(32'hbad901af),
	.w4(32'hbb26f771),
	.w5(32'hbb0a9d88),
	.w6(32'hbb568800),
	.w7(32'hbb83d03b),
	.w8(32'hbb2acca5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf68bbb),
	.w1(32'h3b893f05),
	.w2(32'h3a8cd26b),
	.w3(32'hba33d66a),
	.w4(32'h3b26bf5d),
	.w5(32'h3b6333cd),
	.w6(32'h39f2eb45),
	.w7(32'h392b0432),
	.w8(32'hba84b6ba),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf6204),
	.w1(32'h3b9d1a56),
	.w2(32'h39eb7121),
	.w3(32'h3a92887f),
	.w4(32'h3a9fa4f6),
	.w5(32'h3add0a5f),
	.w6(32'hbb36e3fd),
	.w7(32'hbb25c44c),
	.w8(32'hbbb7a447),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c2b2d),
	.w1(32'hb64ded2f),
	.w2(32'hb9aa2743),
	.w3(32'hbb62f119),
	.w4(32'h3a014f7c),
	.w5(32'hba994571),
	.w6(32'hba6ef795),
	.w7(32'hba788d71),
	.w8(32'h3a3e369f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa825a),
	.w1(32'h3b3e086a),
	.w2(32'h3b587957),
	.w3(32'h3ab9a0d1),
	.w4(32'h3aa8a548),
	.w5(32'h3b3a9148),
	.w6(32'h396069c8),
	.w7(32'h3b09d3fd),
	.w8(32'hba73d887),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2baf73),
	.w1(32'h3a8a20ef),
	.w2(32'h3b11f589),
	.w3(32'h3b38d79a),
	.w4(32'h39240ddb),
	.w5(32'h3a229f0f),
	.w6(32'hba330b49),
	.w7(32'hb9b9aed4),
	.w8(32'h361bed73),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f2fc9),
	.w1(32'h3bba3534),
	.w2(32'h3c420de7),
	.w3(32'hba800028),
	.w4(32'h3b51abd3),
	.w5(32'h3c278c1c),
	.w6(32'h3bac4146),
	.w7(32'h3c2158e6),
	.w8(32'h3bfcc7e7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c192ee9),
	.w1(32'hb9ff87cd),
	.w2(32'hbac909d0),
	.w3(32'h3c14dc94),
	.w4(32'h3add7f73),
	.w5(32'hba11f8fb),
	.w6(32'hbb0d621a),
	.w7(32'hbaa81eb2),
	.w8(32'h3a99ffdb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f55d),
	.w1(32'h3a60695a),
	.w2(32'hbb3d2c41),
	.w3(32'h3b9ac78f),
	.w4(32'h3a89a21d),
	.w5(32'hbac1e7d8),
	.w6(32'hbac206e4),
	.w7(32'hbb0ba654),
	.w8(32'hbac08e3e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b947f),
	.w1(32'hb937c527),
	.w2(32'hba9ae211),
	.w3(32'hba5265c1),
	.w4(32'h3b0b37f9),
	.w5(32'h3a4c8a3c),
	.w6(32'hba9efdbc),
	.w7(32'hba68dc5f),
	.w8(32'hbb18ce06),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4c4ac),
	.w1(32'h3adedd33),
	.w2(32'hbb518f49),
	.w3(32'h3939e897),
	.w4(32'h3b3b6b42),
	.w5(32'h3af455bd),
	.w6(32'hbb4b7c15),
	.w7(32'hbb62cb57),
	.w8(32'hbb839c63),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae505ef),
	.w1(32'h3bdecb33),
	.w2(32'h3c4bf85b),
	.w3(32'hbb6f496b),
	.w4(32'h3b72e337),
	.w5(32'h3c2eda84),
	.w6(32'h3bc1b83f),
	.w7(32'h3c250cbc),
	.w8(32'h3bd9618a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078e92),
	.w1(32'hbb4b8c69),
	.w2(32'h3b03bb79),
	.w3(32'h3c023e7d),
	.w4(32'hbab1b729),
	.w5(32'h3a6c2dd2),
	.w6(32'h3786ca6c),
	.w7(32'hb9b9bd23),
	.w8(32'h38caf4a5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5f4fa),
	.w1(32'hbb73ba46),
	.w2(32'hbb847b46),
	.w3(32'hbb155543),
	.w4(32'h3ab3dd73),
	.w5(32'hba9be77b),
	.w6(32'hbaf14bfd),
	.w7(32'hbb05f585),
	.w8(32'h3a381c31),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6e95),
	.w1(32'hbaac7dcd),
	.w2(32'h38c9de24),
	.w3(32'hbb191997),
	.w4(32'hbb22de23),
	.w5(32'h3adb6161),
	.w6(32'hbb23c6fa),
	.w7(32'h3a5fa8a1),
	.w8(32'hbb4826bf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e2ec),
	.w1(32'hbbb22218),
	.w2(32'hbb82b090),
	.w3(32'hba3781f4),
	.w4(32'hbb7adc2b),
	.w5(32'hbbaf1426),
	.w6(32'hbabb3b79),
	.w7(32'hba23cb3a),
	.w8(32'h39274eb6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d18a0),
	.w1(32'hba2c249a),
	.w2(32'hba1f0ff4),
	.w3(32'hbb2481e9),
	.w4(32'hbb28e7a8),
	.w5(32'hbb71c737),
	.w6(32'hbb2bbec7),
	.w7(32'hbab1ce1a),
	.w8(32'hbae38ff1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7122f),
	.w1(32'h397bcd52),
	.w2(32'hbbae300e),
	.w3(32'hbb8d4567),
	.w4(32'hbb985137),
	.w5(32'hbbb9d48c),
	.w6(32'hbbd5e151),
	.w7(32'hbbb3853e),
	.w8(32'hbb81b6b6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43689e),
	.w1(32'h3b027113),
	.w2(32'h3920ff99),
	.w3(32'hbbe2fe96),
	.w4(32'h38b5b962),
	.w5(32'h39597ad6),
	.w6(32'h3ab59478),
	.w7(32'h3acffee8),
	.w8(32'h39947ea1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10adad),
	.w1(32'hb9a0600a),
	.w2(32'h3b88c5a0),
	.w3(32'h3a8ef8f2),
	.w4(32'hbb5c41d9),
	.w5(32'h3ac63a0d),
	.w6(32'h3b1d019e),
	.w7(32'h3adf7f57),
	.w8(32'h3b0d4761),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2796a7),
	.w1(32'hbb7e7760),
	.w2(32'hba19cc29),
	.w3(32'h3aef3b31),
	.w4(32'hba8c959d),
	.w5(32'hba633db1),
	.w6(32'hbbab689a),
	.w7(32'hbb350054),
	.w8(32'h3bf42020),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07ca62),
	.w1(32'hb900e04b),
	.w2(32'h3ac5681a),
	.w3(32'h3bddbed8),
	.w4(32'h3a531965),
	.w5(32'h3aacf4ca),
	.w6(32'hb8bcc658),
	.w7(32'h39a1690e),
	.w8(32'hbb00e776),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08b0a6),
	.w1(32'h3b2c96a5),
	.w2(32'h39f0f77f),
	.w3(32'hbb0d25b5),
	.w4(32'h3b2b764a),
	.w5(32'h3b2986ad),
	.w6(32'hbb1c3244),
	.w7(32'hbb25f36d),
	.w8(32'hbb492ba1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30ac9f),
	.w1(32'hba98e7f6),
	.w2(32'hbad24e5e),
	.w3(32'h3aa3bc09),
	.w4(32'h3b098849),
	.w5(32'hbb2fd1ac),
	.w6(32'hbad3cdba),
	.w7(32'hbaf8b16a),
	.w8(32'h3ad79e3e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c67999),
	.w1(32'h3b87fc8b),
	.w2(32'h3b702cae),
	.w3(32'h3aa3f2c6),
	.w4(32'h3b2be29c),
	.w5(32'h3b556076),
	.w6(32'h3b02df3b),
	.w7(32'h3ac0abae),
	.w8(32'hbaa390ce),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8b29),
	.w1(32'hbaa05f88),
	.w2(32'hbb0bd61c),
	.w3(32'hba0359a1),
	.w4(32'hbb929304),
	.w5(32'hbb8f3dcd),
	.w6(32'hba333740),
	.w7(32'hbb624506),
	.w8(32'hbabc0819),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348f17),
	.w1(32'hba26d82d),
	.w2(32'hb934f856),
	.w3(32'hbb6fbf4f),
	.w4(32'h39ad4429),
	.w5(32'hba31b2cd),
	.w6(32'hb9f95428),
	.w7(32'hba3421b6),
	.w8(32'hbb17d56d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15215f),
	.w1(32'hbb682b55),
	.w2(32'hba5583a7),
	.w3(32'hba8b81f4),
	.w4(32'h3a8659b8),
	.w5(32'h3a7a494b),
	.w6(32'h3adc654b),
	.w7(32'h3a3b3793),
	.w8(32'h3b3c9865),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07beab),
	.w1(32'hbb94a442),
	.w2(32'hbb5ac327),
	.w3(32'h3b3cd19c),
	.w4(32'hbb82c381),
	.w5(32'hbb8f6fca),
	.w6(32'hbb6521f8),
	.w7(32'hbb349f28),
	.w8(32'h3a097fe9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8170c),
	.w1(32'h3a144818),
	.w2(32'h3af4645f),
	.w3(32'hbb26e764),
	.w4(32'h3ab5bfca),
	.w5(32'h3b32f1ee),
	.w6(32'h3ad0c62a),
	.w7(32'h3b1b24ab),
	.w8(32'h3b5cee1c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55bccb),
	.w1(32'hbaa31189),
	.w2(32'h3b00d572),
	.w3(32'h3b7667a8),
	.w4(32'hba1f68b9),
	.w5(32'h3a165367),
	.w6(32'h3aae287d),
	.w7(32'hb80add1e),
	.w8(32'h3a874bc3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b9c4e),
	.w1(32'hbb36b06b),
	.w2(32'hbbcac0ef),
	.w3(32'hba7f9e88),
	.w4(32'hbb689afb),
	.w5(32'hbb8b4468),
	.w6(32'hbb21966e),
	.w7(32'hbba1db6c),
	.w8(32'hbb7866a7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c35da),
	.w1(32'hba87c7a2),
	.w2(32'hba381766),
	.w3(32'hbb8788ce),
	.w4(32'hbabc8202),
	.w5(32'hba5731a8),
	.w6(32'hbac818c6),
	.w7(32'hba881caf),
	.w8(32'hba84d6a7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b3ea6),
	.w1(32'h3c2b1dd3),
	.w2(32'h3b561c5c),
	.w3(32'hba327dd6),
	.w4(32'h3c1092de),
	.w5(32'h3bd00a6f),
	.w6(32'h3be852f3),
	.w7(32'h3a7d6481),
	.w8(32'hbbdce43b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8a855),
	.w1(32'hbacba4f4),
	.w2(32'hba67610b),
	.w3(32'hbb04f6fa),
	.w4(32'hbb02bd5a),
	.w5(32'hbaec400f),
	.w6(32'hbb43e233),
	.w7(32'hbaf1562f),
	.w8(32'h3a8123d8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca864e),
	.w1(32'h3abae82c),
	.w2(32'h3b8006f2),
	.w3(32'hba4650a8),
	.w4(32'h3a8fbff3),
	.w5(32'h3b1b062d),
	.w6(32'h3a887284),
	.w7(32'h3ba7dca3),
	.w8(32'hbb2bc838),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d2d35),
	.w1(32'hba6b5bbd),
	.w2(32'hbb0dfb12),
	.w3(32'hbb1f13e6),
	.w4(32'hbb827c36),
	.w5(32'hbb382368),
	.w6(32'hbb2e0227),
	.w7(32'hbb3bb67d),
	.w8(32'hbb304158),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a90c9),
	.w1(32'h3bde150e),
	.w2(32'h3c8aa62c),
	.w3(32'hbb39823b),
	.w4(32'h3b20efb3),
	.w5(32'h3c574cf9),
	.w6(32'h3b687fbe),
	.w7(32'h3c43e160),
	.w8(32'h3b8a1ea8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ee5a),
	.w1(32'hba701f4d),
	.w2(32'h3ae81cbf),
	.w3(32'h3bc3a981),
	.w4(32'h3a541d7d),
	.w5(32'h3ae15da0),
	.w6(32'h389e4269),
	.w7(32'h3984845a),
	.w8(32'h39b847db),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc8949),
	.w1(32'hbbac8a33),
	.w2(32'hbb834179),
	.w3(32'h3b2a889a),
	.w4(32'hbb3ea19f),
	.w5(32'hbb56af1a),
	.w6(32'hbb3adacd),
	.w7(32'hbb0a93f9),
	.w8(32'hbb0e805f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fe876),
	.w1(32'hba5ba69c),
	.w2(32'hbb298f0a),
	.w3(32'hbb65d025),
	.w4(32'hba776a3e),
	.w5(32'hbb474aa2),
	.w6(32'h3ac461dd),
	.w7(32'hba7dfe4d),
	.w8(32'h39833b72),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07caa0),
	.w1(32'h3a427857),
	.w2(32'h3a99209d),
	.w3(32'hba941b6b),
	.w4(32'h39780803),
	.w5(32'hbabb0a68),
	.w6(32'hbb3b2de6),
	.w7(32'h38ae3bb3),
	.w8(32'h39e8d5cb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89849b),
	.w1(32'h39c55be6),
	.w2(32'h39b77e42),
	.w3(32'hba157845),
	.w4(32'hb94d9d8f),
	.w5(32'hba084fab),
	.w6(32'hb9d4544e),
	.w7(32'hba4a915e),
	.w8(32'hb890f98e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946d29b),
	.w1(32'h3845e68f),
	.w2(32'hbadf0f3d),
	.w3(32'hb9d04bb2),
	.w4(32'hb90a2f79),
	.w5(32'h3a4e9cdb),
	.w6(32'hbaec9458),
	.w7(32'hbb15d0cc),
	.w8(32'hbbb0f8c0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9368aa),
	.w1(32'hbbb8ca5d),
	.w2(32'hbb9c94ed),
	.w3(32'hbb208ed1),
	.w4(32'hbb9f0619),
	.w5(32'hbb9d3d2e),
	.w6(32'hbbd61636),
	.w7(32'hbbc0f675),
	.w8(32'hbbccb513),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb05e),
	.w1(32'h3b119e90),
	.w2(32'h3b81229e),
	.w3(32'hbbc929a0),
	.w4(32'h3afdf0eb),
	.w5(32'h3b8f3596),
	.w6(32'h3aa92051),
	.w7(32'h3b5f02e0),
	.w8(32'h3905b2cc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93d31),
	.w1(32'h3a860e46),
	.w2(32'h3b6e1e56),
	.w3(32'hbb0aeda4),
	.w4(32'h3ae85419),
	.w5(32'h3bb488cf),
	.w6(32'h3b08087a),
	.w7(32'h3a66eff3),
	.w8(32'hbb0924e2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a10e8),
	.w1(32'h3b078552),
	.w2(32'h3aca6b11),
	.w3(32'h399c4dd6),
	.w4(32'hb9d48ef4),
	.w5(32'hba924799),
	.w6(32'hbaa6e617),
	.w7(32'h39d002f5),
	.w8(32'hbb168462),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e2f5),
	.w1(32'hbb30c4e5),
	.w2(32'hbb074153),
	.w3(32'hba3b77c0),
	.w4(32'hbb018d23),
	.w5(32'h3ac627da),
	.w6(32'hbaf80198),
	.w7(32'hbab85ae3),
	.w8(32'h3aea154f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9264ac),
	.w1(32'hbbbb758c),
	.w2(32'h398b0d13),
	.w3(32'h39aac210),
	.w4(32'hbbb0dcb8),
	.w5(32'hb9931a45),
	.w6(32'hbb9f2181),
	.w7(32'h3a879ae1),
	.w8(32'h3b0ce334),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a7e0f),
	.w1(32'hbadac5b2),
	.w2(32'hbae8894f),
	.w3(32'hba195b0e),
	.w4(32'hbaee9924),
	.w5(32'hbb094a34),
	.w6(32'hbad98539),
	.w7(32'hbb04336c),
	.w8(32'hbb045495),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9b87e),
	.w1(32'hbab51bab),
	.w2(32'hbb3b1c77),
	.w3(32'hbb1eb50c),
	.w4(32'hbb76e488),
	.w5(32'hbb9072bb),
	.w6(32'hbb3329ab),
	.w7(32'hbb0aedf2),
	.w8(32'h3984185e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284077),
	.w1(32'h3ab9f253),
	.w2(32'h393749cd),
	.w3(32'hbad0ee54),
	.w4(32'hbac19abf),
	.w5(32'hbaefbf0a),
	.w6(32'h39c6407d),
	.w7(32'hba7d1ea3),
	.w8(32'hbb134e61),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77d4ae),
	.w1(32'hb9a94b3d),
	.w2(32'h3b124d9c),
	.w3(32'hbb8f429b),
	.w4(32'hb9f597f3),
	.w5(32'h38ce6aa2),
	.w6(32'h3b03fca6),
	.w7(32'h3b936487),
	.w8(32'h3b87d24c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83eff2),
	.w1(32'hbacb699a),
	.w2(32'hbbcae288),
	.w3(32'h3aaa5eed),
	.w4(32'hbaf106ae),
	.w5(32'hbbd0c9c2),
	.w6(32'hbb50c539),
	.w7(32'hbba9215c),
	.w8(32'hbaf2e85a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c633d),
	.w1(32'h3a2e2a08),
	.w2(32'h3abd3af8),
	.w3(32'hbb110592),
	.w4(32'hb9c3ee7b),
	.w5(32'h3a1b2692),
	.w6(32'h378505ab),
	.w7(32'h39b3e922),
	.w8(32'h3901c7b0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa14fee),
	.w1(32'h3b058a29),
	.w2(32'h3abbb4f7),
	.w3(32'h3a8cfea4),
	.w4(32'h3a4a4091),
	.w5(32'h3a06c251),
	.w6(32'h3a27f887),
	.w7(32'h3a0bac9d),
	.w8(32'h3ae96e39),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f7965),
	.w1(32'hbb7af796),
	.w2(32'hbb4f4cd6),
	.w3(32'h3b010b6a),
	.w4(32'hbaf7490a),
	.w5(32'hbbaaec9b),
	.w6(32'hbb5f55d8),
	.w7(32'hbb8617bc),
	.w8(32'hbb05141a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ecf29),
	.w1(32'hbbb7e881),
	.w2(32'hbb8e411e),
	.w3(32'hbb8c645a),
	.w4(32'hbbd053dc),
	.w5(32'hbbfc8f82),
	.w6(32'hbaf28335),
	.w7(32'h39a17639),
	.w8(32'hba98d2f8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe37e),
	.w1(32'hbb13b669),
	.w2(32'h3b8b510f),
	.w3(32'hbb58ac6e),
	.w4(32'hbb6c9726),
	.w5(32'hb98676f9),
	.w6(32'hbaade6dc),
	.w7(32'hb88aae33),
	.w8(32'h3a7bc101),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac82f8b),
	.w1(32'h391521bb),
	.w2(32'hbb467592),
	.w3(32'h39d999c3),
	.w4(32'hba898b6c),
	.w5(32'hbb8e2b51),
	.w6(32'hbb1a84f1),
	.w7(32'hbb00f7b0),
	.w8(32'hbb172cad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab81ba),
	.w1(32'h3a9f2a3f),
	.w2(32'h3ad41dcc),
	.w3(32'hbb708436),
	.w4(32'hba5f34b8),
	.w5(32'hb89c67a4),
	.w6(32'h3ac096bd),
	.w7(32'h3b72965f),
	.w8(32'h3b6c27f4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44c9b6),
	.w1(32'h3b86b1c6),
	.w2(32'h3b5cef97),
	.w3(32'h3aaf39d9),
	.w4(32'h3b3e3b85),
	.w5(32'h3ba9e820),
	.w6(32'h3b979eeb),
	.w7(32'h3b1d745d),
	.w8(32'hbad9b58a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7923dd),
	.w1(32'h3ae41e98),
	.w2(32'h3acccd47),
	.w3(32'h3a762eb7),
	.w4(32'hb969a0f0),
	.w5(32'h3b679551),
	.w6(32'h3aefedfd),
	.w7(32'h3af8aecd),
	.w8(32'hb9017b3f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375026bb),
	.w1(32'h3b0b502f),
	.w2(32'h3b154713),
	.w3(32'h3bb56069),
	.w4(32'hba6ccf07),
	.w5(32'hba6ccc96),
	.w6(32'h3a9291ba),
	.w7(32'h3ab2f3e3),
	.w8(32'h39c0e03a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a864b8c),
	.w1(32'hbb7be2b8),
	.w2(32'h3b0a88eb),
	.w3(32'h3a301d8e),
	.w4(32'hbb4fe099),
	.w5(32'h3b3aac6c),
	.w6(32'hbb57ca2f),
	.w7(32'h3ab8a19a),
	.w8(32'hba60ba44),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854512),
	.w1(32'h3b33356b),
	.w2(32'h391e85d9),
	.w3(32'hb9b60a33),
	.w4(32'h3abb407a),
	.w5(32'h3ab22f1d),
	.w6(32'h3a85cc0f),
	.w7(32'hba02f081),
	.w8(32'hbbb536be),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a88e),
	.w1(32'h3ae2d742),
	.w2(32'h3b67e74e),
	.w3(32'hbb90b9e8),
	.w4(32'h3b8b5f07),
	.w5(32'h3bbcfc27),
	.w6(32'h3a8967fe),
	.w7(32'h3aa35dbb),
	.w8(32'h3b069db3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1f408),
	.w1(32'hbb5dc6f3),
	.w2(32'hbb268492),
	.w3(32'h3b49151a),
	.w4(32'hbb046720),
	.w5(32'hbb00f22b),
	.w6(32'hbb81bc47),
	.w7(32'hbb009e54),
	.w8(32'h39103996),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8940ca),
	.w1(32'h39855756),
	.w2(32'hb9644882),
	.w3(32'hb9d020ee),
	.w4(32'hb8fdeda7),
	.w5(32'h39d7b4cb),
	.w6(32'hba40d6e9),
	.w7(32'hbb096acf),
	.w8(32'hb9acb515),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba123735),
	.w1(32'h3ae399e8),
	.w2(32'h3b16a31b),
	.w3(32'hba8be83a),
	.w4(32'h3a952839),
	.w5(32'h3b30de01),
	.w6(32'hb9cec7f3),
	.w7(32'h3a2fab4a),
	.w8(32'hbb9b5c07),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53d65c),
	.w1(32'h3b96333e),
	.w2(32'h3b44d2b3),
	.w3(32'hbb23be8f),
	.w4(32'h3b31bb8f),
	.w5(32'hba1633e0),
	.w6(32'h3ae64bf0),
	.w7(32'h3ad6e456),
	.w8(32'hbb3f9a1c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be10dd),
	.w1(32'h3aaa660b),
	.w2(32'h3b053e2d),
	.w3(32'h3a855cb6),
	.w4(32'h3922db5a),
	.w5(32'h3ac3e8ef),
	.w6(32'h3b18dc6d),
	.w7(32'h3af8652e),
	.w8(32'h3997b3da),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fde75),
	.w1(32'h3a9740af),
	.w2(32'h3b2080d1),
	.w3(32'h3a3791a5),
	.w4(32'hbadd2a8b),
	.w5(32'h3a8219f4),
	.w6(32'h3a471041),
	.w7(32'h3b437474),
	.w8(32'h3a1b79d0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6f49),
	.w1(32'h3b3b62c7),
	.w2(32'h3b88b452),
	.w3(32'h3b2f5604),
	.w4(32'h3b72e1a9),
	.w5(32'h3b4524f6),
	.w6(32'h3b147ad9),
	.w7(32'h3b271c97),
	.w8(32'hbb85e743),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed4c2),
	.w1(32'hb80eb7dc),
	.w2(32'h3b3c5f13),
	.w3(32'hbb104737),
	.w4(32'hb9c720bc),
	.w5(32'h3aaa4a62),
	.w6(32'h3a8a6ae0),
	.w7(32'h388b6f5d),
	.w8(32'h3aad4ac4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975e0ee),
	.w1(32'h3b31293e),
	.w2(32'h3b40a04a),
	.w3(32'hbb5aac89),
	.w4(32'h3b3352fe),
	.w5(32'hba41fe13),
	.w6(32'h3a010750),
	.w7(32'h3a91707d),
	.w8(32'hbb0996a6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375fdcc3),
	.w1(32'hbb27a26f),
	.w2(32'hbb14bef6),
	.w3(32'h3ab3f0dd),
	.w4(32'hbb045189),
	.w5(32'hbb0a5993),
	.w6(32'h3b0b83dc),
	.w7(32'h3a5de863),
	.w8(32'h3aa349c9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac17954),
	.w1(32'h3a9a76ad),
	.w2(32'hba9337d9),
	.w3(32'h3a67f8f5),
	.w4(32'h3b0675d0),
	.w5(32'h3a6949f4),
	.w6(32'hb9697e29),
	.w7(32'hbb27b82b),
	.w8(32'hbb8dbcbb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61c86c),
	.w1(32'hba3b3f41),
	.w2(32'hbaaec295),
	.w3(32'hba7f60b4),
	.w4(32'hbb92ded3),
	.w5(32'hbbbd312e),
	.w6(32'h3a9b56ad),
	.w7(32'h3ad0ce30),
	.w8(32'h3b83191d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a71e),
	.w1(32'hb9cc1761),
	.w2(32'hb9f4c605),
	.w3(32'hbb57456c),
	.w4(32'h3a11780d),
	.w5(32'h3a59e201),
	.w6(32'hbad4fbf8),
	.w7(32'hbaff34da),
	.w8(32'hbb44d18a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9e1f),
	.w1(32'h3a0bbba2),
	.w2(32'h3b56d928),
	.w3(32'h395cefd7),
	.w4(32'h3b03378e),
	.w5(32'h3a8fadf7),
	.w6(32'h3ac3b856),
	.w7(32'h3ab85e1b),
	.w8(32'h3b125122),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399918c5),
	.w1(32'h3a149894),
	.w2(32'h3985e527),
	.w3(32'hbae5243a),
	.w4(32'h3b48f685),
	.w5(32'h3b848545),
	.w6(32'hbb012d98),
	.w7(32'hbb1ed72f),
	.w8(32'hba19d0a0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa28de4),
	.w1(32'hbad6d1d0),
	.w2(32'hbaea904b),
	.w3(32'h39c1c8d5),
	.w4(32'hbaad63ec),
	.w5(32'hbb06f129),
	.w6(32'h3545060b),
	.w7(32'hbb0722e7),
	.w8(32'hbad91fc8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05cb98),
	.w1(32'hbab8253a),
	.w2(32'hba56cb28),
	.w3(32'hbb0e453f),
	.w4(32'hba824ab4),
	.w5(32'hba0a4203),
	.w6(32'hba43bd44),
	.w7(32'hb9db1293),
	.w8(32'hba90ce6d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0c847),
	.w1(32'h3a335dad),
	.w2(32'hb9df9991),
	.w3(32'hba5c7d71),
	.w4(32'h3b1417d7),
	.w5(32'hb9f375e3),
	.w6(32'h3a3aaf10),
	.w7(32'hba5b882d),
	.w8(32'h38d0db25),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9cf4d),
	.w1(32'hbab377d5),
	.w2(32'h381ce351),
	.w3(32'h3a7589ea),
	.w4(32'h3a803b39),
	.w5(32'h3a0ec987),
	.w6(32'hbb2fd847),
	.w7(32'hba0022c8),
	.w8(32'hbafc662d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56b6f7),
	.w1(32'hbb8491f5),
	.w2(32'hbb8316e3),
	.w3(32'h38f0509a),
	.w4(32'hbb72eb06),
	.w5(32'hbb5b3a70),
	.w6(32'hbb86d51b),
	.w7(32'hbb77f191),
	.w8(32'hba4670e4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00993b),
	.w1(32'hbb0a3eee),
	.w2(32'hbaa5d4ba),
	.w3(32'hba1cea6d),
	.w4(32'h3a423750),
	.w5(32'hba4d3867),
	.w6(32'h384b7b2c),
	.w7(32'hbb0dec3d),
	.w8(32'h39d1a2db),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d1fc9),
	.w1(32'hbb421d02),
	.w2(32'h3ab6a8a6),
	.w3(32'hb8d503f1),
	.w4(32'h3ae080f6),
	.w5(32'h3b8e191e),
	.w6(32'hbb3cbb26),
	.w7(32'h390b8492),
	.w8(32'h390c90c9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecdfc2),
	.w1(32'hb9a756d7),
	.w2(32'h3ad91d2b),
	.w3(32'h3b35dadc),
	.w4(32'h3b1294fb),
	.w5(32'h3b3a98c4),
	.w6(32'hbaa87a42),
	.w7(32'h3accee54),
	.w8(32'h3b43569f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be38d),
	.w1(32'h3a105524),
	.w2(32'h3a331877),
	.w3(32'h3bc0ce0f),
	.w4(32'hba44feb2),
	.w5(32'hbb3c50e5),
	.w6(32'hb9e13ff0),
	.w7(32'hb9be345e),
	.w8(32'hb93df0cb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e6f19),
	.w1(32'h3b35a5e6),
	.w2(32'h3b2c8b78),
	.w3(32'hba253323),
	.w4(32'hbab6eb94),
	.w5(32'h39a8a212),
	.w6(32'h3b4f7c15),
	.w7(32'h3b50ba87),
	.w8(32'hbb75bc9f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a2378),
	.w1(32'hb914afea),
	.w2(32'hbb5340e7),
	.w3(32'hbbca57a3),
	.w4(32'hbacffcb4),
	.w5(32'hba2e7464),
	.w6(32'hb992997c),
	.w7(32'hbb2dddfb),
	.w8(32'hb714ac85),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293a21),
	.w1(32'h39c1a8c5),
	.w2(32'h399ca396),
	.w3(32'hbb868fae),
	.w4(32'h397c153d),
	.w5(32'hbb5f56c6),
	.w6(32'h3b00a3b2),
	.w7(32'h38e0f5d4),
	.w8(32'hbaa6a155),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0372fc),
	.w1(32'h3b97e515),
	.w2(32'h3b81a655),
	.w3(32'hb96a74da),
	.w4(32'h39865250),
	.w5(32'h3abff0bb),
	.w6(32'h382fe119),
	.w7(32'h384a78ba),
	.w8(32'h38c741cd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb4cbb),
	.w1(32'h3a95354c),
	.w2(32'h3b9a2791),
	.w3(32'hba1c82ff),
	.w4(32'h3b970062),
	.w5(32'h3bc2d5d8),
	.w6(32'h3a450edb),
	.w7(32'h3b899d48),
	.w8(32'h393d5ec2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18cf76),
	.w1(32'h3a2b89ad),
	.w2(32'h3c227f74),
	.w3(32'h3ad8e097),
	.w4(32'hbb1defba),
	.w5(32'h3be59106),
	.w6(32'hbad9dd44),
	.w7(32'h3bb9cc30),
	.w8(32'h3ab3af4b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8655bd),
	.w1(32'hb937e2cb),
	.w2(32'hbae556d2),
	.w3(32'h3b2e18ed),
	.w4(32'hbb09bbb7),
	.w5(32'hba7c129b),
	.w6(32'hb9d65bc5),
	.w7(32'hbab15a7e),
	.w8(32'hbacb0f03),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b28f),
	.w1(32'hbab65ff0),
	.w2(32'h3a62eebb),
	.w3(32'h39a435fd),
	.w4(32'hbb07a9d5),
	.w5(32'hbac87627),
	.w6(32'hbb828e57),
	.w7(32'hbaaf5f12),
	.w8(32'h392dccfd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f92be),
	.w1(32'hba60634d),
	.w2(32'hbb944434),
	.w3(32'h3a255495),
	.w4(32'hb8bf1d1e),
	.w5(32'hbb8368c5),
	.w6(32'hb8edecdf),
	.w7(32'hbb15cc57),
	.w8(32'h3aaee258),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13cae1),
	.w1(32'hbb99bbf6),
	.w2(32'hbc008cd5),
	.w3(32'h3a169139),
	.w4(32'hbb448994),
	.w5(32'hbbc16f8a),
	.w6(32'hbbb276e7),
	.w7(32'hbbf13d12),
	.w8(32'hbbb2a686),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaea8d),
	.w1(32'hbb1d07a8),
	.w2(32'hbb1cd11b),
	.w3(32'hbb9366a1),
	.w4(32'hbb03c4c6),
	.w5(32'h3a608643),
	.w6(32'h3b4417e4),
	.w7(32'h3b13eaf3),
	.w8(32'h3ab33ca7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c86b),
	.w1(32'h3b941d83),
	.w2(32'h3b85c44e),
	.w3(32'h3af82f93),
	.w4(32'h3b67f34c),
	.w5(32'h3b382087),
	.w6(32'h3b850554),
	.w7(32'h3b7894d6),
	.w8(32'h3b1d3f00),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13b509),
	.w1(32'hbb35e203),
	.w2(32'h3ade5831),
	.w3(32'h3b11eecf),
	.w4(32'h3a3d5dbb),
	.w5(32'hb9e18e62),
	.w6(32'hbb21a02e),
	.w7(32'hbaa79120),
	.w8(32'hbb4cd25c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080247),
	.w1(32'hb9dc56d5),
	.w2(32'hba0e8638),
	.w3(32'hbb780242),
	.w4(32'hbb3de44e),
	.w5(32'hbaa6e238),
	.w6(32'hbb3d3ee7),
	.w7(32'hba970b04),
	.w8(32'hba6a01f2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fea44),
	.w1(32'h3b18ec2d),
	.w2(32'h38418188),
	.w3(32'hb9d2d3fc),
	.w4(32'h3b25c149),
	.w5(32'h3b0cb24a),
	.w6(32'h3908e24f),
	.w7(32'hba49c17b),
	.w8(32'hbb8e5c19),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cbec),
	.w1(32'hbb8c46a6),
	.w2(32'hbbf2916d),
	.w3(32'hbb1dca3d),
	.w4(32'hbb52ebef),
	.w5(32'hbbdc4eab),
	.w6(32'hbba56279),
	.w7(32'hbbe5a8fc),
	.w8(32'hbb9d6622),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f65aa),
	.w1(32'hba827349),
	.w2(32'hbacadc74),
	.w3(32'hbba377d6),
	.w4(32'hba4ad4be),
	.w5(32'hba1f1e4e),
	.w6(32'hba81c965),
	.w7(32'hbacc0b69),
	.w8(32'hbb349045),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec221),
	.w1(32'h38e9895f),
	.w2(32'h398688c3),
	.w3(32'hbabd5e46),
	.w4(32'hbb1f3e66),
	.w5(32'h3aae4576),
	.w6(32'hb95ff275),
	.w7(32'h3b3091fe),
	.w8(32'h3a5e6ef8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f82986),
	.w1(32'hbb3f03d7),
	.w2(32'hbb88b3ed),
	.w3(32'hba51df96),
	.w4(32'hba3367e0),
	.w5(32'hbbbb0c26),
	.w6(32'hba850b8d),
	.w7(32'hbb490492),
	.w8(32'hbb38797f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb666372),
	.w1(32'h3a7b3d07),
	.w2(32'h3ad6632e),
	.w3(32'hbb22315d),
	.w4(32'h3a5023cb),
	.w5(32'h3af71cd8),
	.w6(32'hb99f3af5),
	.w7(32'hb95afadc),
	.w8(32'hbb6d6de0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514488),
	.w1(32'h3b2d980d),
	.w2(32'hbac433ca),
	.w3(32'hbb2c205f),
	.w4(32'hb91487ce),
	.w5(32'hbb7ab6cd),
	.w6(32'h3b0635a1),
	.w7(32'h3b2473a1),
	.w8(32'hb9ca7677),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7be5d),
	.w1(32'h3a963cc7),
	.w2(32'h3b745de2),
	.w3(32'hba410d6d),
	.w4(32'h3b033aef),
	.w5(32'h3a02a50f),
	.w6(32'h3aa456f1),
	.w7(32'h39ab17d2),
	.w8(32'h3a1190a5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2b832),
	.w1(32'hb980e293),
	.w2(32'hba3151ce),
	.w3(32'h3b3fad1f),
	.w4(32'h395b7f06),
	.w5(32'hba300bf3),
	.w6(32'hb9928145),
	.w7(32'hba1944fe),
	.w8(32'h396d73c6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a682f68),
	.w1(32'hbb300290),
	.w2(32'hbaba8851),
	.w3(32'h3a2cdcc4),
	.w4(32'hbb75247b),
	.w5(32'hb8b0c6bc),
	.w6(32'hbb318437),
	.w7(32'h3a9d3eb8),
	.w8(32'hba9b3559),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f2d57),
	.w1(32'hbb53fd15),
	.w2(32'h3b09136f),
	.w3(32'hbb13ad97),
	.w4(32'h39276f74),
	.w5(32'h3ad79980),
	.w6(32'hba0748d0),
	.w7(32'h3a5b5574),
	.w8(32'hbae9ef35),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba975c5b),
	.w1(32'hbb246abd),
	.w2(32'hbb36a441),
	.w3(32'h38b431f2),
	.w4(32'hbb746021),
	.w5(32'hbbab1b9b),
	.w6(32'hbb28953b),
	.w7(32'hb9c07863),
	.w8(32'hba047367),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eef9c),
	.w1(32'h3a13ffce),
	.w2(32'hbad72577),
	.w3(32'hbba722d1),
	.w4(32'h3a84e306),
	.w5(32'hb9a629e8),
	.w6(32'hb9d36e91),
	.w7(32'h3a185a8a),
	.w8(32'hb8fb3e80),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d1136),
	.w1(32'h3bfd9f7a),
	.w2(32'h3b0b5c3a),
	.w3(32'h3a33d99e),
	.w4(32'hbac74e99),
	.w5(32'hbc9c60a4),
	.w6(32'h3b9a4a88),
	.w7(32'h3c601521),
	.w8(32'h3c7f82a9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule