module layer_8_featuremap_192(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd9724),
	.w1(32'hbc355340),
	.w2(32'hbb0ab0b5),
	.w3(32'h3bc8742f),
	.w4(32'hbbdc6a10),
	.w5(32'hbbb573ab),
	.w6(32'hbc02310d),
	.w7(32'hbb83c91d),
	.w8(32'h3b06790c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c05ba),
	.w1(32'h3a96350f),
	.w2(32'h3bac8a77),
	.w3(32'h3bba9767),
	.w4(32'h3975ada4),
	.w5(32'h3b909e12),
	.w6(32'h39ae2fa7),
	.w7(32'hbae0b234),
	.w8(32'hbba1f04c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c8ca),
	.w1(32'h3bb74d84),
	.w2(32'h3bd476d1),
	.w3(32'hb9fdb263),
	.w4(32'h3c150a30),
	.w5(32'h3c348425),
	.w6(32'hbb028890),
	.w7(32'hbb411504),
	.w8(32'hba8b417e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5506),
	.w1(32'hbbea48ad),
	.w2(32'hbc6bb438),
	.w3(32'h3b748b2d),
	.w4(32'h3bf10c20),
	.w5(32'h3c5d5ee6),
	.w6(32'hbc1a3377),
	.w7(32'h3c769507),
	.w8(32'h3cb59c84),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514286),
	.w1(32'hbb4ac389),
	.w2(32'hbb3a6913),
	.w3(32'h3a5a258b),
	.w4(32'h3afdedb7),
	.w5(32'h3a1aa957),
	.w6(32'hbb81552d),
	.w7(32'hba8ce6df),
	.w8(32'hb8713531),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c05ae1),
	.w1(32'hbad47f93),
	.w2(32'hbc0d4ac7),
	.w3(32'hbbc54a54),
	.w4(32'hbbd18d37),
	.w5(32'h3ac39b45),
	.w6(32'hbc249b81),
	.w7(32'hbaaf17c6),
	.w8(32'h3a76153d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0120ae),
	.w1(32'hbb802a7b),
	.w2(32'hbc212d21),
	.w3(32'hbc41f272),
	.w4(32'h3a95a962),
	.w5(32'hbbd1e2ed),
	.w6(32'hba2ed9ad),
	.w7(32'h3b59e39f),
	.w8(32'h3bc322dd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08e2f),
	.w1(32'hbb00820d),
	.w2(32'hbae3a5d1),
	.w3(32'hbbc2ccd3),
	.w4(32'hbbab21eb),
	.w5(32'hbbbeda20),
	.w6(32'h3b66126e),
	.w7(32'h3b8f6dea),
	.w8(32'h3bd217e7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab513fc),
	.w1(32'hbb8b6db6),
	.w2(32'hbbd82915),
	.w3(32'hbaf8f22c),
	.w4(32'h3bdb62da),
	.w5(32'hb8d142a0),
	.w6(32'h3bc99131),
	.w7(32'h3c5f7ae3),
	.w8(32'h3c9c69f5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8645ee),
	.w1(32'hbcc9ebf1),
	.w2(32'hbbbf0e5a),
	.w3(32'hbbb22d5c),
	.w4(32'hbd2258e7),
	.w5(32'hbcf94310),
	.w6(32'hbbb63c33),
	.w7(32'h3c589a03),
	.w8(32'h3c901153),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f3dd4),
	.w1(32'h3cbcdf58),
	.w2(32'h3ca7ff35),
	.w3(32'hbb0ee6c6),
	.w4(32'h3c1c027c),
	.w5(32'h3cbce444),
	.w6(32'h3bcce8ee),
	.w7(32'h3b118991),
	.w8(32'hbc761c83),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aea64),
	.w1(32'hb9b85e3e),
	.w2(32'h3bd2f6c6),
	.w3(32'h3c098ea2),
	.w4(32'hbc71bf55),
	.w5(32'hbb9f1c3a),
	.w6(32'hb9f401f6),
	.w7(32'h3b90408e),
	.w8(32'hbc51f050),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb859155),
	.w1(32'hbba436c0),
	.w2(32'h3ce0b4f5),
	.w3(32'h3ad057e9),
	.w4(32'hbcbc6168),
	.w5(32'hbc566ab4),
	.w6(32'h3ae8b0af),
	.w7(32'h3ca8d0e1),
	.w8(32'h3c95908a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d084cb1),
	.w1(32'hb968b439),
	.w2(32'h3b9bc480),
	.w3(32'h3c304f2f),
	.w4(32'hbc02cc39),
	.w5(32'h3a3a8840),
	.w6(32'hbc4ce7ef),
	.w7(32'hbc597f90),
	.w8(32'hbba9df7d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891783),
	.w1(32'hbbb0661e),
	.w2(32'hbc533086),
	.w3(32'h3bcd887b),
	.w4(32'h3a9ee807),
	.w5(32'hbbfe36bc),
	.w6(32'h3add8072),
	.w7(32'h3b27c1bf),
	.w8(32'h3c20d758),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa33871),
	.w1(32'hb9047451),
	.w2(32'h3c312acc),
	.w3(32'hbbcfa43a),
	.w4(32'h3af92781),
	.w5(32'h3b80bc46),
	.w6(32'h3be0b447),
	.w7(32'h3b9a7f9f),
	.w8(32'h3b5a4770),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c9656),
	.w1(32'hbc10874a),
	.w2(32'hbc3a4df3),
	.w3(32'h3c2ed000),
	.w4(32'hbb632fe7),
	.w5(32'hbc30bbae),
	.w6(32'hbb36e23d),
	.w7(32'hbbb672dc),
	.w8(32'hbaab6a7f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2598e5),
	.w1(32'hbbf28127),
	.w2(32'hbadbe68d),
	.w3(32'hbbd4e8b9),
	.w4(32'hbba64076),
	.w5(32'hba7cf983),
	.w6(32'hba942074),
	.w7(32'hbb8aaa24),
	.w8(32'hbc1e2247),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a017b),
	.w1(32'h3c9519e3),
	.w2(32'h3cd28453),
	.w3(32'hba1b36f7),
	.w4(32'hbc7d7930),
	.w5(32'hbbf86604),
	.w6(32'h3c0e793c),
	.w7(32'h3c1c613e),
	.w8(32'h3b64a859),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58e218),
	.w1(32'hba9c0166),
	.w2(32'hbc265c17),
	.w3(32'h3bac40c8),
	.w4(32'h3b5b5177),
	.w5(32'hbc043cfa),
	.w6(32'h3b4e5ec9),
	.w7(32'h3b2fd8ca),
	.w8(32'h3c010d1d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c7b31),
	.w1(32'hbca7f08d),
	.w2(32'hbcea9ca0),
	.w3(32'hbc005e9c),
	.w4(32'hbca31dd4),
	.w5(32'hbce37864),
	.w6(32'hbc0f0170),
	.w7(32'hbacdc471),
	.w8(32'hba5b153d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe742e9),
	.w1(32'h3bc85a8d),
	.w2(32'hbb8ee1d9),
	.w3(32'hbc313382),
	.w4(32'h3afc4f11),
	.w5(32'hb9085a7d),
	.w6(32'h3bfc5e60),
	.w7(32'h3bd298e2),
	.w8(32'h3a919196),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a6e06),
	.w1(32'hbba7faa3),
	.w2(32'hbc5fe114),
	.w3(32'h3bb7984c),
	.w4(32'hbc40b814),
	.w5(32'hbc344549),
	.w6(32'hbb81579e),
	.w7(32'hbb3ddc11),
	.w8(32'hbacc564f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1920d),
	.w1(32'h3b8fc893),
	.w2(32'hbac3c2e8),
	.w3(32'h3bcd0266),
	.w4(32'h3baf3341),
	.w5(32'h3a8ee9a4),
	.w6(32'h3c08403e),
	.w7(32'h3b827ea2),
	.w8(32'hbad17165),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3870),
	.w1(32'h3c27e62a),
	.w2(32'h3b10cea5),
	.w3(32'h3bbc7908),
	.w4(32'h3b965cd2),
	.w5(32'h3c0c7d53),
	.w6(32'hbc1170b3),
	.w7(32'hbc4dd819),
	.w8(32'hbc28aa93),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6ad7),
	.w1(32'h3bb6fc45),
	.w2(32'h3ae25291),
	.w3(32'hbb8ba9cb),
	.w4(32'h3b91f562),
	.w5(32'h3b9906c9),
	.w6(32'hbba3b19f),
	.w7(32'hbc8c8a59),
	.w8(32'hbc67461f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cd517),
	.w1(32'h3b02157f),
	.w2(32'hbc3e07f9),
	.w3(32'hbbf9f65f),
	.w4(32'h3bf3329a),
	.w5(32'h3c634797),
	.w6(32'h3b04500e),
	.w7(32'hbbc27772),
	.w8(32'hbc264276),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c664f),
	.w1(32'hbc82680d),
	.w2(32'hbd050b6a),
	.w3(32'hb99f795b),
	.w4(32'hbc135cf8),
	.w5(32'hbca8bf9f),
	.w6(32'hbc41e4c7),
	.w7(32'hbb8d0e33),
	.w8(32'h3bea0f43),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0affb7),
	.w1(32'hbb5a55b9),
	.w2(32'h3bcd5518),
	.w3(32'hbc89407a),
	.w4(32'hb9fcadc2),
	.w5(32'h3c6b3a4a),
	.w6(32'hbb94c18f),
	.w7(32'hbad9d972),
	.w8(32'hbc14baee),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa30b4),
	.w1(32'hbad9e499),
	.w2(32'hbb28e466),
	.w3(32'h3ba033c8),
	.w4(32'hbb0e2c1c),
	.w5(32'hbaeaa564),
	.w6(32'hbae5979a),
	.w7(32'hba81788a),
	.w8(32'h3bddcd45),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d882a),
	.w1(32'hbc2f1444),
	.w2(32'h3c4d06d3),
	.w3(32'h3c06384a),
	.w4(32'hbcb5f5ec),
	.w5(32'hbc8b23b2),
	.w6(32'hba8aeb5c),
	.w7(32'h3bc28f54),
	.w8(32'hb8a1eb86),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c664478),
	.w1(32'h3c56b279),
	.w2(32'h3c60b703),
	.w3(32'h3b099f52),
	.w4(32'hbad9bc52),
	.w5(32'h3c32a91e),
	.w6(32'hbb9efe6c),
	.w7(32'hbc300771),
	.w8(32'hbc839524),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb9ad8),
	.w1(32'hbbd59eda),
	.w2(32'hbc89461b),
	.w3(32'h3b406fde),
	.w4(32'hbb945f8c),
	.w5(32'hba16d023),
	.w6(32'hbc6bb603),
	.w7(32'hbc898c08),
	.w8(32'hbc491584),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d07d),
	.w1(32'hbb8f9a8c),
	.w2(32'hbc2ad59e),
	.w3(32'hbbe9f79f),
	.w4(32'hbbd29022),
	.w5(32'hbc4f0a77),
	.w6(32'h3a95791a),
	.w7(32'hba15c9c0),
	.w8(32'hbbbe174e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caa834),
	.w1(32'hbb849317),
	.w2(32'h3bcecc45),
	.w3(32'hbbf54e52),
	.w4(32'hbc5f6381),
	.w5(32'hbbc3eeb8),
	.w6(32'hbc040ce5),
	.w7(32'hbb5b37af),
	.w8(32'hbb26009e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd527),
	.w1(32'h3b36024e),
	.w2(32'hbba7f01a),
	.w3(32'hb91ff1ab),
	.w4(32'hba9bfdd8),
	.w5(32'h3ba59188),
	.w6(32'h3bea2cc7),
	.w7(32'h3b047b63),
	.w8(32'hbae80093),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e2149),
	.w1(32'h3c14520a),
	.w2(32'hbb87881f),
	.w3(32'h3b4c90c0),
	.w4(32'h3ca823e8),
	.w5(32'h3c4d00c3),
	.w6(32'hbb45c9c9),
	.w7(32'hbc6589ac),
	.w8(32'hbc50566c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8246f9),
	.w1(32'hbb92d59d),
	.w2(32'hbbf22fae),
	.w3(32'hbb02c025),
	.w4(32'h3a6ae776),
	.w5(32'hbbda094e),
	.w6(32'h3b239e91),
	.w7(32'h3bd73a5d),
	.w8(32'h3c626644),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb89983),
	.w1(32'hba76d64a),
	.w2(32'h3c64b781),
	.w3(32'hbbbe10b4),
	.w4(32'h3b733e90),
	.w5(32'h3b6d6dd1),
	.w6(32'hba2a8c3c),
	.w7(32'h3c48586b),
	.w8(32'h3ad1240c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab00d5b),
	.w1(32'hbb502ec5),
	.w2(32'hbbd0c218),
	.w3(32'h3b51cc71),
	.w4(32'h3b29df41),
	.w5(32'hbb02aa4e),
	.w6(32'hbb72b073),
	.w7(32'hbb161018),
	.w8(32'hbad4eeea),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e561c),
	.w1(32'h38b0664e),
	.w2(32'h3b232302),
	.w3(32'hbb6c35c1),
	.w4(32'hbb86dc84),
	.w5(32'hba87be33),
	.w6(32'hbaf8bca2),
	.w7(32'hbabb8986),
	.w8(32'hbb45ac40),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e64074),
	.w1(32'hbae40d83),
	.w2(32'h3c16d5ea),
	.w3(32'hbaf44fde),
	.w4(32'hbcaa47d8),
	.w5(32'hbccf5615),
	.w6(32'h3c893ba1),
	.w7(32'h3c6975d7),
	.w8(32'h3b76e08d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baafeff),
	.w1(32'h3c6d8bde),
	.w2(32'hbb7301be),
	.w3(32'hbbfa8e04),
	.w4(32'h3c922f28),
	.w5(32'h3c71cc7c),
	.w6(32'h3a98bc28),
	.w7(32'hbc711739),
	.w8(32'hbc43e8f2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca19e5b),
	.w1(32'hbbeaa750),
	.w2(32'h3bc70f2a),
	.w3(32'h3bbadc06),
	.w4(32'hbb616a48),
	.w5(32'h3b0b8c10),
	.w6(32'hbb146885),
	.w7(32'h3ad99831),
	.w8(32'hbc6bacff),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38facc),
	.w1(32'hbc29b40a),
	.w2(32'hbc7bd697),
	.w3(32'h3bda3f81),
	.w4(32'hbaee2925),
	.w5(32'hbc036a9d),
	.w6(32'hbbb00d54),
	.w7(32'hbc479df1),
	.w8(32'hbb7fd9f2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b9983),
	.w1(32'h3b845dd9),
	.w2(32'hbb810045),
	.w3(32'hb69e0227),
	.w4(32'h3bbb8fe9),
	.w5(32'hbb6dfb54),
	.w6(32'h3c019239),
	.w7(32'h3b8079a0),
	.w8(32'h3c075abe),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3941a),
	.w1(32'hbb70accd),
	.w2(32'hbc82db58),
	.w3(32'h3aab9b44),
	.w4(32'h3ba8da2e),
	.w5(32'hbae1d159),
	.w6(32'hbb81bd65),
	.w7(32'hbc37117b),
	.w8(32'hbbc3769e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d37f),
	.w1(32'hbb5c2e1a),
	.w2(32'hbbc9ab54),
	.w3(32'hbb905a16),
	.w4(32'h3ae8a769),
	.w5(32'h3abd861b),
	.w6(32'h3c366f67),
	.w7(32'hbbdcb7c9),
	.w8(32'hbba671e6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e81dc),
	.w1(32'hba9a5efb),
	.w2(32'hba9ee6d7),
	.w3(32'h3bad113d),
	.w4(32'hba100f70),
	.w5(32'hba7c0658),
	.w6(32'h3a6591e0),
	.w7(32'hbc2a653e),
	.w8(32'hbbc061b8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac800c2),
	.w1(32'h3b24f60d),
	.w2(32'h3bf27f7f),
	.w3(32'h3a87a338),
	.w4(32'hbc0782fd),
	.w5(32'h3c5b585d),
	.w6(32'h3988843d),
	.w7(32'hbc503ec7),
	.w8(32'hbc0db4e8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85c0a9),
	.w1(32'hbb9640dc),
	.w2(32'hbb8e12d0),
	.w3(32'hbb9fc7e6),
	.w4(32'hba761c7a),
	.w5(32'h3b7fd6ee),
	.w6(32'hbb014f31),
	.w7(32'h3b54f268),
	.w8(32'hba5493a7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3884),
	.w1(32'h3bd2f953),
	.w2(32'h3c49dccc),
	.w3(32'h399869e3),
	.w4(32'hbc4e8c60),
	.w5(32'hbc64c462),
	.w6(32'h3c6700c5),
	.w7(32'h3c5c9c48),
	.w8(32'h3c2890dc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cfa3a),
	.w1(32'hbb7cf0fa),
	.w2(32'hbb018821),
	.w3(32'hbbde663b),
	.w4(32'h3837382c),
	.w5(32'h3b0122c0),
	.w6(32'hbb34f4af),
	.w7(32'hbb0a5d5e),
	.w8(32'hb9bcb408),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41091),
	.w1(32'hbaad625c),
	.w2(32'hbaca34bb),
	.w3(32'hbabbe361),
	.w4(32'hbb6e5971),
	.w5(32'hbc21db30),
	.w6(32'h3b282abd),
	.w7(32'h3b39ae9f),
	.w8(32'h3b0644cc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84317d),
	.w1(32'hbc5962be),
	.w2(32'hbc441ef9),
	.w3(32'hba3d597f),
	.w4(32'h3b8775ad),
	.w5(32'hbb7a1aec),
	.w6(32'hbb7dfae8),
	.w7(32'hbac98d02),
	.w8(32'hbb20d673),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dee78),
	.w1(32'hbac4927a),
	.w2(32'hbb6d669a),
	.w3(32'hbbbf7e66),
	.w4(32'h3a1a7fc4),
	.w5(32'hbb801adf),
	.w6(32'h3a0a4d0d),
	.w7(32'hbba1eb59),
	.w8(32'hbc011ffa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01cf11),
	.w1(32'h3c576ec3),
	.w2(32'hba56a4bb),
	.w3(32'hbba13558),
	.w4(32'h3c71e91c),
	.w5(32'h3cb90648),
	.w6(32'hbbc0d6a7),
	.w7(32'hbc6fbf69),
	.w8(32'hbc83ab3b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d82fc),
	.w1(32'h3b79d8c2),
	.w2(32'hbbdaacc3),
	.w3(32'h3c3f5b13),
	.w4(32'h3c62ec32),
	.w5(32'h3c396174),
	.w6(32'hbb5603df),
	.w7(32'hbc3f8686),
	.w8(32'hbc80dfd0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d1040),
	.w1(32'hbb25dac0),
	.w2(32'hbbad5ff9),
	.w3(32'h3b57e26c),
	.w4(32'hbb4ff818),
	.w5(32'hbbf2e63c),
	.w6(32'hba0b0113),
	.w7(32'hbb49cb5e),
	.w8(32'hbbc81cc6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa029e),
	.w1(32'h3bb470bd),
	.w2(32'h3b29ab03),
	.w3(32'hbbbac6a6),
	.w4(32'h3bd54ba2),
	.w5(32'h3c013f9d),
	.w6(32'hbb6f1b84),
	.w7(32'hbb329471),
	.w8(32'h3af9d5f5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a340293),
	.w1(32'h3b34757f),
	.w2(32'hbbc7d420),
	.w3(32'h3b08d3a3),
	.w4(32'h3cb5e703),
	.w5(32'h3c950faa),
	.w6(32'hbc0783b5),
	.w7(32'hbbbd4d54),
	.w8(32'h39386a0d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b33d2),
	.w1(32'h3c57d4ca),
	.w2(32'hbc8dbb2b),
	.w3(32'hbb7bef8a),
	.w4(32'h3cb31aa0),
	.w5(32'h3c255469),
	.w6(32'h3b8c3829),
	.w7(32'hbc21aede),
	.w8(32'h3a91fb59),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa4a32),
	.w1(32'h3bbf175e),
	.w2(32'h3c29ad98),
	.w3(32'hbc421b5f),
	.w4(32'hbb66ff00),
	.w5(32'h3b49af7a),
	.w6(32'h3bb9d6af),
	.w7(32'h3c7087df),
	.w8(32'h3c3b4dd8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd31b52),
	.w1(32'h3b992890),
	.w2(32'h3ba1962d),
	.w3(32'h3bf5ee4d),
	.w4(32'h3aad3cf0),
	.w5(32'h3adbff06),
	.w6(32'h3b5f5001),
	.w7(32'h3b03ccc2),
	.w8(32'hbb4cb8b8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884ee0d),
	.w1(32'h39e46382),
	.w2(32'h3b3b9909),
	.w3(32'hbabd82b2),
	.w4(32'hbb8a5a0c),
	.w5(32'hbb0855c0),
	.w6(32'h3b52ab01),
	.w7(32'h3a47c261),
	.w8(32'hbb8fa03d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f903),
	.w1(32'hbb2f6918),
	.w2(32'hb8ef6c5d),
	.w3(32'h3a9f733f),
	.w4(32'hbad0e965),
	.w5(32'hba1eb34c),
	.w6(32'h39508bba),
	.w7(32'hbb947b1a),
	.w8(32'hbb8f9c29),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d54c),
	.w1(32'h3be2dd84),
	.w2(32'h3ae3cb5e),
	.w3(32'h3afa7d01),
	.w4(32'h3c13029c),
	.w5(32'h3c0e304c),
	.w6(32'hbb8e89af),
	.w7(32'hbb982e62),
	.w8(32'hbbe80387),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024f1b),
	.w1(32'hbbedda79),
	.w2(32'hbc81c08d),
	.w3(32'h3a1e3ae7),
	.w4(32'hba7cd98b),
	.w5(32'hbc00bd9a),
	.w6(32'h3ba3dc74),
	.w7(32'h3adf93fd),
	.w8(32'h3b129b97),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997696),
	.w1(32'hbb9aadc3),
	.w2(32'hbc86b8cd),
	.w3(32'hbbf4997e),
	.w4(32'hbc805dec),
	.w5(32'hbc3d7de4),
	.w6(32'hbbcc5081),
	.w7(32'hbcd715a3),
	.w8(32'hbc32ef65),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7c752),
	.w1(32'h39fd3d2e),
	.w2(32'hbbdb7aae),
	.w3(32'hbb89f3ca),
	.w4(32'h3b56fb64),
	.w5(32'h3c67c5c3),
	.w6(32'hbb7a859f),
	.w7(32'hbbc01aca),
	.w8(32'hbbe3f2eb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab437),
	.w1(32'hbbf87171),
	.w2(32'hbb16ec05),
	.w3(32'h3b8150a9),
	.w4(32'hbc1c3f9f),
	.w5(32'hbc9d4b74),
	.w6(32'h3c6bba39),
	.w7(32'h3cafd301),
	.w8(32'h3c96d235),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c263514),
	.w1(32'h3bb4f169),
	.w2(32'h3b727767),
	.w3(32'hbbcad532),
	.w4(32'h3bfef16b),
	.w5(32'h3c2d2e17),
	.w6(32'hbb6dcaeb),
	.w7(32'hbb4984e8),
	.w8(32'h3acb3966),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d317),
	.w1(32'h3bb1b967),
	.w2(32'h3bfd7033),
	.w3(32'h3bbc5a2b),
	.w4(32'h3bdca5f1),
	.w5(32'h3bd54922),
	.w6(32'hbb1f6d18),
	.w7(32'hbc7df768),
	.w8(32'hbc2fc3bb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e21f7a),
	.w1(32'hbc00c26b),
	.w2(32'hbc167018),
	.w3(32'h3bb13ee4),
	.w4(32'hb98b87f2),
	.w5(32'h3890ed5e),
	.w6(32'hbc0378de),
	.w7(32'hbc1d18b1),
	.w8(32'h3b785b63),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c342b0f),
	.w1(32'h3c580db4),
	.w2(32'hba345204),
	.w3(32'h3c5ef942),
	.w4(32'h3bf6b74c),
	.w5(32'hbbfa3850),
	.w6(32'h3c371460),
	.w7(32'h3ba959eb),
	.w8(32'hbac9cd8b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c9ebe),
	.w1(32'hba47da98),
	.w2(32'hba8ba411),
	.w3(32'hbc88e8ec),
	.w4(32'hba434f3b),
	.w5(32'hbbf7b4f9),
	.w6(32'h3a418fa1),
	.w7(32'h3bdef012),
	.w8(32'h3c18a2f9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a079364),
	.w1(32'hbc060f22),
	.w2(32'hbb3b2cad),
	.w3(32'h39b26271),
	.w4(32'hbb200164),
	.w5(32'h3bee363f),
	.w6(32'hbc24dc16),
	.w7(32'hbc307c60),
	.w8(32'hbb9f9267),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ed784),
	.w1(32'h3b155d08),
	.w2(32'hbaf3502e),
	.w3(32'h3c09f16b),
	.w4(32'h3ba81db1),
	.w5(32'h3b53479c),
	.w6(32'hbba69cd7),
	.w7(32'hbc0473c7),
	.w8(32'hbbf85790),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b9e1d),
	.w1(32'hbc624d85),
	.w2(32'h3c07f4ff),
	.w3(32'hbabe1e67),
	.w4(32'hbcdcc07b),
	.w5(32'hbc509c75),
	.w6(32'h3b3a651e),
	.w7(32'h3bf4b255),
	.w8(32'h3c0b1817),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c639afc),
	.w1(32'hbbacddc7),
	.w2(32'hbba89af8),
	.w3(32'h3c2452ba),
	.w4(32'hbbefe4a5),
	.w5(32'hbb28fcc5),
	.w6(32'hbbab3d67),
	.w7(32'h3b8b1d02),
	.w8(32'hbac95330),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d8915),
	.w1(32'hbad7d95e),
	.w2(32'hbba84424),
	.w3(32'h3bdb473b),
	.w4(32'h3bcd9deb),
	.w5(32'h3c859f19),
	.w6(32'hbc5fc947),
	.w7(32'hbc3e3ef5),
	.w8(32'hbc278746),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036084),
	.w1(32'hbc29e888),
	.w2(32'hbcad7d76),
	.w3(32'h3b8820a4),
	.w4(32'hbba993d3),
	.w5(32'hbb87dd0b),
	.w6(32'hbbddf5a4),
	.w7(32'hbcc50bc1),
	.w8(32'hbbafd3c1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf5794),
	.w1(32'hba9756c3),
	.w2(32'hbb7c693a),
	.w3(32'hbc08478c),
	.w4(32'hbbed8372),
	.w5(32'hbc5109df),
	.w6(32'hb9c5e185),
	.w7(32'h3aeebf36),
	.w8(32'hbbb38550),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dbbf5),
	.w1(32'hbb239c05),
	.w2(32'hba194aca),
	.w3(32'hbb111076),
	.w4(32'hbba19537),
	.w5(32'hbb07a91e),
	.w6(32'h3b30c2e6),
	.w7(32'h3bed9657),
	.w8(32'h3c2e0777),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834a47),
	.w1(32'hba2eb52d),
	.w2(32'h3b753bda),
	.w3(32'h3b1acc02),
	.w4(32'h3c05b9d0),
	.w5(32'h3bf5c7b1),
	.w6(32'hbc01a6b8),
	.w7(32'hbc5caf45),
	.w8(32'hbc9333c6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89d1b5),
	.w1(32'hbbf6912a),
	.w2(32'hbbca0cf5),
	.w3(32'h3c3f7857),
	.w4(32'hbc574869),
	.w5(32'hbc8a9633),
	.w6(32'hbc41b318),
	.w7(32'hbbb908f8),
	.w8(32'h39d26a19),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf83138),
	.w1(32'hbc6b69dd),
	.w2(32'h3bb5ae52),
	.w3(32'h3c06ddc7),
	.w4(32'hbceac163),
	.w5(32'hbca882c6),
	.w6(32'h3c280788),
	.w7(32'h3caf1225),
	.w8(32'h3ca0574f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c742c9d),
	.w1(32'h3c8f9cbc),
	.w2(32'hbbc7edf3),
	.w3(32'hbb1c22d0),
	.w4(32'h3c404b25),
	.w5(32'h3bfb2f88),
	.w6(32'h3a184974),
	.w7(32'hbc371cf2),
	.w8(32'hbb5fc5f2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb3c9b),
	.w1(32'hbbc5faa1),
	.w2(32'h3c3686e9),
	.w3(32'hbc4bc76a),
	.w4(32'hbcc6acfb),
	.w5(32'hbc4db665),
	.w6(32'hbb103b8c),
	.w7(32'h3bdbe212),
	.w8(32'h3be224ad),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca082e4),
	.w1(32'h3bd421d7),
	.w2(32'h3c59e50c),
	.w3(32'h3b8a2633),
	.w4(32'h3bfadb1a),
	.w5(32'h3c735a9a),
	.w6(32'hbb66bb55),
	.w7(32'hbc0a1e91),
	.w8(32'h3bb3e385),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b489c93),
	.w1(32'h3b43b0f5),
	.w2(32'h3b9c1ca3),
	.w3(32'hb9787b13),
	.w4(32'h3c0b920b),
	.w5(32'h3b3b156b),
	.w6(32'hbbff6c79),
	.w7(32'hbb12777c),
	.w8(32'hbb912de5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ae86),
	.w1(32'hbc10c483),
	.w2(32'hbc3986f2),
	.w3(32'hbb1a8a36),
	.w4(32'hbbac54ed),
	.w5(32'hbc7d10ab),
	.w6(32'hbbd91fc1),
	.w7(32'hbc1e7bec),
	.w8(32'h379caa49),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4033),
	.w1(32'hba0a8da4),
	.w2(32'h38a951a8),
	.w3(32'hbc370b52),
	.w4(32'hbb8e8723),
	.w5(32'hbb93b889),
	.w6(32'hb8b94645),
	.w7(32'h39dfe15b),
	.w8(32'hbb2c9b5a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96558bf),
	.w1(32'hb9fdad94),
	.w2(32'h3a4e1c40),
	.w3(32'hbbc6abc2),
	.w4(32'hbaf8db3e),
	.w5(32'hba843ef3),
	.w6(32'h38f4f359),
	.w7(32'hbb5a434c),
	.w8(32'hbbd498c8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b717e),
	.w1(32'hbb31ca29),
	.w2(32'hbbd79310),
	.w3(32'h389dbf3f),
	.w4(32'h3c970655),
	.w5(32'h3c80bdb1),
	.w6(32'hbbfab419),
	.w7(32'hbc8ab843),
	.w8(32'hbbe988ca),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0133a),
	.w1(32'hbaaf1ab0),
	.w2(32'h3bb4e24f),
	.w3(32'h3bc0507b),
	.w4(32'h3bbfed00),
	.w5(32'h3c29a16c),
	.w6(32'hbba48539),
	.w7(32'hb83852e6),
	.w8(32'h3b2b6c3c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1fba9),
	.w1(32'hb92653a1),
	.w2(32'hbadf453c),
	.w3(32'h3c381e3e),
	.w4(32'hbbe90153),
	.w5(32'h3b2ba79a),
	.w6(32'h394b99f9),
	.w7(32'hbb2c9ce3),
	.w8(32'hba3a14fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20743c),
	.w1(32'h3b2a9004),
	.w2(32'h3bb49ccd),
	.w3(32'h3bd44bb7),
	.w4(32'hbb1ae4fe),
	.w5(32'h3ae3975d),
	.w6(32'h39a1aa4f),
	.w7(32'h3b8e993e),
	.w8(32'h3aaf5de0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b7ff3),
	.w1(32'hbbca2b97),
	.w2(32'h3b9cac23),
	.w3(32'h3ab2276f),
	.w4(32'h3b1454ad),
	.w5(32'h3b85512d),
	.w6(32'h3bac8180),
	.w7(32'h3bb6dd86),
	.w8(32'h3b46320b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56475b),
	.w1(32'h3b158a52),
	.w2(32'hbc5c2a7a),
	.w3(32'h3ae85548),
	.w4(32'h3c976ab4),
	.w5(32'h3c9f7bdc),
	.w6(32'hbbddbbf2),
	.w7(32'hbcc89e68),
	.w8(32'hbc4d6d90),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a8b19),
	.w1(32'h39ccaef0),
	.w2(32'h3c21896c),
	.w3(32'h3ba29ff0),
	.w4(32'hbc256b65),
	.w5(32'hbb443540),
	.w6(32'h3ae99f3c),
	.w7(32'hbbaaef04),
	.w8(32'hbca28e6a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad86e8f),
	.w1(32'hbb940c3b),
	.w2(32'h3a8a9cf1),
	.w3(32'hbae2516a),
	.w4(32'hbc05698b),
	.w5(32'h3b4ef76e),
	.w6(32'h39c219ec),
	.w7(32'h3b06cc72),
	.w8(32'h383059be),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba842d4f),
	.w1(32'hbc00c05d),
	.w2(32'hbc8b3f89),
	.w3(32'hbb27ce95),
	.w4(32'h38b6895c),
	.w5(32'hbad6a3d9),
	.w6(32'hbae6fe3f),
	.w7(32'hbc00f037),
	.w8(32'hbae8d07f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc856),
	.w1(32'hbc6d3d0c),
	.w2(32'h3aca3d9c),
	.w3(32'hbba58e3d),
	.w4(32'hbc29acea),
	.w5(32'hbba5c84e),
	.w6(32'hbc0c80a5),
	.w7(32'hbb0deef2),
	.w8(32'hbb0b7631),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ac4f),
	.w1(32'h3b980ec9),
	.w2(32'h3b07b7fb),
	.w3(32'hbbe26eb5),
	.w4(32'hbad2d021),
	.w5(32'hba12ca09),
	.w6(32'h3c1fc0a7),
	.w7(32'h3b5b037d),
	.w8(32'h39df61f8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6e33),
	.w1(32'hba77a14b),
	.w2(32'hbc084a76),
	.w3(32'h3b88730d),
	.w4(32'h3b4a2b2a),
	.w5(32'hbb714315),
	.w6(32'h3bcbb4ac),
	.w7(32'h39dc5127),
	.w8(32'h3bd27560),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bc465),
	.w1(32'hbbe6174a),
	.w2(32'h3c599471),
	.w3(32'h3b5504b0),
	.w4(32'hbb42b4c2),
	.w5(32'h3beea67e),
	.w6(32'hbb73fb3b),
	.w7(32'h3c276f73),
	.w8(32'h3b1422e9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eadd9),
	.w1(32'h3c3a536b),
	.w2(32'hbbfb7637),
	.w3(32'h3bb5b533),
	.w4(32'h3ca3cb9e),
	.w5(32'h3c7427cd),
	.w6(32'hbb4c448b),
	.w7(32'hbcc4c69c),
	.w8(32'hbce0f06d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce32dac),
	.w1(32'h3c3ef9a3),
	.w2(32'h3c771891),
	.w3(32'h3aea6391),
	.w4(32'h3c12f9a1),
	.w5(32'h3c31f754),
	.w6(32'h3c5be96d),
	.w7(32'h3c9cc9ea),
	.w8(32'h3cbfa110),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b39c3),
	.w1(32'hb7e013ae),
	.w2(32'h3bdc8cb3),
	.w3(32'h3c56794a),
	.w4(32'hbb4d93d4),
	.w5(32'h3afda847),
	.w6(32'hb9bd08d0),
	.w7(32'h390b11fa),
	.w8(32'hbb6fda1f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb6134),
	.w1(32'hbbfced6b),
	.w2(32'hbc0ddc41),
	.w3(32'h3b6fd08e),
	.w4(32'h3c20c16a),
	.w5(32'hb71ecf59),
	.w6(32'hbb08818f),
	.w7(32'hbc06c412),
	.w8(32'h3975ff44),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5efc2),
	.w1(32'h3b07415c),
	.w2(32'h3973c6c8),
	.w3(32'hbaca14ab),
	.w4(32'hb9bb89b5),
	.w5(32'hb93cc2ad),
	.w6(32'h39c068e0),
	.w7(32'h3a1d3bd2),
	.w8(32'hbb2b3063),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2430a9),
	.w1(32'h3b857955),
	.w2(32'h3c2029aa),
	.w3(32'hbafdb725),
	.w4(32'h3b8f8677),
	.w5(32'h3c23e42f),
	.w6(32'h3bd37ba9),
	.w7(32'h3bfcf9ac),
	.w8(32'h3bbb3c94),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b1454),
	.w1(32'h3cbfb143),
	.w2(32'h3cb86e71),
	.w3(32'h3bd39117),
	.w4(32'h3c88e7d8),
	.w5(32'h3c8e9381),
	.w6(32'h3a343473),
	.w7(32'hbc4345cb),
	.w8(32'hbc684245),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d2ba8),
	.w1(32'hbc0fedb4),
	.w2(32'h3c403723),
	.w3(32'h3c11301e),
	.w4(32'hbd02946b),
	.w5(32'hbcb80504),
	.w6(32'h3b8353c8),
	.w7(32'h3c27679d),
	.w8(32'h3b8d5cdb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8556d7),
	.w1(32'h3b0108d4),
	.w2(32'h3c0535c6),
	.w3(32'hba7e662e),
	.w4(32'hbae8deb0),
	.w5(32'h3ba1b35e),
	.w6(32'h3a082a5b),
	.w7(32'h3aa9e394),
	.w8(32'hbb43a0cd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aacdd),
	.w1(32'h3c5ad550),
	.w2(32'h3bd34db0),
	.w3(32'h3b8616cf),
	.w4(32'h3cf03c35),
	.w5(32'h3c9bf506),
	.w6(32'h3bba80f0),
	.w7(32'hbb4d7db4),
	.w8(32'h3ba85d6e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388abca6),
	.w1(32'h3be25070),
	.w2(32'hb9c1fe11),
	.w3(32'hbaf7793e),
	.w4(32'h3b890261),
	.w5(32'h3bcffa05),
	.w6(32'h3bc82896),
	.w7(32'h3bfb455b),
	.w8(32'h3b932107),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dd16c),
	.w1(32'h3c883d95),
	.w2(32'h3c992e65),
	.w3(32'h3ba135cf),
	.w4(32'hbb8eba62),
	.w5(32'h3cce7f41),
	.w6(32'hbc505ed6),
	.w7(32'hbc096ca4),
	.w8(32'hbc195969),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0766dd),
	.w1(32'h3bb3236e),
	.w2(32'h3b03c1db),
	.w3(32'h3c6cc99c),
	.w4(32'h3a863bd6),
	.w5(32'hbbbc336b),
	.w6(32'h3c1709e1),
	.w7(32'h3be085e9),
	.w8(32'h3a81caa7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0986e),
	.w1(32'hbc862579),
	.w2(32'hbca14bb9),
	.w3(32'hbc21b2ec),
	.w4(32'hbc603f44),
	.w5(32'hbbf4b23d),
	.w6(32'hbba6607a),
	.w7(32'hbca94e0f),
	.w8(32'hbc5fd49e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d374e),
	.w1(32'hbb135008),
	.w2(32'h3bc6c1b5),
	.w3(32'h3a58f7c2),
	.w4(32'h3b8e0897),
	.w5(32'h3b8c4985),
	.w6(32'hbb22350c),
	.w7(32'hbb6bfadd),
	.w8(32'hbc241017),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ca59b),
	.w1(32'h3b380c36),
	.w2(32'h3b38265c),
	.w3(32'h3ab7c012),
	.w4(32'h39146dc8),
	.w5(32'h3b51ad0c),
	.w6(32'h3b56383d),
	.w7(32'h3b0376ca),
	.w8(32'hbb6a20a8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74b489),
	.w1(32'h3c30f0a6),
	.w2(32'h3b9ee530),
	.w3(32'hba4b11fe),
	.w4(32'h3ba7df9c),
	.w5(32'h3bedd68b),
	.w6(32'h3c37c0e9),
	.w7(32'h3c0b60b6),
	.w8(32'h3bbe3500),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c013e3a),
	.w1(32'h3c2b90c8),
	.w2(32'h3baaa079),
	.w3(32'h3beac1fe),
	.w4(32'h3c7afe62),
	.w5(32'h3c0b5ac9),
	.w6(32'hbc2f141a),
	.w7(32'hbba48f1a),
	.w8(32'hbbff7954),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0436ff),
	.w1(32'h3af11279),
	.w2(32'h3ab2eaab),
	.w3(32'h3b6f94f2),
	.w4(32'hb9c8c6e5),
	.w5(32'h3b348239),
	.w6(32'h3abfd5bf),
	.w7(32'hba8565fc),
	.w8(32'hbb68e28f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9cabd),
	.w1(32'hbb481c34),
	.w2(32'hbb033da2),
	.w3(32'h3b8ea804),
	.w4(32'h39b964b6),
	.w5(32'hb970d114),
	.w6(32'h39259a41),
	.w7(32'hba41926e),
	.w8(32'h38cff1a9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1489e4),
	.w1(32'hbb934b26),
	.w2(32'h3c2f7da2),
	.w3(32'h394f4784),
	.w4(32'hbc84d8d2),
	.w5(32'hbb83569e),
	.w6(32'hbbdf2154),
	.w7(32'h3abd8c72),
	.w8(32'hbc160c49),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule