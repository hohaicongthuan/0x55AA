module layer_10_featuremap_383(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb203ed4),
	.w1(32'hbafcbaa7),
	.w2(32'hbae67a7b),
	.w3(32'hbb83da36),
	.w4(32'hbbb017c8),
	.w5(32'hbb8635e2),
	.w6(32'hbb9a4524),
	.w7(32'hbaf35007),
	.w8(32'h3a383de0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb02443),
	.w1(32'hbae0e0c7),
	.w2(32'hba9e6861),
	.w3(32'hbb8533c7),
	.w4(32'h3bda3c08),
	.w5(32'h3afca03f),
	.w6(32'hb99537ea),
	.w7(32'h3ad42c57),
	.w8(32'hbb795d3a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc651654),
	.w1(32'h3b912484),
	.w2(32'h3bd055c1),
	.w3(32'hbc365735),
	.w4(32'h3c099b4d),
	.w5(32'h3b3f74df),
	.w6(32'hbc8651a1),
	.w7(32'h3b64586b),
	.w8(32'hbba68425),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cf231),
	.w1(32'hbb185787),
	.w2(32'h3b969d4e),
	.w3(32'h3c097c5b),
	.w4(32'h3c319935),
	.w5(32'h3c277be9),
	.w6(32'hbb435669),
	.w7(32'h3afecba3),
	.w8(32'h380185ba),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19ecb8),
	.w1(32'h3ae241be),
	.w2(32'h3aed1deb),
	.w3(32'h3a504b9f),
	.w4(32'h3ac42398),
	.w5(32'hba06057e),
	.w6(32'hbbb94bd5),
	.w7(32'h394e191b),
	.w8(32'hbb09dde3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40bed6),
	.w1(32'hb98706e3),
	.w2(32'h3a6f2181),
	.w3(32'h3b6dbc4d),
	.w4(32'hbac96032),
	.w5(32'h3be7a08e),
	.w6(32'hba993547),
	.w7(32'hba29f25a),
	.w8(32'h3b9f0df5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4eb9f),
	.w1(32'hbb258bc2),
	.w2(32'hbc0daeb9),
	.w3(32'h3ae3c658),
	.w4(32'hbb8d459f),
	.w5(32'hbc1fb97e),
	.w6(32'h3a360ef6),
	.w7(32'hbbe66cf8),
	.w8(32'hbb9727c6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4cd16),
	.w1(32'h3aaa2c10),
	.w2(32'hbbdf2c64),
	.w3(32'hbc1345e4),
	.w4(32'h3c23f9d4),
	.w5(32'h3b860b2a),
	.w6(32'hba532cc2),
	.w7(32'h3b9016f6),
	.w8(32'h3b4e8a97),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3d3b0),
	.w1(32'hbbae2bbc),
	.w2(32'hbb9013a5),
	.w3(32'h3c419e2f),
	.w4(32'hbb5c3f70),
	.w5(32'hbb24ea52),
	.w6(32'h3c43aac8),
	.w7(32'hbbad0ddd),
	.w8(32'hb8ebb87c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc759e3),
	.w1(32'h3ca02d83),
	.w2(32'h3c46ee8a),
	.w3(32'hbc4b00b4),
	.w4(32'h3bd8d85a),
	.w5(32'hbbdd9a3c),
	.w6(32'hbc30d9ca),
	.w7(32'h3b305a18),
	.w8(32'hbbd54529),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be72c66),
	.w1(32'h3c121048),
	.w2(32'h3c399f53),
	.w3(32'hbc05dd05),
	.w4(32'hbb34fd6e),
	.w5(32'hbbaa9020),
	.w6(32'hbba333a6),
	.w7(32'hbc0b359f),
	.w8(32'hbc2080cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfad183),
	.w1(32'h3ae200f4),
	.w2(32'h3b9ecadc),
	.w3(32'h3888cd42),
	.w4(32'h3ac4cc17),
	.w5(32'h3baba908),
	.w6(32'hbc0dc150),
	.w7(32'hb9c4ccf7),
	.w8(32'h3a98ddbb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0daed2),
	.w1(32'h3c4369d9),
	.w2(32'h3c00c943),
	.w3(32'h3b5a79ab),
	.w4(32'h3c8869ef),
	.w5(32'h3c8bbb14),
	.w6(32'hba918fd2),
	.w7(32'h3bacfdf0),
	.w8(32'hb769d550),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba969c0d),
	.w1(32'h3a59f176),
	.w2(32'hbb10a28a),
	.w3(32'hbbad452b),
	.w4(32'hbb145597),
	.w5(32'hbbfbebfd),
	.w6(32'hbc52d4a0),
	.w7(32'hbbe31ebf),
	.w8(32'hbbbe7cab),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ebf8e),
	.w1(32'hbb112aa4),
	.w2(32'h3b342be6),
	.w3(32'hbb1cc27c),
	.w4(32'hbc6220ad),
	.w5(32'hbbf5d806),
	.w6(32'hbafc2b88),
	.w7(32'hbc429d34),
	.w8(32'hbbf61aa3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b5bc),
	.w1(32'h395c1335),
	.w2(32'hbb119a33),
	.w3(32'h3b89055e),
	.w4(32'h39bb913f),
	.w5(32'hbb2268d9),
	.w6(32'hbbbaab50),
	.w7(32'hbb20900d),
	.w8(32'hbb5c209b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e1b56),
	.w1(32'hbb95a3cc),
	.w2(32'h3ac4d508),
	.w3(32'hbb2c66ef),
	.w4(32'hbc0fc2bc),
	.w5(32'h3a28ce8b),
	.w6(32'hbb4e987e),
	.w7(32'hbc5efef1),
	.w8(32'hbbbd91ff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf33a33),
	.w1(32'h3bddd61d),
	.w2(32'hbbcbda41),
	.w3(32'h3b3be965),
	.w4(32'h3bfecc88),
	.w5(32'hbbe5677b),
	.w6(32'hbbee07e7),
	.w7(32'hba8330fc),
	.w8(32'hbbef007f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbddb67),
	.w1(32'h3b8a8769),
	.w2(32'h3b8d0a57),
	.w3(32'hbc3ead86),
	.w4(32'h3a5817d9),
	.w5(32'h3b726fa7),
	.w6(32'hbc5c37c2),
	.w7(32'hba7a4943),
	.w8(32'h3ab7f0ab),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ab06f),
	.w1(32'hba12982e),
	.w2(32'hb9cbfc28),
	.w3(32'hb9a16232),
	.w4(32'h3a29ebcd),
	.w5(32'h393d7ed9),
	.w6(32'hbaa9db6c),
	.w7(32'h3a6532b1),
	.w8(32'hbb271278),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83380),
	.w1(32'h3c026b89),
	.w2(32'h3b593a79),
	.w3(32'h3bfe5018),
	.w4(32'h3c068ad4),
	.w5(32'h3b960b65),
	.w6(32'h3a1c9400),
	.w7(32'h3b8d76e1),
	.w8(32'hbb35cac6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9902d0c),
	.w1(32'hbaf6c209),
	.w2(32'h3a773fe3),
	.w3(32'hbbb30634),
	.w4(32'hbb077d13),
	.w5(32'h3b631cc6),
	.w6(32'hbc0c952e),
	.w7(32'h390c5b42),
	.w8(32'hb90a41ac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e418),
	.w1(32'h3bf80b7b),
	.w2(32'h3c082cd8),
	.w3(32'h3be6ca88),
	.w4(32'h3b9364c7),
	.w5(32'h39bc6d25),
	.w6(32'hb981c0c6),
	.w7(32'h39eed70f),
	.w8(32'hbb9fdfc9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101449),
	.w1(32'h3b62e81a),
	.w2(32'h3c226976),
	.w3(32'hba8ddd03),
	.w4(32'h3bc703ce),
	.w5(32'h3c612b4b),
	.w6(32'hba9734be),
	.w7(32'hbbfbb526),
	.w8(32'hbb687f47),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee4f6),
	.w1(32'hbb7cbdcf),
	.w2(32'hbb139cd1),
	.w3(32'hbb1e31ec),
	.w4(32'hbad09001),
	.w5(32'hbb4ee22a),
	.w6(32'hbc3a20fe),
	.w7(32'h3b785eef),
	.w8(32'h3b40965b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f8088),
	.w1(32'h3c1dda5a),
	.w2(32'h3be0eedc),
	.w3(32'hb9ad4efd),
	.w4(32'h3c035543),
	.w5(32'h3bf43791),
	.w6(32'h3a001eb3),
	.w7(32'h3b5e4e7b),
	.w8(32'hb9296354),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be25a95),
	.w1(32'h3b75c41e),
	.w2(32'hbb41929e),
	.w3(32'h3b128a9d),
	.w4(32'hbb308f67),
	.w5(32'hbc0ea960),
	.w6(32'h3a987b95),
	.w7(32'h3bded2e3),
	.w8(32'h3bb9d673),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf7ede),
	.w1(32'hbb815c70),
	.w2(32'hbab91e3a),
	.w3(32'hbad35ee5),
	.w4(32'h3ad08327),
	.w5(32'h3a422ed6),
	.w6(32'h3b9fe73c),
	.w7(32'hbae8a336),
	.w8(32'h3b519d00),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c31c),
	.w1(32'h3b3dca7c),
	.w2(32'h3addf539),
	.w3(32'hbb1d3af7),
	.w4(32'h3b1a0020),
	.w5(32'hbbc976a1),
	.w6(32'hbb4c8035),
	.w7(32'hba96584d),
	.w8(32'hbb2cd67b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710da4),
	.w1(32'h3b4b9b78),
	.w2(32'h399a72ba),
	.w3(32'hbb2d5a9b),
	.w4(32'h3c5a2f22),
	.w5(32'h3b9d368b),
	.w6(32'hbb37f3f6),
	.w7(32'h3c413b8d),
	.w8(32'h3c0cd815),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a386952),
	.w1(32'h394c2abe),
	.w2(32'h3b5acd40),
	.w3(32'hbbcee4bb),
	.w4(32'h3b5d7eb3),
	.w5(32'h3af3dabe),
	.w6(32'h3a966789),
	.w7(32'h3a910f30),
	.w8(32'h3b11f04b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45e5a3),
	.w1(32'h3af3dfda),
	.w2(32'h393e2bda),
	.w3(32'h3bbbc1b3),
	.w4(32'h3a99f23f),
	.w5(32'hbb27abf3),
	.w6(32'h3ad327ea),
	.w7(32'h3b931e85),
	.w8(32'h39aba8a1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4ba36),
	.w1(32'h3b9af8c2),
	.w2(32'hbb851b96),
	.w3(32'hbbc320f8),
	.w4(32'h3be92ecf),
	.w5(32'hbabc66a8),
	.w6(32'hbbb1299a),
	.w7(32'h3bec413e),
	.w8(32'h3c2078af),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3c72f),
	.w1(32'hbbc13686),
	.w2(32'hbb256bfc),
	.w3(32'hbb80484c),
	.w4(32'hbbdb6461),
	.w5(32'hba993323),
	.w6(32'h3c0476e3),
	.w7(32'hbbb1fd7a),
	.w8(32'h3b9cf05f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7926d),
	.w1(32'h3a98f403),
	.w2(32'hbc0c0d9b),
	.w3(32'hba6ed0f3),
	.w4(32'h3c30ad36),
	.w5(32'hba5fe3b4),
	.w6(32'h3b35fb49),
	.w7(32'h3c444e52),
	.w8(32'h3c428258),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5547),
	.w1(32'h3c0d15e2),
	.w2(32'h3b763cf9),
	.w3(32'h3af35842),
	.w4(32'h3c383cfd),
	.w5(32'h3b5c25da),
	.w6(32'h3c3f1aea),
	.w7(32'h3a42f7d9),
	.w8(32'hbb9a47d1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0864e6),
	.w1(32'h3c0e26e1),
	.w2(32'h3c5bd15e),
	.w3(32'hbc51444c),
	.w4(32'h3c5a72d2),
	.w5(32'h3cae71ce),
	.w6(32'hbc34c961),
	.w7(32'h3c3cf1d9),
	.w8(32'h3ca0ad9f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd8dab),
	.w1(32'hbb035849),
	.w2(32'hbb73d134),
	.w3(32'h3c1bb5fd),
	.w4(32'hbadf1dec),
	.w5(32'hbc6d9e75),
	.w6(32'h3c886fb4),
	.w7(32'h3c0691a0),
	.w8(32'hbc1d61ad),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b365c),
	.w1(32'hbb1dcbb4),
	.w2(32'h3c0ff220),
	.w3(32'hbc88af55),
	.w4(32'hbc836ec6),
	.w5(32'hbc4490d6),
	.w6(32'hbc53855e),
	.w7(32'hbc486956),
	.w8(32'hbc34f0ce),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c488284),
	.w1(32'h3c46648c),
	.w2(32'hb982776c),
	.w3(32'h3c05ecc4),
	.w4(32'h3c73d743),
	.w5(32'hbb92d3f9),
	.w6(32'h3a3cb94b),
	.w7(32'h3c6bcd09),
	.w8(32'h3a874600),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba427bd1),
	.w1(32'h3c3841a2),
	.w2(32'h3c7c4d27),
	.w3(32'hbbd32592),
	.w4(32'h3c07ebe5),
	.w5(32'h3bec14ed),
	.w6(32'hbb7dd459),
	.w7(32'h3c1ac13a),
	.w8(32'h3c3ce8dd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84199a),
	.w1(32'h3b8f4374),
	.w2(32'h3a739d42),
	.w3(32'h3c8feb00),
	.w4(32'hbbb420fb),
	.w5(32'hbc1993b1),
	.w6(32'h3c380cd2),
	.w7(32'hbb91ca94),
	.w8(32'hbbe5b47f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adab08f),
	.w1(32'h3b837e35),
	.w2(32'h3bb59a3b),
	.w3(32'h3b985243),
	.w4(32'h3c5db1bf),
	.w5(32'h3c5354cc),
	.w6(32'h3af5dd48),
	.w7(32'h3bbbd8a0),
	.w8(32'h3be6115f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4e17f),
	.w1(32'hbb14e8e7),
	.w2(32'h3b14c3f5),
	.w3(32'h3b504109),
	.w4(32'hba8f8785),
	.w5(32'h3a2eed8f),
	.w6(32'hbc13275b),
	.w7(32'hbb861989),
	.w8(32'hbb464ee9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d7547),
	.w1(32'h3b56a632),
	.w2(32'h3ad015be),
	.w3(32'hbae34995),
	.w4(32'h3b0c8db6),
	.w5(32'h3bac0407),
	.w6(32'h399a32cd),
	.w7(32'h3b1ab39c),
	.w8(32'h3b337c77),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c23f63),
	.w1(32'h3ba772cd),
	.w2(32'h3b21ca79),
	.w3(32'hba8f1b5a),
	.w4(32'h3a854e5f),
	.w5(32'h3b35a752),
	.w6(32'hbaf80e5a),
	.w7(32'h3a88f3fa),
	.w8(32'h3ab7c914),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba74688),
	.w1(32'h3ba19915),
	.w2(32'h3c1e780e),
	.w3(32'h3ab5ffe0),
	.w4(32'hbad6ccb3),
	.w5(32'h3acafcd2),
	.w6(32'h387c0276),
	.w7(32'hbc4d1540),
	.w8(32'hbc75b79d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becc43f),
	.w1(32'h3cb39d80),
	.w2(32'h3c708fd2),
	.w3(32'hbc17f066),
	.w4(32'h3c91e0d5),
	.w5(32'h3bfe3b4c),
	.w6(32'hbce4cba7),
	.w7(32'h3c866aa2),
	.w8(32'h3c32f614),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28af97),
	.w1(32'hbb2346bc),
	.w2(32'hba194906),
	.w3(32'h3bfb5fba),
	.w4(32'hbaa35f40),
	.w5(32'h3acfcd47),
	.w6(32'h3c38a6b6),
	.w7(32'hba85dcee),
	.w8(32'h3b8fc818),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0aa70),
	.w1(32'h3a834e83),
	.w2(32'h3be54b8a),
	.w3(32'hbbc764b9),
	.w4(32'hbbdf0bf8),
	.w5(32'h3ac571e1),
	.w6(32'hbb7ee93f),
	.w7(32'hbacd27c9),
	.w8(32'h3bba59dd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19923d),
	.w1(32'hbb09fc5b),
	.w2(32'h39653074),
	.w3(32'h3c2fac38),
	.w4(32'hba1a80ca),
	.w5(32'hb92950fa),
	.w6(32'h3be18593),
	.w7(32'hbb43be06),
	.w8(32'hba630200),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6247c9),
	.w1(32'h39f0fef4),
	.w2(32'hba9b8709),
	.w3(32'h3a4b7f84),
	.w4(32'hbb199a34),
	.w5(32'hbbb573da),
	.w6(32'hbb7cbdc8),
	.w7(32'hb949b11d),
	.w8(32'hbbfc56bc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb281573),
	.w1(32'h3a27eb60),
	.w2(32'h3a8f3f6b),
	.w3(32'hbb72e8c6),
	.w4(32'h3af30f6b),
	.w5(32'h3bca1a22),
	.w6(32'hbaf9518f),
	.w7(32'h3ba9a35d),
	.w8(32'h3c9fc59b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099080),
	.w1(32'h3bc9ce86),
	.w2(32'hbbf6b7e7),
	.w3(32'h3c29fed5),
	.w4(32'h3c878803),
	.w5(32'h3aab1c97),
	.w6(32'h3c52c873),
	.w7(32'h3c498ca7),
	.w8(32'h3c409ca1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc434398),
	.w1(32'h3c22b18a),
	.w2(32'h3a35bbcf),
	.w3(32'hbc2f809b),
	.w4(32'h3c507c7f),
	.w5(32'hbbe7b59a),
	.w6(32'h3a23fc6f),
	.w7(32'h3c82c828),
	.w8(32'h3ae46200),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36cf9),
	.w1(32'h3b262e07),
	.w2(32'hbafc53b3),
	.w3(32'hbb6e1437),
	.w4(32'h3c50bdd6),
	.w5(32'h3bbafe4c),
	.w6(32'h392cd761),
	.w7(32'h3be3894b),
	.w8(32'h3adf2738),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1122),
	.w1(32'hbb04fbd5),
	.w2(32'hba8c26e2),
	.w3(32'hbc68d1d8),
	.w4(32'hbb03f3ec),
	.w5(32'h3a97dd5c),
	.w6(32'hbc8fad88),
	.w7(32'hbb497f11),
	.w8(32'hba4d2d42),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29213),
	.w1(32'h3a4d1838),
	.w2(32'hba665da5),
	.w3(32'hbbd28978),
	.w4(32'h3ad8a315),
	.w5(32'h3bbf1057),
	.w6(32'hbbc791c8),
	.w7(32'hba89c779),
	.w8(32'h3ada4c81),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1267c0),
	.w1(32'hbb1623b6),
	.w2(32'h3bc2af72),
	.w3(32'hbb8a9789),
	.w4(32'hbb3c7ba9),
	.w5(32'h3c2939b4),
	.w6(32'h3706a040),
	.w7(32'hbbbd5774),
	.w8(32'h3ab40b06),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa99e57),
	.w1(32'h3bab4ea6),
	.w2(32'hbb4535cc),
	.w3(32'h3af86755),
	.w4(32'h3c0cb614),
	.w5(32'h3b4eecac),
	.w6(32'hbb3dd9ea),
	.w7(32'h3b85ebc4),
	.w8(32'h3b142ad8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e12b),
	.w1(32'hbbe5e21e),
	.w2(32'hbb9cd8d3),
	.w3(32'h3a05f6f1),
	.w4(32'hbb9885b3),
	.w5(32'hbb689f39),
	.w6(32'hbb5811f7),
	.w7(32'hbbcea7e5),
	.w8(32'hbc0a89cb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e05d1),
	.w1(32'hbb125bce),
	.w2(32'h39dfaa05),
	.w3(32'h38c0c51b),
	.w4(32'hbb6f6acb),
	.w5(32'hbba7fc1f),
	.w6(32'hbba4f7cb),
	.w7(32'hbbbd8135),
	.w8(32'hbbc4018d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901f7da),
	.w1(32'h3b42f71f),
	.w2(32'hbbeb34eb),
	.w3(32'h3ba79ef3),
	.w4(32'h3c0385fe),
	.w5(32'hbc024fcb),
	.w6(32'hbba03b64),
	.w7(32'h3a74e76a),
	.w8(32'hbc3c021a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02fe8d),
	.w1(32'hbbd30a0f),
	.w2(32'h3a9e93ac),
	.w3(32'hbc61a51a),
	.w4(32'hbbb8e847),
	.w5(32'h3ad81da3),
	.w6(32'hbc808d4d),
	.w7(32'hbb3879bc),
	.w8(32'hb99ea236),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b356174),
	.w1(32'h3bda4859),
	.w2(32'h39d3a31a),
	.w3(32'h3b8b3832),
	.w4(32'h3bd1fed0),
	.w5(32'hbb03d0c1),
	.w6(32'h39bee5c6),
	.w7(32'h3b6e63cd),
	.w8(32'hbb92d1af),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025d31),
	.w1(32'hbb872c99),
	.w2(32'hbb527fd8),
	.w3(32'hbc2129fc),
	.w4(32'hbc3b44ba),
	.w5(32'hbc11c84e),
	.w6(32'hbc15d121),
	.w7(32'hbc1450d0),
	.w8(32'hbbbbc75f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72f0b8),
	.w1(32'hbb7d6366),
	.w2(32'hbc9057f0),
	.w3(32'h3c0d46f3),
	.w4(32'hbb082033),
	.w5(32'hbce82a55),
	.w6(32'hbb01996f),
	.w7(32'hbbf073cc),
	.w8(32'hbc9a5ade),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc157bb),
	.w1(32'h3bb8f427),
	.w2(32'h3a93ebf5),
	.w3(32'hbcb0d880),
	.w4(32'hbaed6fae),
	.w5(32'hbc0ce0d0),
	.w6(32'hbc84452d),
	.w7(32'hbbd70658),
	.w8(32'hbbe02d15),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacedcb1),
	.w1(32'hbb162b4a),
	.w2(32'hbbe72c40),
	.w3(32'hbc1a63b0),
	.w4(32'hbb2e6c12),
	.w5(32'hbc46666c),
	.w6(32'hbc06de3b),
	.w7(32'hbbd04425),
	.w8(32'hbc15f2d7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc256734),
	.w1(32'h3a90dda2),
	.w2(32'h3c2adfe9),
	.w3(32'hbc25ceac),
	.w4(32'hbc09a463),
	.w5(32'h3bb1b795),
	.w6(32'hbb27a066),
	.w7(32'hb993b20e),
	.w8(32'h3c0020cd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01bca2),
	.w1(32'h3bd612d5),
	.w2(32'hbbd6a881),
	.w3(32'h3c6ac9df),
	.w4(32'h3bff711c),
	.w5(32'hbc049275),
	.w6(32'h3ae7b525),
	.w7(32'h3b3d80ee),
	.w8(32'hbb99b9e2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc589b64),
	.w1(32'hbb6161b7),
	.w2(32'h3b73027c),
	.w3(32'hbc0b0d2c),
	.w4(32'hbbc9dbbc),
	.w5(32'hb931e91f),
	.w6(32'hb9b368d4),
	.w7(32'hbac87234),
	.w8(32'h3b9c2b34),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c745),
	.w1(32'hbb368de3),
	.w2(32'h3c50a7ed),
	.w3(32'hbb9d6475),
	.w4(32'hbbe327f8),
	.w5(32'h3c03aad3),
	.w6(32'hbb991c9f),
	.w7(32'hbb387240),
	.w8(32'h3c48a213),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32249a),
	.w1(32'hba37213d),
	.w2(32'hb91bff7f),
	.w3(32'h3bec4b69),
	.w4(32'hbac3d16a),
	.w5(32'hbb523e53),
	.w6(32'h3b466ebf),
	.w7(32'h3b1b565c),
	.w8(32'h3ada1035),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87745f),
	.w1(32'h3a8bfed3),
	.w2(32'hb932b138),
	.w3(32'h3b3c7199),
	.w4(32'hbbaf81e1),
	.w5(32'h3c2ccbac),
	.w6(32'h3aa07cdb),
	.w7(32'hbb139817),
	.w8(32'hbb26c708),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75b85d),
	.w1(32'hbbdb8ec9),
	.w2(32'hbb99ebef),
	.w3(32'hbc015331),
	.w4(32'hbba7d0f3),
	.w5(32'hbb14dcd1),
	.w6(32'hbb89a2f1),
	.w7(32'hbb38c713),
	.w8(32'hbb1f5109),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b9d5),
	.w1(32'h3bb92c05),
	.w2(32'h3b787a9b),
	.w3(32'hbbb40814),
	.w4(32'h3c3ac56c),
	.w5(32'h3b433bfd),
	.w6(32'hbb942718),
	.w7(32'h3ab3aea3),
	.w8(32'h3bb609c7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080ff3),
	.w1(32'hba6db45c),
	.w2(32'h3ac2fe66),
	.w3(32'hbc03b964),
	.w4(32'h3ad35652),
	.w5(32'hbbb35ccb),
	.w6(32'hbbd21d09),
	.w7(32'h3c0a63c4),
	.w8(32'hb9b0b61a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957aa6),
	.w1(32'hbc1e50b6),
	.w2(32'hbc2266a7),
	.w3(32'hbc1c2178),
	.w4(32'hbc457a86),
	.w5(32'hbbaf258c),
	.w6(32'hbb98d467),
	.w7(32'hbc5446a1),
	.w8(32'hbbc87b1f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54a913),
	.w1(32'h3c9d1d53),
	.w2(32'hbb0de028),
	.w3(32'hbbf9d86e),
	.w4(32'h3ced8d2a),
	.w5(32'h3c81fbfe),
	.w6(32'hbc14ff40),
	.w7(32'h3b805851),
	.w8(32'h3ca658c6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf6fef),
	.w1(32'h3c445dc5),
	.w2(32'h3baa5484),
	.w3(32'hbabc93f7),
	.w4(32'h3c2b293d),
	.w5(32'hbbf562f9),
	.w6(32'h3bce1e0e),
	.w7(32'h3c5d8aeb),
	.w8(32'h3b2a8a95),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d4620),
	.w1(32'h38c29636),
	.w2(32'hbc03d2d3),
	.w3(32'h3b8994d7),
	.w4(32'hba46bce9),
	.w5(32'hbb0e2fef),
	.w6(32'h3bd46d46),
	.w7(32'hbb0e851e),
	.w8(32'hbbe4b3db),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30c29),
	.w1(32'h39cdc4c1),
	.w2(32'hbb88a01a),
	.w3(32'hbb7e1885),
	.w4(32'hb89afd94),
	.w5(32'hbb87c02d),
	.w6(32'hbad57f8f),
	.w7(32'h3b928d53),
	.w8(32'h3a8e5a51),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692d4d),
	.w1(32'hbb2c13a0),
	.w2(32'hbb1b93e5),
	.w3(32'hbb572e34),
	.w4(32'hbbd5482e),
	.w5(32'hbba5098d),
	.w6(32'hb9a303f2),
	.w7(32'hba65b729),
	.w8(32'hbb9d5203),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0669f6),
	.w1(32'h3b1aef93),
	.w2(32'hbb50f270),
	.w3(32'hbc0f306b),
	.w4(32'hbab8b5fe),
	.w5(32'hbb302b73),
	.w6(32'hbbe51328),
	.w7(32'h3b13de7f),
	.w8(32'hbbc6a7d3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc311acd),
	.w1(32'hbc1aa3d7),
	.w2(32'hbbec9d26),
	.w3(32'hbc2dbda1),
	.w4(32'hbc3db121),
	.w5(32'hbb399ecb),
	.w6(32'hbb9f2be6),
	.w7(32'hbc5a964c),
	.w8(32'hbaf43f63),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d9fad),
	.w1(32'h3bacc862),
	.w2(32'h3b90dbc4),
	.w3(32'h3be84502),
	.w4(32'h3b0c8750),
	.w5(32'h3b60d73d),
	.w6(32'h3c43fe54),
	.w7(32'h399ae782),
	.w8(32'h3bd261fa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898186),
	.w1(32'hbb48b925),
	.w2(32'h3acdebac),
	.w3(32'h3b82bd7d),
	.w4(32'hbba2462d),
	.w5(32'h3c19397f),
	.w6(32'h3c29ea57),
	.w7(32'hbc0ec90e),
	.w8(32'h3c1a7c69),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9bc71),
	.w1(32'hbacfca15),
	.w2(32'hbb95419a),
	.w3(32'hbac646cb),
	.w4(32'h3ba583c9),
	.w5(32'h3a7712fa),
	.w6(32'h3b790d91),
	.w7(32'h371ecea3),
	.w8(32'hbb172a00),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04ad4),
	.w1(32'hba419f68),
	.w2(32'hbbc466ef),
	.w3(32'hbc3f268a),
	.w4(32'hbba05609),
	.w5(32'h3b904b7e),
	.w6(32'hbc78f177),
	.w7(32'hbc433ec0),
	.w8(32'hbb442f8d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde1373),
	.w1(32'h3a829688),
	.w2(32'h3bafc22c),
	.w3(32'hbb65aeaf),
	.w4(32'h3b98ed55),
	.w5(32'h3ae776ce),
	.w6(32'hbb0417cf),
	.w7(32'h3b6f67e0),
	.w8(32'h3b5a8214),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9fe66),
	.w1(32'h3aaf6700),
	.w2(32'h3b5755dd),
	.w3(32'h3c481158),
	.w4(32'hbb1b9ac7),
	.w5(32'hbbd958d9),
	.w6(32'h3b90a9d8),
	.w7(32'h3b0282da),
	.w8(32'hbb0fbb5d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9077926),
	.w1(32'hbb32b46c),
	.w2(32'h3adf64cc),
	.w3(32'hbc11a581),
	.w4(32'hbc42dcec),
	.w5(32'hbb725242),
	.w6(32'hbb6a847e),
	.w7(32'hbbc69f74),
	.w8(32'hba616d17),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30f3e0),
	.w1(32'h3b95fe82),
	.w2(32'hb8127418),
	.w3(32'hbb3dcb10),
	.w4(32'h3b521bbc),
	.w5(32'hbbf723e5),
	.w6(32'h3aaa5063),
	.w7(32'hba2b9e45),
	.w8(32'hbb11317a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3eef2),
	.w1(32'hbba0b406),
	.w2(32'hbbf4a349),
	.w3(32'h3b20ea20),
	.w4(32'h3bdba51e),
	.w5(32'hbb2664d8),
	.w6(32'h3b1dd37a),
	.w7(32'hbbb8b723),
	.w8(32'h3a9c6748),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63e44),
	.w1(32'h3c0f641e),
	.w2(32'h3c04fdd8),
	.w3(32'hbbf07d3e),
	.w4(32'h3c00a403),
	.w5(32'hba32ecda),
	.w6(32'hbbc4c3a5),
	.w7(32'h3bf4e0ec),
	.w8(32'h3bec090e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351d6a),
	.w1(32'h3a7c94bb),
	.w2(32'hbc01972b),
	.w3(32'hba824133),
	.w4(32'hbadace20),
	.w5(32'hbbc52476),
	.w6(32'h3b3c0cdf),
	.w7(32'hbb2bfbf9),
	.w8(32'hbbe5907e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c3542),
	.w1(32'h3b72e834),
	.w2(32'h3bdeb005),
	.w3(32'h3b5fd56e),
	.w4(32'h3a8249bc),
	.w5(32'h3bc123b3),
	.w6(32'h3a7a3224),
	.w7(32'hba11f5e4),
	.w8(32'h3b122f98),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0600bb),
	.w1(32'hbc264203),
	.w2(32'hbbc9cbe5),
	.w3(32'h3b301dd7),
	.w4(32'hbbf2dae1),
	.w5(32'hba456223),
	.w6(32'h38fdf0ba),
	.w7(32'hbc71c2a6),
	.w8(32'hbafdb2da),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992c3c),
	.w1(32'h3c00b544),
	.w2(32'h3c36b9a1),
	.w3(32'hbb6f7c32),
	.w4(32'hbc2c351c),
	.w5(32'h3b1154e8),
	.w6(32'hbaf8ccd8),
	.w7(32'hbb9930ff),
	.w8(32'hbaaddb86),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22026a),
	.w1(32'hbb6a456a),
	.w2(32'hbaac0dc3),
	.w3(32'h3b74c278),
	.w4(32'h39a3827b),
	.w5(32'hbbc6b7f5),
	.w6(32'h3b9410d9),
	.w7(32'hba94c6d0),
	.w8(32'hbbc79443),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f186a),
	.w1(32'hbb2752ae),
	.w2(32'hb75b93dc),
	.w3(32'hbb98e0ff),
	.w4(32'hbc0b6fd9),
	.w5(32'h3b4796a2),
	.w6(32'h3990e622),
	.w7(32'hbbd9c60c),
	.w8(32'hba56e9d2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7468b),
	.w1(32'h3aeedc50),
	.w2(32'h3b0abfed),
	.w3(32'hbbb33499),
	.w4(32'h3b2316d8),
	.w5(32'h3b940e37),
	.w6(32'hbb52bab8),
	.w7(32'h3b25960b),
	.w8(32'h3b92bfd8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f9c2),
	.w1(32'h3af76710),
	.w2(32'h3b8dd3d0),
	.w3(32'hbb31f724),
	.w4(32'hbba461e5),
	.w5(32'h3b891f39),
	.w6(32'hbac2dbcc),
	.w7(32'hbaf2776a),
	.w8(32'h3a84e63d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254bf9),
	.w1(32'h38aab901),
	.w2(32'hbb2bb0a9),
	.w3(32'hbb88d179),
	.w4(32'h3b587861),
	.w5(32'h3c0e6125),
	.w6(32'h3b3bf437),
	.w7(32'h3b48187b),
	.w8(32'h3b83d3a5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb375),
	.w1(32'hbba8a7c8),
	.w2(32'hbb1f1b89),
	.w3(32'hbc5bb128),
	.w4(32'hbb52909c),
	.w5(32'h3a8752ee),
	.w6(32'hbc1bd3ce),
	.w7(32'hbb0ee574),
	.w8(32'hb924fe2b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf49592),
	.w1(32'hbba1bbdf),
	.w2(32'hbbfbc099),
	.w3(32'h3aebc7b1),
	.w4(32'hbbc311bb),
	.w5(32'hbbd4639e),
	.w6(32'h3b184706),
	.w7(32'hbbd63e0f),
	.w8(32'hbc1dcae7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265503),
	.w1(32'h3b5fa4d8),
	.w2(32'h3c0c86a3),
	.w3(32'hbbdb7943),
	.w4(32'hbbaffd4a),
	.w5(32'hbbf75f8a),
	.w6(32'hbb48c328),
	.w7(32'hbb350718),
	.w8(32'hbb424df7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b4a6b),
	.w1(32'h3b1bcd82),
	.w2(32'h3a7ef1ac),
	.w3(32'h3c5028c5),
	.w4(32'hbb8fbc46),
	.w5(32'h3bbde00d),
	.w6(32'hba6e561b),
	.w7(32'hbb4b2332),
	.w8(32'h3a84f19e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3034dc),
	.w1(32'h3ba18ddc),
	.w2(32'h3aef4924),
	.w3(32'h3b9eaa0f),
	.w4(32'h3c01f424),
	.w5(32'h3c3b1571),
	.w6(32'h3b544c26),
	.w7(32'h3a9abcfc),
	.w8(32'h3c2a9111),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb951),
	.w1(32'hbc055bda),
	.w2(32'h3927b8f6),
	.w3(32'hbbc1dcc3),
	.w4(32'hbbb3f5b6),
	.w5(32'h3a0bd2b5),
	.w6(32'h3aad44ab),
	.w7(32'hbb586a38),
	.w8(32'hbb777e15),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb4f1),
	.w1(32'hba6c1f5f),
	.w2(32'hbac1b8d0),
	.w3(32'h3aaec2a4),
	.w4(32'hbb07d90d),
	.w5(32'hbba93025),
	.w6(32'hbbc75f8e),
	.w7(32'h3b99c23e),
	.w8(32'hbb2a72d6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ef58e),
	.w1(32'hbbd1500d),
	.w2(32'hba836d64),
	.w3(32'h3c03e651),
	.w4(32'hbc166b44),
	.w5(32'hbbb1c422),
	.w6(32'h3c05eb4c),
	.w7(32'hbbc4f59d),
	.w8(32'hbbec4ba1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0c686),
	.w1(32'hbb39ddf0),
	.w2(32'h3bd70baa),
	.w3(32'hbad69c68),
	.w4(32'hb61fff5c),
	.w5(32'h3ba999f0),
	.w6(32'h3a9b5603),
	.w7(32'h3bf3b27c),
	.w8(32'h3bc31a59),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde8a63),
	.w1(32'h3bd3e09a),
	.w2(32'hb9e0fc01),
	.w3(32'h3bbd7ebd),
	.w4(32'hb9585927),
	.w5(32'hbc22e04f),
	.w6(32'h399791c6),
	.w7(32'h38d6f11c),
	.w8(32'hbbacbcf9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eb5ad),
	.w1(32'hba4402fb),
	.w2(32'hb780fd68),
	.w3(32'h3bf209a7),
	.w4(32'hba5f3bed),
	.w5(32'h3ba8850f),
	.w6(32'h397fb37c),
	.w7(32'hba7d2cc4),
	.w8(32'h3b0d967f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c31e),
	.w1(32'hbaacd159),
	.w2(32'h3bb1f8c8),
	.w3(32'h39bd2b07),
	.w4(32'hbb456cda),
	.w5(32'h3b771fd6),
	.w6(32'h39eabe5a),
	.w7(32'hbb6af75c),
	.w8(32'h3ad2cd9b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a75d),
	.w1(32'h3bdd9708),
	.w2(32'h3a2a9347),
	.w3(32'hbc48285e),
	.w4(32'h3bf456ae),
	.w5(32'hbc0fe599),
	.w6(32'hbb75c415),
	.w7(32'h3c328cfb),
	.w8(32'h399d9557),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd1dcd),
	.w1(32'hbb93403a),
	.w2(32'h3b2b7005),
	.w3(32'hbb8a22a8),
	.w4(32'hbbe6517a),
	.w5(32'h3b031065),
	.w6(32'hbac0a0c3),
	.w7(32'hbaee0af1),
	.w8(32'h3bd36e1f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c856),
	.w1(32'h3ba640a5),
	.w2(32'h3c0d6fee),
	.w3(32'hbc25ed09),
	.w4(32'h3b94d960),
	.w5(32'h3c48a0ea),
	.w6(32'hbbbac75b),
	.w7(32'h3b841472),
	.w8(32'h3c2f67c7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2877f),
	.w1(32'h3b184e26),
	.w2(32'hb9b5178b),
	.w3(32'h3b3e9d1b),
	.w4(32'h3abe0ce0),
	.w5(32'hb9790839),
	.w6(32'h3b01f05b),
	.w7(32'h3ab69535),
	.w8(32'h3aa46aa9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e98b1),
	.w1(32'hbb70c475),
	.w2(32'hb9abf52f),
	.w3(32'hbbe3c0db),
	.w4(32'hb9bb2233),
	.w5(32'h3b4ffe17),
	.w6(32'hbbf278b8),
	.w7(32'h3b9ee627),
	.w8(32'h3bcbe714),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1f35),
	.w1(32'h395ebeb5),
	.w2(32'hbb04095f),
	.w3(32'h3c1affd4),
	.w4(32'h3b800e82),
	.w5(32'hbb1ffa08),
	.w6(32'h3c108857),
	.w7(32'h3c082a62),
	.w8(32'h39b4f5ba),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3577e),
	.w1(32'hbc545027),
	.w2(32'hbbe449b7),
	.w3(32'hbbefc977),
	.w4(32'hbc8b90ab),
	.w5(32'hbc08fca4),
	.w6(32'hbae7a998),
	.w7(32'hbc71be59),
	.w8(32'hbc274eba),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7c34f),
	.w1(32'hbb8fe9cd),
	.w2(32'h3bb422d6),
	.w3(32'hbb3321af),
	.w4(32'hbbd010eb),
	.w5(32'h3b95a721),
	.w6(32'hbb19429c),
	.w7(32'hbb9ea4f1),
	.w8(32'h38e2db5f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5808f8),
	.w1(32'hbb5beef5),
	.w2(32'hbb972399),
	.w3(32'hbaf5272b),
	.w4(32'hb9bc2691),
	.w5(32'hba02f1d7),
	.w6(32'hba29fd6a),
	.w7(32'h3aea04ed),
	.w8(32'hbaa62a22),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75ae26),
	.w1(32'hbbce3246),
	.w2(32'hbae353db),
	.w3(32'hbc25f10a),
	.w4(32'h3c829384),
	.w5(32'h3afbf21c),
	.w6(32'hbc0d2085),
	.w7(32'h3afa9d6a),
	.w8(32'h3b6c458a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfa72f),
	.w1(32'h3a9d50d5),
	.w2(32'hbb694aa2),
	.w3(32'hbacf2285),
	.w4(32'hbbbec01e),
	.w5(32'h3bc859fc),
	.w6(32'h3b3e2c19),
	.w7(32'hbbc84f6d),
	.w8(32'hbbcfd58f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d02de8),
	.w1(32'h3c77712a),
	.w2(32'h3b4adffa),
	.w3(32'hbbde0f40),
	.w4(32'h3cddeb20),
	.w5(32'h3b99bcf0),
	.w6(32'hbc24ca67),
	.w7(32'h3c9c248a),
	.w8(32'h3b503867),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9d4e),
	.w1(32'hbb20180b),
	.w2(32'h3a83ebe2),
	.w3(32'h3c40416c),
	.w4(32'h3ae26e9e),
	.w5(32'h3af06bc2),
	.w6(32'h3c152de1),
	.w7(32'h3b3a5680),
	.w8(32'h3a9e77fd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0c4d),
	.w1(32'h3aebe812),
	.w2(32'hbb6223c5),
	.w3(32'h3c044d75),
	.w4(32'h3b29d884),
	.w5(32'h3a9c81e9),
	.w6(32'h3bbd11f2),
	.w7(32'hba174854),
	.w8(32'h3b3bca49),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2675e),
	.w1(32'h3a98e90b),
	.w2(32'h3b336ab8),
	.w3(32'hbb1017d0),
	.w4(32'h3ad4d1be),
	.w5(32'h3ad10e66),
	.w6(32'hba206484),
	.w7(32'h3bfa6572),
	.w8(32'h3bde919d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8859),
	.w1(32'hba63722c),
	.w2(32'h3a72f1aa),
	.w3(32'h3bc27257),
	.w4(32'h3621e5cc),
	.w5(32'h3b661bca),
	.w6(32'hba6fa54f),
	.w7(32'hbaf0c231),
	.w8(32'hbb7b46a4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b750),
	.w1(32'hbb804579),
	.w2(32'h3958f4f6),
	.w3(32'h3af7de56),
	.w4(32'hbc2a4bd6),
	.w5(32'hbc077869),
	.w6(32'h39eb3010),
	.w7(32'hbba9328b),
	.w8(32'hbb553bf1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaab30),
	.w1(32'h3b76a835),
	.w2(32'h3b7305e4),
	.w3(32'h3a5f9feb),
	.w4(32'h3c12ccf1),
	.w5(32'h3a9d936e),
	.w6(32'hbb632115),
	.w7(32'h3ad789f8),
	.w8(32'h3a2f595c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182fbe),
	.w1(32'h3b44a09a),
	.w2(32'hb8f5ddf8),
	.w3(32'hbbecdfa3),
	.w4(32'h3b2bafda),
	.w5(32'hbc8661ae),
	.w6(32'hba69b510),
	.w7(32'h3ac657ed),
	.w8(32'hbc2e923e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bcddb),
	.w1(32'h3b5102af),
	.w2(32'h3beb347f),
	.w3(32'h3ac23cef),
	.w4(32'h3ab394cd),
	.w5(32'h3b9ce471),
	.w6(32'h3b129c5e),
	.w7(32'h3bf3c0c0),
	.w8(32'h3c1c0ff1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4b32),
	.w1(32'hbafa9ae8),
	.w2(32'hba8db808),
	.w3(32'h3b9b8e8e),
	.w4(32'hbb9c7f42),
	.w5(32'h396cab63),
	.w6(32'h3b4d562b),
	.w7(32'hbc300b59),
	.w8(32'hbb98cbf4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7660ac),
	.w1(32'h391cdfb4),
	.w2(32'h3bdafdb7),
	.w3(32'h39c2a176),
	.w4(32'hbc0ab336),
	.w5(32'h3b933139),
	.w6(32'hbb03dba9),
	.w7(32'hbb9f9cbd),
	.w8(32'hbb893729),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66462b),
	.w1(32'hbb8083e0),
	.w2(32'hbbf98b8a),
	.w3(32'h3b44870b),
	.w4(32'hb9c4d48b),
	.w5(32'h3a0032c1),
	.w6(32'h3b12bbd6),
	.w7(32'hbb82d8a3),
	.w8(32'hbbdb4f65),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9370b9),
	.w1(32'hbb027239),
	.w2(32'hbc600ccd),
	.w3(32'hbb4c49ce),
	.w4(32'h39e80da8),
	.w5(32'hbbecf9b4),
	.w6(32'hbbbd07ff),
	.w7(32'h3b389f2c),
	.w8(32'hbc278b83),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0970),
	.w1(32'h3beb5fb6),
	.w2(32'hbb430cd6),
	.w3(32'hbbe70e99),
	.w4(32'h38f9ad4d),
	.w5(32'h369b1710),
	.w6(32'hbc10959b),
	.w7(32'h3b0124e6),
	.w8(32'hbac34c79),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7c531),
	.w1(32'h3950d802),
	.w2(32'hbbac1e19),
	.w3(32'hbb93b870),
	.w4(32'hba3e485e),
	.w5(32'hbbe4a20f),
	.w6(32'h397d4be2),
	.w7(32'h3b63b49b),
	.w8(32'hbbfae6cf),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb187910),
	.w1(32'h3b6698c8),
	.w2(32'hbc17d813),
	.w3(32'hbc068a5e),
	.w4(32'h3ba04148),
	.w5(32'hbc3f1cf3),
	.w6(32'hbb2cc8cd),
	.w7(32'h3ba5e4f6),
	.w8(32'hbc2caf6d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb86204),
	.w1(32'hbb51099d),
	.w2(32'hbbbbc3da),
	.w3(32'hbbeb2893),
	.w4(32'hbb20fef2),
	.w5(32'hbb831b1e),
	.w6(32'hbb586f0c),
	.w7(32'hbc26bb27),
	.w8(32'hbab7a384),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5e58),
	.w1(32'h3c415bf5),
	.w2(32'h3bf28fd6),
	.w3(32'hbc2319d0),
	.w4(32'h3c35d6c7),
	.w5(32'hb9a29a70),
	.w6(32'hbba0e834),
	.w7(32'h3ba4ada7),
	.w8(32'hb88e1aa7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc0e18),
	.w1(32'h3a87b3ed),
	.w2(32'hbb6b0d0a),
	.w3(32'h3ba5d265),
	.w4(32'h3b1a20c5),
	.w5(32'hbb20346d),
	.w6(32'h3c0cd5cd),
	.w7(32'h3c1831d3),
	.w8(32'hbb993221),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3111a6),
	.w1(32'hbb7dbae4),
	.w2(32'hbbdb1d24),
	.w3(32'hbbcdc7f7),
	.w4(32'hbba77da5),
	.w5(32'hbbc735e2),
	.w6(32'hbbc5261e),
	.w7(32'hbbb1d8b4),
	.w8(32'hbc11415c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc327611),
	.w1(32'hbb8cc3f4),
	.w2(32'hbbdc8f7f),
	.w3(32'hbc67a5f4),
	.w4(32'hbb93463d),
	.w5(32'hbbb940b7),
	.w6(32'hbad6ef81),
	.w7(32'hbbd8affb),
	.w8(32'hbc063647),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be7ca),
	.w1(32'h3b9c21ec),
	.w2(32'hbc3e00d0),
	.w3(32'h3a71aa2f),
	.w4(32'h3c0f5cd0),
	.w5(32'hbc5dfcfe),
	.w6(32'hbc03be51),
	.w7(32'h3c25a307),
	.w8(32'hbc7e1b53),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cef8e),
	.w1(32'h3afc1773),
	.w2(32'h3ba6c655),
	.w3(32'hbc2d6cd9),
	.w4(32'h3bb6098d),
	.w5(32'h3c2960a8),
	.w6(32'hbbcaf963),
	.w7(32'hbb2da40a),
	.w8(32'h3a7b0938),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12b068),
	.w1(32'hbc134e35),
	.w2(32'h3bf34d6e),
	.w3(32'h3ba3af57),
	.w4(32'hbc941d3b),
	.w5(32'hbb899003),
	.w6(32'hbbf30341),
	.w7(32'hbc247703),
	.w8(32'h3ba5c92e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e9822),
	.w1(32'hbaa2b1da),
	.w2(32'h3be49259),
	.w3(32'hbb1e6883),
	.w4(32'h3c0190dd),
	.w5(32'h3c10383a),
	.w6(32'h3bd37f23),
	.w7(32'h3ba264dd),
	.w8(32'h3c06a259),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04fa75),
	.w1(32'h3ad77ee4),
	.w2(32'hbb6cf976),
	.w3(32'h3be8d3a2),
	.w4(32'hbb2c1149),
	.w5(32'hbbcb508c),
	.w6(32'h3b17f604),
	.w7(32'h39c6ba31),
	.w8(32'hbbbc69be),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c54a3),
	.w1(32'hb98c109e),
	.w2(32'hbb972a0c),
	.w3(32'hba927b6a),
	.w4(32'hbb6436de),
	.w5(32'hbbf3ef85),
	.w6(32'h3aa96e38),
	.w7(32'hbb6ff90d),
	.w8(32'hbb173890),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b542247),
	.w1(32'hbbbfcff6),
	.w2(32'hbb2053fa),
	.w3(32'hb9d7b58b),
	.w4(32'hbb60dfc1),
	.w5(32'hbbde0ac4),
	.w6(32'h3ab046e6),
	.w7(32'h3af7212c),
	.w8(32'h3b4990c6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59a868),
	.w1(32'hba4dad9c),
	.w2(32'h3c57bf12),
	.w3(32'h3c7100f6),
	.w4(32'h3cb4fe79),
	.w5(32'h3c264868),
	.w6(32'h3bb42813),
	.w7(32'h3b13e456),
	.w8(32'hbba7b674),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837c54),
	.w1(32'hbc3d7df8),
	.w2(32'hbc38455b),
	.w3(32'hbbd6b1b9),
	.w4(32'hbc203eee),
	.w5(32'hbba3eacd),
	.w6(32'hbc133aa3),
	.w7(32'hbc517bf8),
	.w8(32'hbc1e419d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e8b3),
	.w1(32'h3add5ba2),
	.w2(32'h3a3a4497),
	.w3(32'hbb5c75fd),
	.w4(32'h3b969647),
	.w5(32'hbb54029b),
	.w6(32'hbb3e75bd),
	.w7(32'hbb8ace2a),
	.w8(32'hbb8901b6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9dd22),
	.w1(32'hbb9bb28b),
	.w2(32'hbb4c3cb3),
	.w3(32'hbbcccb1a),
	.w4(32'hbbeffb88),
	.w5(32'h3ac0c898),
	.w6(32'h39fdf4e7),
	.w7(32'hbbe7e754),
	.w8(32'hb99e6491),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b99c),
	.w1(32'h3a1a58cd),
	.w2(32'h3b151bf6),
	.w3(32'hbb37a56b),
	.w4(32'h3b1cd4d3),
	.w5(32'h3c07b667),
	.w6(32'hbaf8c818),
	.w7(32'hbbb48a97),
	.w8(32'h3b81f5c2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbe247),
	.w1(32'hb9bbeb79),
	.w2(32'hbb23bd5e),
	.w3(32'h3b2dd395),
	.w4(32'hbab0f9c1),
	.w5(32'hbbeb72d9),
	.w6(32'hba82d85c),
	.w7(32'hba58bd19),
	.w8(32'h39f24bb9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb475),
	.w1(32'h3c1bc704),
	.w2(32'hbb9747e2),
	.w3(32'h3adc131c),
	.w4(32'h3bb73346),
	.w5(32'hbc87864f),
	.w6(32'h3a7a7b11),
	.w7(32'h3c114dd0),
	.w8(32'hbb01ed54),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11aeb1),
	.w1(32'h3b3fd283),
	.w2(32'h3900d234),
	.w3(32'hbb1e6639),
	.w4(32'hbb6acf58),
	.w5(32'hbbaf3ca5),
	.w6(32'h3bdede38),
	.w7(32'hbb3ddced),
	.w8(32'h3b3fb2c9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2255d6),
	.w1(32'hbae0b6fa),
	.w2(32'h3c37e6fc),
	.w3(32'h3b11acdb),
	.w4(32'hbbde1d9c),
	.w5(32'h3c9f17f1),
	.w6(32'h3b79fc40),
	.w7(32'hbb076f30),
	.w8(32'h3bc0edc8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacfb38),
	.w1(32'hbbe0acdd),
	.w2(32'hbb3e3e8a),
	.w3(32'h3b5f8c85),
	.w4(32'hbc0ae28f),
	.w5(32'hba5b214c),
	.w6(32'h3ad88adf),
	.w7(32'hbc0e8b86),
	.w8(32'hbb55a5a0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf05a9b),
	.w1(32'h3c3ffd9b),
	.w2(32'hbb43a7d0),
	.w3(32'hbb855bea),
	.w4(32'h3c133643),
	.w5(32'hbc875910),
	.w6(32'hbaf34a6b),
	.w7(32'h3be29fdd),
	.w8(32'hbb8535a1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba60e06),
	.w1(32'h3a7006be),
	.w2(32'h3b1b5e0b),
	.w3(32'h3c00729c),
	.w4(32'h3afa9fcc),
	.w5(32'hbc133e20),
	.w6(32'h3c146b7c),
	.w7(32'h3aae39f7),
	.w8(32'hbba4f582),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40e885),
	.w1(32'h3bfa02ac),
	.w2(32'hbafcb9c7),
	.w3(32'h3c1e5c69),
	.w4(32'h3c1ae6f9),
	.w5(32'h3bbb74a4),
	.w6(32'h3b91f8ff),
	.w7(32'h39cede0b),
	.w8(32'h3aa42aa5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ece2),
	.w1(32'hbbb8d786),
	.w2(32'hbbdf28bd),
	.w3(32'hbb75cd10),
	.w4(32'hbbcd2cac),
	.w5(32'hbb358d16),
	.w6(32'hb815a5cb),
	.w7(32'hbb9b6e0f),
	.w8(32'hbb856ab3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362c5f),
	.w1(32'h3a03db64),
	.w2(32'h3b4ef922),
	.w3(32'hbbdad407),
	.w4(32'hba944c5b),
	.w5(32'h3c676526),
	.w6(32'hbb53e685),
	.w7(32'h3a1a27cb),
	.w8(32'h3bfd7fb4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b716d),
	.w1(32'h3c98192d),
	.w2(32'h3c7948b8),
	.w3(32'hbc27b819),
	.w4(32'h3ca5e429),
	.w5(32'hbbf60816),
	.w6(32'hbc02d15e),
	.w7(32'h3cac64c7),
	.w8(32'h3b6e55a4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77a183),
	.w1(32'hb7902ffd),
	.w2(32'h3af7b30f),
	.w3(32'h3c3744f5),
	.w4(32'h3b1c4131),
	.w5(32'h3ab3291a),
	.w6(32'h3c209ec9),
	.w7(32'h3bad1746),
	.w8(32'h3b041915),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2533d8),
	.w1(32'h3b1f1e40),
	.w2(32'hbbd62fb7),
	.w3(32'h3b38151d),
	.w4(32'h3ae7109a),
	.w5(32'hbc49c34d),
	.w6(32'hba5889c2),
	.w7(32'h3b071bb7),
	.w8(32'hbb9aa01d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802641),
	.w1(32'h3bc2e1ab),
	.w2(32'h3b3e7e38),
	.w3(32'hb95ca65a),
	.w4(32'h38040bc0),
	.w5(32'h3b7d6d72),
	.w6(32'hbb94213b),
	.w7(32'hbbfc6f05),
	.w8(32'hbb519e5f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec66a),
	.w1(32'h3b8b843f),
	.w2(32'hbb6298a5),
	.w3(32'hb92fc4c2),
	.w4(32'h38caeb51),
	.w5(32'hbbeae760),
	.w6(32'hbbdedd59),
	.w7(32'h3b90985d),
	.w8(32'h3a338759),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9795f),
	.w1(32'hbb42f78b),
	.w2(32'hbbc6a384),
	.w3(32'h3c038e88),
	.w4(32'hbb89ad5e),
	.w5(32'hbc534c97),
	.w6(32'h3b3382ea),
	.w7(32'hbc124961),
	.w8(32'hbbfaf3e8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc418),
	.w1(32'hbb1fef3d),
	.w2(32'hbb02cbfe),
	.w3(32'hbc2a35b5),
	.w4(32'hbbeb7b5a),
	.w5(32'hbbff411f),
	.w6(32'hbc1bf04b),
	.w7(32'hbc14647c),
	.w8(32'hbb3cca76),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991e995),
	.w1(32'h3c1edbf0),
	.w2(32'hbb46de83),
	.w3(32'hbbc86ee3),
	.w4(32'h3c81087f),
	.w5(32'hbb9a2d18),
	.w6(32'hbb2ff33c),
	.w7(32'h3c3450a4),
	.w8(32'hbae0c148),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafed9c2),
	.w1(32'h3b378105),
	.w2(32'h3c39fa0e),
	.w3(32'hb95c1115),
	.w4(32'hbb243b60),
	.w5(32'h3c211181),
	.w6(32'hbb85e3a1),
	.w7(32'h3bcf1389),
	.w8(32'h3cb5eaa6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18de6a),
	.w1(32'hb8b17031),
	.w2(32'hbad224df),
	.w3(32'h3b1b75a8),
	.w4(32'hbb6e1cd8),
	.w5(32'hbc0c7dbf),
	.w6(32'h3c18d544),
	.w7(32'hbbda5b66),
	.w8(32'h3a09e1f6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eba60),
	.w1(32'hba80f023),
	.w2(32'hb995fb30),
	.w3(32'hbb10f59a),
	.w4(32'hbb7c6b86),
	.w5(32'hbbebd751),
	.w6(32'h3b2f49dc),
	.w7(32'hbabdefe1),
	.w8(32'h3a85be3c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080c31),
	.w1(32'hbba31c72),
	.w2(32'h3ae72439),
	.w3(32'hb9d72997),
	.w4(32'hbbe22e20),
	.w5(32'hba6061a4),
	.w6(32'h3b1fae5f),
	.w7(32'hbb9b8cb8),
	.w8(32'h3b540eba),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca9d7),
	.w1(32'h3ba038e0),
	.w2(32'h3bdde7ca),
	.w3(32'hbb939cd1),
	.w4(32'hbb157248),
	.w5(32'h3b6c0984),
	.w6(32'hbb19361b),
	.w7(32'h3b0d65fa),
	.w8(32'h3b05a91f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b0b8),
	.w1(32'hbb6f5d88),
	.w2(32'hbb3ce037),
	.w3(32'hbaf1b2ea),
	.w4(32'hbbf25819),
	.w5(32'h3b5c2ab4),
	.w6(32'h3b17f22c),
	.w7(32'hbb861b5a),
	.w8(32'hbb52e7df),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1af5bc),
	.w1(32'hbbc69715),
	.w2(32'hbabb1e1a),
	.w3(32'hba67635a),
	.w4(32'hbc407621),
	.w5(32'hba6d005a),
	.w6(32'h39bf177b),
	.w7(32'hbbaa4437),
	.w8(32'hbb8b192c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca6ca2),
	.w1(32'h39436f0f),
	.w2(32'h3bf8e885),
	.w3(32'h3a4929f7),
	.w4(32'hbb7742c2),
	.w5(32'h3c804303),
	.w6(32'h3ad4456e),
	.w7(32'h3ad708aa),
	.w8(32'h3c0d7d32),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5432),
	.w1(32'h3c4df7a0),
	.w2(32'h3ba03219),
	.w3(32'h3ac745c2),
	.w4(32'h3c37e43d),
	.w5(32'h3b9e0476),
	.w6(32'hbb13835f),
	.w7(32'h3b29c64f),
	.w8(32'hbb2e4aee),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3779c),
	.w1(32'hbc0746de),
	.w2(32'h3c05c081),
	.w3(32'h3c5d1077),
	.w4(32'hbb955e57),
	.w5(32'hbaf51c2c),
	.w6(32'h3a534eda),
	.w7(32'hbb8e59ab),
	.w8(32'h36be76ba),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ae159),
	.w1(32'hbbe77832),
	.w2(32'h3ba7f4db),
	.w3(32'h3b7e9fcf),
	.w4(32'hbb30ba13),
	.w5(32'h3c15e22b),
	.w6(32'hbb914565),
	.w7(32'hbb8fc90a),
	.w8(32'h3b86e61a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93de5),
	.w1(32'h3a164baa),
	.w2(32'hba93926b),
	.w3(32'h3a2175e0),
	.w4(32'hba0f6268),
	.w5(32'hbae0e6a4),
	.w6(32'hba6559f3),
	.w7(32'hbb3cf136),
	.w8(32'hba6f70bc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ef31),
	.w1(32'hbb8e7f3f),
	.w2(32'hbb9f31a0),
	.w3(32'hbbbe1722),
	.w4(32'hbb91a33c),
	.w5(32'h39a3debb),
	.w6(32'hbb076383),
	.w7(32'hbb5aef3f),
	.w8(32'hbbd51ea8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd4a3),
	.w1(32'h3c553003),
	.w2(32'h3b1c36ea),
	.w3(32'hbb3206b4),
	.w4(32'h3c037f9c),
	.w5(32'hbc1a5f80),
	.w6(32'hbba0d9b5),
	.w7(32'h3c455161),
	.w8(32'hbb41b13a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97611a),
	.w1(32'h3b879cd3),
	.w2(32'h3c51e639),
	.w3(32'hbb1c9bd3),
	.w4(32'hbb2185a2),
	.w5(32'h3bf5391f),
	.w6(32'h3ae88e60),
	.w7(32'hbbb28898),
	.w8(32'h3bc3c007),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b182a08),
	.w1(32'hbb87c155),
	.w2(32'hbbd42b48),
	.w3(32'hbbf26ed2),
	.w4(32'h3bb6c260),
	.w5(32'hbbc70b76),
	.w6(32'hbb20e61f),
	.w7(32'h3aef1974),
	.w8(32'hbb3aa88b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389858fc),
	.w1(32'hbc03812d),
	.w2(32'h3aa3070c),
	.w3(32'hb9a81f53),
	.w4(32'hbc54930d),
	.w5(32'hbbff8345),
	.w6(32'h39e78e34),
	.w7(32'hbbf1b76d),
	.w8(32'h3b9ee65e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52038c),
	.w1(32'h3c67b1ca),
	.w2(32'h3b594916),
	.w3(32'hbc448d44),
	.w4(32'h3cbeccd4),
	.w5(32'hba3343a3),
	.w6(32'hbbd37310),
	.w7(32'h3ca496e0),
	.w8(32'h38c59b3b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c117047),
	.w1(32'h3a154f3a),
	.w2(32'hbb9befa7),
	.w3(32'h3c0ae96b),
	.w4(32'h3b458b00),
	.w5(32'hbba0af5d),
	.w6(32'hbab7aacb),
	.w7(32'h3ae6f207),
	.w8(32'hba15d7fc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad1736),
	.w1(32'hba64001e),
	.w2(32'hba4a535f),
	.w3(32'hbb8ea67e),
	.w4(32'hba48089a),
	.w5(32'h3a27011e),
	.w6(32'hba00d0ae),
	.w7(32'hb522373e),
	.w8(32'h3a6565ee),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5f171),
	.w1(32'h3b1bc6f6),
	.w2(32'h3b666b4e),
	.w3(32'hbb7fb891),
	.w4(32'h3b4eb694),
	.w5(32'h3aafc811),
	.w6(32'hbb3dd637),
	.w7(32'hba133813),
	.w8(32'h3a6cb35c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4c740),
	.w1(32'h3b39d9d3),
	.w2(32'hba491e55),
	.w3(32'h3b71311b),
	.w4(32'h3ba3dc4f),
	.w5(32'h3ba1bdac),
	.w6(32'h3a7d5928),
	.w7(32'h3b6c89ce),
	.w8(32'h3b6e5837),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d8998),
	.w1(32'h3be0fa78),
	.w2(32'h3bafba9a),
	.w3(32'h3a85297e),
	.w4(32'h3bca1818),
	.w5(32'h3b968cb2),
	.w6(32'h3af9418b),
	.w7(32'h3bbe3b07),
	.w8(32'h3b87b695),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84f8b7),
	.w1(32'hbbd5d5fb),
	.w2(32'hba9fc4fb),
	.w3(32'hbb1db1dc),
	.w4(32'hbbaaec1c),
	.w5(32'hbb02bc0e),
	.w6(32'h3aa5bf54),
	.w7(32'hbbc0f680),
	.w8(32'h39b9bfde),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2195da),
	.w1(32'hbbc17c1c),
	.w2(32'hbb947540),
	.w3(32'hbb511c93),
	.w4(32'hbbdbc5fc),
	.w5(32'hbba42627),
	.w6(32'h3a31bc87),
	.w7(32'hbb992ce0),
	.w8(32'hba177b48),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09278),
	.w1(32'hbbbba7a2),
	.w2(32'hbb8a563f),
	.w3(32'hbbbce325),
	.w4(32'hbb69260e),
	.w5(32'hbb85ad63),
	.w6(32'h3b81433e),
	.w7(32'h38c7a453),
	.w8(32'hbb538d25),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ee8b),
	.w1(32'h395612c8),
	.w2(32'h38bfd49a),
	.w3(32'h3b6b2556),
	.w4(32'hbaa61eb8),
	.w5(32'hbadd1658),
	.w6(32'h3b31bfa9),
	.w7(32'h3b0c393a),
	.w8(32'hbab3f6d8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda6923),
	.w1(32'h39e6de9a),
	.w2(32'hba773fb0),
	.w3(32'hbb608d9b),
	.w4(32'hbb141d6c),
	.w5(32'hbbd54298),
	.w6(32'hba91238a),
	.w7(32'h3b2d93ac),
	.w8(32'hbaf6aebc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f5867),
	.w1(32'h3b8d86a0),
	.w2(32'hbab0a4d4),
	.w3(32'h3a028464),
	.w4(32'hb8e3110a),
	.w5(32'hbb36c3b8),
	.w6(32'hb99fe406),
	.w7(32'hbb4be9af),
	.w8(32'hbb907589),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e299b),
	.w1(32'h3b871228),
	.w2(32'h3bbb4084),
	.w3(32'hbbace16a),
	.w4(32'h3c109583),
	.w5(32'h3b34d0d7),
	.w6(32'hbc2165c8),
	.w7(32'h3c1a1c65),
	.w8(32'h3ba317df),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40e0ca),
	.w1(32'hbb770c63),
	.w2(32'hbb0b6798),
	.w3(32'hba84060c),
	.w4(32'hbb6d2710),
	.w5(32'hbb0d497a),
	.w6(32'h3ab2b314),
	.w7(32'hbbbe7137),
	.w8(32'hbb5c2893),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95522a),
	.w1(32'h397e41ef),
	.w2(32'h3af6849a),
	.w3(32'hbb5f32ff),
	.w4(32'h3a08ab5b),
	.w5(32'hba2ee869),
	.w6(32'hbb4bcc21),
	.w7(32'h3b02048a),
	.w8(32'h3b4cb6dc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb4b29),
	.w1(32'h3b680c25),
	.w2(32'h3baf8143),
	.w3(32'h3a90262a),
	.w4(32'hbb94b21a),
	.w5(32'h3abcb3c3),
	.w6(32'h3b036dcf),
	.w7(32'hbc15b2ea),
	.w8(32'hbaf4caa7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1a231),
	.w1(32'h3c1886d9),
	.w2(32'h3b849872),
	.w3(32'hbadef175),
	.w4(32'h3b475715),
	.w5(32'h3b730018),
	.w6(32'hbb8a64f1),
	.w7(32'h3a80bfe3),
	.w8(32'hba9f6ce7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d13c6),
	.w1(32'h3a6f7814),
	.w2(32'hbb02ced4),
	.w3(32'hbb8b0da6),
	.w4(32'hbad98735),
	.w5(32'h3a530015),
	.w6(32'hbb47ddf7),
	.w7(32'h3a1c7891),
	.w8(32'hbba3b467),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f790c),
	.w1(32'h3a09cf40),
	.w2(32'h3b1f203d),
	.w3(32'hb8632419),
	.w4(32'h3a67de94),
	.w5(32'h3b57e25e),
	.w6(32'hbbca717d),
	.w7(32'h3a96bbd1),
	.w8(32'h3a28e3b8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0f669),
	.w1(32'hbb65f0da),
	.w2(32'hbb913732),
	.w3(32'hbc026725),
	.w4(32'hbc0c1473),
	.w5(32'hbbc784a6),
	.w6(32'hbbb58288),
	.w7(32'hbb0df4a5),
	.w8(32'hbb8faef8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a198290),
	.w1(32'hbb6342ee),
	.w2(32'hbb3d04cd),
	.w3(32'hbbd284df),
	.w4(32'hbb82aa80),
	.w5(32'hbbb92d21),
	.w6(32'hbbec82cd),
	.w7(32'hbbe06df9),
	.w8(32'hbb85ff8a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc62e88),
	.w1(32'h3ab2cec9),
	.w2(32'h3a7ef62b),
	.w3(32'hbae22123),
	.w4(32'hb9a83719),
	.w5(32'h3bde19df),
	.w6(32'hbaa5e9c1),
	.w7(32'hbb8bbea5),
	.w8(32'hbb30f070),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02e8ee),
	.w1(32'h3a3ab471),
	.w2(32'h3b36e3ea),
	.w3(32'hbbe19fef),
	.w4(32'h3b430079),
	.w5(32'h3c14848e),
	.w6(32'hbc0aec0b),
	.w7(32'h39cb7f4d),
	.w8(32'h3b1c0dce),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a4f33),
	.w1(32'h3b3aae4e),
	.w2(32'h3ad8299f),
	.w3(32'h3a9a70ea),
	.w4(32'h3a2d1ad5),
	.w5(32'h3b8bc2e0),
	.w6(32'h39b86f58),
	.w7(32'hbafcca5a),
	.w8(32'h3a4d0184),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71011c),
	.w1(32'h3ae16d8c),
	.w2(32'hbb048cd6),
	.w3(32'h3b391f83),
	.w4(32'hb9220fc0),
	.w5(32'hbc16bfa3),
	.w6(32'h38f64e0c),
	.w7(32'hb9677c4b),
	.w8(32'hbb35e3a4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1059e1),
	.w1(32'h3c413e9b),
	.w2(32'h3c06808c),
	.w3(32'hba0a71a9),
	.w4(32'h3c272bea),
	.w5(32'h3b428188),
	.w6(32'hb98b72a2),
	.w7(32'h3c0a7afa),
	.w8(32'h3ba1a0ed),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25dafe),
	.w1(32'h3ba9b31e),
	.w2(32'h3b93489e),
	.w3(32'h3ad9f28b),
	.w4(32'h3a49280c),
	.w5(32'h3ae30309),
	.w6(32'h3afe9b67),
	.w7(32'h3b14f5ae),
	.w8(32'h39ec6867),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22bbbe),
	.w1(32'hbbc472f1),
	.w2(32'hba5e8973),
	.w3(32'hbac85551),
	.w4(32'hbbcbb7e8),
	.w5(32'h3b1548e0),
	.w6(32'hbb65af8f),
	.w7(32'hbb08bcfe),
	.w8(32'h3760adb5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592771),
	.w1(32'h3b235951),
	.w2(32'hbb0341ce),
	.w3(32'h3b9b730a),
	.w4(32'hba7ede44),
	.w5(32'hbadb3fc9),
	.w6(32'h3a956472),
	.w7(32'hb915042e),
	.w8(32'hbb597d4f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97cde),
	.w1(32'h3c2bad81),
	.w2(32'h3bf119e5),
	.w3(32'hbab59640),
	.w4(32'h3c0ae6ee),
	.w5(32'h3be7f70a),
	.w6(32'h3a7ddd6c),
	.w7(32'h3b9b9c92),
	.w8(32'h3b5af358),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad59dc),
	.w1(32'h3b4c194e),
	.w2(32'hbb943c4f),
	.w3(32'hbba062b1),
	.w4(32'h3a4dff29),
	.w5(32'h3ae0dc3f),
	.w6(32'hbad83b13),
	.w7(32'hbad3ca55),
	.w8(32'hba687e41),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba036b7),
	.w1(32'h3bdc0867),
	.w2(32'h3aa4dd4c),
	.w3(32'h3b6fbe26),
	.w4(32'h3a5159bb),
	.w5(32'h3ad33e5b),
	.w6(32'h3bb58641),
	.w7(32'hbad06fc6),
	.w8(32'h3b1c3019),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45e693),
	.w1(32'h3c176c9d),
	.w2(32'h3bc39720),
	.w3(32'hbb42bd88),
	.w4(32'h3bd90aec),
	.w5(32'h3b75d193),
	.w6(32'hbb000acf),
	.w7(32'h3ba17c3d),
	.w8(32'h3bb1cfa0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaae2f6),
	.w1(32'h3b8e47aa),
	.w2(32'hb9db4b41),
	.w3(32'h3a73aaf8),
	.w4(32'h3b3bf073),
	.w5(32'h3a25ccdc),
	.w6(32'h3bab13e7),
	.w7(32'h3ac6e3c7),
	.w8(32'hb9c4e6e8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52cff1),
	.w1(32'h3b893a84),
	.w2(32'h3c83b63e),
	.w3(32'hbab327ba),
	.w4(32'h3b0388a0),
	.w5(32'h3c6ccb55),
	.w6(32'hbb7ca209),
	.w7(32'h3ac63e63),
	.w8(32'h3bdfa65d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58c45a),
	.w1(32'h3bacf1f5),
	.w2(32'hbb7cbca9),
	.w3(32'h3c217e28),
	.w4(32'h3bd1d1a9),
	.w5(32'h3a4e635c),
	.w6(32'h3983c140),
	.w7(32'h3ba0a3e7),
	.w8(32'hbb2cf262),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25f614),
	.w1(32'hbb5e23b7),
	.w2(32'hbbae4ab3),
	.w3(32'h3c270882),
	.w4(32'hbb9a99ae),
	.w5(32'hbc0420ef),
	.w6(32'h3c5acd36),
	.w7(32'hbb68b709),
	.w8(32'hbac7bd62),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3b6e2),
	.w1(32'h3b63c327),
	.w2(32'hbb9b5046),
	.w3(32'hbb5606b0),
	.w4(32'h3abcfe68),
	.w5(32'hbb8724b2),
	.w6(32'hbc089967),
	.w7(32'hbac5c1a4),
	.w8(32'hbb3c7c1a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74a3ec),
	.w1(32'h3aa30393),
	.w2(32'h3bb3489d),
	.w3(32'h3a17ee8e),
	.w4(32'h3bbfdead),
	.w5(32'h3c1a60e9),
	.w6(32'hba3a8849),
	.w7(32'h3bac0d8a),
	.w8(32'h3bb428dc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab637ee),
	.w1(32'hbb1cf682),
	.w2(32'hbab59271),
	.w3(32'hbb2bc4ed),
	.w4(32'hbb5dade6),
	.w5(32'h39a33f71),
	.w6(32'hbb562f89),
	.w7(32'hbb75360a),
	.w8(32'hba92a44b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a304a37),
	.w1(32'hbafc1115),
	.w2(32'h3aa70fcf),
	.w3(32'h3a34618d),
	.w4(32'h3a21beac),
	.w5(32'hba85a6fa),
	.w6(32'h3af1a6d8),
	.w7(32'hbb80f7a9),
	.w8(32'hbb144575),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76c80a),
	.w1(32'h3b412f14),
	.w2(32'hb9ae9f7d),
	.w3(32'hba90a6af),
	.w4(32'hbb79b956),
	.w5(32'hbbaaf1d8),
	.w6(32'hb9276fc7),
	.w7(32'hbc1f6e5c),
	.w8(32'hbbc982d4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907364e),
	.w1(32'hba0f7bfc),
	.w2(32'h3b603f4b),
	.w3(32'h3b76e6fe),
	.w4(32'hba6a9604),
	.w5(32'h3c115186),
	.w6(32'h3adae081),
	.w7(32'hbab83ca9),
	.w8(32'h39170a9a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03095),
	.w1(32'hbaceef04),
	.w2(32'hbbee86f4),
	.w3(32'h3c1a266a),
	.w4(32'h3b093f2b),
	.w5(32'hbba34c22),
	.w6(32'h3a62b7ba),
	.w7(32'hbb1347b9),
	.w8(32'hbbd0c831),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510954),
	.w1(32'h3b6d469a),
	.w2(32'hbaf20973),
	.w3(32'h3b197925),
	.w4(32'h3baefec7),
	.w5(32'hb848eb0b),
	.w6(32'hbb861967),
	.w7(32'hb9965842),
	.w8(32'hbb93fb92),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f7cb7),
	.w1(32'hbc3661fe),
	.w2(32'h3bb0b1c4),
	.w3(32'hbade1c7f),
	.w4(32'hbc33838e),
	.w5(32'h3b335f42),
	.w6(32'hbb921066),
	.w7(32'hbc7a6a19),
	.w8(32'hbadf947d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846d5a),
	.w1(32'hbb9cfa62),
	.w2(32'hbb978df1),
	.w3(32'h3b9ba590),
	.w4(32'hbb84d60a),
	.w5(32'hbc0e0042),
	.w6(32'h3b96134a),
	.w7(32'hbba232ba),
	.w8(32'hbbd21a84),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bd177),
	.w1(32'hba841fd0),
	.w2(32'hbb66286d),
	.w3(32'hbb8242f2),
	.w4(32'h3a971837),
	.w5(32'hbb3348ef),
	.w6(32'hbb4fbf5c),
	.w7(32'h3aec9887),
	.w8(32'hba83657e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0ed57),
	.w1(32'h3ac40e2f),
	.w2(32'h39e27139),
	.w3(32'hbb1fcfcf),
	.w4(32'h3bb60fc9),
	.w5(32'h3b271193),
	.w6(32'hbb450475),
	.w7(32'h3a45956b),
	.w8(32'h3a823258),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1956e),
	.w1(32'h3b78bee7),
	.w2(32'hbb9610a6),
	.w3(32'hbb92cb43),
	.w4(32'hba0d8d21),
	.w5(32'hbb561307),
	.w6(32'hbb8e5b85),
	.w7(32'hbbcc4117),
	.w8(32'hbc01ca56),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4ce6),
	.w1(32'h3ab8c21b),
	.w2(32'h3a60d9bf),
	.w3(32'h3af40db7),
	.w4(32'hba0386e4),
	.w5(32'hbaca27ad),
	.w6(32'hbb3392c0),
	.w7(32'hba4e24c6),
	.w8(32'hbba26d47),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8d81f),
	.w1(32'h3c39edcc),
	.w2(32'h3c8bbd7a),
	.w3(32'hba372860),
	.w4(32'h3bb0a0de),
	.w5(32'h3c921a5c),
	.w6(32'h3a30387b),
	.w7(32'h3bf5e889),
	.w8(32'h3c906870),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70b14c),
	.w1(32'hbb1edf1a),
	.w2(32'hb9567ba7),
	.w3(32'h3c70d563),
	.w4(32'hbad3b561),
	.w5(32'hbb1d2216),
	.w6(32'h3c7c828a),
	.w7(32'hb98376f0),
	.w8(32'hbadf795e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad6f1),
	.w1(32'hbc09dd2d),
	.w2(32'h3a553cab),
	.w3(32'h3b856794),
	.w4(32'hbbf49ce5),
	.w5(32'h39bb7b03),
	.w6(32'h3b40b77e),
	.w7(32'hbb641188),
	.w8(32'h39432a44),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35e308),
	.w1(32'hbbb21ef5),
	.w2(32'hbb659148),
	.w3(32'h3b11e9c8),
	.w4(32'hbbb2ea1e),
	.w5(32'hbb62e534),
	.w6(32'h3b18f6e2),
	.w7(32'hbb77d6ab),
	.w8(32'hbbcc5057),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4fa51),
	.w1(32'hbbbd4775),
	.w2(32'hbbe702d5),
	.w3(32'hbbe97165),
	.w4(32'hbb077c43),
	.w5(32'hbc15c275),
	.w6(32'hbc5b4d51),
	.w7(32'hbb4c57ef),
	.w8(32'hbbcbbb93),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099360),
	.w1(32'h3a896767),
	.w2(32'h3a820e2b),
	.w3(32'hbbc3dfd1),
	.w4(32'hba8b384c),
	.w5(32'hbb8407e5),
	.w6(32'hbb9d6908),
	.w7(32'hbbfa298d),
	.w8(32'hbbd106a8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef586c),
	.w1(32'hbaeadd4e),
	.w2(32'hbbc1662d),
	.w3(32'hbb3c7c6e),
	.w4(32'hbaebdf6b),
	.w5(32'hbba2928c),
	.w6(32'hbc2b1d0a),
	.w7(32'hbbb1b8df),
	.w8(32'hbb8640f9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d55f4),
	.w1(32'h3bf6a9ab),
	.w2(32'h3b901a52),
	.w3(32'h3baf8af6),
	.w4(32'h3b598270),
	.w5(32'h3af5dc04),
	.w6(32'h3a5ead52),
	.w7(32'h398c51ae),
	.w8(32'h3a816e84),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc33fe4),
	.w1(32'hba7a1b71),
	.w2(32'h3aeb167c),
	.w3(32'h3bf8963e),
	.w4(32'hbb62291d),
	.w5(32'h3ac947c9),
	.w6(32'h3bb2bf8a),
	.w7(32'hbb8e92f3),
	.w8(32'hbb96f27a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule