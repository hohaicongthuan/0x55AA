module layer_8_featuremap_110(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4814d),
	.w1(32'h3b5c97f9),
	.w2(32'hbc0e0660),
	.w3(32'h3b30b16e),
	.w4(32'hbc2a9e66),
	.w5(32'hbb652a99),
	.w6(32'hbaea72a2),
	.w7(32'hbbf951c6),
	.w8(32'hbb8166b5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1b082),
	.w1(32'h38286be9),
	.w2(32'hbb996937),
	.w3(32'hbc04a171),
	.w4(32'hba360012),
	.w5(32'h3ca9e3d8),
	.w6(32'hba67f07d),
	.w7(32'hbb36457d),
	.w8(32'h3c8124c0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895a56),
	.w1(32'h3a32f19f),
	.w2(32'h3ccbd64b),
	.w3(32'h3c1d20e4),
	.w4(32'h3c36d37c),
	.w5(32'h3b650242),
	.w6(32'h3bc6cf2a),
	.w7(32'h3c867cca),
	.w8(32'hba39caee),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f580),
	.w1(32'hbbed3bda),
	.w2(32'hbcc64abc),
	.w3(32'h3babe8d7),
	.w4(32'h3a85eac2),
	.w5(32'hbb0c356a),
	.w6(32'hbc62ac13),
	.w7(32'hbc55054f),
	.w8(32'hbc8c1950),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06de86),
	.w1(32'h3b7e882d),
	.w2(32'hbaacaa5e),
	.w3(32'hba8870c7),
	.w4(32'hbb02e4dc),
	.w5(32'hba8ade1d),
	.w6(32'hbc0428c0),
	.w7(32'hbb5e8d0a),
	.w8(32'h3bc16dd2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833ea8),
	.w1(32'hbb39b4f1),
	.w2(32'hbc99e6d5),
	.w3(32'hbc361533),
	.w4(32'hb97899af),
	.w5(32'h3a551b1a),
	.w6(32'hbba39466),
	.w7(32'h3c228cce),
	.w8(32'h3bf3c782),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72600d),
	.w1(32'h382ff412),
	.w2(32'hbc1f171d),
	.w3(32'hbb2a1a49),
	.w4(32'h3bc32f46),
	.w5(32'hbb8e36af),
	.w6(32'h3c499bc2),
	.w7(32'hbbfe23eb),
	.w8(32'hbb589c98),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ba49f),
	.w1(32'h3bd4188f),
	.w2(32'h3c88390b),
	.w3(32'hbc1f3143),
	.w4(32'h3c8713d3),
	.w5(32'h3ca1775f),
	.w6(32'hbc0d46d1),
	.w7(32'h3d0ba900),
	.w8(32'h3d40173f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a39ca),
	.w1(32'h3b13cb33),
	.w2(32'h3bcc2c97),
	.w3(32'hbb96d2fc),
	.w4(32'hbbe39fc3),
	.w5(32'h3bd4e9db),
	.w6(32'h3b0ac264),
	.w7(32'hbc31fe16),
	.w8(32'h3bb4d04a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13b54),
	.w1(32'h3b2b8c47),
	.w2(32'h3c7f8ae1),
	.w3(32'hbc6a62d7),
	.w4(32'h3b941bb9),
	.w5(32'h398b628d),
	.w6(32'hbc384282),
	.w7(32'h3a576c94),
	.w8(32'hbcfc1c00),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00923d),
	.w1(32'h3bb5551f),
	.w2(32'h3cb7cc62),
	.w3(32'h3beb51db),
	.w4(32'h3b02da28),
	.w5(32'h3a0404a3),
	.w6(32'h3b7fbd9d),
	.w7(32'h3c1b4d9c),
	.w8(32'h3c73fbbc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad7716),
	.w1(32'hbc790bdc),
	.w2(32'hbbbfc5ac),
	.w3(32'h3a8d3948),
	.w4(32'hba60ce82),
	.w5(32'hbb1e274c),
	.w6(32'hbc8d23de),
	.w7(32'hba20c1ee),
	.w8(32'hbba437ad),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e2c8),
	.w1(32'hbc04dc2b),
	.w2(32'h3b6b2657),
	.w3(32'hbc83e403),
	.w4(32'h3af4c947),
	.w5(32'h3b477a58),
	.w6(32'hbc95fd7a),
	.w7(32'h3b63c7a7),
	.w8(32'h3c50dd03),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fbec2),
	.w1(32'hbac68ecd),
	.w2(32'hbb37de77),
	.w3(32'hbb2d10ce),
	.w4(32'hbb1a9a10),
	.w5(32'hbbac6ebd),
	.w6(32'hb9a4f8ec),
	.w7(32'hbb8b714e),
	.w8(32'h3a59e768),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b973229),
	.w1(32'h39bbee5d),
	.w2(32'hbaa65523),
	.w3(32'h3681f5b6),
	.w4(32'hbb4872a9),
	.w5(32'hbb71724e),
	.w6(32'h3b00a047),
	.w7(32'hbafa2080),
	.w8(32'hbb051293),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6c65),
	.w1(32'h3b12e03a),
	.w2(32'hb9c70aa3),
	.w3(32'h391d444a),
	.w4(32'h3af0fc27),
	.w5(32'h3ba2de30),
	.w6(32'h3aa509e7),
	.w7(32'h3bbe71a3),
	.w8(32'hbc67c772),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272150),
	.w1(32'hbb0e31a3),
	.w2(32'h3afc2205),
	.w3(32'hbc00117d),
	.w4(32'h3b43322f),
	.w5(32'h3c897af3),
	.w6(32'h3c5d9d88),
	.w7(32'h3a8d8d6d),
	.w8(32'h3d317d8f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b3457),
	.w1(32'h3c1c9550),
	.w2(32'hbb6c9cab),
	.w3(32'hbc88717a),
	.w4(32'hbc31b3d6),
	.w5(32'hbc0a1b31),
	.w6(32'hbb7cdc68),
	.w7(32'h3b389749),
	.w8(32'hbb956b95),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445a76),
	.w1(32'h3c272f50),
	.w2(32'h3ca1b638),
	.w3(32'hbb2b4060),
	.w4(32'h39a775c8),
	.w5(32'h3a90f49a),
	.w6(32'hbd314cb1),
	.w7(32'h3b52c7d4),
	.w8(32'h3bf42784),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bdc13),
	.w1(32'hbb92723e),
	.w2(32'h3a2e994a),
	.w3(32'hbc85be98),
	.w4(32'h3b34c443),
	.w5(32'hbc5ebeea),
	.w6(32'hbcc7844d),
	.w7(32'h3ba4ac59),
	.w8(32'hbcb7760d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008924),
	.w1(32'h3b83a417),
	.w2(32'hbbbe51b7),
	.w3(32'hbbc46ff1),
	.w4(32'hbaa9aadf),
	.w5(32'hbc1e341c),
	.w6(32'h3c89d384),
	.w7(32'h3c5a3130),
	.w8(32'hbd17e6e5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc697b34),
	.w1(32'hb96a3ae4),
	.w2(32'hbc29836e),
	.w3(32'h3c2fdf13),
	.w4(32'h3c176bdc),
	.w5(32'h3b2fc823),
	.w6(32'h3c46a8bc),
	.w7(32'h3b871961),
	.w8(32'h3d2e54e2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43f2d),
	.w1(32'h3aa01be7),
	.w2(32'h3cbe1a28),
	.w3(32'hbc00a631),
	.w4(32'hbc042178),
	.w5(32'hbb997c8a),
	.w6(32'hbcc38f7d),
	.w7(32'h3c56cd7d),
	.w8(32'hbbde4127),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde8303),
	.w1(32'hbbacfbc9),
	.w2(32'h3b8cc046),
	.w3(32'hbaa5041c),
	.w4(32'hbb505427),
	.w5(32'hbc2b800d),
	.w6(32'hbaf5ef06),
	.w7(32'h3b1ca60f),
	.w8(32'hbc09694d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc315e74),
	.w1(32'hbc3e4481),
	.w2(32'hbaa67294),
	.w3(32'hbc16fd3f),
	.w4(32'hbad4b009),
	.w5(32'h3b60ecc3),
	.w6(32'hbc1d284a),
	.w7(32'h3aedab94),
	.w8(32'hbadcd61e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc2c2),
	.w1(32'h3b373d4d),
	.w2(32'hbb859a2d),
	.w3(32'hbb58ee79),
	.w4(32'hbbdb23b1),
	.w5(32'hbc237c07),
	.w6(32'h3afc69da),
	.w7(32'hbc7ca2eb),
	.w8(32'h3bc42fe6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce233b8),
	.w1(32'hbc567513),
	.w2(32'h3bc6593e),
	.w3(32'hbc639ef8),
	.w4(32'hbbb97855),
	.w5(32'hba272955),
	.w6(32'hbc4032dc),
	.w7(32'h3b20e904),
	.w8(32'hbc9c7985),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8821d7),
	.w1(32'h3cf36127),
	.w2(32'h3d3163e4),
	.w3(32'h3c86d548),
	.w4(32'hbaa4f543),
	.w5(32'h3b0a28b8),
	.w6(32'hbd248ba3),
	.w7(32'hbc3f0e51),
	.w8(32'h3ce0d3fd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c106a46),
	.w1(32'h3b1a66d6),
	.w2(32'h3c344445),
	.w3(32'hbc2cbb95),
	.w4(32'hbbcb159c),
	.w5(32'hbcc8b192),
	.w6(32'hbc565111),
	.w7(32'hbb37b766),
	.w8(32'h3d0376c7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301f5e),
	.w1(32'hbbfab076),
	.w2(32'hbb4d1358),
	.w3(32'h3c20f792),
	.w4(32'hbba1454c),
	.w5(32'h3b8cb33c),
	.w6(32'hbbed5e21),
	.w7(32'h3c7f7f75),
	.w8(32'hbd4a4cf5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1687fa),
	.w1(32'hb80f16bf),
	.w2(32'h3b1b3424),
	.w3(32'hbc3382cf),
	.w4(32'h3b65f42c),
	.w5(32'h3b97b4b7),
	.w6(32'h3c6ae246),
	.w7(32'h3b193648),
	.w8(32'h3bb39a6a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395149a2),
	.w1(32'h3a9b3e66),
	.w2(32'h3a0f0a2b),
	.w3(32'hbb9a43ea),
	.w4(32'h3b7234bc),
	.w5(32'h3b279495),
	.w6(32'hba9dfbc8),
	.w7(32'hbbe7ec95),
	.w8(32'hbc0f83bf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac9f23),
	.w1(32'h3a75364e),
	.w2(32'hbc49eede),
	.w3(32'hbc15a9d7),
	.w4(32'hb9239146),
	.w5(32'h3bd3c32c),
	.w6(32'h3c710bb9),
	.w7(32'hbbf56bc7),
	.w8(32'h3c5e8061),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e15d6),
	.w1(32'hbad368ed),
	.w2(32'h3af6a803),
	.w3(32'h3bcdb95e),
	.w4(32'hbaa994c2),
	.w5(32'h3c2a49d9),
	.w6(32'hbc7c0c69),
	.w7(32'hbbce74ba),
	.w8(32'hbbc1faf4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4e1bf),
	.w1(32'h3c02f4d4),
	.w2(32'hbb512ef6),
	.w3(32'hbb433df2),
	.w4(32'h3ba77a9a),
	.w5(32'hbb746628),
	.w6(32'h3bfe95d7),
	.w7(32'h3beeecee),
	.w8(32'hbbe9260d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66bd00),
	.w1(32'h3c3ffbdd),
	.w2(32'h3b2e4d2a),
	.w3(32'h3bb3c023),
	.w4(32'hbabe107f),
	.w5(32'hbcbfa5a4),
	.w6(32'h3b13e1e2),
	.w7(32'h3c699bbd),
	.w8(32'hbca7dcf9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cb9ba),
	.w1(32'hbbd1459d),
	.w2(32'h3be164a0),
	.w3(32'h3a2ba1ec),
	.w4(32'h3b598c74),
	.w5(32'hbbd5b9a4),
	.w6(32'hbbf71484),
	.w7(32'hb987e4b3),
	.w8(32'h3c9607cd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34086),
	.w1(32'h3be60ba1),
	.w2(32'h3b3f5ad3),
	.w3(32'hbb83272a),
	.w4(32'hbb9f1a43),
	.w5(32'hbba9f940),
	.w6(32'hbc761745),
	.w7(32'hbb507510),
	.w8(32'h3b821e79),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984871),
	.w1(32'h3ac5bce6),
	.w2(32'h3c95945e),
	.w3(32'h3acd34b0),
	.w4(32'h3bcc3765),
	.w5(32'h3b8a0e35),
	.w6(32'hb8bbec9e),
	.w7(32'hba52dc76),
	.w8(32'h3d1416c7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9a18e),
	.w1(32'h3cdd72ca),
	.w2(32'h3b849fe8),
	.w3(32'hbcdbb063),
	.w4(32'h3bb16406),
	.w5(32'h3a9ad794),
	.w6(32'h3c22e787),
	.w7(32'h3bf75811),
	.w8(32'hbb27647a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd15c34e),
	.w1(32'hbc68c03e),
	.w2(32'hbc8d055a),
	.w3(32'hbd417c92),
	.w4(32'hbd1451a5),
	.w5(32'hbd036f6b),
	.w6(32'hbd646904),
	.w7(32'hbd12712a),
	.w8(32'hbd31bd96),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca94e9d),
	.w1(32'hbb50a3b2),
	.w2(32'h3c526dfd),
	.w3(32'hbc20cc2c),
	.w4(32'hbc4ee62a),
	.w5(32'hbba02965),
	.w6(32'hbbe61e5e),
	.w7(32'h3cd84ac3),
	.w8(32'hbd2255f8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a6017),
	.w1(32'h3bb5fa4a),
	.w2(32'hb92caa9e),
	.w3(32'h3c9df415),
	.w4(32'hbafab537),
	.w5(32'hbba18320),
	.w6(32'h3c05a230),
	.w7(32'hba9b24f9),
	.w8(32'hbb635ce3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700bc52),
	.w1(32'hbc78c5b9),
	.w2(32'hbbd7c0c2),
	.w3(32'h3acf9ae6),
	.w4(32'hbc02529b),
	.w5(32'hbc1fae33),
	.w6(32'hbc4aecd0),
	.w7(32'hbbd4d478),
	.w8(32'h3ba28424),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab01243),
	.w1(32'h3b0ef94f),
	.w2(32'h3a119b9d),
	.w3(32'hbbb7e22c),
	.w4(32'h3c338bf3),
	.w5(32'hbb648fd1),
	.w6(32'hbc1147be),
	.w7(32'hbb78616b),
	.w8(32'h3d61dd3b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc715ec5),
	.w1(32'hbb45cc3b),
	.w2(32'h3c40f093),
	.w3(32'hbc1ecbc8),
	.w4(32'h3c3ec05e),
	.w5(32'hba425e58),
	.w6(32'hbc6f526f),
	.w7(32'h3c8e78f7),
	.w8(32'h3c5e6eac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079c52),
	.w1(32'h3c01d4e2),
	.w2(32'h3a0f7739),
	.w3(32'h3b74f35f),
	.w4(32'hbbcaad7f),
	.w5(32'hbc244a3f),
	.w6(32'h3b319dad),
	.w7(32'h3c3e40a8),
	.w8(32'h3ba4b771),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe2cb4),
	.w1(32'hbbbac1ca),
	.w2(32'hb89147ab),
	.w3(32'hbc213fcc),
	.w4(32'hbaa879ed),
	.w5(32'h3c06c322),
	.w6(32'h3bf0ea62),
	.w7(32'hbc925625),
	.w8(32'h3da6a4fb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99e16),
	.w1(32'h39e1f4e9),
	.w2(32'h3aa1dd18),
	.w3(32'hbc464a94),
	.w4(32'h3aeb8e52),
	.w5(32'h3c31615f),
	.w6(32'hbc3571bb),
	.w7(32'h3c24c599),
	.w8(32'hbc5896c8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79a5e1),
	.w1(32'hbc0d05cc),
	.w2(32'hbcaaea52),
	.w3(32'hbb41dfe3),
	.w4(32'hbcb02151),
	.w5(32'hbbcbfdbe),
	.w6(32'hbc8b94d9),
	.w7(32'hbc2aa687),
	.w8(32'h3ca7cf2b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc61a12),
	.w1(32'hbc55d8ab),
	.w2(32'h3b62988e),
	.w3(32'hbd19beb9),
	.w4(32'h3bee87ae),
	.w5(32'h3c4902a9),
	.w6(32'hbc6d99ac),
	.w7(32'h3c415ee5),
	.w8(32'hbadbeeb0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd91871),
	.w1(32'h3c83d85b),
	.w2(32'hbc388010),
	.w3(32'hbcce5931),
	.w4(32'hbbe97ef7),
	.w5(32'hbbb3aefd),
	.w6(32'hbc90185b),
	.w7(32'hbc436e54),
	.w8(32'h3c00a686),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e79d),
	.w1(32'hbb2bb7a2),
	.w2(32'h3b02d09d),
	.w3(32'h3c5a3a02),
	.w4(32'h3ae5b7c3),
	.w5(32'h3b9ba53f),
	.w6(32'h3c10c60b),
	.w7(32'h3b6c2472),
	.w8(32'hbc7e804c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c0dcc),
	.w1(32'hbb7ed624),
	.w2(32'hbbcc9af8),
	.w3(32'hbc1c2b4d),
	.w4(32'hbbcb38df),
	.w5(32'hbb915d3b),
	.w6(32'h387249f2),
	.w7(32'hbbbe64b3),
	.w8(32'h3b616ebc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb23a60),
	.w1(32'h395de801),
	.w2(32'h3bc00b37),
	.w3(32'hbb1e1fa1),
	.w4(32'h3c3004fc),
	.w5(32'hbc54a6cd),
	.w6(32'hba1312d3),
	.w7(32'hbb0b807f),
	.w8(32'h3c4469d9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc813f43),
	.w1(32'hba31e389),
	.w2(32'hbc1bd0f8),
	.w3(32'h3c7af757),
	.w4(32'h3bdce706),
	.w5(32'h3c48911a),
	.w6(32'hbaa2849c),
	.w7(32'hbc555bb6),
	.w8(32'h3d2dbf93),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803a04),
	.w1(32'hba36ede1),
	.w2(32'h3ba0282a),
	.w3(32'h3c3ee45b),
	.w4(32'hbbeab415),
	.w5(32'hbab510a7),
	.w6(32'hbb22756a),
	.w7(32'hbae4c969),
	.w8(32'hbba6632d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14023b),
	.w1(32'h3c4f1e52),
	.w2(32'h3c682685),
	.w3(32'hbbb93f9b),
	.w4(32'h3bb4c34a),
	.w5(32'hbb884acd),
	.w6(32'hbb590545),
	.w7(32'h3c498731),
	.w8(32'hbb8c56c2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda69ca),
	.w1(32'h3b24511f),
	.w2(32'h3b6e45d9),
	.w3(32'hbc05e082),
	.w4(32'h3bacc3ae),
	.w5(32'h3b47d051),
	.w6(32'hbb2788bc),
	.w7(32'h3bf8d097),
	.w8(32'h3cb65ce6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79c5e8),
	.w1(32'hbb33e8e4),
	.w2(32'hb9c1db96),
	.w3(32'hbc0bde7a),
	.w4(32'hbc84c303),
	.w5(32'hbbf13555),
	.w6(32'hbb8365b2),
	.w7(32'hbc0f5456),
	.w8(32'h3a86e01a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1c31),
	.w1(32'hbc0953df),
	.w2(32'h3b992416),
	.w3(32'h3a6e2375),
	.w4(32'hbc65fb68),
	.w5(32'hbc32803d),
	.w6(32'hbbfdeca7),
	.w7(32'h3b8a7089),
	.w8(32'hbd0e2d3d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b1465),
	.w1(32'hbc35031a),
	.w2(32'hbac43af6),
	.w3(32'h3ba02e3a),
	.w4(32'hbc6c6a0d),
	.w5(32'hbb87723e),
	.w6(32'h3c63f0c6),
	.w7(32'hbbd2f523),
	.w8(32'hbafc76e0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf64a9a),
	.w1(32'hbc3d5277),
	.w2(32'h3bb236ea),
	.w3(32'hbcd79692),
	.w4(32'hbc6db362),
	.w5(32'hbce0f1ce),
	.w6(32'hbccc8a1e),
	.w7(32'hbceff617),
	.w8(32'hbc346f17),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3068b6),
	.w1(32'hbc353e9e),
	.w2(32'h3c7615f7),
	.w3(32'h3a04ce8d),
	.w4(32'h3c39d27c),
	.w5(32'h3bdff41c),
	.w6(32'hbc4c285d),
	.w7(32'h3ad4a7f5),
	.w8(32'h3c833b5a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522e6e),
	.w1(32'h3c9f4288),
	.w2(32'h3842efda),
	.w3(32'hbc98a954),
	.w4(32'hbae0677c),
	.w5(32'hb9467bbf),
	.w6(32'h3c86675f),
	.w7(32'h3b1e4aa5),
	.w8(32'hbbe1fd00),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480a36),
	.w1(32'hbc31f162),
	.w2(32'h3c24edb3),
	.w3(32'h3c11baa2),
	.w4(32'hbaada35d),
	.w5(32'h39477c94),
	.w6(32'hba560dc8),
	.w7(32'h3ab2fd96),
	.w8(32'hb9d9239b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c5ba1),
	.w1(32'h3a7602ef),
	.w2(32'h3a94c81e),
	.w3(32'hbba12703),
	.w4(32'hbc0bb94a),
	.w5(32'h3c2ae888),
	.w6(32'h3af70538),
	.w7(32'h3bbe46f0),
	.w8(32'hbb6e0ae3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b4108),
	.w1(32'h3c21a7e4),
	.w2(32'h3c45379a),
	.w3(32'hbd14daed),
	.w4(32'hbb2084eb),
	.w5(32'h3c23ce69),
	.w6(32'h3beef7ec),
	.w7(32'h3aa3f4d8),
	.w8(32'hbd0f1879),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe318bf),
	.w1(32'hbb844c4e),
	.w2(32'h3a07dfdc),
	.w3(32'h3c37d1a0),
	.w4(32'h393d3a71),
	.w5(32'hbbd76bb6),
	.w6(32'h3cafd84c),
	.w7(32'h3c848a6e),
	.w8(32'h3d01c554),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95810a),
	.w1(32'h3ca0ca08),
	.w2(32'h3bada9bc),
	.w3(32'h3b826f11),
	.w4(32'hbc125a28),
	.w5(32'h3c7ee008),
	.w6(32'h3c8e86d2),
	.w7(32'hbb49b2b6),
	.w8(32'h39b5e37f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f46a5),
	.w1(32'hbc6a1f7e),
	.w2(32'h3c4a64d9),
	.w3(32'hb883c453),
	.w4(32'hbc82769d),
	.w5(32'hbbc73885),
	.w6(32'hbad3d09e),
	.w7(32'h3beb9910),
	.w8(32'hbcf18707),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd77a6),
	.w1(32'hbcb2e628),
	.w2(32'h3ca4fba1),
	.w3(32'h3c123fd4),
	.w4(32'h3b828e32),
	.w5(32'h3d1f71b0),
	.w6(32'h3a487c7d),
	.w7(32'hbb39fa2a),
	.w8(32'h3c14d530),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c4e5c),
	.w1(32'h3c94df9c),
	.w2(32'hbae01f4b),
	.w3(32'hbc780603),
	.w4(32'h3bfd2f31),
	.w5(32'hba8bb3f7),
	.w6(32'hbbbf2433),
	.w7(32'hb6ab3cb5),
	.w8(32'hbc48ed26),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45a8b8),
	.w1(32'hbbc41223),
	.w2(32'hbbb7c9c7),
	.w3(32'hbb5f8bb2),
	.w4(32'h3ba3f034),
	.w5(32'h3b74d750),
	.w6(32'hbbeb9482),
	.w7(32'h3bec1295),
	.w8(32'hbcd05fa8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f977c),
	.w1(32'hba28dc4f),
	.w2(32'hbbb5b8a0),
	.w3(32'h3be7e4a6),
	.w4(32'h3c07c7bf),
	.w5(32'hbbb15b09),
	.w6(32'h3bbffdbc),
	.w7(32'h3c367a37),
	.w8(32'hbc07c462),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824e3f),
	.w1(32'h3bf9c84b),
	.w2(32'h3c08e0ad),
	.w3(32'h3be5907d),
	.w4(32'h3c3eca59),
	.w5(32'h3d13d638),
	.w6(32'h3b923c11),
	.w7(32'hbc17b244),
	.w8(32'h3d2d827c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7a531),
	.w1(32'h3c233c76),
	.w2(32'h3ba62d8c),
	.w3(32'hb921f26c),
	.w4(32'h3af6f2ea),
	.w5(32'h3aa33be6),
	.w6(32'h3b28f976),
	.w7(32'h3be2e704),
	.w8(32'h3b292445),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd72dd1),
	.w1(32'h3b00609d),
	.w2(32'hbab76d94),
	.w3(32'hbc31987e),
	.w4(32'hbbd9565e),
	.w5(32'hbb4c30f1),
	.w6(32'hbc6401d9),
	.w7(32'hbc405e7b),
	.w8(32'hbbdcd2da),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc296ddb),
	.w1(32'hbb14fcad),
	.w2(32'hbb1db50d),
	.w3(32'hbc1cb5ae),
	.w4(32'hbc03db61),
	.w5(32'h3a13209c),
	.w6(32'hbc45136d),
	.w7(32'hbc44e985),
	.w8(32'hbc04c87c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc18c94),
	.w1(32'hbb59124a),
	.w2(32'hbb3a6996),
	.w3(32'hbb513f4a),
	.w4(32'h3b3a5173),
	.w5(32'h3ae5d8b8),
	.w6(32'hbb9e45c3),
	.w7(32'hbbb334f4),
	.w8(32'hbbfd2e1c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0792d6),
	.w1(32'hba5dd102),
	.w2(32'hbbcbbc72),
	.w3(32'hbb1d1332),
	.w4(32'hbbaac05f),
	.w5(32'h3a909d35),
	.w6(32'hbb64a893),
	.w7(32'h3b7aba01),
	.w8(32'hbab47e52),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0981d6),
	.w1(32'hbc0357c3),
	.w2(32'hbaa18149),
	.w3(32'h3a148851),
	.w4(32'h3b15a29d),
	.w5(32'hbb0b42ff),
	.w6(32'h3b591d6d),
	.w7(32'hba3a0c7b),
	.w8(32'hba421267),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9225),
	.w1(32'hba4a8035),
	.w2(32'hbb4a2801),
	.w3(32'hbca3a145),
	.w4(32'hbbb73466),
	.w5(32'hbafcfc5a),
	.w6(32'hbc96edee),
	.w7(32'hbb72acf0),
	.w8(32'hbb23c9ea),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01b964),
	.w1(32'hbc6925bf),
	.w2(32'hba42fc74),
	.w3(32'hbd4580e7),
	.w4(32'hbceee7a7),
	.w5(32'hbccb3931),
	.w6(32'hbd400257),
	.w7(32'hbc259608),
	.w8(32'hbd0e5df0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd22e5b),
	.w1(32'hbc6f3008),
	.w2(32'hbaf5fbfa),
	.w3(32'hbd068d88),
	.w4(32'hbc621b5a),
	.w5(32'hbc59cf3c),
	.w6(32'hbd3504fc),
	.w7(32'hbca91272),
	.w8(32'h38e832c2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50f212),
	.w1(32'h3c4b3c39),
	.w2(32'hbbb62adf),
	.w3(32'hbc4b333e),
	.w4(32'hbbdc2ac6),
	.w5(32'hbc9a70f0),
	.w6(32'hbc018d4a),
	.w7(32'hbb6e0ef8),
	.w8(32'hbbbd1c90),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617a64),
	.w1(32'hbb6a4fbb),
	.w2(32'hbc5c695a),
	.w3(32'hbb8ec7b5),
	.w4(32'hbc605a9e),
	.w5(32'hbc9c9bb6),
	.w6(32'hbc49930d),
	.w7(32'hbc9b12c4),
	.w8(32'hbcd80ec7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad7e2b),
	.w1(32'hbc8f6a0c),
	.w2(32'h3c3a096d),
	.w3(32'hbc02906b),
	.w4(32'h3c14efaf),
	.w5(32'h3c553db4),
	.w6(32'hbccf0acb),
	.w7(32'h3b800940),
	.w8(32'h3b8377de),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d67f),
	.w1(32'hb9ae3f95),
	.w2(32'hbb5497d2),
	.w3(32'hba3af681),
	.w4(32'hbb16b96a),
	.w5(32'hbb122897),
	.w6(32'hba586c29),
	.w7(32'hbbb65f0c),
	.w8(32'hbbbd25ca),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394c7d),
	.w1(32'h39c2a8d9),
	.w2(32'h3c0589fb),
	.w3(32'h39d2c313),
	.w4(32'hbc18f001),
	.w5(32'h387b9290),
	.w6(32'hbb5cc002),
	.w7(32'h3bbc0c2c),
	.w8(32'hbaceca61),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e6e6),
	.w1(32'hbc069f97),
	.w2(32'hbb0a9a1a),
	.w3(32'hbc5e3d64),
	.w4(32'h3b27f1be),
	.w5(32'h3b3a03e4),
	.w6(32'hbbe39007),
	.w7(32'h3a4ad129),
	.w8(32'hbc0e07b9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35a8ed),
	.w1(32'hbb877466),
	.w2(32'h3ab2f3b7),
	.w3(32'h3b6dbf3f),
	.w4(32'hba642077),
	.w5(32'hba69721e),
	.w6(32'hbb2f5de3),
	.w7(32'hb90f7121),
	.w8(32'hba82f03f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb577b7a),
	.w1(32'hbb084def),
	.w2(32'h3b6d87b3),
	.w3(32'hbbd3a36c),
	.w4(32'hbc9a0f8c),
	.w5(32'hbc904641),
	.w6(32'hbc8d5ee0),
	.w7(32'h3c355ebf),
	.w8(32'hbb8aabe9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3010d9),
	.w1(32'hbc60f84d),
	.w2(32'hbc17d9f9),
	.w3(32'hbc9b973e),
	.w4(32'h3aabf630),
	.w5(32'h3c83fb82),
	.w6(32'hbc7cb1a0),
	.w7(32'hbc3b7e11),
	.w8(32'h3cc5e3f8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc647521),
	.w1(32'h39ebdea2),
	.w2(32'hbb9a5231),
	.w3(32'h3a457cf9),
	.w4(32'hbb440a4d),
	.w5(32'hbb40b920),
	.w6(32'h3c28be90),
	.w7(32'hbbb92b49),
	.w8(32'hbbea818f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ffdba),
	.w1(32'hb99df91b),
	.w2(32'h3c15ffa1),
	.w3(32'hbbc34f9a),
	.w4(32'hbbfca380),
	.w5(32'hbbecb10d),
	.w6(32'hbc53b38a),
	.w7(32'hbb8fc132),
	.w8(32'hbb8e8a3e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd59e9),
	.w1(32'h3b395ab1),
	.w2(32'h3c277d26),
	.w3(32'hbcb97c0f),
	.w4(32'h3afec381),
	.w5(32'h3c3c0f2b),
	.w6(32'hbcad6efe),
	.w7(32'h3ba6be68),
	.w8(32'h3cf3d732),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b82a0),
	.w1(32'hb93347eb),
	.w2(32'hbc0d3cbe),
	.w3(32'h3a05271f),
	.w4(32'h3b02c94d),
	.w5(32'h3a8d9906),
	.w6(32'h3bb0420e),
	.w7(32'hbc141a51),
	.w8(32'hbc3ef9dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b31d),
	.w1(32'hbaa51e76),
	.w2(32'h3cd100ff),
	.w3(32'h3af8fe5b),
	.w4(32'h3d077ad5),
	.w5(32'h3c391bac),
	.w6(32'h3a6271ce),
	.w7(32'h3cefa4a0),
	.w8(32'h3c4af674),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1405ac),
	.w1(32'h3afe8634),
	.w2(32'hbb8a8979),
	.w3(32'hbb62ea92),
	.w4(32'hbb92d713),
	.w5(32'h3a2871ba),
	.w6(32'hb98b04e7),
	.w7(32'h3ba445e1),
	.w8(32'h3c7b68b6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12740e),
	.w1(32'h3c6b05f1),
	.w2(32'hbbac002c),
	.w3(32'h3bae84bf),
	.w4(32'hbb87e2fa),
	.w5(32'hba8038b2),
	.w6(32'h3c155916),
	.w7(32'hb92c9b8d),
	.w8(32'hbc4535fb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80d63),
	.w1(32'hbc19100f),
	.w2(32'hbba722bc),
	.w3(32'hbb15f99f),
	.w4(32'hbba834bf),
	.w5(32'hbbf94f63),
	.w6(32'hbbfe4072),
	.w7(32'hbbb3b918),
	.w8(32'hbc334d4f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61f917),
	.w1(32'hb9acd832),
	.w2(32'h3c6f5de8),
	.w3(32'h3aab7c2a),
	.w4(32'h3ab7516e),
	.w5(32'hbb40e3bd),
	.w6(32'hbbcdd172),
	.w7(32'h3ce9ac9a),
	.w8(32'h3abbe407),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb450b6),
	.w1(32'hbc148dbc),
	.w2(32'h3ba5d2bb),
	.w3(32'hbc79e196),
	.w4(32'hbb02f0f4),
	.w5(32'hbb1bf499),
	.w6(32'hbb358326),
	.w7(32'h3c0d2682),
	.w8(32'h3bbbcc75),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd81436),
	.w1(32'h3ac74eac),
	.w2(32'h3c15322e),
	.w3(32'hba09b495),
	.w4(32'h3c3d889a),
	.w5(32'h3bd36bcb),
	.w6(32'h3b9c492a),
	.w7(32'h3bd7f151),
	.w8(32'h3a5a7da7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003251),
	.w1(32'hbbbb2736),
	.w2(32'h3c27f67b),
	.w3(32'hbbf4f16b),
	.w4(32'hbb22347c),
	.w5(32'hbbf8ad22),
	.w6(32'hbba4ef96),
	.w7(32'hbbf35bd8),
	.w8(32'hbba46f54),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b63dd),
	.w1(32'h3abf4073),
	.w2(32'hbc32f8ce),
	.w3(32'hbb2f65c5),
	.w4(32'h3b0b6971),
	.w5(32'hbbb9f913),
	.w6(32'hbb384eac),
	.w7(32'h3c66516f),
	.w8(32'h3c933e45),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb1cfe),
	.w1(32'h3a1bf98f),
	.w2(32'h3b986b58),
	.w3(32'hbbe5eea9),
	.w4(32'h3bb06b0f),
	.w5(32'h3b3bb717),
	.w6(32'hbb8de521),
	.w7(32'h3c37279b),
	.w8(32'h3b081094),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc70d7),
	.w1(32'h3adc52d6),
	.w2(32'hba6a4c00),
	.w3(32'h3b531644),
	.w4(32'hbba23c2b),
	.w5(32'hbc56a5e9),
	.w6(32'h3b856e48),
	.w7(32'h3cd144c4),
	.w8(32'h3b5592fa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840ee5),
	.w1(32'hbabbfc3b),
	.w2(32'h3bb9a027),
	.w3(32'hbc6fd7eb),
	.w4(32'hbc41ebbc),
	.w5(32'h3bcda30b),
	.w6(32'hbbdc3bb9),
	.w7(32'hbc1280ae),
	.w8(32'h3b99e1ba),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5d8c8),
	.w1(32'h3bf5524a),
	.w2(32'hbaba7771),
	.w3(32'h39d3bf86),
	.w4(32'h3a296de6),
	.w5(32'hbad5f672),
	.w6(32'h3bad6b1e),
	.w7(32'h3ccd565a),
	.w8(32'h3c02eda7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3135a2),
	.w1(32'h3c08f377),
	.w2(32'hbc644329),
	.w3(32'hbc54a947),
	.w4(32'hbc2463f2),
	.w5(32'hbbbcfe92),
	.w6(32'h3acc6879),
	.w7(32'h3a9bc72a),
	.w8(32'hbb0a0751),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2ddd2),
	.w1(32'hbbcb1b11),
	.w2(32'h3bb45209),
	.w3(32'hbb80f0a7),
	.w4(32'h3bdb643f),
	.w5(32'hbab84dfc),
	.w6(32'hbb66e195),
	.w7(32'h3b19df61),
	.w8(32'hbaf418b3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f511),
	.w1(32'hbba0e3c4),
	.w2(32'hbb78e62a),
	.w3(32'hbba63979),
	.w4(32'hbbf89aa8),
	.w5(32'hbb940b99),
	.w6(32'hbb8683ce),
	.w7(32'hbc0b27f2),
	.w8(32'hbc6e11d1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2b07),
	.w1(32'hbc3e57c8),
	.w2(32'h3c5e4c81),
	.w3(32'hbb85bbb7),
	.w4(32'hbb792a05),
	.w5(32'hbaf21092),
	.w6(32'hbb971951),
	.w7(32'hbc05ed4c),
	.w8(32'hbc1f3957),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46d961),
	.w1(32'hbc2c0fa6),
	.w2(32'h3c6b770e),
	.w3(32'h3b19948f),
	.w4(32'h3aadbd9b),
	.w5(32'hbb345014),
	.w6(32'hbc4a17e9),
	.w7(32'hbb27ac88),
	.w8(32'h3c543ddc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6958e4),
	.w1(32'h3b3fa83c),
	.w2(32'hbacf853e),
	.w3(32'h3a71f9d5),
	.w4(32'h3b5821e5),
	.w5(32'hbb006206),
	.w6(32'h3b88ee00),
	.w7(32'h3a3422b9),
	.w8(32'hbbcad4a3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd6485),
	.w1(32'hbab6e328),
	.w2(32'h3bdc6925),
	.w3(32'hbbf7b849),
	.w4(32'h3b4df369),
	.w5(32'h3b3326ad),
	.w6(32'hbbeed40e),
	.w7(32'h3b35d8d1),
	.w8(32'h3900b3cd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19393c),
	.w1(32'h39dd6a35),
	.w2(32'hbb519bb4),
	.w3(32'hba33f02d),
	.w4(32'hbb76cfd0),
	.w5(32'h3b375383),
	.w6(32'hbaf120b9),
	.w7(32'h3b69fa88),
	.w8(32'h3c124b83),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef4ded),
	.w1(32'hba9f7fe4),
	.w2(32'h3aa05a20),
	.w3(32'hbba5fe78),
	.w4(32'h3a8ac9a6),
	.w5(32'hbbe951bb),
	.w6(32'hbb613599),
	.w7(32'hbb9b2669),
	.w8(32'hbb864c54),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36c0ef),
	.w1(32'hbbd3e89a),
	.w2(32'hbafc41da),
	.w3(32'hbc63b750),
	.w4(32'hbbfed647),
	.w5(32'hbb8f6009),
	.w6(32'hbc01e23d),
	.w7(32'hbb923ce2),
	.w8(32'hbb96edc4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb209ff4),
	.w1(32'hbb2014aa),
	.w2(32'hbc0bdcce),
	.w3(32'h3b5d615a),
	.w4(32'hbb993d81),
	.w5(32'h39c3d311),
	.w6(32'hb9ba993b),
	.w7(32'hbbba0f4d),
	.w8(32'hbae1b231),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afad443),
	.w1(32'hbbb43625),
	.w2(32'h3b3413e3),
	.w3(32'h3b32608a),
	.w4(32'h3adeb036),
	.w5(32'h3a736780),
	.w6(32'hbb9a3827),
	.w7(32'h3b7cdd02),
	.w8(32'hba9df4e4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88500),
	.w1(32'h3a73ec04),
	.w2(32'h3bbef500),
	.w3(32'h3b4aadbf),
	.w4(32'hbc26223f),
	.w5(32'hbc865d8c),
	.w6(32'h3b787f8e),
	.w7(32'hbacd200c),
	.w8(32'hbbae56d2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6898b),
	.w1(32'hbb07ca67),
	.w2(32'h3b81df74),
	.w3(32'hbc370f8b),
	.w4(32'hbbd48c97),
	.w5(32'hbb2d4775),
	.w6(32'hbc045a82),
	.w7(32'hba1b95d4),
	.w8(32'h3bb13881),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24881a),
	.w1(32'hbb892da0),
	.w2(32'hb8e510a2),
	.w3(32'hbbeb964a),
	.w4(32'hbc2d1bbe),
	.w5(32'hbbe2ea67),
	.w6(32'hbb1dac29),
	.w7(32'hbb6f641a),
	.w8(32'hbbf4dfc3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7526b),
	.w1(32'hbb81c9d2),
	.w2(32'hbca1f29f),
	.w3(32'hbbf83958),
	.w4(32'hbbb72d28),
	.w5(32'hbbe21df9),
	.w6(32'hbbc6cf7c),
	.w7(32'hbc47c65a),
	.w8(32'hbc78de37),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78ee13),
	.w1(32'hbc36dd5e),
	.w2(32'h3b6b6f7a),
	.w3(32'hbc35e8fd),
	.w4(32'h3b124e0f),
	.w5(32'hba06a63c),
	.w6(32'hbc682481),
	.w7(32'h37ef6013),
	.w8(32'h3b65260c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule