module LineBuffer(data_in, data_out, Clk, valid_in, valid_out, Rst);
    parameter DATA_WIDTH = 32;
    parameter COUNTER_WIDTH = 7;
    parameter BUFFER_DEPTH = 97;

    input  Clk, valid_in, Rst;
    input  [DATA_WIDTH - 1:0] data_in;

    output valid_out;
    output reg [DATA_WIDTH - 1:0] data_out;

	reg [DATA_WIDTH - 1:0] Buffer [BUFFER_DEPTH - 1:0];
    reg [COUNTER_WIDTH - 1:0] Counter;
	 
    always @ (posedge Clk or negedge Rst) begin
		if (!Rst) Counter <= 0;
        else begin
            if (valid_in) begin
                if (Counter >= BUFFER_DEPTH) Counter <= Counter;
                else Counter <= Counter + 1;

                data_out <= Buffer[BUFFER_DEPTH - 1];
                
                Buffer[1] <= Buffer[0];
                Buffer[2] <= Buffer[1];
                Buffer[3] <= Buffer[2];
                Buffer[4] <= Buffer[3];
                Buffer[5] <= Buffer[4];
                Buffer[6] <= Buffer[5];
                Buffer[7] <= Buffer[6];
                Buffer[8] <= Buffer[7];
                Buffer[9] <= Buffer[8];
                Buffer[10] <= Buffer[9];
                Buffer[11] <= Buffer[10];
                Buffer[12] <= Buffer[11];
                Buffer[13] <= Buffer[12];
                Buffer[14] <= Buffer[13];
                Buffer[15] <= Buffer[14];
                Buffer[16] <= Buffer[15];
                Buffer[17] <= Buffer[16];
                Buffer[18] <= Buffer[17];
                Buffer[19] <= Buffer[18];
                Buffer[20] <= Buffer[19];
                Buffer[21] <= Buffer[20];
                Buffer[22] <= Buffer[21];
                Buffer[23] <= Buffer[22];
                Buffer[24] <= Buffer[23];
                Buffer[25] <= Buffer[24];
                Buffer[26] <= Buffer[25];
                Buffer[27] <= Buffer[26];
                Buffer[28] <= Buffer[27];
                Buffer[29] <= Buffer[28];
                Buffer[30] <= Buffer[29];
                Buffer[31] <= Buffer[30];
                Buffer[32] <= Buffer[31];
                Buffer[33] <= Buffer[32];
                Buffer[34] <= Buffer[33];
                Buffer[35] <= Buffer[34];
                Buffer[36] <= Buffer[35];
                Buffer[37] <= Buffer[36];
                Buffer[38] <= Buffer[37];
                Buffer[39] <= Buffer[38];
                Buffer[40] <= Buffer[39];
                Buffer[41] <= Buffer[40];
                Buffer[42] <= Buffer[41];
                Buffer[43] <= Buffer[42];
                Buffer[44] <= Buffer[43];
                Buffer[45] <= Buffer[44];
                Buffer[46] <= Buffer[45];
                Buffer[47] <= Buffer[46];
                Buffer[48] <= Buffer[47];
                Buffer[49] <= Buffer[48];
                Buffer[50] <= Buffer[49];
                Buffer[51] <= Buffer[50];
                Buffer[52] <= Buffer[51];
                Buffer[53] <= Buffer[52];
                Buffer[54] <= Buffer[53];
                Buffer[55] <= Buffer[54];
                Buffer[56] <= Buffer[55];
                Buffer[57] <= Buffer[56];
                Buffer[58] <= Buffer[57];
                Buffer[59] <= Buffer[58];
                Buffer[60] <= Buffer[59];
                Buffer[61] <= Buffer[60];
                Buffer[62] <= Buffer[61];
                Buffer[63] <= Buffer[62];
                Buffer[64] <= Buffer[63];
                Buffer[65] <= Buffer[64];
                Buffer[66] <= Buffer[65];
                Buffer[67] <= Buffer[66];
                Buffer[68] <= Buffer[67];
                Buffer[69] <= Buffer[68];
                Buffer[70] <= Buffer[69];
                Buffer[71] <= Buffer[70];
                Buffer[72] <= Buffer[71];
                Buffer[73] <= Buffer[72];
                Buffer[74] <= Buffer[73];
                Buffer[75] <= Buffer[74];
                Buffer[76] <= Buffer[75];
                Buffer[77] <= Buffer[76];
                Buffer[78] <= Buffer[77];
                Buffer[79] <= Buffer[78];
                Buffer[80] <= Buffer[79];
                Buffer[81] <= Buffer[80];
                Buffer[82] <= Buffer[81];
                Buffer[83] <= Buffer[82];
                Buffer[84] <= Buffer[83];
                Buffer[85] <= Buffer[84];
                Buffer[86] <= Buffer[85];
                Buffer[87] <= Buffer[86];
                Buffer[88] <= Buffer[87];
                Buffer[89] <= Buffer[88];
                Buffer[90] <= Buffer[89];
                Buffer[91] <= Buffer[90];
                Buffer[92] <= Buffer[91];
                Buffer[93] <= Buffer[92];
                Buffer[94] <= Buffer[93];
                Buffer[95] <= Buffer[94];
                Buffer[96] <= Buffer[95];
                
                Buffer[0] <= data_in;
            end else begin
                Counter <= Counter;

                Buffer[0] <= Buffer[0];
                Buffer[1] <= Buffer[1];
                Buffer[2] <= Buffer[2];
                Buffer[3] <= Buffer[3];
                Buffer[4] <= Buffer[4];
                Buffer[5] <= Buffer[5];
                Buffer[6] <= Buffer[6];
                Buffer[7] <= Buffer[7];
                Buffer[8] <= Buffer[8];
                Buffer[9] <= Buffer[9];
                Buffer[10] <= Buffer[10];
                Buffer[11] <= Buffer[11];
                Buffer[12] <= Buffer[12];
                Buffer[13] <= Buffer[13];
                Buffer[14] <= Buffer[14];
                Buffer[15] <= Buffer[15];
                Buffer[16] <= Buffer[16];
                Buffer[17] <= Buffer[17];
                Buffer[18] <= Buffer[18];
                Buffer[19] <= Buffer[19];
                Buffer[20] <= Buffer[20];
                Buffer[21] <= Buffer[21];
                Buffer[22] <= Buffer[22];
                Buffer[23] <= Buffer[23];
                Buffer[24] <= Buffer[24];
                Buffer[25] <= Buffer[25];
                Buffer[26] <= Buffer[26];
                Buffer[27] <= Buffer[27];
                Buffer[28] <= Buffer[28];
                Buffer[29] <= Buffer[29];
                Buffer[30] <= Buffer[30];
                Buffer[31] <= Buffer[31];
                Buffer[32] <= Buffer[32];
                Buffer[33] <= Buffer[33];
                Buffer[34] <= Buffer[34];
                Buffer[35] <= Buffer[35];
                Buffer[36] <= Buffer[36];
                Buffer[37] <= Buffer[37];
                Buffer[38] <= Buffer[38];
                Buffer[39] <= Buffer[39];
                Buffer[40] <= Buffer[40];
                Buffer[41] <= Buffer[41];
                Buffer[42] <= Buffer[42];
                Buffer[43] <= Buffer[43];
                Buffer[44] <= Buffer[44];
                Buffer[45] <= Buffer[45];
                Buffer[46] <= Buffer[46];
                Buffer[47] <= Buffer[47];
                Buffer[48] <= Buffer[48];
                Buffer[49] <= Buffer[49];
                Buffer[50] <= Buffer[50];
                Buffer[51] <= Buffer[51];
                Buffer[52] <= Buffer[52];
                Buffer[53] <= Buffer[53];
                Buffer[54] <= Buffer[54];
                Buffer[55] <= Buffer[55];
                Buffer[56] <= Buffer[56];
                Buffer[57] <= Buffer[57];
                Buffer[58] <= Buffer[58];
                Buffer[59] <= Buffer[59];
                Buffer[60] <= Buffer[60];
                Buffer[61] <= Buffer[61];
                Buffer[62] <= Buffer[62];
                Buffer[63] <= Buffer[63];
                Buffer[64] <= Buffer[64];
                Buffer[65] <= Buffer[65];
                Buffer[66] <= Buffer[66];
                Buffer[67] <= Buffer[67];
                Buffer[68] <= Buffer[68];
                Buffer[69] <= Buffer[69];
                Buffer[70] <= Buffer[70];
                Buffer[71] <= Buffer[71];
                Buffer[72] <= Buffer[72];
                Buffer[73] <= Buffer[73];
                Buffer[74] <= Buffer[74];
                Buffer[75] <= Buffer[75];
                Buffer[76] <= Buffer[76];
                Buffer[77] <= Buffer[77];
                Buffer[78] <= Buffer[78];
                Buffer[79] <= Buffer[79];
                Buffer[80] <= Buffer[80];
                Buffer[81] <= Buffer[81];
                Buffer[82] <= Buffer[82];
                Buffer[83] <= Buffer[83];
                Buffer[84] <= Buffer[84];
                Buffer[85] <= Buffer[85];
                Buffer[86] <= Buffer[86];
                Buffer[87] <= Buffer[87];
                Buffer[88] <= Buffer[88];
                Buffer[89] <= Buffer[89];
                Buffer[90] <= Buffer[90];
                Buffer[91] <= Buffer[91];
                Buffer[92] <= Buffer[92];
                Buffer[93] <= Buffer[93];
                Buffer[94] <= Buffer[94];
                Buffer[95] <= Buffer[95];
                Buffer[96] <= Buffer[96];
            end
        end
	end

    assign valid_out = (Counter >= BUFFER_DEPTH) ? 1'b1 : 1'b0;

endmodule