module layer_10_featuremap_273(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abe33),
	.w1(32'hba7a3269),
	.w2(32'h3b0677be),
	.w3(32'hba338c71),
	.w4(32'hba82a85e),
	.w5(32'hbb756475),
	.w6(32'hbb11e0d8),
	.w7(32'h3b5664b5),
	.w8(32'hba340e88),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80dac),
	.w1(32'hbb8268be),
	.w2(32'hbb90b3d0),
	.w3(32'hbae09c59),
	.w4(32'hbbb70641),
	.w5(32'h381e811c),
	.w6(32'hbb68376f),
	.w7(32'hbb7f3e1f),
	.w8(32'h3b5c8332),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed91c),
	.w1(32'hbc98f389),
	.w2(32'hbc09f634),
	.w3(32'hbc26f599),
	.w4(32'hbcb6706b),
	.w5(32'hbb376711),
	.w6(32'hbbc481a0),
	.w7(32'hbcbea067),
	.w8(32'hbb81fc3d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e2c1),
	.w1(32'hb9a3573c),
	.w2(32'hbabfa4ab),
	.w3(32'hbbaf96b5),
	.w4(32'hbc0adc69),
	.w5(32'hba9d8baa),
	.w6(32'h3a0a1de3),
	.w7(32'hbc04ecdd),
	.w8(32'hbbaa322c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834f5c),
	.w1(32'hbc05c5b2),
	.w2(32'hbae8560e),
	.w3(32'hbc1ead45),
	.w4(32'h39f3bdf5),
	.w5(32'h3b184d3b),
	.w6(32'hbb3066d8),
	.w7(32'hbbb37a18),
	.w8(32'h3b2bd611),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfdfdb),
	.w1(32'hbb044fa2),
	.w2(32'hba664227),
	.w3(32'h3b0dd8b5),
	.w4(32'h3a9af755),
	.w5(32'h39fbd743),
	.w6(32'h3ac6f469),
	.w7(32'hba4d347c),
	.w8(32'h3af970ac),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf45fa0),
	.w1(32'h3c47fc4d),
	.w2(32'hbbdf1db3),
	.w3(32'h3b8f5f4c),
	.w4(32'h3c0bd457),
	.w5(32'hbbe29540),
	.w6(32'h3aa864a4),
	.w7(32'h3bf4452f),
	.w8(32'hbbbf8fd8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc5d90),
	.w1(32'h3b1bc7a7),
	.w2(32'hbb0a434f),
	.w3(32'hbbf348cd),
	.w4(32'h3c044c2e),
	.w5(32'hba8e94be),
	.w6(32'hbc1100de),
	.w7(32'hbb02a5e5),
	.w8(32'hba629c4c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b5987),
	.w1(32'hb8aadca8),
	.w2(32'h3ba707a6),
	.w3(32'h3b1daae7),
	.w4(32'h3bb4d438),
	.w5(32'h3b13d316),
	.w6(32'hba4d236c),
	.w7(32'h3b89268c),
	.w8(32'h3b1a9411),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58cd07),
	.w1(32'h39d4ed7e),
	.w2(32'hbbf1cd96),
	.w3(32'h3b1bff2f),
	.w4(32'h3b953537),
	.w5(32'hbbc1132c),
	.w6(32'h3ac4837a),
	.w7(32'h3a656362),
	.w8(32'hbbd6f00e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a7ff),
	.w1(32'hbbd3f6f2),
	.w2(32'hbb9ea726),
	.w3(32'hba91fd40),
	.w4(32'h3a331413),
	.w5(32'hbc03d6ed),
	.w6(32'h3c0f0f63),
	.w7(32'hbb829d0a),
	.w8(32'hbb619c76),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e4037),
	.w1(32'h3d1f6f70),
	.w2(32'h3a009834),
	.w3(32'hbac48c31),
	.w4(32'h3d088780),
	.w5(32'h3bae26a7),
	.w6(32'h3c50060c),
	.w7(32'h3d24d1f0),
	.w8(32'h3c12e741),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63d9ec),
	.w1(32'h3bb182f6),
	.w2(32'hbbc9027f),
	.w3(32'h3c13941c),
	.w4(32'h3bb71c05),
	.w5(32'hbc0d874b),
	.w6(32'h3b5c64e8),
	.w7(32'h3b390c8a),
	.w8(32'hbbcb2c7c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc8c8b),
	.w1(32'h3b994034),
	.w2(32'hbb77d9ae),
	.w3(32'h3a292d5d),
	.w4(32'hbc4f90b0),
	.w5(32'hbb81a3c4),
	.w6(32'h3c87191c),
	.w7(32'hbc1228fd),
	.w8(32'hbb625821),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b021),
	.w1(32'hbae27e67),
	.w2(32'h38cd34ad),
	.w3(32'h3b11709f),
	.w4(32'hbb83d39d),
	.w5(32'hbc70e0c5),
	.w6(32'h3b4fdd04),
	.w7(32'h3aea2c48),
	.w8(32'hbc6d39b9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31edce),
	.w1(32'hbc0d72e6),
	.w2(32'hbc8bed18),
	.w3(32'hbb39227b),
	.w4(32'hbbec9fb4),
	.w5(32'hbc095970),
	.w6(32'hbac42c0b),
	.w7(32'hbbe6a318),
	.w8(32'hbbf43280),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a43526),
	.w1(32'h3a2f7401),
	.w2(32'h3bf9c806),
	.w3(32'hba6d4a88),
	.w4(32'h3b54a0ef),
	.w5(32'h3b102656),
	.w6(32'hbbcc8bc5),
	.w7(32'h3bf366f3),
	.w8(32'h3b9aeed1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cdeaf),
	.w1(32'h3ab1c42a),
	.w2(32'hbc538217),
	.w3(32'h3b0f1971),
	.w4(32'h3aa0a02d),
	.w5(32'hbbf4e979),
	.w6(32'hbb3b6ca3),
	.w7(32'hbc75d826),
	.w8(32'hbc1a43a2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beaa45f),
	.w1(32'hbb34ed57),
	.w2(32'hbc21fd63),
	.w3(32'hbb1fd9ce),
	.w4(32'h3bb4e34a),
	.w5(32'hbbdfcc80),
	.w6(32'hbc1182e2),
	.w7(32'hbafe02c9),
	.w8(32'hbb38673d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f04a1),
	.w1(32'hbc356707),
	.w2(32'hba3dc671),
	.w3(32'hbca544db),
	.w4(32'h3c40c7e2),
	.w5(32'h3bdd8ce9),
	.w6(32'hbc72cc84),
	.w7(32'h3c10fdc3),
	.w8(32'h3c1a384b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb429),
	.w1(32'hbbb92802),
	.w2(32'hbbde432f),
	.w3(32'hbc0b5031),
	.w4(32'h3b4c0743),
	.w5(32'h3ac3c05c),
	.w6(32'hba348160),
	.w7(32'h3a8ab2f5),
	.w8(32'hbad444a2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39860034),
	.w1(32'h38dc2443),
	.w2(32'h3b478166),
	.w3(32'hbb771496),
	.w4(32'hba177a09),
	.w5(32'hbb59f4ad),
	.w6(32'hbc04ce58),
	.w7(32'hbb2822b0),
	.w8(32'hbc1eb0f1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5983f0),
	.w1(32'h3bbb157d),
	.w2(32'hbc535d8d),
	.w3(32'hbc100f0b),
	.w4(32'h3bfd2a61),
	.w5(32'hbcb58b80),
	.w6(32'h3a4c4328),
	.w7(32'h3c183933),
	.w8(32'hbcc63280),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e2c5f),
	.w1(32'hbc64bd29),
	.w2(32'hbc8658a5),
	.w3(32'hbc450de5),
	.w4(32'hbc5076e4),
	.w5(32'h3bb19c4b),
	.w6(32'hbb3799cb),
	.w7(32'hbc41ff87),
	.w8(32'h3c081548),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf25430),
	.w1(32'h3a82ef96),
	.w2(32'h3ce64d6d),
	.w3(32'h3c7f3dc2),
	.w4(32'hbb627f15),
	.w5(32'hbbafc1f8),
	.w6(32'h3c59304a),
	.w7(32'h3c9ca50a),
	.w8(32'hba697164),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb393a14),
	.w1(32'h3adad9e7),
	.w2(32'h3b696ac4),
	.w3(32'h3b89896f),
	.w4(32'h3b7548fe),
	.w5(32'hba4b41fe),
	.w6(32'h38487ad5),
	.w7(32'h3b015c66),
	.w8(32'h3b31142e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f271ce),
	.w1(32'h3b10030e),
	.w2(32'h3bb6af6a),
	.w3(32'h3a978df1),
	.w4(32'h3bc60742),
	.w5(32'h3b3896e0),
	.w6(32'hbb689669),
	.w7(32'hbb2211f7),
	.w8(32'hbaa90b06),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c0742),
	.w1(32'h39b188ee),
	.w2(32'hbbc28481),
	.w3(32'hbc313ff9),
	.w4(32'h3b22a5fa),
	.w5(32'h3ac85c8a),
	.w6(32'hbc2007b2),
	.w7(32'h3bedcbcd),
	.w8(32'h3b0b2501),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d71ade),
	.w1(32'h3cd9398a),
	.w2(32'h3c6db882),
	.w3(32'h3c2abebc),
	.w4(32'hbb20fc67),
	.w5(32'hbbe2e921),
	.w6(32'h3d0477ae),
	.w7(32'h3c6679b8),
	.w8(32'hbbcc4148),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c4cbc),
	.w1(32'hbbcf1931),
	.w2(32'hbbcc87e9),
	.w3(32'hbc1a13ff),
	.w4(32'hbc076576),
	.w5(32'hbc16398b),
	.w6(32'h3c41c5e9),
	.w7(32'hbc37bc6f),
	.w8(32'hbc58e03b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57465c),
	.w1(32'hbc393666),
	.w2(32'hbc5b37c2),
	.w3(32'hbc9dda5b),
	.w4(32'hbc7f19e6),
	.w5(32'hbbe7322b),
	.w6(32'hbb5409e9),
	.w7(32'hbc67b0f7),
	.w8(32'hb9ced1bb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52814),
	.w1(32'hbc032938),
	.w2(32'hbc360712),
	.w3(32'hbc61e5ec),
	.w4(32'hbc51aae6),
	.w5(32'hbab387c4),
	.w6(32'hbc098000),
	.w7(32'hbc0925e1),
	.w8(32'hbaab9279),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dd6b9),
	.w1(32'hbb314c9e),
	.w2(32'h3af07b74),
	.w3(32'hbaa51e2f),
	.w4(32'h3a8fab96),
	.w5(32'h39fa1018),
	.w6(32'hbb280494),
	.w7(32'h3c2404f8),
	.w8(32'h3af72e50),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2118),
	.w1(32'hb9288fda),
	.w2(32'hbb0e3089),
	.w3(32'hbb9e79d3),
	.w4(32'hbc3e4fcb),
	.w5(32'hbc099b3b),
	.w6(32'h3c4cab25),
	.w7(32'hbc54f529),
	.w8(32'hba070fe0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe94b26),
	.w1(32'h39276151),
	.w2(32'h3c272e91),
	.w3(32'h3bf3e514),
	.w4(32'hbaa380a8),
	.w5(32'h3c8a743b),
	.w6(32'h3cc329d6),
	.w7(32'h3c127948),
	.w8(32'h3c3219a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e57b0),
	.w1(32'h3b7bd8c4),
	.w2(32'h3c943a88),
	.w3(32'hbb7c53f8),
	.w4(32'h3bbce96e),
	.w5(32'h390e9c85),
	.w6(32'hbc503151),
	.w7(32'h3c325aac),
	.w8(32'hbb6af59d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbab91b),
	.w1(32'h3c4cf474),
	.w2(32'hbc41a87b),
	.w3(32'hbc8b73c0),
	.w4(32'h39e87cba),
	.w5(32'h3902dd22),
	.w6(32'hbae41a39),
	.w7(32'h3cba0b01),
	.w8(32'hbc663938),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02dae9),
	.w1(32'h3a071b2d),
	.w2(32'hba6d9c8b),
	.w3(32'h3a2cd9d4),
	.w4(32'hbb82a225),
	.w5(32'hbc5eb81f),
	.w6(32'h3b861efb),
	.w7(32'hbaaf62ff),
	.w8(32'hbc93664a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52f913),
	.w1(32'hbb7124e3),
	.w2(32'h3abaf494),
	.w3(32'hbc11310c),
	.w4(32'hbc7a1af1),
	.w5(32'h3ae8ab9f),
	.w6(32'h3ae41758),
	.w7(32'h3a71e0fb),
	.w8(32'h3b704230),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a437f5b),
	.w1(32'hb8aebc0d),
	.w2(32'h3bab33a8),
	.w3(32'h3ae75b02),
	.w4(32'h3b3278c7),
	.w5(32'h3bf7dd3b),
	.w6(32'hbaad6cb0),
	.w7(32'h3b47597d),
	.w8(32'hbbf92436),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8673d0),
	.w1(32'h3ce73090),
	.w2(32'h3cb523b8),
	.w3(32'h3c6aa8c6),
	.w4(32'h3d06b539),
	.w5(32'h3bb712db),
	.w6(32'h3b9ad493),
	.w7(32'h3cc43ebd),
	.w8(32'h3be0b5f9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14440a),
	.w1(32'h3b7404a8),
	.w2(32'h3acf2828),
	.w3(32'h3b7f5fa8),
	.w4(32'h3b4a8a3c),
	.w5(32'hbaa65c5c),
	.w6(32'hb9d30b8f),
	.w7(32'h3a30b829),
	.w8(32'hbb0c3236),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39a7db),
	.w1(32'hbc083c28),
	.w2(32'h3ab036f1),
	.w3(32'hbbf03563),
	.w4(32'hbad2f20b),
	.w5(32'hbb7df6d9),
	.w6(32'hbc0ba8be),
	.w7(32'h3b8c351e),
	.w8(32'h3b4d9d3b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d565),
	.w1(32'hbaced097),
	.w2(32'hbb2dd697),
	.w3(32'hbc4c8713),
	.w4(32'h3b26d2aa),
	.w5(32'hbb9daade),
	.w6(32'hbae81eac),
	.w7(32'h3a5c3f1b),
	.w8(32'hbba39add),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf8768),
	.w1(32'hbbb44c5a),
	.w2(32'hbba5fbb6),
	.w3(32'hbc117279),
	.w4(32'hbc51f5ef),
	.w5(32'hbb8accf2),
	.w6(32'hbc28b1d1),
	.w7(32'hbbf958a0),
	.w8(32'h3a6b59af),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a8c5),
	.w1(32'h3b74cb51),
	.w2(32'h3b360229),
	.w3(32'hbbe87308),
	.w4(32'h3b361e3c),
	.w5(32'hbb86ae64),
	.w6(32'hbc00db4f),
	.w7(32'h3b6aa61c),
	.w8(32'hbb993db5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf76fd),
	.w1(32'h3b878293),
	.w2(32'h3afed30a),
	.w3(32'h3b9cb17c),
	.w4(32'h3b1195eb),
	.w5(32'hbb99c1d7),
	.w6(32'h3c161780),
	.w7(32'hb9991727),
	.w8(32'hbc5656c2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf78bfb),
	.w1(32'h3c1d8c93),
	.w2(32'h3b40f992),
	.w3(32'h3bea80cf),
	.w4(32'h3c939edc),
	.w5(32'h3b910436),
	.w6(32'hbba4dea0),
	.w7(32'h3be32afe),
	.w8(32'hb9dbb8e5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85853c),
	.w1(32'h3b677ac0),
	.w2(32'hba95e45d),
	.w3(32'h3b8fc9a2),
	.w4(32'h3b0e38dc),
	.w5(32'hbb398470),
	.w6(32'hb8d7926b),
	.w7(32'h39fd6f7a),
	.w8(32'hbb993a46),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ee1e),
	.w1(32'hbb3a6653),
	.w2(32'hbb0ab31e),
	.w3(32'hbba20e5b),
	.w4(32'hbb419f57),
	.w5(32'h3ac994e8),
	.w6(32'hbc2e156a),
	.w7(32'hbb7eb0c6),
	.w8(32'hbc090985),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a151d),
	.w1(32'h3b8d9b2a),
	.w2(32'h3a950916),
	.w3(32'h3c331cf7),
	.w4(32'h3b0b8343),
	.w5(32'h3757b267),
	.w6(32'h3cc9d390),
	.w7(32'h3b1d8ead),
	.w8(32'hbb962e98),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad1142),
	.w1(32'h3c329558),
	.w2(32'h3ad881cc),
	.w3(32'hbb348c1c),
	.w4(32'hbb1f6bba),
	.w5(32'hbc7ab59d),
	.w6(32'hbc0d51d7),
	.w7(32'hbb3fad33),
	.w8(32'hbb9ffd83),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad13ec6),
	.w1(32'h3b3815e5),
	.w2(32'hbbdbd075),
	.w3(32'hba5e892b),
	.w4(32'h3c27d5fd),
	.w5(32'h3b6e6cc4),
	.w6(32'h3cfe6292),
	.w7(32'h3b8afe86),
	.w8(32'hbbd34735),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35ae9c),
	.w1(32'h3c6f1551),
	.w2(32'h3bf451d3),
	.w3(32'h3c73548e),
	.w4(32'h3ccaaa04),
	.w5(32'h3c0a95e7),
	.w6(32'h3ad33d09),
	.w7(32'h3d0671df),
	.w8(32'h3c3e6cf3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd71a7f),
	.w1(32'hbc213eae),
	.w2(32'h3c171977),
	.w3(32'hbca18cf8),
	.w4(32'h3c8dc19a),
	.w5(32'hbc16b5cc),
	.w6(32'hbcd07831),
	.w7(32'h3cbb46ac),
	.w8(32'hbb2b1222),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8701fc),
	.w1(32'h3be25eaf),
	.w2(32'hbaddc5cc),
	.w3(32'h3a8b59b8),
	.w4(32'hbc40897f),
	.w5(32'h3b92aab4),
	.w6(32'h3ccad0d9),
	.w7(32'hbc27286c),
	.w8(32'hbc5b4a6a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c7bab),
	.w1(32'h3c8b7874),
	.w2(32'h3c1cdf26),
	.w3(32'h3c260ed8),
	.w4(32'h3b3085e9),
	.w5(32'hbb8de3eb),
	.w6(32'h3b2941b2),
	.w7(32'hbbe5abaa),
	.w8(32'hbbf12535),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a80aa),
	.w1(32'hbb7452b2),
	.w2(32'hbac85463),
	.w3(32'h3ba8be9a),
	.w4(32'h3bcd5c9d),
	.w5(32'hbad890af),
	.w6(32'h3c88f56f),
	.w7(32'h3b040b12),
	.w8(32'hbb3c9194),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0adf3f),
	.w1(32'hb8dd75d1),
	.w2(32'hbb07d743),
	.w3(32'hbba041da),
	.w4(32'hbac83bd1),
	.w5(32'h39867967),
	.w6(32'hbc1ff21f),
	.w7(32'hbb18a3ef),
	.w8(32'hbc25bbff),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35a84),
	.w1(32'hbc34701e),
	.w2(32'hbb97ab6d),
	.w3(32'hbbc511fc),
	.w4(32'h3ba6475f),
	.w5(32'hbb77736b),
	.w6(32'hbc65b55b),
	.w7(32'hbb7ab1c3),
	.w8(32'hbb26fba9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1052),
	.w1(32'hbba4d9dd),
	.w2(32'hbb95b73f),
	.w3(32'hbaa624d6),
	.w4(32'hbbbb9515),
	.w5(32'hbbf0e3b7),
	.w6(32'hba8c6ab6),
	.w7(32'hbbadd545),
	.w8(32'hbba9b3f8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca2b0),
	.w1(32'hbb17b449),
	.w2(32'h3b387d5d),
	.w3(32'hba9c6ac0),
	.w4(32'hbae7392c),
	.w5(32'hbbfe928a),
	.w6(32'hbc11de2e),
	.w7(32'hbb6e00c1),
	.w8(32'hbbd1cb5e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeebc9),
	.w1(32'hbb348046),
	.w2(32'h39c070e8),
	.w3(32'hbbf33f6b),
	.w4(32'hbc27112d),
	.w5(32'h3bc20204),
	.w6(32'h3aee50a1),
	.w7(32'hbba63a9b),
	.w8(32'h38684f9c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58bd8d),
	.w1(32'h3cb16a55),
	.w2(32'h3cd824df),
	.w3(32'h3caf4f57),
	.w4(32'h3c5ed9ec),
	.w5(32'hbc26c374),
	.w6(32'h3c1e1cfd),
	.w7(32'h3cda37ae),
	.w8(32'hbbf149b9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71ae1c),
	.w1(32'hbc5120c1),
	.w2(32'hbb8ab4fe),
	.w3(32'hbc86712c),
	.w4(32'hbc384e7e),
	.w5(32'h396b4a13),
	.w6(32'h3bcf2a0c),
	.w7(32'hbbe37fb4),
	.w8(32'h3994c1ba),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80cc5c),
	.w1(32'h3ac58acc),
	.w2(32'hbb923336),
	.w3(32'hbb6af65f),
	.w4(32'h3c5236bd),
	.w5(32'hbb41cab9),
	.w6(32'h3bde4edf),
	.w7(32'h3ca9c73d),
	.w8(32'h397497ce),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1c2a4),
	.w1(32'hbc02dc18),
	.w2(32'hbc8b0fa7),
	.w3(32'h3b888285),
	.w4(32'h3b2d1270),
	.w5(32'h3b83ed29),
	.w6(32'h3c1b8f4f),
	.w7(32'h3bc52d29),
	.w8(32'h3b7cc744),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02f98f),
	.w1(32'h3c123561),
	.w2(32'h3c36c9da),
	.w3(32'hbb824dfa),
	.w4(32'h3c19623c),
	.w5(32'h3be92520),
	.w6(32'hbc447208),
	.w7(32'hbb88a2cb),
	.w8(32'hbba4683c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b338c),
	.w1(32'hbcab56c7),
	.w2(32'h3c897624),
	.w3(32'hbcb996cd),
	.w4(32'h3c64cf0d),
	.w5(32'hbbcf0bdb),
	.w6(32'hbc7d807a),
	.w7(32'h3bfa662f),
	.w8(32'hbbe23522),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d7e93),
	.w1(32'hbaa85c83),
	.w2(32'h3ba5210b),
	.w3(32'hbc0b04f7),
	.w4(32'hbb5d7ac5),
	.w5(32'hbc749d00),
	.w6(32'hbcba771d),
	.w7(32'hbb2db4fd),
	.w8(32'hbc624c6b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dec5b),
	.w1(32'hbbd65fdd),
	.w2(32'h3bab30a0),
	.w3(32'hbb4fce6f),
	.w4(32'h3bc768e4),
	.w5(32'h3b52e46b),
	.w6(32'hbc3aabc5),
	.w7(32'h3bae338e),
	.w8(32'h3c11a2e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9e239),
	.w1(32'hbc13c01d),
	.w2(32'h3a9ebc47),
	.w3(32'hbb625a50),
	.w4(32'hbb870153),
	.w5(32'hbba78b9e),
	.w6(32'hbbe52814),
	.w7(32'hbb9f75f7),
	.w8(32'hbac550b2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22271f),
	.w1(32'h3b6826a7),
	.w2(32'hbb1f3514),
	.w3(32'hbaf33172),
	.w4(32'hbc0b231d),
	.w5(32'h3c149d44),
	.w6(32'hbc1e2d47),
	.w7(32'hbc2dc8b9),
	.w8(32'h3bfba9a2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768bc9),
	.w1(32'hba39c615),
	.w2(32'h3b23a823),
	.w3(32'h3bd4908d),
	.w4(32'hb920a21c),
	.w5(32'h3a07844e),
	.w6(32'h3c1e5759),
	.w7(32'h38a08875),
	.w8(32'h3a90e171),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39176c32),
	.w1(32'hbaf864c6),
	.w2(32'hbb6122f2),
	.w3(32'h3ab00879),
	.w4(32'h3a13f8cf),
	.w5(32'hb9478aa9),
	.w6(32'h3c4bd27c),
	.w7(32'h3b0b0d15),
	.w8(32'h38cefc87),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34dd43),
	.w1(32'h3b3a8e6a),
	.w2(32'hbc047bb7),
	.w3(32'h3abfa489),
	.w4(32'hba29e472),
	.w5(32'hba10897b),
	.w6(32'h3bcdff70),
	.w7(32'hbb22416c),
	.w8(32'h3b3b02fc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46c0fe),
	.w1(32'h3c9f5f6a),
	.w2(32'hbb10dc42),
	.w3(32'h3ba6bb2d),
	.w4(32'h3cd92669),
	.w5(32'hbc10dfbb),
	.w6(32'h3c7e5959),
	.w7(32'h3cb48328),
	.w8(32'hbbd4e4ae),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a2b5),
	.w1(32'hbb883148),
	.w2(32'hba3e496a),
	.w3(32'hbc21c73e),
	.w4(32'hbc1cac47),
	.w5(32'hbb955c12),
	.w6(32'h39aabac7),
	.w7(32'hbb2666ad),
	.w8(32'hb993d1ad),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b572d67),
	.w1(32'hbbc45684),
	.w2(32'hbb477da0),
	.w3(32'h3af1d848),
	.w4(32'hbb4e19f7),
	.w5(32'h3b22c566),
	.w6(32'hbb910263),
	.w7(32'hbc02d911),
	.w8(32'hba651758),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39507d2d),
	.w1(32'h3b2bfbb9),
	.w2(32'hba727c97),
	.w3(32'h3b8a5fa5),
	.w4(32'h3b5f610c),
	.w5(32'hba1f801a),
	.w6(32'h3bbe5bac),
	.w7(32'h3bb72824),
	.w8(32'hbb9c46e7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae56941),
	.w1(32'hba94ef34),
	.w2(32'h3b91e53b),
	.w3(32'hbc280695),
	.w4(32'h3befefcc),
	.w5(32'h3bc21ad9),
	.w6(32'hbc47edea),
	.w7(32'h3be7f4c1),
	.w8(32'h3c03b3a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c69d99),
	.w1(32'h3b87c54b),
	.w2(32'hbbe28970),
	.w3(32'hba9c5bc2),
	.w4(32'h3b1aa9e9),
	.w5(32'hbb9fcdef),
	.w6(32'hbb69dc7b),
	.w7(32'hbb7fdf01),
	.w8(32'hbb641557),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad48478),
	.w1(32'hbbb83a6e),
	.w2(32'hbbec174a),
	.w3(32'hbc32f96f),
	.w4(32'hbbfb10c9),
	.w5(32'hba6b1436),
	.w6(32'h3c0f4a55),
	.w7(32'hbb4735e4),
	.w8(32'h3b281893),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab97500),
	.w1(32'hbba3bb4e),
	.w2(32'hbaae88f7),
	.w3(32'hbb4298cb),
	.w4(32'hbc04ff67),
	.w5(32'h3c0e0f5b),
	.w6(32'h3c568136),
	.w7(32'hbc0031c3),
	.w8(32'h3bc59678),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa86e3),
	.w1(32'h3aa85650),
	.w2(32'hbb1c4fb3),
	.w3(32'hbbc86579),
	.w4(32'hbb7ecb18),
	.w5(32'hbbff9ddb),
	.w6(32'h3b2f66b1),
	.w7(32'h3a2fc58a),
	.w8(32'hb5ed1953),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc380c),
	.w1(32'hbc412511),
	.w2(32'hbc041cef),
	.w3(32'hbafbb60d),
	.w4(32'hbad6e359),
	.w5(32'h3bba0ed0),
	.w6(32'h3bfa00ed),
	.w7(32'h3b0274ea),
	.w8(32'h3c7d7fbb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d85c5),
	.w1(32'hbc8873b5),
	.w2(32'h3b196bf1),
	.w3(32'hbc941b42),
	.w4(32'hbc0d0d57),
	.w5(32'hbbd2584c),
	.w6(32'hbc77e6e5),
	.w7(32'hba305b6b),
	.w8(32'hbbd7a3d8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc781ff6),
	.w1(32'hbc093a43),
	.w2(32'hbc1fc8d6),
	.w3(32'hbc177fea),
	.w4(32'hb9e06ce6),
	.w5(32'h3aed8257),
	.w6(32'hbbb532d2),
	.w7(32'h3b579056),
	.w8(32'h3a6c0703),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b379301),
	.w1(32'h3b485c6f),
	.w2(32'h3b8009bc),
	.w3(32'hbb22ca4d),
	.w4(32'hbb6be3a7),
	.w5(32'h3c218592),
	.w6(32'hbb8f4409),
	.w7(32'hbb5644ab),
	.w8(32'h3b8fcbda),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb930b9),
	.w1(32'h3cc77011),
	.w2(32'hbc5270c6),
	.w3(32'h3cdca0df),
	.w4(32'hb9887ea1),
	.w5(32'hbbc8824c),
	.w6(32'h3cfcd1a4),
	.w7(32'hbc614fe8),
	.w8(32'hbc357fe1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bad95),
	.w1(32'hb9755fa5),
	.w2(32'hbbf99391),
	.w3(32'hba8c7074),
	.w4(32'h3ab72555),
	.w5(32'h3ba681a7),
	.w6(32'h3b6f3d09),
	.w7(32'h3b0a87eb),
	.w8(32'h3c8021e1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6812be),
	.w1(32'h3c11d201),
	.w2(32'hbbf228fd),
	.w3(32'h3c6488b2),
	.w4(32'h3c16e74a),
	.w5(32'hbc150d92),
	.w6(32'h3cc50038),
	.w7(32'hb8ebe080),
	.w8(32'hbc837e97),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa82a2),
	.w1(32'hbb326161),
	.w2(32'h3a28fbb7),
	.w3(32'hbc48d217),
	.w4(32'hbb812be0),
	.w5(32'h3b3832fe),
	.w6(32'hbbf08dd7),
	.w7(32'h3b92048e),
	.w8(32'h3b6029ca),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28731a),
	.w1(32'h3c691c46),
	.w2(32'hbc68a4b8),
	.w3(32'h3c84f6fa),
	.w4(32'hbc425c6d),
	.w5(32'hbc4a47ac),
	.w6(32'h3cbfa03f),
	.w7(32'hbc4b8827),
	.w8(32'hbc742c8e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4972f),
	.w1(32'hbbf45955),
	.w2(32'hbc2686c8),
	.w3(32'hbadab142),
	.w4(32'hbc154cbd),
	.w5(32'hbc019b0e),
	.w6(32'hba7d7138),
	.w7(32'hbbd51864),
	.w8(32'hbc3d224a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac381e1),
	.w1(32'hbbf04bfc),
	.w2(32'hbba34fe9),
	.w3(32'hbb8a5b28),
	.w4(32'h3b52f87f),
	.w5(32'h39bd7aad),
	.w6(32'hbbc25837),
	.w7(32'hba493839),
	.w8(32'hbb3fa1ba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29d563),
	.w1(32'hbba1c8c3),
	.w2(32'hbb245437),
	.w3(32'h3a0733eb),
	.w4(32'hbba33925),
	.w5(32'hbbfd8f39),
	.w6(32'hbc74d102),
	.w7(32'hbb957f26),
	.w8(32'hbb8c2021),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43f38),
	.w1(32'hbb32358a),
	.w2(32'hbcb973e7),
	.w3(32'h3baea9da),
	.w4(32'hbc3d11b6),
	.w5(32'hbb59fec1),
	.w6(32'h3ab84b27),
	.w7(32'hbc8df9a3),
	.w8(32'hbbb0a880),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952984),
	.w1(32'h393f9d1c),
	.w2(32'hbc127ff0),
	.w3(32'hba317be8),
	.w4(32'h3afc9423),
	.w5(32'hba1dc36b),
	.w6(32'h3b9b0d6c),
	.w7(32'h3c1228db),
	.w8(32'hbb049d1f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d98e),
	.w1(32'h3c7945ae),
	.w2(32'hbbc50509),
	.w3(32'hbc692325),
	.w4(32'hbb31c969),
	.w5(32'hbbc7ff16),
	.w6(32'hbc4eff44),
	.w7(32'hbc3688c7),
	.w8(32'hbc8a308e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ab96),
	.w1(32'h3b8309d4),
	.w2(32'hbab2cd9c),
	.w3(32'hbbaa6c9d),
	.w4(32'h38a4a9c1),
	.w5(32'hbb8123ca),
	.w6(32'h3b0751be),
	.w7(32'h3b37602b),
	.w8(32'hbbb66a0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14eaca),
	.w1(32'h3b2dd4f0),
	.w2(32'hb946e4f9),
	.w3(32'hbb8b477f),
	.w4(32'hbb892d88),
	.w5(32'hbb893ff3),
	.w6(32'hba30430e),
	.w7(32'hbb3aa476),
	.w8(32'hbb729e4d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79bd74),
	.w1(32'h3baab7a2),
	.w2(32'hbc5fbe81),
	.w3(32'hbbf57022),
	.w4(32'h3aa1a820),
	.w5(32'hbb287e9e),
	.w6(32'hbb13cf39),
	.w7(32'h3b2d832e),
	.w8(32'hbbc24f84),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77dd0e),
	.w1(32'h3aa78ee1),
	.w2(32'h3a1405e8),
	.w3(32'h39fc7c36),
	.w4(32'h3a755704),
	.w5(32'hba59c7fa),
	.w6(32'h3ad1192e),
	.w7(32'h3a9d08ef),
	.w8(32'hbb34f905),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe25d72),
	.w1(32'h3a2969fa),
	.w2(32'hbc2cc34c),
	.w3(32'hbb161e34),
	.w4(32'hbbb23bd6),
	.w5(32'hbc0d2fce),
	.w6(32'hbc3d7f87),
	.w7(32'hbb83b5fc),
	.w8(32'hbc0b0a81),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846e42),
	.w1(32'h3a2ce187),
	.w2(32'h3a0eb1d6),
	.w3(32'hbab57449),
	.w4(32'h3ab8b38d),
	.w5(32'h3b158807),
	.w6(32'hbb03908d),
	.w7(32'h3b48f2e1),
	.w8(32'h3b01117d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba591e18),
	.w1(32'h3a8f8551),
	.w2(32'h38ed475b),
	.w3(32'hba0be754),
	.w4(32'hb9cf2f18),
	.w5(32'h399c4117),
	.w6(32'hba6f517d),
	.w7(32'hb9fb57d0),
	.w8(32'h374fa601),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f06f),
	.w1(32'h3b269b39),
	.w2(32'h3a47582b),
	.w3(32'h39d05962),
	.w4(32'hba55ef09),
	.w5(32'hbb96e64c),
	.w6(32'h3b116a9c),
	.w7(32'h39fb5457),
	.w8(32'hbb45d2b6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ceaf),
	.w1(32'h39c40f81),
	.w2(32'hbb28dfed),
	.w3(32'hb9fd8a3f),
	.w4(32'h3b939e7c),
	.w5(32'hbb608b75),
	.w6(32'hbb2584a3),
	.w7(32'h3a975ec6),
	.w8(32'hbbab1927),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0dfa),
	.w1(32'hba626c76),
	.w2(32'hbaa9457a),
	.w3(32'hbb4f8d6f),
	.w4(32'hbb2fb221),
	.w5(32'hbb15388b),
	.w6(32'hbad60c18),
	.w7(32'hbad93c97),
	.w8(32'hbb3acee1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208748),
	.w1(32'hbb0ba54b),
	.w2(32'h3a3d4095),
	.w3(32'hbab62f60),
	.w4(32'hbad2c953),
	.w5(32'hba845eac),
	.w6(32'hb960e08c),
	.w7(32'h3b020a47),
	.w8(32'h39b3b4be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d56bc3),
	.w1(32'hb9b4b521),
	.w2(32'h364ff43e),
	.w3(32'hba4aff8b),
	.w4(32'hbaeb0246),
	.w5(32'hbb89a128),
	.w6(32'h3ac295a3),
	.w7(32'h370786d6),
	.w8(32'hbba34b5a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed819e),
	.w1(32'h3bc3323a),
	.w2(32'h3ae1d77e),
	.w3(32'hbb8f4817),
	.w4(32'h3a8d6d10),
	.w5(32'hbb23c3e5),
	.w6(32'hbc054e1a),
	.w7(32'hbbf3e102),
	.w8(32'hbbf0fb8f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95bcf6),
	.w1(32'hbb0d6594),
	.w2(32'hbc10da93),
	.w3(32'hba99d0d0),
	.w4(32'hbb244818),
	.w5(32'hbbc0932d),
	.w6(32'hbb978801),
	.w7(32'hbb11ce59),
	.w8(32'hbbb20105),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939fb94),
	.w1(32'h3ad98ce5),
	.w2(32'hba836d58),
	.w3(32'h3a28243a),
	.w4(32'hbb09ac86),
	.w5(32'hbb01ff05),
	.w6(32'h3ae4dfc7),
	.w7(32'hbaf70f90),
	.w8(32'hbb142e23),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921aedb),
	.w1(32'h3a821c9b),
	.w2(32'h3a5f27fd),
	.w3(32'h39bb4551),
	.w4(32'h38018079),
	.w5(32'hba6e7f59),
	.w6(32'h39a6fbef),
	.w7(32'h39a1d090),
	.w8(32'hba141dbc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9923a8),
	.w1(32'hbb0f59d4),
	.w2(32'hbb0cd14a),
	.w3(32'hbab61771),
	.w4(32'hba85c6a5),
	.w5(32'hbb090f27),
	.w6(32'hbabb454d),
	.w7(32'hba867b8e),
	.w8(32'hbb66cbf9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b6e92),
	.w1(32'hba32a18d),
	.w2(32'h3a910d18),
	.w3(32'h3ac07e29),
	.w4(32'hb9855381),
	.w5(32'hbab8b68c),
	.w6(32'h3a27b961),
	.w7(32'hb99bacae),
	.w8(32'hba2a1732),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca21a9),
	.w1(32'hb9429d8b),
	.w2(32'hba632944),
	.w3(32'hba88ca26),
	.w4(32'hb9d8a5e0),
	.w5(32'h39ebb52d),
	.w6(32'hb9f2825f),
	.w7(32'hbada07e0),
	.w8(32'h3ad136fe),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919589f),
	.w1(32'hbaf73a9e),
	.w2(32'hba0d9b26),
	.w3(32'hbb33aa34),
	.w4(32'h39ff5572),
	.w5(32'hbb42a241),
	.w6(32'hbad6bf57),
	.w7(32'h3a2dd767),
	.w8(32'hbaf1ca1a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c01ae),
	.w1(32'h3a323e39),
	.w2(32'h3a1163e1),
	.w3(32'h3a09d962),
	.w4(32'h3a60587a),
	.w5(32'hba49e074),
	.w6(32'h3a15ccff),
	.w7(32'h3a0797af),
	.w8(32'hba93c8d7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf7abd),
	.w1(32'h3b063aef),
	.w2(32'hbb00bdc2),
	.w3(32'h3a0fa1ce),
	.w4(32'h3b798401),
	.w5(32'h3accc39a),
	.w6(32'h3a0850ab),
	.w7(32'h3ae76286),
	.w8(32'hba511fbf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b032c3),
	.w1(32'hbb6a316a),
	.w2(32'hbb08792d),
	.w3(32'hba92ca30),
	.w4(32'hbc1a55bd),
	.w5(32'hbc0b4734),
	.w6(32'h3b39c819),
	.w7(32'hbb76b3c8),
	.w8(32'hbbf3135d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f15d4),
	.w1(32'hba58ba99),
	.w2(32'hbaa12462),
	.w3(32'hba0c8738),
	.w4(32'h3a93a6f9),
	.w5(32'hb9634495),
	.w6(32'hbaa5a766),
	.w7(32'h3a587ec0),
	.w8(32'h3a638c09),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81fbd6),
	.w1(32'h39810da9),
	.w2(32'h3973b0b4),
	.w3(32'h3a0b13a1),
	.w4(32'hb91aef4e),
	.w5(32'hb9a8129f),
	.w6(32'h3a00edb3),
	.w7(32'hb8260730),
	.w8(32'hba435736),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea406e),
	.w1(32'hb97c2322),
	.w2(32'h39f914a2),
	.w3(32'hba3982e0),
	.w4(32'hba6e8479),
	.w5(32'hba88ba83),
	.w6(32'hba3ad2be),
	.w7(32'hb9cce408),
	.w8(32'hba44aefb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d2848),
	.w1(32'hbaf9d39d),
	.w2(32'hbaca0278),
	.w3(32'hba7b27e6),
	.w4(32'hb9c22ef8),
	.w5(32'h396d0dba),
	.w6(32'hba6588f5),
	.w7(32'hba6af463),
	.w8(32'h39336014),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a6aa),
	.w1(32'h3c8e7881),
	.w2(32'h3b847b9a),
	.w3(32'h3b1bc017),
	.w4(32'h3bc56be1),
	.w5(32'hbb95039a),
	.w6(32'hbc0ec5d6),
	.w7(32'hbb237c45),
	.w8(32'hbc2b69c2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39065a8b),
	.w1(32'h3ab10775),
	.w2(32'hbbb72b18),
	.w3(32'h3b093039),
	.w4(32'h3ba598c6),
	.w5(32'hbb771e32),
	.w6(32'hbb21f708),
	.w7(32'h3a57b8e3),
	.w8(32'hbbc282f6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cce250),
	.w1(32'hbaa84c5a),
	.w2(32'hbb85163b),
	.w3(32'hb818c34f),
	.w4(32'hbaa50724),
	.w5(32'hbabaf4fe),
	.w6(32'h3aac2ba4),
	.w7(32'hb9c58b66),
	.w8(32'hbaabb885),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af73172),
	.w1(32'h3b17c23b),
	.w2(32'hba245db5),
	.w3(32'hbb3d1dd6),
	.w4(32'h39f30d8a),
	.w5(32'hbaa3e7a7),
	.w6(32'hbadfa4d8),
	.w7(32'hbb4411ae),
	.w8(32'hbb4f6bf8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51d40c),
	.w1(32'hb92966e0),
	.w2(32'hba5f6f80),
	.w3(32'hb9430f9d),
	.w4(32'h38d2f3d0),
	.w5(32'hb9c86105),
	.w6(32'hb99919dc),
	.w7(32'h3a2e8c95),
	.w8(32'hbb7a7e6d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c9b43e),
	.w1(32'h39e5f097),
	.w2(32'hba7321ed),
	.w3(32'hb9e5be5e),
	.w4(32'h3a0429fc),
	.w5(32'hbb4a030d),
	.w6(32'hbb35c841),
	.w7(32'hbb3c6547),
	.w8(32'hbb9fe1f2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37b6b),
	.w1(32'hba7c1f36),
	.w2(32'hba9f1af4),
	.w3(32'hbac759db),
	.w4(32'hbacea6e0),
	.w5(32'hbb76e00a),
	.w6(32'h39a2d1af),
	.w7(32'h398ba879),
	.w8(32'hbb0106a7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2094da),
	.w1(32'h3b885172),
	.w2(32'hbc093d70),
	.w3(32'h3b8c8897),
	.w4(32'h3be93edb),
	.w5(32'h39f202ed),
	.w6(32'h3a5e2aad),
	.w7(32'h3ba8762e),
	.w8(32'hbb6e94cb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39693ea1),
	.w1(32'h3afbb7a9),
	.w2(32'h3a844f9f),
	.w3(32'h399f4608),
	.w4(32'hbb482d9b),
	.w5(32'hbb87c2e4),
	.w6(32'h3b3a9b61),
	.w7(32'hbaf1dd33),
	.w8(32'hbba4b9bc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a680bc1),
	.w1(32'hba457028),
	.w2(32'hbba0c0bc),
	.w3(32'h39325c56),
	.w4(32'hba2d6564),
	.w5(32'hbba002ba),
	.w6(32'hba1172b5),
	.w7(32'hba348229),
	.w8(32'hbbbf3404),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f861a),
	.w1(32'h3b39b650),
	.w2(32'hbbadf561),
	.w3(32'hb7ca097a),
	.w4(32'h3b8fa645),
	.w5(32'hb9b538a0),
	.w6(32'hba15937f),
	.w7(32'h3aa7d603),
	.w8(32'hbb57cf9a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b84939),
	.w1(32'h3b4a17f4),
	.w2(32'h3a9be7da),
	.w3(32'hbb274278),
	.w4(32'hbb249913),
	.w5(32'hbb36f9e2),
	.w6(32'hb8e897dd),
	.w7(32'hbb23764e),
	.w8(32'hbb8828c5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d43763),
	.w1(32'h3968c03b),
	.w2(32'hbb6b9759),
	.w3(32'h3ab1e2bf),
	.w4(32'h3b27753f),
	.w5(32'hbb086d5a),
	.w6(32'h3aeac6d5),
	.w7(32'h3b03e37c),
	.w8(32'hbb5bb31a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a427a0e),
	.w1(32'h3a341316),
	.w2(32'hb9c0cfc9),
	.w3(32'h3839f5b4),
	.w4(32'h3a50a090),
	.w5(32'hb9bbcee0),
	.w6(32'hba73182e),
	.w7(32'h3a5b4c5d),
	.w8(32'hbaf5e65f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c2cf8),
	.w1(32'h3ac78534),
	.w2(32'hbb5c05d1),
	.w3(32'h38a6e8c6),
	.w4(32'hbb25149c),
	.w5(32'hbb354548),
	.w6(32'h39ad243d),
	.w7(32'hbaaeb595),
	.w8(32'hbba2e724),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5925f),
	.w1(32'h3a4fc9e8),
	.w2(32'h3aa62476),
	.w3(32'h3a8f3e1f),
	.w4(32'h3a82ea59),
	.w5(32'hba243cd1),
	.w6(32'hba08e36f),
	.w7(32'hb9d77116),
	.w8(32'hbb3ba75a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de4f5),
	.w1(32'hb88f09a1),
	.w2(32'h394c5940),
	.w3(32'h3a2a87d8),
	.w4(32'h38f8e0d2),
	.w5(32'hba257a04),
	.w6(32'hb96f36ed),
	.w7(32'h3819832e),
	.w8(32'hbae512a1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63aab1),
	.w1(32'hbad21506),
	.w2(32'hbad63a7e),
	.w3(32'h3989c75b),
	.w4(32'hba06c14b),
	.w5(32'hba2d6c3a),
	.w6(32'hb9bc3a6b),
	.w7(32'hba84e297),
	.w8(32'hba8676ca),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f1b5d),
	.w1(32'hb9404cdf),
	.w2(32'hba92e5b8),
	.w3(32'h39203e1e),
	.w4(32'hba5b023f),
	.w5(32'hb9d52733),
	.w6(32'h3903fb8b),
	.w7(32'hba96fda8),
	.w8(32'hba474bb1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf6aab),
	.w1(32'h3a4d9d15),
	.w2(32'hbac615e9),
	.w3(32'hbb3e8698),
	.w4(32'hbb00a726),
	.w5(32'hbb26af06),
	.w6(32'h3a7e3f22),
	.w7(32'hb92a4f45),
	.w8(32'hbb892870),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92b141),
	.w1(32'h3970ea51),
	.w2(32'hba9d97b2),
	.w3(32'h3a8713bd),
	.w4(32'h3ad81a48),
	.w5(32'hbad4cf79),
	.w6(32'hbac7629f),
	.w7(32'hb8bf1f8e),
	.w8(32'hbb6654a0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950b146),
	.w1(32'hb786df6b),
	.w2(32'hb6f0bbc0),
	.w3(32'h39aa9755),
	.w4(32'h39ef4444),
	.w5(32'h39d84125),
	.w6(32'hba456359),
	.w7(32'h39b21d40),
	.w8(32'h3a6c8a42),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a043c94),
	.w1(32'hb90f3fbc),
	.w2(32'hbba80113),
	.w3(32'h3a4a12be),
	.w4(32'h3b475b9e),
	.w5(32'hbac5055c),
	.w6(32'hba5798b9),
	.w7(32'h3acc5fbd),
	.w8(32'hbaf2ad8f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a100ec5),
	.w1(32'h39e12bcf),
	.w2(32'hb9aa7393),
	.w3(32'hba2672a2),
	.w4(32'h3980f756),
	.w5(32'hba3555ff),
	.w6(32'hba58b755),
	.w7(32'hb9bb44d4),
	.w8(32'hbb337bb8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3172b7),
	.w1(32'h3b5e92e0),
	.w2(32'hbbe4c86f),
	.w3(32'h3b141aab),
	.w4(32'h3b6d6dd2),
	.w5(32'hb9ae4c0a),
	.w6(32'h3a8d8f58),
	.w7(32'h3b0e0a2d),
	.w8(32'hbb4ece1a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc551ab),
	.w1(32'hb9e5df7e),
	.w2(32'h3ab23358),
	.w3(32'hbc0598a4),
	.w4(32'hbbc9b7fb),
	.w5(32'hbbc96635),
	.w6(32'hbb6e8f39),
	.w7(32'h3b3def42),
	.w8(32'hbb5c7d02),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817a0a),
	.w1(32'hbb343949),
	.w2(32'hbaa6b0fb),
	.w3(32'hba9229ef),
	.w4(32'hbb37a914),
	.w5(32'hbb850341),
	.w6(32'hb95d99b7),
	.w7(32'hbaed00da),
	.w8(32'hbbaa1498),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba378cf5),
	.w1(32'hbaa24f58),
	.w2(32'h38dd9f34),
	.w3(32'hba8501f1),
	.w4(32'h3a0713c0),
	.w5(32'hbb5aa527),
	.w6(32'hba95f621),
	.w7(32'hb9c584ae),
	.w8(32'hbb4ef332),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c49d6),
	.w1(32'hbabf3af3),
	.w2(32'hbb0ef875),
	.w3(32'hbb91337c),
	.w4(32'hbb1d80a9),
	.w5(32'hbb31ac53),
	.w6(32'hbb6489e8),
	.w7(32'hbaf0aa70),
	.w8(32'hbad48af7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9965c94),
	.w1(32'hb9db69e6),
	.w2(32'hba8bb2e4),
	.w3(32'hbafca761),
	.w4(32'hbb2a9391),
	.w5(32'hbb823685),
	.w6(32'hba3b9912),
	.w7(32'h38777797),
	.w8(32'hbb5b8f12),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237df6),
	.w1(32'hba9d5d03),
	.w2(32'hba4a4b69),
	.w3(32'hbafa16db),
	.w4(32'hbb081f5e),
	.w5(32'hbb26539c),
	.w6(32'h3824a83e),
	.w7(32'hb9818440),
	.w8(32'hbad1f5a7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9089c85),
	.w1(32'h3ac8d157),
	.w2(32'hbaa127d3),
	.w3(32'h3a3ea59f),
	.w4(32'h39e69268),
	.w5(32'h3a802db9),
	.w6(32'h366b6d18),
	.w7(32'hba87f01c),
	.w8(32'hba83189e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80ad09),
	.w1(32'hbac4475c),
	.w2(32'h3a1a9b37),
	.w3(32'h3ab520f3),
	.w4(32'hba27f743),
	.w5(32'hbabe94fe),
	.w6(32'h3b1dbeea),
	.w7(32'h3b01f6f0),
	.w8(32'hba9c65d5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb937),
	.w1(32'h3b9e7410),
	.w2(32'hbb32c8ef),
	.w3(32'h3ae3dc94),
	.w4(32'h3b962f76),
	.w5(32'hbab6df59),
	.w6(32'h3a70e143),
	.w7(32'h3b2d5dcc),
	.w8(32'hbb97be0a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62ce56),
	.w1(32'h3aa7f1b4),
	.w2(32'hba9a54bd),
	.w3(32'h3b1399d4),
	.w4(32'h3b1ba1ba),
	.w5(32'h3998e2c3),
	.w6(32'h3a993cff),
	.w7(32'h3a9e8284),
	.w8(32'h3a45a243),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba655570),
	.w1(32'hba0512bf),
	.w2(32'h3b4e5ac2),
	.w3(32'hbb42b78a),
	.w4(32'hbaebcff2),
	.w5(32'hbb44e1ab),
	.w6(32'hbb618980),
	.w7(32'hbb248d2a),
	.w8(32'hbacf31ff),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9a3c2),
	.w1(32'hb9d62180),
	.w2(32'hba14502d),
	.w3(32'hb9a0beb7),
	.w4(32'hb8e30a3a),
	.w5(32'hb96884f8),
	.w6(32'hb9efe720),
	.w7(32'hba211c40),
	.w8(32'h39164f35),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c7f9),
	.w1(32'h3b31e087),
	.w2(32'hba4720f8),
	.w3(32'h3b5eba79),
	.w4(32'h3b90b5ef),
	.w5(32'hb989ba42),
	.w6(32'h39cfa030),
	.w7(32'hb9ada245),
	.w8(32'hbb92d969),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2ff0f),
	.w1(32'hbb1dd813),
	.w2(32'h39bfae25),
	.w3(32'hbb43e65f),
	.w4(32'hbab53a51),
	.w5(32'h3949d46e),
	.w6(32'hbaeb1d0d),
	.w7(32'hba332ecf),
	.w8(32'h37eb22fe),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d82a5f),
	.w1(32'hb9ae5505),
	.w2(32'hbac37285),
	.w3(32'hb96d785a),
	.w4(32'h3a6b0fe6),
	.w5(32'hbacf5fdd),
	.w6(32'hba330e50),
	.w7(32'hba6719ae),
	.w8(32'hbaa0d12b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dcc55),
	.w1(32'hba8b542b),
	.w2(32'hba9435f2),
	.w3(32'hb9bd9f29),
	.w4(32'hbb3386d7),
	.w5(32'hbb0a4d70),
	.w6(32'h3a43a914),
	.w7(32'hbac3d2ab),
	.w8(32'hbb194d34),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f6a92),
	.w1(32'h3c092ac6),
	.w2(32'hbae6c036),
	.w3(32'h39a2dc26),
	.w4(32'h3ba5e225),
	.w5(32'hb953d538),
	.w6(32'hbbb6ac76),
	.w7(32'hbb41cc24),
	.w8(32'hbbbb1a45),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad99877),
	.w1(32'hbb078079),
	.w2(32'hbabeb98e),
	.w3(32'hbabc7100),
	.w4(32'hb88cd617),
	.w5(32'h3a591c0c),
	.w6(32'hba20b2bb),
	.w7(32'hb98dadc2),
	.w8(32'h3a6d4529),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5287d9),
	.w1(32'h3a550b65),
	.w2(32'h3b574347),
	.w3(32'hbae59f0b),
	.w4(32'hbb2c36a8),
	.w5(32'hbb2b4bd0),
	.w6(32'h3a2e71bb),
	.w7(32'h39e42cfe),
	.w8(32'hbb9aece4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad412a5),
	.w1(32'h38be8b41),
	.w2(32'h3a9551f0),
	.w3(32'hbb176fe7),
	.w4(32'hba4a3516),
	.w5(32'hba3bab38),
	.w6(32'hbb2719e1),
	.w7(32'hb7f1c3f0),
	.w8(32'h3a48cfd5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad5e06),
	.w1(32'hbb5f963a),
	.w2(32'hbb5b4296),
	.w3(32'hbb7d367d),
	.w4(32'hba68e3a0),
	.w5(32'hbaaf1462),
	.w6(32'hbbbfd6c3),
	.w7(32'hb99228f9),
	.w8(32'hbabe2113),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5baa6),
	.w1(32'h3ad19318),
	.w2(32'hba9a6fdd),
	.w3(32'h3b0a5c61),
	.w4(32'hba0d807f),
	.w5(32'hbb2073a1),
	.w6(32'h3b68d3d5),
	.w7(32'h39b93c30),
	.w8(32'hbb7a34f4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70fe53),
	.w1(32'h3a075386),
	.w2(32'hbb416214),
	.w3(32'h3a2257ad),
	.w4(32'h3b870c4e),
	.w5(32'hbab97f71),
	.w6(32'hbb006840),
	.w7(32'h3a728c1b),
	.w8(32'hbb44124d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33a191),
	.w1(32'h3983863f),
	.w2(32'h399cad82),
	.w3(32'h394a7886),
	.w4(32'h3a60fa53),
	.w5(32'hba6ec687),
	.w6(32'h39ed3963),
	.w7(32'h39dd7699),
	.w8(32'hb9892008),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaada3b),
	.w1(32'hbad6a107),
	.w2(32'hbb4f4716),
	.w3(32'hbb0f5d48),
	.w4(32'hbb0dbd05),
	.w5(32'hbb5b6bb0),
	.w6(32'hbb5322b3),
	.w7(32'hbaf2b874),
	.w8(32'hbb2b18bb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d275b),
	.w1(32'hbaa2edfc),
	.w2(32'hb9a6124b),
	.w3(32'hba7994bf),
	.w4(32'h3a0bd4ae),
	.w5(32'hbab4fb2c),
	.w6(32'hb9d698a0),
	.w7(32'hb6d5fa55),
	.w8(32'hbac2b541),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad93334),
	.w1(32'h3a062a76),
	.w2(32'h39a99aec),
	.w3(32'h3ad4b697),
	.w4(32'h3a285495),
	.w5(32'h3a435f2d),
	.w6(32'h39f39207),
	.w7(32'h3a98561f),
	.w8(32'hba3aa48d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821cc8),
	.w1(32'h3a0ad63a),
	.w2(32'hb9a0ef80),
	.w3(32'h3a77b5dc),
	.w4(32'hbaae0316),
	.w5(32'hba72313b),
	.w6(32'h3a49de51),
	.w7(32'hbaa6ed28),
	.w8(32'hba8f8f1d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b358460),
	.w1(32'hbabe6cef),
	.w2(32'hbba07e68),
	.w3(32'hb932abdc),
	.w4(32'hbb4461c7),
	.w5(32'hbbc189e9),
	.w6(32'hbab8ff15),
	.w7(32'hba5159d3),
	.w8(32'hbbed87aa),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dbe39),
	.w1(32'hbb27eec8),
	.w2(32'hb9a5e1ae),
	.w3(32'h39a0aa2e),
	.w4(32'h3a36090e),
	.w5(32'h3949d688),
	.w6(32'hbac16f01),
	.w7(32'h3a151148),
	.w8(32'hb995ae58),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c1e77),
	.w1(32'hba3c22ae),
	.w2(32'hb91f6769),
	.w3(32'h3903efe0),
	.w4(32'hba9d2f4e),
	.w5(32'hba63e2f3),
	.w6(32'hb6a86760),
	.w7(32'hba5da195),
	.w8(32'hba1b9f4a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f781),
	.w1(32'h3a43d944),
	.w2(32'hb94b4558),
	.w3(32'hbafca496),
	.w4(32'hbb0c0085),
	.w5(32'hbb36160c),
	.w6(32'hbac9910a),
	.w7(32'hbb453099),
	.w8(32'hbb1a45da),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80e7a),
	.w1(32'h389f8882),
	.w2(32'hbc1b1617),
	.w3(32'hbbd0ad64),
	.w4(32'hbb1f3d66),
	.w5(32'hbbcf2b30),
	.w6(32'hb8a7d1e8),
	.w7(32'h38f841e0),
	.w8(32'hbbffd001),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e8822),
	.w1(32'h3b935e29),
	.w2(32'hbb7ed971),
	.w3(32'hbb979ac2),
	.w4(32'h398a9d9f),
	.w5(32'h3b2a669f),
	.w6(32'hbb39875c),
	.w7(32'h3a56f028),
	.w8(32'h38df32e7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b3c3),
	.w1(32'hbb026070),
	.w2(32'hba4e49e1),
	.w3(32'hba5cd433),
	.w4(32'h395514cf),
	.w5(32'h3a3f3431),
	.w6(32'hba5aa0a0),
	.w7(32'hb70e4e7c),
	.w8(32'h3a8005ff),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a9e3b),
	.w1(32'h3b9bb158),
	.w2(32'hbb5e977b),
	.w3(32'h3b976d04),
	.w4(32'h3c156ad0),
	.w5(32'hbb197378),
	.w6(32'hbb2de735),
	.w7(32'h3987d407),
	.w8(32'hbc0e8961),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d55d5),
	.w1(32'hbbbabf19),
	.w2(32'h3ad63cfc),
	.w3(32'hbad8dd24),
	.w4(32'hbaeb71a5),
	.w5(32'hbba5f080),
	.w6(32'hb9b5d200),
	.w7(32'h3b8ad92a),
	.w8(32'hbb565aa4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11f98d),
	.w1(32'h3b06e595),
	.w2(32'hbadf7719),
	.w3(32'h3a6e1ba0),
	.w4(32'h3b3a78a8),
	.w5(32'h39dbcbfd),
	.w6(32'h3a7ae897),
	.w7(32'h3b07005f),
	.w8(32'h38e533bf),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71a89f4),
	.w1(32'h38e74210),
	.w2(32'h39a0abde),
	.w3(32'hba3ce885),
	.w4(32'hb99e4092),
	.w5(32'hba2bf633),
	.w6(32'hbaceeee8),
	.w7(32'hbaa95302),
	.w8(32'hb9b5514b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377c4cee),
	.w1(32'h38d0fc1a),
	.w2(32'hb89e6d7c),
	.w3(32'hba3d0abe),
	.w4(32'h39d8ce7a),
	.w5(32'hb97fd4ec),
	.w6(32'hbace4f5f),
	.w7(32'hb9c4f98b),
	.w8(32'hba8bcd82),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95fee2),
	.w1(32'hb92ddf9e),
	.w2(32'h39275664),
	.w3(32'hb8f5c59a),
	.w4(32'hb9966e35),
	.w5(32'hbac08782),
	.w6(32'hba9e1f95),
	.w7(32'hba62dd8b),
	.w8(32'hbae3ea24),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edced2),
	.w1(32'h3bcf17b9),
	.w2(32'hb9b9e309),
	.w3(32'hba457a75),
	.w4(32'h3b82b8ea),
	.w5(32'h3ac5e37e),
	.w6(32'hba9d7ea8),
	.w7(32'h3b7ab4cc),
	.w8(32'hbaeb94ed),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17fcc1),
	.w1(32'h3b10a12d),
	.w2(32'hb9ac2346),
	.w3(32'h3a7ac320),
	.w4(32'h3acf543e),
	.w5(32'h39d4593a),
	.w6(32'hbac662db),
	.w7(32'hbb1666c3),
	.w8(32'hba8fc8df),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb6b08),
	.w1(32'hb83bdc48),
	.w2(32'hba3c3edf),
	.w3(32'hbb1ae1d7),
	.w4(32'hbb3b31b7),
	.w5(32'hbb8120f5),
	.w6(32'hba939662),
	.w7(32'hbb2577b8),
	.w8(32'hbb85e148),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c1fb1),
	.w1(32'h39cc8278),
	.w2(32'hba121f5c),
	.w3(32'hba050702),
	.w4(32'hba965d2d),
	.w5(32'hbaf646db),
	.w6(32'hb986db41),
	.w7(32'hba07df39),
	.w8(32'hbb14dadf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba893c5d),
	.w1(32'h39d31368),
	.w2(32'hbb80b465),
	.w3(32'h38f431c2),
	.w4(32'h3b4a5b05),
	.w5(32'hba016035),
	.w6(32'hbb0f5007),
	.w7(32'hb92a60e1),
	.w8(32'hbb674ace),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5bb16),
	.w1(32'h3a4a15fb),
	.w2(32'h3a623eeb),
	.w3(32'hbb794ed1),
	.w4(32'hba18e2fc),
	.w5(32'hba6ad2aa),
	.w6(32'hbad62ca5),
	.w7(32'hba3fb61a),
	.w8(32'hb9cc25a4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15866e),
	.w1(32'h3a2946d1),
	.w2(32'h39b7546d),
	.w3(32'h3a810eb3),
	.w4(32'hb9974f95),
	.w5(32'hb8a0dbdf),
	.w6(32'h3a38ca7b),
	.w7(32'hb9c9fb14),
	.w8(32'h39d9e557),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39247b48),
	.w1(32'hbb91c179),
	.w2(32'hbbd788d2),
	.w3(32'hbb7e1a49),
	.w4(32'hbb803ec9),
	.w5(32'hbbefa41a),
	.w6(32'hbbd087f6),
	.w7(32'hbb8382b4),
	.w8(32'hbbdb8d9a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa85a3),
	.w1(32'hba2f5737),
	.w2(32'hba6a8d6f),
	.w3(32'hb9977994),
	.w4(32'h3a3e50bc),
	.w5(32'hb985fbc0),
	.w6(32'hb93a86a0),
	.w7(32'h3a40e412),
	.w8(32'hba0e9e5a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1ac20),
	.w1(32'h3b051837),
	.w2(32'hbb1ee026),
	.w3(32'h389dd794),
	.w4(32'h3ac49eea),
	.w5(32'hbb36aa87),
	.w6(32'hba9aa1da),
	.w7(32'h38d52f12),
	.w8(32'hbb4bfe96),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1934e0),
	.w1(32'h394716f1),
	.w2(32'hba52da47),
	.w3(32'hbb2ccfb4),
	.w4(32'hbb9cd758),
	.w5(32'hbbb2023a),
	.w6(32'h3a011ac7),
	.w7(32'hbab1ae63),
	.w8(32'hbbb69932),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d130),
	.w1(32'h39ad717b),
	.w2(32'hbab1ee44),
	.w3(32'hbb3045d4),
	.w4(32'hbad0ba02),
	.w5(32'hbb29c0dc),
	.w6(32'hb94797b0),
	.w7(32'h39120ab4),
	.w8(32'hbb3c1f32),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf13af),
	.w1(32'hb94ad4b4),
	.w2(32'hbad3302f),
	.w3(32'hba754992),
	.w4(32'hbabe51ea),
	.w5(32'h3a26d4b1),
	.w6(32'hb9a0aee8),
	.w7(32'hbad4f626),
	.w8(32'hb9d9a1b4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6772fb),
	.w1(32'hb91b4adc),
	.w2(32'h3b31b155),
	.w3(32'hbae52ec8),
	.w4(32'hbb216ee5),
	.w5(32'hbb902c09),
	.w6(32'hbaa07411),
	.w7(32'hba989005),
	.w8(32'hbb36cd55),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae121e1),
	.w1(32'hb9898a70),
	.w2(32'hbb890fa8),
	.w3(32'h3a16a245),
	.w4(32'h3accd909),
	.w5(32'hba183cb4),
	.w6(32'hbaa616c2),
	.w7(32'hba80b82b),
	.w8(32'hbb346001),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00477),
	.w1(32'h3b1b1d2d),
	.w2(32'hb9f27773),
	.w3(32'h3ab2008d),
	.w4(32'h3b180b6c),
	.w5(32'hbb755ce1),
	.w6(32'hba9ad54c),
	.w7(32'h39a62020),
	.w8(32'hbb63b2db),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4dee),
	.w1(32'hb9b99ef4),
	.w2(32'hba688f5c),
	.w3(32'hbabbb716),
	.w4(32'hba90ff62),
	.w5(32'h3a330f8f),
	.w6(32'hba653b26),
	.w7(32'hba6fc854),
	.w8(32'h3a4e7cfc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cd1ff),
	.w1(32'hba0dbad1),
	.w2(32'hb9baaea1),
	.w3(32'h3a08a8d8),
	.w4(32'h39ea140c),
	.w5(32'h3a8fa59e),
	.w6(32'h392aecbc),
	.w7(32'h3925f706),
	.w8(32'h3b23689d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a6ea),
	.w1(32'h3c527c01),
	.w2(32'h3bacfb1c),
	.w3(32'hbb0c8dc6),
	.w4(32'h3b9e3e15),
	.w5(32'hbb9eb4a8),
	.w6(32'hba1b41df),
	.w7(32'hbb5b1742),
	.w8(32'hbc1f84a2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da712),
	.w1(32'h3b8177d5),
	.w2(32'hba9bcaf5),
	.w3(32'h39d07ce9),
	.w4(32'h3a707517),
	.w5(32'hbb030114),
	.w6(32'hbb8a2ae4),
	.w7(32'hbba4fffa),
	.w8(32'hbbe481a7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45bc64),
	.w1(32'h3a4cc262),
	.w2(32'hbab9e4d7),
	.w3(32'hbb833e3f),
	.w4(32'hbb4397f7),
	.w5(32'hbb924e4f),
	.w6(32'h372ed5c2),
	.w7(32'hba5a74df),
	.w8(32'hbb9b92d9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b0d09),
	.w1(32'h3a892719),
	.w2(32'hbc3dec3c),
	.w3(32'h398fc82d),
	.w4(32'h3b875bed),
	.w5(32'hba308876),
	.w6(32'h3ba6c156),
	.w7(32'h3c16baab),
	.w8(32'hbbcc292f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccd4f0),
	.w1(32'hbad759c5),
	.w2(32'hbabb8e13),
	.w3(32'h38b33e53),
	.w4(32'hb9781d7f),
	.w5(32'hbafb3790),
	.w6(32'hbac86d39),
	.w7(32'hbb183b22),
	.w8(32'hbb3dfdd6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaea50f),
	.w1(32'hbacd1528),
	.w2(32'hbb4214f1),
	.w3(32'hba93fcaa),
	.w4(32'hba8c5c67),
	.w5(32'hbb6cd8bb),
	.w6(32'hbb2d9e20),
	.w7(32'hbb74f9dd),
	.w8(32'hbb670b07),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb811355),
	.w1(32'h3cbb5362),
	.w2(32'h3ab8f89d),
	.w3(32'hbc0f4fd2),
	.w4(32'h3c669c4e),
	.w5(32'h3aef3d24),
	.w6(32'hbc491db2),
	.w7(32'h3c04dc87),
	.w8(32'hbc1c6854),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b882603),
	.w1(32'h3b839347),
	.w2(32'hbb8cbf61),
	.w3(32'h3b7f7255),
	.w4(32'h3c0d350a),
	.w5(32'hbb1f936d),
	.w6(32'hbb4e9d5d),
	.w7(32'h3a1e0e8d),
	.w8(32'hbbdebcf5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5837f),
	.w1(32'h3aa29684),
	.w2(32'hbbb0d574),
	.w3(32'hbac14e51),
	.w4(32'hb9955ce5),
	.w5(32'h39d21599),
	.w6(32'hba7d3760),
	.w7(32'hbacac751),
	.w8(32'hbb9a1ccd),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44fd28),
	.w1(32'hba9d1560),
	.w2(32'hba9b5624),
	.w3(32'hbb783b4f),
	.w4(32'hbbad54c6),
	.w5(32'hbb83ec2f),
	.w6(32'hba804611),
	.w7(32'hbb17997f),
	.w8(32'hbb529e6d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12c77),
	.w1(32'hbb41058c),
	.w2(32'hbb2e5285),
	.w3(32'hbac3333c),
	.w4(32'hbbbfaf62),
	.w5(32'hbbe97876),
	.w6(32'h3a88f08e),
	.w7(32'hbb36864d),
	.w8(32'hbbd4dce5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba935cd5),
	.w1(32'hba5d2520),
	.w2(32'hb9b5aa7a),
	.w3(32'hbaddba52),
	.w4(32'hba20c83e),
	.w5(32'h3a40013d),
	.w6(32'hba375bb4),
	.w7(32'h38e864ab),
	.w8(32'hbab0b02f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8788f5),
	.w1(32'hbb05e91b),
	.w2(32'h39f0b5b7),
	.w3(32'h39a35225),
	.w4(32'hb9196dd7),
	.w5(32'hbab44511),
	.w6(32'hb9f08f28),
	.w7(32'h3ac00475),
	.w8(32'hba315fd7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d761e),
	.w1(32'h3a780d33),
	.w2(32'hbacbe8d0),
	.w3(32'h3a9326eb),
	.w4(32'h3b2fcd2c),
	.w5(32'hbadd4259),
	.w6(32'hbadcc63a),
	.w7(32'h39957474),
	.w8(32'hbb4c2268),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9390a7),
	.w1(32'h3a19ac69),
	.w2(32'hba0c356e),
	.w3(32'hb9377680),
	.w4(32'h3a472beb),
	.w5(32'hbaaef577),
	.w6(32'hba3a10ce),
	.w7(32'h392d5a5b),
	.w8(32'hbb310dff),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc3bdd),
	.w1(32'h3bba1865),
	.w2(32'h3bbd9f7c),
	.w3(32'h3b1d774d),
	.w4(32'h3c1ab2fa),
	.w5(32'hbc0b151b),
	.w6(32'hb9d4a88e),
	.w7(32'h3c1572a6),
	.w8(32'hbbe5c55d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bec8bd),
	.w1(32'h3c015563),
	.w2(32'hbad3225d),
	.w3(32'hbbc1729c),
	.w4(32'h3b1134c9),
	.w5(32'hbc8263a4),
	.w6(32'hbbd402e0),
	.w7(32'hbb3d129c),
	.w8(32'hbcb25107),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21881c),
	.w1(32'hb9c0be9d),
	.w2(32'h3c086009),
	.w3(32'hb9e42151),
	.w4(32'h3c1d7e17),
	.w5(32'hbb3cee67),
	.w6(32'h3b22c2b7),
	.w7(32'h3c6368b2),
	.w8(32'h3bcd5e08),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c1d6),
	.w1(32'hbb958bb3),
	.w2(32'h3b326a26),
	.w3(32'hbb04bd9a),
	.w4(32'hbacef42a),
	.w5(32'h3b140052),
	.w6(32'hba8ca23d),
	.w7(32'h3b83a697),
	.w8(32'h3ac651a8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6795bf),
	.w1(32'h3bcd3a6d),
	.w2(32'hbc53d371),
	.w3(32'h3ab3c7cb),
	.w4(32'h3a227738),
	.w5(32'h3a0592a0),
	.w6(32'hbabd3725),
	.w7(32'hbba2a0d8),
	.w8(32'h3a12db03),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf7e55),
	.w1(32'h3acdf0b4),
	.w2(32'hbb5f6d9b),
	.w3(32'hbbd7b7ee),
	.w4(32'h38a0894d),
	.w5(32'hbbc481fe),
	.w6(32'hbbe38968),
	.w7(32'hbba6b05b),
	.w8(32'hbc04ec29),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9034),
	.w1(32'hbb9da05b),
	.w2(32'h3bf46c2f),
	.w3(32'h39210171),
	.w4(32'h3c8c4c04),
	.w5(32'hba5f1b98),
	.w6(32'hbb9525b8),
	.w7(32'h3c5bb1c0),
	.w8(32'hbb4b952e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d6afe),
	.w1(32'h3bb105cf),
	.w2(32'hba8ac2d9),
	.w3(32'h3b1de52f),
	.w4(32'h3ba7953d),
	.w5(32'hbb84b851),
	.w6(32'h3b2a38fd),
	.w7(32'h3b95db72),
	.w8(32'hbc352f2c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7aaf),
	.w1(32'hbb8fc3a2),
	.w2(32'h3be97ca3),
	.w3(32'hbbdb0f6d),
	.w4(32'hba645240),
	.w5(32'hbb70b145),
	.w6(32'hbc1a5984),
	.w7(32'hbaf62291),
	.w8(32'hbb999074),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63343f),
	.w1(32'h3bf58d4e),
	.w2(32'h3c164e37),
	.w3(32'h3bfa311c),
	.w4(32'h3c1ae2d9),
	.w5(32'hbbe62b32),
	.w6(32'h3bcc10e4),
	.w7(32'h3c2a207e),
	.w8(32'hbc0eb546),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d6e7),
	.w1(32'hbbe5bedb),
	.w2(32'h3aab859e),
	.w3(32'hbbc8acc9),
	.w4(32'h3bf4158e),
	.w5(32'hbb712b53),
	.w6(32'hbc01e4dd),
	.w7(32'h3b9f0be3),
	.w8(32'hbbb2bab8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82af55),
	.w1(32'h3b27c904),
	.w2(32'hbb336c1b),
	.w3(32'hbb0ef5f4),
	.w4(32'hbbd403d8),
	.w5(32'hba4947e3),
	.w6(32'h3a8a9fd6),
	.w7(32'h3a0bb653),
	.w8(32'h3b07172f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36a26e),
	.w1(32'h3c6a1277),
	.w2(32'h3c00fac2),
	.w3(32'hbb2b7105),
	.w4(32'hbbb66d9d),
	.w5(32'h3bb762a8),
	.w6(32'h3bc57a53),
	.w7(32'h3b10e5a1),
	.w8(32'h3bae0620),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2ed8f),
	.w1(32'hbba7633b),
	.w2(32'hbbd31557),
	.w3(32'hb92a9489),
	.w4(32'h3b029e88),
	.w5(32'h3b1caec6),
	.w6(32'h3a5781cb),
	.w7(32'h3bda06ca),
	.w8(32'h391c3975),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baccbb9),
	.w1(32'h3a1bc579),
	.w2(32'hbc10ba77),
	.w3(32'h399bf704),
	.w4(32'hbbac7d8c),
	.w5(32'hbb3978f9),
	.w6(32'hbb1cb3f0),
	.w7(32'hbc192151),
	.w8(32'hbae1eacf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06a6e3),
	.w1(32'hbbbdfbde),
	.w2(32'hbc043b5b),
	.w3(32'h3987f648),
	.w4(32'h3bec1041),
	.w5(32'h3b2b2255),
	.w6(32'h389d6d71),
	.w7(32'h3bf038e1),
	.w8(32'hbbb35220),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b99ea),
	.w1(32'h3adf049c),
	.w2(32'h3b589875),
	.w3(32'h3bf74dad),
	.w4(32'h3b96ab4b),
	.w5(32'h3a826b15),
	.w6(32'h3b86c421),
	.w7(32'h3ba12ecd),
	.w8(32'h3b2748ed),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0689d),
	.w1(32'hbb708f19),
	.w2(32'h3aa3cc32),
	.w3(32'hb91a8760),
	.w4(32'hbb18c99f),
	.w5(32'hbb4f4dea),
	.w6(32'hbb4f01b1),
	.w7(32'hba6bf027),
	.w8(32'hbc12cb71),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69b4a),
	.w1(32'hb9a4a563),
	.w2(32'h3bf2c274),
	.w3(32'hba4cd5e6),
	.w4(32'h3b067c42),
	.w5(32'hbb140f7f),
	.w6(32'h3986efc1),
	.w7(32'h3bd0477e),
	.w8(32'hbba75546),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecb6ff),
	.w1(32'hbbbd3381),
	.w2(32'h3a97aa20),
	.w3(32'h3a435923),
	.w4(32'h3ba2e1a2),
	.w5(32'hbb4d7a7b),
	.w6(32'hbbb8c79a),
	.w7(32'h3b311ba2),
	.w8(32'hbb8fdd5e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bec1d),
	.w1(32'hbb51b20f),
	.w2(32'hbb62c3b1),
	.w3(32'hbae01adb),
	.w4(32'h3b155b71),
	.w5(32'hbbc93b86),
	.w6(32'hbbc8f38b),
	.w7(32'h3b2dc2cb),
	.w8(32'hbbda9b74),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a88a8),
	.w1(32'hba9b3b98),
	.w2(32'h3a70f863),
	.w3(32'hbc0564c7),
	.w4(32'hba387692),
	.w5(32'h3a8cbefb),
	.w6(32'hbbe7a383),
	.w7(32'hbaf2e2fa),
	.w8(32'hbb146044),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34ab71),
	.w1(32'h396e5838),
	.w2(32'hbb11806b),
	.w3(32'h3b97c078),
	.w4(32'hbb03a80e),
	.w5(32'h3a7f5e28),
	.w6(32'h3a8a9e4e),
	.w7(32'hbbdbd92e),
	.w8(32'h3af976cb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb279f2),
	.w1(32'hb9b288d4),
	.w2(32'hbbf20b3d),
	.w3(32'hbbd19d06),
	.w4(32'hbc1d01b0),
	.w5(32'hb9a4a273),
	.w6(32'hbb0f5148),
	.w7(32'hbc49d4a5),
	.w8(32'h3b73d389),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a692ce0),
	.w1(32'hbb7451be),
	.w2(32'hbbe7c8fe),
	.w3(32'h3ba56a11),
	.w4(32'hba319213),
	.w5(32'h3bf22a45),
	.w6(32'hbb057cb5),
	.w7(32'hba805ca4),
	.w8(32'h3bbe78b5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15dd5c),
	.w1(32'h3b96dd25),
	.w2(32'hbb6a0984),
	.w3(32'h3915ffcb),
	.w4(32'hbbdd173e),
	.w5(32'hbad0b0d1),
	.w6(32'h3a969d62),
	.w7(32'hbbf52d2f),
	.w8(32'h3b024c07),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228917),
	.w1(32'hbb5c81f8),
	.w2(32'hbb7279e5),
	.w3(32'hb9ba891b),
	.w4(32'hbbdb351f),
	.w5(32'h3869182e),
	.w6(32'hbae73b59),
	.w7(32'hbba140fb),
	.w8(32'h3b6e64ba),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bb793),
	.w1(32'hbb4dfe6c),
	.w2(32'hbc03d3ef),
	.w3(32'hb97bba0e),
	.w4(32'h3be652f5),
	.w5(32'hbc413d78),
	.w6(32'hbb83bbbb),
	.w7(32'h3aaeba2e),
	.w8(32'hbc850b5a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0521d5),
	.w1(32'h3b8c52b5),
	.w2(32'h3c4f36e0),
	.w3(32'h3bf23400),
	.w4(32'h3c061d63),
	.w5(32'hbb2f37b0),
	.w6(32'h3c3d37ea),
	.w7(32'h3c99051b),
	.w8(32'hba9df905),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aec6a7),
	.w1(32'h389e33ee),
	.w2(32'hbae85850),
	.w3(32'hbc528a38),
	.w4(32'hbb9bba10),
	.w5(32'hbbb0dd1c),
	.w6(32'hbbdcc956),
	.w7(32'hbc161bd0),
	.w8(32'hbbbca92d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule