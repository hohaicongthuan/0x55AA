module layer_8_featuremap_77(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5b96),
	.w1(32'hbaa5ea05),
	.w2(32'hbacef906),
	.w3(32'hbbcb0ecd),
	.w4(32'hbc0705e6),
	.w5(32'hbbfcc951),
	.w6(32'hbb80c727),
	.w7(32'hbbfa3684),
	.w8(32'hbc22f2de),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8756fa),
	.w1(32'h3bc34abf),
	.w2(32'h3aafed9a),
	.w3(32'h3a72d626),
	.w4(32'h3ac80ff8),
	.w5(32'hbafb3e5a),
	.w6(32'h3b84bf6a),
	.w7(32'h3a2b985e),
	.w8(32'hbb4e5ff6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf871),
	.w1(32'h3b73a624),
	.w2(32'h3b7578a9),
	.w3(32'h3ac270dc),
	.w4(32'h393aeaaa),
	.w5(32'hb97bd027),
	.w6(32'h3ba498c4),
	.w7(32'h3b8bb99b),
	.w8(32'hb8602f7d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88fbb4),
	.w1(32'hbb2dffc8),
	.w2(32'hbab22575),
	.w3(32'hbb33c12b),
	.w4(32'hbb56b009),
	.w5(32'hba39136b),
	.w6(32'hbbffea7f),
	.w7(32'hbbdf04de),
	.w8(32'hb9136165),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3b1b),
	.w1(32'h3b981151),
	.w2(32'h3b12c8ec),
	.w3(32'hb9aa2118),
	.w4(32'h3a3afd7b),
	.w5(32'hbb1cf704),
	.w6(32'h3b4f8221),
	.w7(32'h3ad1e028),
	.w8(32'h3b8836b4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6ed3),
	.w1(32'h3c25795a),
	.w2(32'h3c24f6ab),
	.w3(32'h3b61a51e),
	.w4(32'h3bea3472),
	.w5(32'h3bd06caf),
	.w6(32'h3c1ba533),
	.w7(32'h3c4be390),
	.w8(32'h3bf65c5e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cfb33),
	.w1(32'h3bc27a85),
	.w2(32'h3b846ce6),
	.w3(32'hb8467112),
	.w4(32'h3b325818),
	.w5(32'h3af9a401),
	.w6(32'h3bb2ac9b),
	.w7(32'h3b6f3e23),
	.w8(32'h3a8143bc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967243),
	.w1(32'h3ba147d9),
	.w2(32'h3b006c77),
	.w3(32'hbb696d9b),
	.w4(32'hbb5b59e3),
	.w5(32'hbb855aaa),
	.w6(32'h39382735),
	.w7(32'hba70ef33),
	.w8(32'h3ad4a37f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf155),
	.w1(32'h3b94ff7f),
	.w2(32'hba5dfe1e),
	.w3(32'h3904a150),
	.w4(32'hbabee1fc),
	.w5(32'hbb1a5cb3),
	.w6(32'h3b3d71dc),
	.w7(32'hbb63f672),
	.w8(32'hbc06d116),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afab9d5),
	.w1(32'hb8a4130a),
	.w2(32'hba1e321e),
	.w3(32'h3b6c149f),
	.w4(32'h3b5cdb29),
	.w5(32'h3bd83831),
	.w6(32'hbb1479d4),
	.w7(32'hbb169e0f),
	.w8(32'hb8822a64),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf724c),
	.w1(32'hbbb72348),
	.w2(32'hba56dd27),
	.w3(32'hbc10ab6a),
	.w4(32'hbc5f8fcb),
	.w5(32'hbc076401),
	.w6(32'hbbdb648f),
	.w7(32'hbb839003),
	.w8(32'hbb390744),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131c46),
	.w1(32'h39bedf44),
	.w2(32'hb897a8bd),
	.w3(32'hbb82c8f9),
	.w4(32'hbb59fec4),
	.w5(32'hbb33ec7b),
	.w6(32'h3a8edfef),
	.w7(32'h392a0561),
	.w8(32'h39e31c4b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6aa46),
	.w1(32'h3bca2424),
	.w2(32'h3b406bac),
	.w3(32'h3a1a56b1),
	.w4(32'h3a8a2fa0),
	.w5(32'h3b01e4e5),
	.w6(32'h3b3e2d1b),
	.w7(32'h3990901d),
	.w8(32'h3c242d0f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd0894),
	.w1(32'h3bc426a3),
	.w2(32'h3bc022e6),
	.w3(32'h3b3d5b32),
	.w4(32'h3aab49dd),
	.w5(32'h3a2600ac),
	.w6(32'h3bda424f),
	.w7(32'h3becb174),
	.w8(32'h3b8c1a19),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b04c),
	.w1(32'h3b82fcbd),
	.w2(32'h3b55bd03),
	.w3(32'h3aed5468),
	.w4(32'h3b0897f9),
	.w5(32'h3a5dcbb7),
	.w6(32'h3b6dc614),
	.w7(32'h3b81277e),
	.w8(32'h3a8c23b4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a785c0a),
	.w1(32'h3a3b98e6),
	.w2(32'hb94737c1),
	.w3(32'hb95e4e8f),
	.w4(32'hba9cb844),
	.w5(32'hb9de6500),
	.w6(32'h399633cc),
	.w7(32'hb8930f03),
	.w8(32'h3b01ad30),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58235b),
	.w1(32'hbb838b30),
	.w2(32'hbb1d7d8e),
	.w3(32'h3b8569d8),
	.w4(32'h3c037cd1),
	.w5(32'h3c3e37c9),
	.w6(32'h3ba320e5),
	.w7(32'h3b2de3f9),
	.w8(32'h3ac6f807),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaae2da),
	.w1(32'h3a100eaf),
	.w2(32'h3ae07fde),
	.w3(32'hbbc8d51b),
	.w4(32'hbbd93146),
	.w5(32'hbb0a6845),
	.w6(32'h3875ec5f),
	.w7(32'h3a4076e8),
	.w8(32'h3b14af98),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3888ae),
	.w1(32'hbb9aa216),
	.w2(32'h3c1685af),
	.w3(32'hbc46b5b9),
	.w4(32'hbca148ba),
	.w5(32'hbc1d3269),
	.w6(32'h3b6a3c9f),
	.w7(32'h3b49424f),
	.w8(32'h3c6c1a21),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac76a4),
	.w1(32'hba5e54e6),
	.w2(32'h3b7d8b85),
	.w3(32'hbc282658),
	.w4(32'hbc10c7bc),
	.w5(32'hbc16cf96),
	.w6(32'h3966960e),
	.w7(32'h38af1359),
	.w8(32'hbb52ec07),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6100f7),
	.w1(32'hba1ba5b5),
	.w2(32'h3a62e3ea),
	.w3(32'h3aaad0c2),
	.w4(32'h39e0d694),
	.w5(32'hba1af241),
	.w6(32'h3a445c9d),
	.w7(32'h3a0deac0),
	.w8(32'h3c0fafd3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c263470),
	.w1(32'h3c4b5f37),
	.w2(32'h3c39382d),
	.w3(32'h3bd7ccb9),
	.w4(32'h3c190c86),
	.w5(32'h3c18072c),
	.w6(32'h3c2061c7),
	.w7(32'h3c3192f3),
	.w8(32'h3aa3a833),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c1a1c),
	.w1(32'hbc0c0647),
	.w2(32'hbc218e59),
	.w3(32'h385abbf9),
	.w4(32'hbc9502f9),
	.w5(32'hbcb458c6),
	.w6(32'hbc1a29d4),
	.w7(32'hbcabbf95),
	.w8(32'hbc7e04e1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d59f8),
	.w1(32'hbb22e3e9),
	.w2(32'hbb33627b),
	.w3(32'hbbe70c21),
	.w4(32'hbbb3a9ec),
	.w5(32'hbbd8d97d),
	.w6(32'hba83f2e1),
	.w7(32'hbb871795),
	.w8(32'hbb9be3bb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae80eaf),
	.w1(32'hbb7d8726),
	.w2(32'hbb015a04),
	.w3(32'hba23f0a6),
	.w4(32'hbb1cc616),
	.w5(32'hb9872c27),
	.w6(32'hbb2fcc5d),
	.w7(32'hba8c138b),
	.w8(32'hba9e1499),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7054b2),
	.w1(32'hba8d1bc7),
	.w2(32'hbac21fac),
	.w3(32'hbb9b52e7),
	.w4(32'hbc1a7fae),
	.w5(32'hbc57f17e),
	.w6(32'hbbfc1017),
	.w7(32'hbc2fd701),
	.w8(32'hbc36abc4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad410ed),
	.w1(32'hbb5311e5),
	.w2(32'hbb394d24),
	.w3(32'hba16d017),
	.w4(32'hbb1f505c),
	.w5(32'hbac4fbb0),
	.w6(32'hbb2e8b51),
	.w7(32'hbb4c2ca9),
	.w8(32'hba58ca64),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdafdfaa),
	.w1(32'hbcc858db),
	.w2(32'hbc31de59),
	.w3(32'hbc44bbc0),
	.w4(32'h3b93aa6c),
	.w5(32'hbd3d199d),
	.w6(32'hbda46663),
	.w7(32'hbd2ae7b4),
	.w8(32'hbb1b082e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23e1f3),
	.w1(32'h3ba161d9),
	.w2(32'h3ae712fb),
	.w3(32'hbb90ed64),
	.w4(32'hbaf4515d),
	.w5(32'hbb257cc8),
	.w6(32'h3b0bb992),
	.w7(32'h3a8cc8b0),
	.w8(32'hbab2e6b3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f6cd4),
	.w1(32'h39f0c390),
	.w2(32'hbabb0648),
	.w3(32'hb9739964),
	.w4(32'h38b62296),
	.w5(32'hbabceed4),
	.w6(32'h39f87704),
	.w7(32'hb9378704),
	.w8(32'hbacd83e3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e43bf),
	.w1(32'hbb9903d8),
	.w2(32'hbb363636),
	.w3(32'hbbdeef1a),
	.w4(32'hbba1738f),
	.w5(32'hbb377f9d),
	.w6(32'hbb30fdd1),
	.w7(32'hbaf61914),
	.w8(32'hbaea22d2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f28e9),
	.w1(32'hba64d6e3),
	.w2(32'hba07e601),
	.w3(32'h3b071b8c),
	.w4(32'h3b333ed4),
	.w5(32'h3a76364b),
	.w6(32'h3a15aa9d),
	.w7(32'h3ad384fe),
	.w8(32'h39905558),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16f28d),
	.w1(32'h3abee53c),
	.w2(32'hbaceb7e4),
	.w3(32'hbaa02567),
	.w4(32'hb9a3bec9),
	.w5(32'hbb261b40),
	.w6(32'hbb6dc9df),
	.w7(32'hbb8e348b),
	.w8(32'hbb1e3306),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0012ec),
	.w1(32'hbb0cd51d),
	.w2(32'h39098700),
	.w3(32'h39cff8e6),
	.w4(32'h3ac44f33),
	.w5(32'h3a479f79),
	.w6(32'hbba4c531),
	.w7(32'hba3704f3),
	.w8(32'h3c066aec),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcb6b6),
	.w1(32'h3bebef2c),
	.w2(32'h3bf91cea),
	.w3(32'h3b6192cc),
	.w4(32'h3b92d632),
	.w5(32'h3b4b3843),
	.w6(32'h3c3140f1),
	.w7(32'h3c4ef9d6),
	.w8(32'h3bd18c96),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57e17c),
	.w1(32'hb93a104d),
	.w2(32'h3aa7b165),
	.w3(32'hbc19f8f9),
	.w4(32'hbc0972f0),
	.w5(32'hbbcb7ed1),
	.w6(32'hb98373bf),
	.w7(32'hbb43a110),
	.w8(32'hbb244346),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332b7c),
	.w1(32'hbb232337),
	.w2(32'hba8e7877),
	.w3(32'hbac28986),
	.w4(32'hbadcfb5a),
	.w5(32'hb95e0063),
	.w6(32'hbb137089),
	.w7(32'hba624bbe),
	.w8(32'hbb3feedd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c1390),
	.w1(32'hbacd5343),
	.w2(32'hbba54c30),
	.w3(32'h389ebb89),
	.w4(32'hba32d9cc),
	.w5(32'hbba1eeb8),
	.w6(32'h3a07d9dd),
	.w7(32'hbaaa4599),
	.w8(32'h3b97700b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddaf59),
	.w1(32'h3c02a44e),
	.w2(32'h3bb6dd04),
	.w3(32'h3b57ce50),
	.w4(32'h3b94bafa),
	.w5(32'h3a74dfd8),
	.w6(32'h3bca1537),
	.w7(32'h3bce5f4e),
	.w8(32'hbaa7397a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d96ac),
	.w1(32'h39f340d4),
	.w2(32'hb8c1183f),
	.w3(32'h3a02a4a1),
	.w4(32'h3a3d1150),
	.w5(32'h3910edc0),
	.w6(32'hba512708),
	.w7(32'hba7c7fe7),
	.w8(32'hba7b6d24),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18abc4),
	.w1(32'hbc0961bd),
	.w2(32'hbbeb26e6),
	.w3(32'hbc8f50bd),
	.w4(32'hbc94a7d9),
	.w5(32'hbc9c3540),
	.w6(32'hbc91fc84),
	.w7(32'hbc7e7343),
	.w8(32'hbc5305c6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9394a7f),
	.w1(32'hb8e6ca89),
	.w2(32'h3b82905c),
	.w3(32'hba335da5),
	.w4(32'hb7d8e76e),
	.w5(32'h3b45faa5),
	.w6(32'h3aa4905e),
	.w7(32'h3b3151c6),
	.w8(32'h3bb9b6e2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba101cbb),
	.w1(32'h398632fb),
	.w2(32'h3a1e5ece),
	.w3(32'hb98b48d9),
	.w4(32'h3a7405da),
	.w5(32'h3a22da9f),
	.w6(32'hb8328d4c),
	.w7(32'h391f8a9a),
	.w8(32'h3ad5d373),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf81f0a),
	.w1(32'hbb357fc8),
	.w2(32'hbb0353fe),
	.w3(32'hbb8572b8),
	.w4(32'hbba8f1fd),
	.w5(32'hbbb1d3cf),
	.w6(32'hbb9b7943),
	.w7(32'hbb94899b),
	.w8(32'hbb82a2fe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67371c),
	.w1(32'h3ab8614a),
	.w2(32'h3b9e9b38),
	.w3(32'hbacdf5d0),
	.w4(32'hbb4d8f53),
	.w5(32'hba35f4f5),
	.w6(32'h39d08500),
	.w7(32'h3ac196af),
	.w8(32'h3ba6df35),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fecc),
	.w1(32'hb9ef0bba),
	.w2(32'h3b0fa7b8),
	.w3(32'hbb406371),
	.w4(32'hba14790e),
	.w5(32'h3b19f420),
	.w6(32'hbb2da793),
	.w7(32'h3a1667a0),
	.w8(32'h3b0b7aaa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629a10),
	.w1(32'hbb43ecb8),
	.w2(32'hbb15c113),
	.w3(32'hba81b4b9),
	.w4(32'hbad5ddc4),
	.w5(32'hbaa2fb59),
	.w6(32'hba8a5c00),
	.w7(32'hba10aace),
	.w8(32'h39242f20),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273379),
	.w1(32'h3aec2fc1),
	.w2(32'h3b80d25a),
	.w3(32'h3a8da425),
	.w4(32'hbb1ab7df),
	.w5(32'hbb6e0d8c),
	.w6(32'h3a92cc67),
	.w7(32'hba8247f1),
	.w8(32'h3a80b3a2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14e91b),
	.w1(32'hba39b8a0),
	.w2(32'h3ada8834),
	.w3(32'hba8e9c7c),
	.w4(32'hba39cb10),
	.w5(32'h3b01ce13),
	.w6(32'h3ad7b98d),
	.w7(32'h3b18d991),
	.w8(32'h3b716411),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99bd2a),
	.w1(32'hbafda2b5),
	.w2(32'hbac4626c),
	.w3(32'hbb7930b2),
	.w4(32'hbbe55745),
	.w5(32'hbbbb22e7),
	.w6(32'hbb968501),
	.w7(32'hbb8d9e78),
	.w8(32'hbb70afcc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c388480),
	.w1(32'h3c24ea90),
	.w2(32'h3ae2b96d),
	.w3(32'h3c4004c0),
	.w4(32'h3c2f7abb),
	.w5(32'h3aaf7875),
	.w6(32'h3c31b95d),
	.w7(32'h3c01ae4f),
	.w8(32'h3af53151),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ddfa6),
	.w1(32'h3a4b79e0),
	.w2(32'h3c0bcbac),
	.w3(32'hbba2556b),
	.w4(32'hbc12a972),
	.w5(32'hbb062ee4),
	.w6(32'h3be5838d),
	.w7(32'h3b4878fc),
	.w8(32'h3c26eae2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f6e4c),
	.w1(32'hba5f177b),
	.w2(32'hb9c6738e),
	.w3(32'hbb679021),
	.w4(32'hbbf57d7f),
	.w5(32'hbbb99f8a),
	.w6(32'hbb06a9d9),
	.w7(32'hbbcb09ba),
	.w8(32'hbbd24fee),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba132cef),
	.w1(32'hbb179203),
	.w2(32'hb9e01880),
	.w3(32'hbb3e61cc),
	.w4(32'hbba6c7bf),
	.w5(32'hbad5381b),
	.w6(32'h3a0be816),
	.w7(32'hbaaaf3e5),
	.w8(32'h3afdbddc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfa233),
	.w1(32'hbb106dc4),
	.w2(32'hbaf210ea),
	.w3(32'hba43532c),
	.w4(32'hba40979a),
	.w5(32'hba49caa7),
	.w6(32'hbacaf432),
	.w7(32'hbac9b18c),
	.w8(32'hb8a49d3c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb651ae1),
	.w1(32'hbb26252e),
	.w2(32'hbad4cdc8),
	.w3(32'h392c9d98),
	.w4(32'hbc004180),
	.w5(32'hbc11952e),
	.w6(32'hbb92de40),
	.w7(32'hbb5015c5),
	.w8(32'hba9add5d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40625d),
	.w1(32'h3af70689),
	.w2(32'h3b890c40),
	.w3(32'h3a7d1088),
	.w4(32'h3b2c2186),
	.w5(32'h3b69acef),
	.w6(32'h3b3bf4de),
	.w7(32'h3b257b52),
	.w8(32'h3a01c697),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823aa65),
	.w1(32'h39bb5df9),
	.w2(32'h3b7f186b),
	.w3(32'hbbc1fae7),
	.w4(32'hbbe26294),
	.w5(32'hba83451d),
	.w6(32'hbb58c1e4),
	.w7(32'hbaa81d61),
	.w8(32'h3b396f35),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1465db),
	.w1(32'h3a96c378),
	.w2(32'h3a582332),
	.w3(32'hba903e35),
	.w4(32'hba0d4b4e),
	.w5(32'hba8952c6),
	.w6(32'hba05cae5),
	.w7(32'hbaae09c7),
	.w8(32'h3902b151),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a719d91),
	.w1(32'h39832b83),
	.w2(32'hba0dd39b),
	.w3(32'hba63013d),
	.w4(32'hbafca28d),
	.w5(32'hbb064e73),
	.w6(32'hbadb7390),
	.w7(32'hbacabfc7),
	.w8(32'hba7471dd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ca485),
	.w1(32'hbae22ec2),
	.w2(32'h393839bd),
	.w3(32'h3a8d924d),
	.w4(32'h3ac22c9e),
	.w5(32'h3a030bdd),
	.w6(32'hbae0df38),
	.w7(32'hbb06c3d6),
	.w8(32'h39539b1f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ed358),
	.w1(32'hb98c5f01),
	.w2(32'hba110c63),
	.w3(32'h3a22aeb6),
	.w4(32'h39bab9ed),
	.w5(32'h39477f44),
	.w6(32'h39647316),
	.w7(32'h3920ec2d),
	.w8(32'h395b226f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee35d9),
	.w1(32'hb9b6b7ed),
	.w2(32'h3ab7e974),
	.w3(32'hbbfc222f),
	.w4(32'hbbd9efb8),
	.w5(32'hbb914f72),
	.w6(32'hbb686f22),
	.w7(32'hbab73378),
	.w8(32'hb85537b0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade5c3b),
	.w1(32'hbacd6eb8),
	.w2(32'hbb292700),
	.w3(32'hb9d26185),
	.w4(32'hbba146a3),
	.w5(32'hbb3dbc4e),
	.w6(32'hb96a9270),
	.w7(32'hbafb1b1c),
	.w8(32'hbaf3ec3c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f9e0f),
	.w1(32'hbb0b3be4),
	.w2(32'hbb5a0fe5),
	.w3(32'hbaa7cc78),
	.w4(32'hbb48a97d),
	.w5(32'hbb9aae21),
	.w6(32'hbac1b5b9),
	.w7(32'hbb80e36a),
	.w8(32'hbbb4d692),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28dc7c),
	.w1(32'hba264f06),
	.w2(32'h3aa0e780),
	.w3(32'hbb733b43),
	.w4(32'hbb94dac0),
	.w5(32'hbb5247d7),
	.w6(32'hbb550a68),
	.w7(32'hbb647867),
	.w8(32'hba9d29a6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803eff),
	.w1(32'h3b806990),
	.w2(32'h3b5bf5c6),
	.w3(32'h3ad73ce2),
	.w4(32'h3a76c86d),
	.w5(32'hb9a38cb1),
	.w6(32'h3b3787fb),
	.w7(32'h3b2f8a25),
	.w8(32'hb8c60970),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf27974),
	.w1(32'h3a89f28f),
	.w2(32'h3b2f649c),
	.w3(32'h39f223b2),
	.w4(32'h3a2e8dfe),
	.w5(32'h3a4642f6),
	.w6(32'hb9d90bef),
	.w7(32'h3b17237f),
	.w8(32'h3b6a3543),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d099f8),
	.w1(32'h381509dd),
	.w2(32'h383a87e2),
	.w3(32'h397e44ca),
	.w4(32'h38253688),
	.w5(32'h390a75d7),
	.w6(32'hb8f64770),
	.w7(32'hb9153886),
	.w8(32'hba8be551),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca70d),
	.w1(32'hbb7031c2),
	.w2(32'hb9185896),
	.w3(32'hbb93de16),
	.w4(32'hbc4e6980),
	.w5(32'hbc65937a),
	.w6(32'hbbb61877),
	.w7(32'hbbdef317),
	.w8(32'hbb39b351),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b24e4),
	.w1(32'h394c0ec0),
	.w2(32'hb6dafdb2),
	.w3(32'hb55f983d),
	.w4(32'h389ebfb5),
	.w5(32'h37069ccd),
	.w6(32'h395093ef),
	.w7(32'h386566dc),
	.w8(32'h36eda272),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32652b),
	.w1(32'hbb0aa2d6),
	.w2(32'hba890670),
	.w3(32'hbb9cd80b),
	.w4(32'hbba906a9),
	.w5(32'hbb9c5a07),
	.w6(32'hbb7ee89c),
	.w7(32'hbb9f5a3d),
	.w8(32'hbb8b4d8c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38425fae),
	.w1(32'hb78bc6a1),
	.w2(32'hb70b025f),
	.w3(32'hb9bb279f),
	.w4(32'hb99a0828),
	.w5(32'hb8617ff1),
	.w6(32'hb8eb532a),
	.w7(32'hb95d4901),
	.w8(32'hbac89403),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad38ef1),
	.w1(32'h3b7b80b2),
	.w2(32'hba975b23),
	.w3(32'h3b5fb602),
	.w4(32'h3b605403),
	.w5(32'h3a3f6faf),
	.w6(32'hbb1bf1fd),
	.w7(32'hb956460c),
	.w8(32'hbaaf79fd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d68f4a),
	.w1(32'hb91b6600),
	.w2(32'hb9977fad),
	.w3(32'hb917b79b),
	.w4(32'hb9a496ad),
	.w5(32'hb994dfb6),
	.w6(32'hb931a66c),
	.w7(32'hb93b19b8),
	.w8(32'h38a6f15f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162645),
	.w1(32'hb8e2a491),
	.w2(32'hbae24a34),
	.w3(32'hba210f63),
	.w4(32'hba193971),
	.w5(32'hbaef1217),
	.w6(32'hbb2c4a31),
	.w7(32'hbb94623a),
	.w8(32'hbb91cc53),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35484eb6),
	.w1(32'hb8c709f9),
	.w2(32'hb8a0cd06),
	.w3(32'hb9133b83),
	.w4(32'hb94dada0),
	.w5(32'hb926206f),
	.w6(32'h370366d0),
	.w7(32'hb86dcb11),
	.w8(32'hbaae17ce),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b95f),
	.w1(32'hbb874e16),
	.w2(32'hba61f54a),
	.w3(32'hbbcf6ee9),
	.w4(32'hbc2ba048),
	.w5(32'hbc27cd83),
	.w6(32'hbc1748af),
	.w7(32'hbc1b1155),
	.w8(32'hbbd82fbc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9922535),
	.w1(32'h3a01c4d8),
	.w2(32'h3b049567),
	.w3(32'hbaba319e),
	.w4(32'hb8dfa90b),
	.w5(32'h3823f077),
	.w6(32'hb94217b2),
	.w7(32'h3ad34c4a),
	.w8(32'h3b8371b6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7821e74),
	.w1(32'hb9a2a228),
	.w2(32'h38929439),
	.w3(32'hb77d695d),
	.w4(32'hb8e02b8e),
	.w5(32'h381b5719),
	.w6(32'h3750c779),
	.w7(32'hb8f3933d),
	.w8(32'hb881bde2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba327d8f),
	.w1(32'h388d6d75),
	.w2(32'hba7c809c),
	.w3(32'h3a61efc2),
	.w4(32'h3a22b283),
	.w5(32'hba8696f8),
	.w6(32'h37197271),
	.w7(32'h378b5007),
	.w8(32'hb8917c96),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934ef79),
	.w1(32'h3a441927),
	.w2(32'h3ad69a1b),
	.w3(32'hbb24e87c),
	.w4(32'hbb0841fb),
	.w5(32'hba048d89),
	.w6(32'hba4a85cf),
	.w7(32'hba1766a5),
	.w8(32'hb970f976),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01bdd6),
	.w1(32'h3adc57a1),
	.w2(32'h3b8a35a0),
	.w3(32'hbbb52a69),
	.w4(32'hbbeea56d),
	.w5(32'hbbbb5b98),
	.w6(32'hbbc84263),
	.w7(32'hbbb8054b),
	.w8(32'hbb99b1df),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c692d),
	.w1(32'hbb5210bf),
	.w2(32'hbba56db5),
	.w3(32'hbc3f7317),
	.w4(32'hbc0318d8),
	.w5(32'hbc128c5a),
	.w6(32'hbc280aa0),
	.w7(32'hbbdfc163),
	.w8(32'hbb149fae),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb707ccf),
	.w1(32'hbb819937),
	.w2(32'hbb308455),
	.w3(32'hbc27d972),
	.w4(32'hbc81953a),
	.w5(32'hbc915e8c),
	.w6(32'hbc529727),
	.w7(32'hbc761319),
	.w8(32'hbc6bfa91),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2287e2),
	.w1(32'hba80d34b),
	.w2(32'h3a917c28),
	.w3(32'hbbcf4f2d),
	.w4(32'hbc0358d6),
	.w5(32'hbc18385b),
	.w6(32'hbae360f4),
	.w7(32'hbba0e9fd),
	.w8(32'hbbf5bb0a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4fd68),
	.w1(32'h39085c8d),
	.w2(32'h39b87051),
	.w3(32'h3a00ee4e),
	.w4(32'h39ba3370),
	.w5(32'h3a1fe347),
	.w6(32'h39d3c88a),
	.w7(32'h38963be8),
	.w8(32'hb9bcc956),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c8150),
	.w1(32'hba3b9af9),
	.w2(32'hb92f1219),
	.w3(32'hb9a2426e),
	.w4(32'hb9f36867),
	.w5(32'hb92e698e),
	.w6(32'hb9f92725),
	.w7(32'hb94d251e),
	.w8(32'hb97dbfa4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39591933),
	.w1(32'h3969ae67),
	.w2(32'h376249e9),
	.w3(32'h39f12401),
	.w4(32'hb95fe64e),
	.w5(32'hb7f951b3),
	.w6(32'h384cd448),
	.w7(32'h38dbcaac),
	.w8(32'h39cfd6f0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e30382),
	.w1(32'hbafffe6c),
	.w2(32'hbb6876bd),
	.w3(32'hbb0f0513),
	.w4(32'hbb4a45e9),
	.w5(32'hbb47465d),
	.w6(32'hbb212e77),
	.w7(32'hbbbaa376),
	.w8(32'hbbd5caac),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8628d),
	.w1(32'h3a279d24),
	.w2(32'h3979a843),
	.w3(32'hba879a29),
	.w4(32'hba995225),
	.w5(32'hba94ea99),
	.w6(32'hb99becf8),
	.w7(32'hb8461c29),
	.w8(32'hba8349e2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9639c),
	.w1(32'hba9d1254),
	.w2(32'hbac47984),
	.w3(32'hb838bc8f),
	.w4(32'hba3496dc),
	.w5(32'hba6807a4),
	.w6(32'hba7eb3f4),
	.w7(32'hbabf56ae),
	.w8(32'hbb241fb6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39474aa9),
	.w1(32'h3a049ab9),
	.w2(32'h3a32b282),
	.w3(32'hbb4b42b9),
	.w4(32'hbb34ffe5),
	.w5(32'hbaf25374),
	.w6(32'hba8d1e1c),
	.w7(32'hb9c4740f),
	.w8(32'h3a80b3f1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ed008),
	.w1(32'hb9a6a9e3),
	.w2(32'h3a17468a),
	.w3(32'hbb2ec86e),
	.w4(32'hbb2e8da9),
	.w5(32'hbad9bdf4),
	.w6(32'hbafa0481),
	.w7(32'hbab1490d),
	.w8(32'hb980085b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa34485),
	.w1(32'hb9c0eca1),
	.w2(32'h3a71cef0),
	.w3(32'h390cc98a),
	.w4(32'h3a3ac254),
	.w5(32'h39ffc7bd),
	.w6(32'h380fae9d),
	.w7(32'h3a95f00b),
	.w8(32'h3a82bdba),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb821d062),
	.w1(32'h39722764),
	.w2(32'h3b848e00),
	.w3(32'hbb06c7ec),
	.w4(32'hbb1b66e6),
	.w5(32'h3a38cec4),
	.w6(32'hbae9f2a1),
	.w7(32'hbb0732a9),
	.w8(32'h3a7d4dc0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cfa33),
	.w1(32'h39bf3737),
	.w2(32'hba915797),
	.w3(32'hbb489725),
	.w4(32'hbb4cbd69),
	.w5(32'hbbd01dbb),
	.w6(32'h38944322),
	.w7(32'hbb99392b),
	.w8(32'hbbc4ba63),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a68a2c),
	.w1(32'hba876222),
	.w2(32'hbaa696c6),
	.w3(32'hba6c2770),
	.w4(32'hbae17161),
	.w5(32'hbab621c2),
	.w6(32'h3a4389e7),
	.w7(32'h3a4b21ff),
	.w8(32'hbaa39f41),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba242d38),
	.w1(32'hb9e8501a),
	.w2(32'hba050063),
	.w3(32'hba6976c9),
	.w4(32'hba395432),
	.w5(32'hba70739f),
	.w6(32'hba4c30c0),
	.w7(32'hba1afac6),
	.w8(32'hb9cf2573),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c2932),
	.w1(32'hba278ab2),
	.w2(32'hb96e613d),
	.w3(32'hb9e646e0),
	.w4(32'hb9f1d43f),
	.w5(32'hb92ccaa9),
	.w6(32'hb9c58a34),
	.w7(32'hb9542768),
	.w8(32'hb9b7f561),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872ef4b),
	.w1(32'hb9cccca1),
	.w2(32'hb95478ac),
	.w3(32'h39899237),
	.w4(32'hb99c8a36),
	.w5(32'hb982707d),
	.w6(32'hb9282558),
	.w7(32'hb9dbff73),
	.w8(32'hb99e73a0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f5ed6),
	.w1(32'hbac9c41d),
	.w2(32'hbb4a1be3),
	.w3(32'h39b4b77c),
	.w4(32'hba74e365),
	.w5(32'hbb33f40b),
	.w6(32'hbafcc162),
	.w7(32'hbb3f856b),
	.w8(32'hbba75df9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc57c4),
	.w1(32'hba5b9303),
	.w2(32'hba8a90bc),
	.w3(32'hba33e5da),
	.w4(32'hba81ca43),
	.w5(32'hbacfea88),
	.w6(32'hba714cb2),
	.w7(32'hbaa60cf0),
	.w8(32'h390851e8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a676e80),
	.w1(32'h3b15953e),
	.w2(32'h3b6cd030),
	.w3(32'hba1e818f),
	.w4(32'h3ab09573),
	.w5(32'h3b480d10),
	.w6(32'h3b2b92b1),
	.w7(32'h3b30d057),
	.w8(32'h3b995fe4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f82452),
	.w1(32'hb9e0f0df),
	.w2(32'hba1d2ca7),
	.w3(32'hb9ce3e0b),
	.w4(32'hb98f69c8),
	.w5(32'hb8adb9f3),
	.w6(32'hb8c54692),
	.w7(32'h38f0b6bc),
	.w8(32'h3b66bbf4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878739),
	.w1(32'h3b8c8d93),
	.w2(32'h3b95a8ab),
	.w3(32'hbae59aa7),
	.w4(32'hbb89a0b3),
	.w5(32'hbbb16033),
	.w6(32'hbb02b574),
	.w7(32'hbb938745),
	.w8(32'hb9a62c70),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83e391),
	.w1(32'hbb5d1615),
	.w2(32'h3bd8884a),
	.w3(32'h3b53bcb8),
	.w4(32'hbbd999b9),
	.w5(32'hbaaa96e6),
	.w6(32'hbbc30e42),
	.w7(32'hbaf9e12e),
	.w8(32'hbbec09a4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05c1a2),
	.w1(32'h3b0dda35),
	.w2(32'h3b265a46),
	.w3(32'h3aa83ff3),
	.w4(32'h3a06134f),
	.w5(32'h399de50f),
	.w6(32'h3ac9b547),
	.w7(32'h3b1d4959),
	.w8(32'hbafd79fb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c77e2),
	.w1(32'h3b260c1e),
	.w2(32'hba20fbed),
	.w3(32'hbb10f1ef),
	.w4(32'hba79ebd1),
	.w5(32'hbb412d93),
	.w6(32'h3a2872f7),
	.w7(32'hba5f27f7),
	.w8(32'h3986b73f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d224),
	.w1(32'h3c4566c2),
	.w2(32'h3b668c65),
	.w3(32'h3b89adf0),
	.w4(32'h3bcc4291),
	.w5(32'hb9f12fe5),
	.w6(32'h3b4ae2c3),
	.w7(32'hbbb81140),
	.w8(32'hbb7efecc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab07e6b),
	.w1(32'h3c275204),
	.w2(32'h3bd4dbc4),
	.w3(32'h3ba61370),
	.w4(32'h3c36c315),
	.w5(32'h3bf2943c),
	.w6(32'h3b7579b3),
	.w7(32'h3b8cf120),
	.w8(32'h3ba8f742),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71edc4),
	.w1(32'h3c2def2c),
	.w2(32'h3bcfc46f),
	.w3(32'hbb1499f3),
	.w4(32'h3b47fa79),
	.w5(32'h3a992137),
	.w6(32'h3bc2a0cc),
	.w7(32'h3acaefba),
	.w8(32'h3b8fbf2e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58a84b),
	.w1(32'hbbb3b75f),
	.w2(32'hbb9cde2f),
	.w3(32'h3ad3f664),
	.w4(32'hba9c4a2f),
	.w5(32'hbb155739),
	.w6(32'hbb8885ef),
	.w7(32'hbabd3c66),
	.w8(32'h3870c249),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dd893),
	.w1(32'h3c0ac3b0),
	.w2(32'h3b3c51c9),
	.w3(32'h3a1a4e34),
	.w4(32'h3b1cb2bf),
	.w5(32'hba20400e),
	.w6(32'h3b2f6ef3),
	.w7(32'hba71900e),
	.w8(32'h39f096a0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa73146),
	.w1(32'h3acafa84),
	.w2(32'h3a4bbb49),
	.w3(32'h37a14ab6),
	.w4(32'hb90dd9c0),
	.w5(32'hba0e4956),
	.w6(32'h3a390ed7),
	.w7(32'hba114be2),
	.w8(32'h3a3bd424),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d432),
	.w1(32'h3b72950f),
	.w2(32'h3accaba0),
	.w3(32'h3b58ec37),
	.w4(32'h3b184799),
	.w5(32'h392eb514),
	.w6(32'h3ad085f8),
	.w7(32'hb9afbcb0),
	.w8(32'h393f055f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b321dd9),
	.w1(32'hbc13c339),
	.w2(32'hbc4c81ca),
	.w3(32'hba6a6ec4),
	.w4(32'hbb90049f),
	.w5(32'hbc3f227b),
	.w6(32'hbc20a12e),
	.w7(32'hbc306b37),
	.w8(32'h3af9cc58),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77f898),
	.w1(32'h3aaef53f),
	.w2(32'h391f6d27),
	.w3(32'hbb8a23af),
	.w4(32'hbb0860bf),
	.w5(32'hbb3c290a),
	.w6(32'hba9f7f1c),
	.w7(32'hbac4753f),
	.w8(32'h3a71e8db),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989ef42),
	.w1(32'h3bc71c76),
	.w2(32'h3c26d319),
	.w3(32'hbb0942dd),
	.w4(32'h3b89d014),
	.w5(32'h3bb97f58),
	.w6(32'h3be866cb),
	.w7(32'h3c2d0ae6),
	.w8(32'hb90a898f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954080c),
	.w1(32'hbaabb23c),
	.w2(32'hbb8370ab),
	.w3(32'hba6864ec),
	.w4(32'hbbbca5af),
	.w5(32'hbbf7811d),
	.w6(32'hb955a1d8),
	.w7(32'hbb725dcc),
	.w8(32'hbb724e3c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c1362),
	.w1(32'h3a91a0a8),
	.w2(32'hb6fcfa33),
	.w3(32'hba9f80c8),
	.w4(32'hbab4f43e),
	.w5(32'h3a99857c),
	.w6(32'hbad8222a),
	.w7(32'hbb191d2e),
	.w8(32'hba2e58d6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30b505),
	.w1(32'h3b22e899),
	.w2(32'h3b9e21a6),
	.w3(32'h3bf18fb0),
	.w4(32'h3ba41c61),
	.w5(32'h3b6a18e5),
	.w6(32'h3bd1ea7b),
	.w7(32'h3b1a64fe),
	.w8(32'hbad460f5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ee9a8),
	.w1(32'hbb030e8b),
	.w2(32'h39d0d68b),
	.w3(32'hbb0a1fb3),
	.w4(32'hbb1e868b),
	.w5(32'hb9f8ed3a),
	.w6(32'hba88181a),
	.w7(32'h382e644b),
	.w8(32'h3b339f5a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63a70f),
	.w1(32'h3b5ad17d),
	.w2(32'h3a89a9dc),
	.w3(32'h3b38d046),
	.w4(32'h3b3a9625),
	.w5(32'h3abb7d3a),
	.w6(32'h3a3e823e),
	.w7(32'h39b4fb88),
	.w8(32'hbaa701b6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d23cf),
	.w1(32'hba799fc4),
	.w2(32'hbab558c9),
	.w3(32'h3b03c1b2),
	.w4(32'h3bc5bcc9),
	.w5(32'h3b0a831a),
	.w6(32'hb8f0a634),
	.w7(32'hbb0b37a7),
	.w8(32'h3b474eca),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd960),
	.w1(32'h3c71090a),
	.w2(32'h3b92c7d4),
	.w3(32'h3a6bca86),
	.w4(32'h3addc034),
	.w5(32'hbb8cc302),
	.w6(32'h3c338943),
	.w7(32'h3a9be49c),
	.w8(32'h3a31c999),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e11165),
	.w1(32'h3bc1bb70),
	.w2(32'h3abde3ab),
	.w3(32'hb9f37745),
	.w4(32'h3b72f74b),
	.w5(32'h3a42bda2),
	.w6(32'h3b44b371),
	.w7(32'hba1ba5db),
	.w8(32'hbacb1695),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c6eb),
	.w1(32'hbbc3fbc9),
	.w2(32'hbb649e15),
	.w3(32'hbbc3793a),
	.w4(32'hbadf8c23),
	.w5(32'h39636f70),
	.w6(32'hb9d89b49),
	.w7(32'hbab1344c),
	.w8(32'h3bf84d0e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule