module layer_8_featuremap_67(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bf0e2),
	.w1(32'h3bcf5c28),
	.w2(32'h3bee12ef),
	.w3(32'hbc2062bd),
	.w4(32'h3a9bd1f4),
	.w5(32'h3b304451),
	.w6(32'hbc1ded0f),
	.w7(32'hbbc91450),
	.w8(32'hbc0a9564),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74daca),
	.w1(32'h3af54d35),
	.w2(32'h3b88cf72),
	.w3(32'hbb0af452),
	.w4(32'hbab47557),
	.w5(32'hb9d9d7e2),
	.w6(32'h3a1f1deb),
	.w7(32'h3aaf94ba),
	.w8(32'hbb023729),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85213a),
	.w1(32'hb9f50dfe),
	.w2(32'h3a17410f),
	.w3(32'h3b1a5d86),
	.w4(32'hba21edb7),
	.w5(32'hba04dc5d),
	.w6(32'h3b983998),
	.w7(32'h3b90b979),
	.w8(32'h3af3643f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab04372),
	.w1(32'hbbdc17eb),
	.w2(32'hbb944ea8),
	.w3(32'hbbf6386f),
	.w4(32'hb9a4d075),
	.w5(32'hba9e85a3),
	.w6(32'hbc731442),
	.w7(32'hbc3f478e),
	.w8(32'hbb707e47),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1442a6),
	.w1(32'h3bfc2d2a),
	.w2(32'h3c2c34cd),
	.w3(32'h38a4daf7),
	.w4(32'h3b72aa01),
	.w5(32'h3bfb933c),
	.w6(32'h3b1d12a2),
	.w7(32'h3ba09c88),
	.w8(32'h3bfe3bdd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f2b2),
	.w1(32'hbbae4b4f),
	.w2(32'hbb89ed55),
	.w3(32'h3c064ff4),
	.w4(32'h3be22473),
	.w5(32'h3c112edc),
	.w6(32'h3bb8d483),
	.w7(32'h3c086600),
	.w8(32'h3afa5120),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025d15),
	.w1(32'hba314969),
	.w2(32'h3afab125),
	.w3(32'hbb86d575),
	.w4(32'hbb549b12),
	.w5(32'hba31e9b8),
	.w6(32'hbae2257f),
	.w7(32'hb9016941),
	.w8(32'h3a34f7c5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdce368),
	.w1(32'h3bf3e4c6),
	.w2(32'h3c0e3178),
	.w3(32'h3bac7b76),
	.w4(32'h3c0b6dfa),
	.w5(32'h3c1ee30f),
	.w6(32'h3aaa3f67),
	.w7(32'h3ac2267e),
	.w8(32'hbb32301d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa47e5),
	.w1(32'h3bfa1294),
	.w2(32'h3c412913),
	.w3(32'hba57b2c7),
	.w4(32'h3793e8e2),
	.w5(32'h3b5bbbc6),
	.w6(32'h3a989ed8),
	.w7(32'h3b427f91),
	.w8(32'h3b95bc22),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ce5bb),
	.w1(32'h3c1f502a),
	.w2(32'hba445c53),
	.w3(32'hbc04f1ff),
	.w4(32'hbb7c1675),
	.w5(32'h3b0da911),
	.w6(32'hbb3c3bd7),
	.w7(32'hbbc3d376),
	.w8(32'hbb59a103),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf881),
	.w1(32'h3be21833),
	.w2(32'h3bed3a2e),
	.w3(32'hbb783504),
	.w4(32'h3be6ae50),
	.w5(32'h3c229c00),
	.w6(32'hbc3c825b),
	.w7(32'hbc11baa3),
	.w8(32'hbbc998f9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6ec7),
	.w1(32'h3bcd6888),
	.w2(32'h3bc5f570),
	.w3(32'hbc0c1aa9),
	.w4(32'hbb7d92ac),
	.w5(32'hb973dafa),
	.w6(32'hbc05c916),
	.w7(32'hbb9dc7a2),
	.w8(32'hbb944af8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a7ad),
	.w1(32'hbac53726),
	.w2(32'h3a6b3d94),
	.w3(32'hbb876a5c),
	.w4(32'hbbc2e97d),
	.w5(32'hbb694774),
	.w6(32'h3a2f97b7),
	.w7(32'h3a6b55e2),
	.w8(32'h3ade82c7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23a2a2),
	.w1(32'h3aa38aeb),
	.w2(32'h3b9c98fe),
	.w3(32'h3ad98ee7),
	.w4(32'h3b217ed8),
	.w5(32'h3bcd14e8),
	.w6(32'h3b6e19e7),
	.w7(32'h3bbfe649),
	.w8(32'h3ac26d5e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39033073),
	.w1(32'h3a809f1a),
	.w2(32'h3b20488c),
	.w3(32'h38db4c27),
	.w4(32'h3a43cf28),
	.w5(32'h3b53295d),
	.w6(32'h3ade401e),
	.w7(32'h3b14e38d),
	.w8(32'hba1ded25),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cb747),
	.w1(32'h3a8f90cd),
	.w2(32'h3a522855),
	.w3(32'hbab8c9a5),
	.w4(32'hba88a3e7),
	.w5(32'hb9f812d5),
	.w6(32'hb914179b),
	.w7(32'hb9e751f1),
	.w8(32'h3a1e8b78),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6170f4),
	.w1(32'hba97a83d),
	.w2(32'hbb26a657),
	.w3(32'h3c073a2f),
	.w4(32'h3c151c1f),
	.w5(32'h3bc9d768),
	.w6(32'h3aff439c),
	.w7(32'h3af482a7),
	.w8(32'hbad76a19),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2339b9),
	.w1(32'h3ba4589a),
	.w2(32'h3bd8e7eb),
	.w3(32'hbb0b3207),
	.w4(32'hba2c84fb),
	.w5(32'h3ad9330b),
	.w6(32'hbb30eb4a),
	.w7(32'h3acdcda3),
	.w8(32'hbb9208b6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d033c59),
	.w1(32'h3d293a81),
	.w2(32'h3c3e0461),
	.w3(32'hbc735bbf),
	.w4(32'h3cc141a5),
	.w5(32'h3b6ec50e),
	.w6(32'hbcb23fa3),
	.w7(32'hbcc29ced),
	.w8(32'hbd02093d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47f32e),
	.w1(32'h3c04abe2),
	.w2(32'hbb610344),
	.w3(32'h3ab22259),
	.w4(32'hbb4efa8c),
	.w5(32'hbc160591),
	.w6(32'hbbb2bcc3),
	.w7(32'hbb9a0a96),
	.w8(32'hbc2976f9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf05dfc),
	.w1(32'hbb2eeee8),
	.w2(32'h39a0c2dd),
	.w3(32'hbc04cf31),
	.w4(32'hbb887bb3),
	.w5(32'hb9e32828),
	.w6(32'h3b8c5acf),
	.w7(32'h388bf0d2),
	.w8(32'hbbef19b0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e322),
	.w1(32'hbb71f1e9),
	.w2(32'h3a17699f),
	.w3(32'hbb14a3c9),
	.w4(32'hbb8fc834),
	.w5(32'hb9816ef6),
	.w6(32'h3b6b022a),
	.w7(32'h3b135579),
	.w8(32'h3a692f4e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6d41a),
	.w1(32'h3c45ef3a),
	.w2(32'h3b8a4ce9),
	.w3(32'hbc7dc8a0),
	.w4(32'h3c0046c7),
	.w5(32'h3bf98928),
	.w6(32'hbcd433f1),
	.w7(32'hbcaf5edf),
	.w8(32'hbcb925b1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3319ce),
	.w1(32'hbc074a2b),
	.w2(32'h3b7fdc70),
	.w3(32'hbc24be1f),
	.w4(32'hbb8aa00c),
	.w5(32'h3b30707b),
	.w6(32'hbb0f292c),
	.w7(32'h3ac49ae4),
	.w8(32'hbb8fa476),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974feb),
	.w1(32'hbb42006f),
	.w2(32'hbbabe061),
	.w3(32'hbb825439),
	.w4(32'hbb34cff6),
	.w5(32'hbb623908),
	.w6(32'hbb535014),
	.w7(32'hbb808950),
	.w8(32'h3b814394),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c838f),
	.w1(32'h3c445836),
	.w2(32'h3bfa1e0a),
	.w3(32'hbbce06d5),
	.w4(32'h3b68da3a),
	.w5(32'h3b78149c),
	.w6(32'hbc84975e),
	.w7(32'hbc082cd0),
	.w8(32'hbc03c609),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90188a),
	.w1(32'hba199b34),
	.w2(32'h39c3182a),
	.w3(32'h3a53bda1),
	.w4(32'hba8f207b),
	.w5(32'hba1ad146),
	.w6(32'h3aaf34b3),
	.w7(32'h3b612437),
	.w8(32'hba268e24),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d925806),
	.w1(32'h3d9b6522),
	.w2(32'h3c81ac8e),
	.w3(32'hbd4f76fa),
	.w4(32'h3c9d4677),
	.w5(32'h3d5cc6fc),
	.w6(32'hbd1358bb),
	.w7(32'hbdcade6e),
	.w8(32'hbdd866b9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9396),
	.w1(32'h3c22d9fe),
	.w2(32'h3bed969d),
	.w3(32'hbbe14778),
	.w4(32'h3b629433),
	.w5(32'h3aff6d42),
	.w6(32'hbbda181d),
	.w7(32'hbc2140b5),
	.w8(32'hbbcc5dbc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c545dd),
	.w1(32'hba74e5da),
	.w2(32'h3adcdcf1),
	.w3(32'hb9c1514c),
	.w4(32'hba442f90),
	.w5(32'h3a6a285e),
	.w6(32'hba066181),
	.w7(32'h38736964),
	.w8(32'hbb77b3e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c12908),
	.w1(32'h3b14db85),
	.w2(32'hbbccbdef),
	.w3(32'hbaf5d0b0),
	.w4(32'hba6f8453),
	.w5(32'h3a8b5e50),
	.w6(32'hbb742ace),
	.w7(32'hbbd7697c),
	.w8(32'hbae2d755),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801a64),
	.w1(32'hba04ec3b),
	.w2(32'h3afa4d78),
	.w3(32'hbb7dbe55),
	.w4(32'hbb68fffc),
	.w5(32'hbb8077d3),
	.w6(32'hba7e48ea),
	.w7(32'h3a713b3e),
	.w8(32'h386692b5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad78a9e),
	.w1(32'h3b35aa1f),
	.w2(32'h3aff0d91),
	.w3(32'hbb5d3174),
	.w4(32'h3ac6082d),
	.w5(32'h3b543f1d),
	.w6(32'h3b2509ba),
	.w7(32'hbacdbb3a),
	.w8(32'h3b00de54),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10207f),
	.w1(32'hba8114bc),
	.w2(32'hbb5ede71),
	.w3(32'hba37f8e4),
	.w4(32'h39e6758e),
	.w5(32'h3b2b5d3d),
	.w6(32'h3b007fd6),
	.w7(32'hb8726a2c),
	.w8(32'h3b682f0f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575b94),
	.w1(32'hbc3ceadf),
	.w2(32'hbb68c934),
	.w3(32'hbbd2205f),
	.w4(32'hbbf5f6de),
	.w5(32'hbaa706c3),
	.w6(32'h3bee9ee6),
	.w7(32'h3c05beb6),
	.w8(32'hbb4d301c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e4dd9),
	.w1(32'h3c2e91d0),
	.w2(32'h3c409e22),
	.w3(32'hbc32af8c),
	.w4(32'h3aae321a),
	.w5(32'h3b809f3d),
	.w6(32'hbc047742),
	.w7(32'hbb964a7a),
	.w8(32'hbc3499e7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18282b),
	.w1(32'hbb4dad5b),
	.w2(32'hbb7dda22),
	.w3(32'hbb40d116),
	.w4(32'hbb4174e6),
	.w5(32'hbb990ef7),
	.w6(32'hbb255055),
	.w7(32'hbb74b203),
	.w8(32'hbad965ac),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8865b4),
	.w1(32'h3b124f6b),
	.w2(32'h3c03697f),
	.w3(32'h3a1edafa),
	.w4(32'hb9e42901),
	.w5(32'h3b504b2e),
	.w6(32'h399a1078),
	.w7(32'h3b0bd771),
	.w8(32'h3bb172d1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e418b),
	.w1(32'h3b1c6fc1),
	.w2(32'h3ba50c40),
	.w3(32'h398f9c4f),
	.w4(32'h3ab7045f),
	.w5(32'h3bdcbb7e),
	.w6(32'h3b82e25e),
	.w7(32'h3ba0d3ef),
	.w8(32'hbb114069),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0633),
	.w1(32'hbb744e53),
	.w2(32'hbb735bca),
	.w3(32'hbb800213),
	.w4(32'hbb93fa9a),
	.w5(32'hbb8f15bf),
	.w6(32'hbb45b382),
	.w7(32'hbb45d057),
	.w8(32'h39c5510f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0094a9),
	.w1(32'h3b911307),
	.w2(32'hbc1958d0),
	.w3(32'hba89fb25),
	.w4(32'h3b665c8e),
	.w5(32'hb99df6a8),
	.w6(32'hbcb9411e),
	.w7(32'hbc961ec1),
	.w8(32'hbc827ba9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fc76e),
	.w1(32'h3afa8a1c),
	.w2(32'hbacbfe70),
	.w3(32'h3a3299a7),
	.w4(32'h3b0091ef),
	.w5(32'hbb1b670d),
	.w6(32'h39c6fd70),
	.w7(32'hbb57cca5),
	.w8(32'hbb964eaa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775a31),
	.w1(32'hbac83070),
	.w2(32'hbadaa1f7),
	.w3(32'hb8101e6d),
	.w4(32'hba5c82d6),
	.w5(32'hba8674dc),
	.w6(32'h3a8d4b60),
	.w7(32'h3831f36b),
	.w8(32'hba72ca19),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93c1d),
	.w1(32'h3a1339a1),
	.w2(32'hba9fed3d),
	.w3(32'hba9114f8),
	.w4(32'h3b6d3bc5),
	.w5(32'h3b868eb6),
	.w6(32'hbc15c9c6),
	.w7(32'hbbf3fe70),
	.w8(32'hbbaa03a2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9c68),
	.w1(32'h3be5d7da),
	.w2(32'hbb448424),
	.w3(32'h3b43759b),
	.w4(32'h3c53e799),
	.w5(32'h3ba79557),
	.w6(32'hbc5dfdcf),
	.w7(32'hbc3be036),
	.w8(32'hbc5bea2a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac69f6c),
	.w1(32'hbac302cc),
	.w2(32'hbb6ef928),
	.w3(32'hbb803aba),
	.w4(32'hbb834e46),
	.w5(32'hbbbd8394),
	.w6(32'hba50e9b2),
	.w7(32'hbbc53ec0),
	.w8(32'hbbda5bdf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77525c1),
	.w1(32'h37184101),
	.w2(32'h372555c4),
	.w3(32'hb73a6355),
	.w4(32'h37151aa1),
	.w5(32'h36ec32b1),
	.w6(32'hb7141390),
	.w7(32'h3781475a),
	.w8(32'h37e5bd81),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba321249),
	.w1(32'h3a9556a9),
	.w2(32'hbba81ce1),
	.w3(32'hbbc4a6c9),
	.w4(32'h3b61a4cc),
	.w5(32'hbafc4076),
	.w6(32'hbc1f820e),
	.w7(32'hbc6f09f8),
	.w8(32'hbc96799e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95417f5),
	.w1(32'hba0b2dbf),
	.w2(32'hbb0522ea),
	.w3(32'hb884c484),
	.w4(32'hba0c8f23),
	.w5(32'hba402954),
	.w6(32'hba824797),
	.w7(32'hbaae2672),
	.w8(32'hbadac9e5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba451e75),
	.w1(32'h3a548238),
	.w2(32'hbaca93e8),
	.w3(32'hbb6acd4a),
	.w4(32'h3b9fd4fc),
	.w5(32'h3aee81a6),
	.w6(32'hbc8e20d6),
	.w7(32'hbc44f9cf),
	.w8(32'hbb9b9f4f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba3985),
	.w1(32'hbad1bb46),
	.w2(32'hba975633),
	.w3(32'h3b890a81),
	.w4(32'hbbebba8d),
	.w5(32'hbbf19749),
	.w6(32'h3c6220af),
	.w7(32'h3992650a),
	.w8(32'hbbb5eea5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92cdf6),
	.w1(32'h3c8cfab6),
	.w2(32'hbc3101b3),
	.w3(32'h3cc2606c),
	.w4(32'h3d17dba9),
	.w5(32'h3c5dc217),
	.w6(32'hbcd93c08),
	.w7(32'hbc443b83),
	.w8(32'hbca5a824),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c005db7),
	.w1(32'h3c2ab388),
	.w2(32'h3bc8ab53),
	.w3(32'h3ba1fb4b),
	.w4(32'h3c08398e),
	.w5(32'h3beba0e9),
	.w6(32'hbbc14d82),
	.w7(32'hbb733ec7),
	.w8(32'hbaebff17),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cb5f0),
	.w1(32'h39fdc6c0),
	.w2(32'h3b1d7c16),
	.w3(32'hbbd8ea34),
	.w4(32'hbbb5d0ef),
	.w5(32'hbc07872b),
	.w6(32'hbab129b3),
	.w7(32'h3a8a0354),
	.w8(32'hba9dbb44),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e0f83),
	.w1(32'h38ee939b),
	.w2(32'h38d2fc40),
	.w3(32'hb703a040),
	.w4(32'h3877354d),
	.w5(32'h38ba45d2),
	.w6(32'h37a50220),
	.w7(32'h388a1690),
	.w8(32'h38b85462),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19d7f1),
	.w1(32'h3b881409),
	.w2(32'h3a8cb86a),
	.w3(32'hbc9d797c),
	.w4(32'hbc021b3a),
	.w5(32'hbb326040),
	.w6(32'hbb6fdebc),
	.w7(32'hbc87c37e),
	.w8(32'hbc84d4e1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74a22),
	.w1(32'hbb9330a2),
	.w2(32'hbb0f3afb),
	.w3(32'hbb7c9daf),
	.w4(32'hbbb0d225),
	.w5(32'hbb986903),
	.w6(32'hbab89bf6),
	.w7(32'hbb27f1cd),
	.w8(32'hbb3e73be),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd90dfe),
	.w1(32'h3c02cea3),
	.w2(32'h3a9639a2),
	.w3(32'h3c5729a2),
	.w4(32'h3c82ea15),
	.w5(32'h3bda4ed4),
	.w6(32'hbbc3a47c),
	.w7(32'hbaa0ece4),
	.w8(32'hbb6d852d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4634),
	.w1(32'h3b6e924e),
	.w2(32'hbb183a5e),
	.w3(32'h3abc4acf),
	.w4(32'h3bdf851c),
	.w5(32'h3bb65fc7),
	.w6(32'hbb957ad9),
	.w7(32'hbbaacf38),
	.w8(32'hbba86bb0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59856),
	.w1(32'hbbf881fa),
	.w2(32'hbc1652c7),
	.w3(32'hbb9e0d98),
	.w4(32'hbb414edc),
	.w5(32'hbb8dc95d),
	.w6(32'hbc2ff1be),
	.w7(32'hbbc81539),
	.w8(32'hbc08ea68),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6014),
	.w1(32'h3a2b1ecf),
	.w2(32'h39d27066),
	.w3(32'h3a5c228f),
	.w4(32'h3a4c75a8),
	.w5(32'h3a0ce26e),
	.w6(32'h3a06dd3f),
	.w7(32'h3a3292d5),
	.w8(32'h3a041825),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848abe9),
	.w1(32'hba129480),
	.w2(32'hba5a45db),
	.w3(32'hb89fd218),
	.w4(32'hb9c36d49),
	.w5(32'hba0aae6b),
	.w6(32'hba213312),
	.w7(32'hba8945a3),
	.w8(32'hba580f59),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4df04d),
	.w1(32'h3c2160ad),
	.w2(32'h3b4c2058),
	.w3(32'hbbcbfaf1),
	.w4(32'hbb31c661),
	.w5(32'hbb89ff2a),
	.w6(32'hbc236f04),
	.w7(32'hbc6ba628),
	.w8(32'hbc37b79b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4484),
	.w1(32'hbabc3543),
	.w2(32'hbb106879),
	.w3(32'h3ae248bd),
	.w4(32'h3b0ebb79),
	.w5(32'hba3960a8),
	.w6(32'hb94f0b16),
	.w7(32'h3aca0ced),
	.w8(32'hbac33b92),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007ef9),
	.w1(32'hbaa77a45),
	.w2(32'hba6290ba),
	.w3(32'hbaed9731),
	.w4(32'hba516b3c),
	.w5(32'hba2edf2b),
	.w6(32'hbb5a4d7e),
	.w7(32'hbb0b993a),
	.w8(32'hbb202d77),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59f711),
	.w1(32'h3bb19c67),
	.w2(32'h3b9e57b7),
	.w3(32'h3abc85bd),
	.w4(32'h3baa0deb),
	.w5(32'h3b938e94),
	.w6(32'h3a2621b6),
	.w7(32'hba86795d),
	.w8(32'hbb1d338a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6beea2),
	.w1(32'h3a242b6b),
	.w2(32'hbabc00e6),
	.w3(32'h3bb64f5a),
	.w4(32'h3b8f9177),
	.w5(32'h3b6bf52b),
	.w6(32'h3b561ffc),
	.w7(32'h3b0071b1),
	.w8(32'h3a4e2f69),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cce97),
	.w1(32'hba75bc50),
	.w2(32'hbb2f58b0),
	.w3(32'hbc299429),
	.w4(32'hbc1db311),
	.w5(32'hbc2a2a36),
	.w6(32'hbaed7922),
	.w7(32'hbc0f9755),
	.w8(32'hbc3757e8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a066250),
	.w1(32'h399ad713),
	.w2(32'h354dab45),
	.w3(32'h39b5b328),
	.w4(32'h39701793),
	.w5(32'hb9409378),
	.w6(32'h385a6c21),
	.w7(32'h381dab4c),
	.w8(32'hb952217c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc7e32),
	.w1(32'h3b0db76c),
	.w2(32'hbbfea545),
	.w3(32'hbb887a20),
	.w4(32'h3cc2352b),
	.w5(32'h3cbd6e1e),
	.w6(32'hbcb9aff0),
	.w7(32'hbc8d9075),
	.w8(32'hbcfeab1b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5d9d8),
	.w1(32'hb80717c0),
	.w2(32'h38240fff),
	.w3(32'h39169aad),
	.w4(32'hb6beb303),
	.w5(32'h37aa0c03),
	.w6(32'h3960795a),
	.w7(32'h38cc182f),
	.w8(32'h38f69c14),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16afa1),
	.w1(32'h3ba739f5),
	.w2(32'h3b54aedb),
	.w3(32'hbb4c766f),
	.w4(32'h3a6c13d9),
	.w5(32'h3a9629df),
	.w6(32'hbbc4fa21),
	.w7(32'hbba58673),
	.w8(32'hbbc2b282),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386606de),
	.w1(32'hb9138790),
	.w2(32'hb986c0fe),
	.w3(32'hb8df914b),
	.w4(32'hb9a6b15c),
	.w5(32'hb98483c1),
	.w6(32'hb91be661),
	.w7(32'hb9de5edc),
	.w8(32'hb9bedadb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1132),
	.w1(32'h3ba5619a),
	.w2(32'h3bd45add),
	.w3(32'hbc526e20),
	.w4(32'hbc4bcbd3),
	.w5(32'hbb9b3a44),
	.w6(32'hbb966849),
	.w7(32'hbbeccc57),
	.w8(32'hbbc6e548),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb776c5bd),
	.w1(32'h383f0d07),
	.w2(32'h37cfd66b),
	.w3(32'hb85766c5),
	.w4(32'hb6d5aa13),
	.w5(32'hb7765cb1),
	.w6(32'h36b63b66),
	.w7(32'h37eae5a8),
	.w8(32'h3791aa47),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce101f),
	.w1(32'h3be196f7),
	.w2(32'h3bba6c02),
	.w3(32'h3b56bed3),
	.w4(32'h3bb3957b),
	.w5(32'h3bd4d965),
	.w6(32'hba77f667),
	.w7(32'hba7db874),
	.w8(32'h39e1125a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de7733),
	.w1(32'h390dc316),
	.w2(32'h39099c07),
	.w3(32'hb63911e4),
	.w4(32'h37fa191d),
	.w5(32'h37ec64b2),
	.w6(32'hb6fa43c0),
	.w7(32'hb6a94cc9),
	.w8(32'hb7c69e3c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20f56a),
	.w1(32'h3c8058fe),
	.w2(32'h3bde74de),
	.w3(32'hbb71b197),
	.w4(32'h3c1df4ca),
	.w5(32'h3c0bb3ad),
	.w6(32'hbc2745db),
	.w7(32'hbc2e3d32),
	.w8(32'hbc631f8e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83de8a),
	.w1(32'hbad76e86),
	.w2(32'hbb3737ac),
	.w3(32'hbbb6981f),
	.w4(32'hbbb5fba3),
	.w5(32'hbb515e0d),
	.w6(32'h3a956cda),
	.w7(32'hbba255eb),
	.w8(32'hbb7f7719),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2711b),
	.w1(32'hb90a46dc),
	.w2(32'hb7b3d80c),
	.w3(32'h3a11b693),
	.w4(32'h39b7daf0),
	.w5(32'h3922a26b),
	.w6(32'h3a34fa3f),
	.w7(32'hb927c043),
	.w8(32'h3996e2c9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37059105),
	.w1(32'hb75e9062),
	.w2(32'hb94c8e60),
	.w3(32'h387cac8b),
	.w4(32'h38c4b36f),
	.w5(32'h36cf8b3b),
	.w6(32'hb8b9e719),
	.w7(32'hb7a5ad7a),
	.w8(32'hb8f2e6f0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf74efa),
	.w1(32'hbbcbf5fb),
	.w2(32'hbc21cecc),
	.w3(32'h3b92b5ca),
	.w4(32'h3bc9aca6),
	.w5(32'h3b25d3dc),
	.w6(32'hbb10966d),
	.w7(32'h3af5caef),
	.w8(32'hba914d86),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f676a),
	.w1(32'h3bb4e96f),
	.w2(32'hba8a49ca),
	.w3(32'hbb8a7cf5),
	.w4(32'h3b62ddf3),
	.w5(32'hba8458ac),
	.w6(32'hbc5b6375),
	.w7(32'hbc8424d6),
	.w8(32'hbc850acf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ac9e),
	.w1(32'hbc5fba8a),
	.w2(32'hbc97b6a4),
	.w3(32'hbc01907d),
	.w4(32'hbbf0a663),
	.w5(32'hbcbbfcca),
	.w6(32'hbcc14397),
	.w7(32'hbc974f4c),
	.w8(32'hbcbd4033),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40ddeb),
	.w1(32'h3c7e0e54),
	.w2(32'h3c300269),
	.w3(32'hbb15258a),
	.w4(32'h3c552bdb),
	.w5(32'h3c484298),
	.w6(32'hbcc2c2fc),
	.w7(32'hbcaa750f),
	.w8(32'hbc9fc369),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98d0d0),
	.w1(32'h3adca4f7),
	.w2(32'hbb11009d),
	.w3(32'hba55bb84),
	.w4(32'h3c208680),
	.w5(32'h3bb4ea43),
	.w6(32'hbc86ecea),
	.w7(32'hbbdfaf6b),
	.w8(32'hbb213cdd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba3a59),
	.w1(32'hb8ab8330),
	.w2(32'h37104bcf),
	.w3(32'hb9fae3a7),
	.w4(32'hb955381c),
	.w5(32'hb989f9a9),
	.w6(32'hb9977a6b),
	.w7(32'h38708c34),
	.w8(32'h38919ab0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e09d7),
	.w1(32'hb80c8286),
	.w2(32'hb62d6b70),
	.w3(32'hb8bbd50d),
	.w4(32'hb7b5ce87),
	.w5(32'hb795390e),
	.w6(32'hb83a7d90),
	.w7(32'h37ab723c),
	.w8(32'h3834efa6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad60e),
	.w1(32'hb9410c17),
	.w2(32'hb9858796),
	.w3(32'hb91c0d49),
	.w4(32'hb8bb16be),
	.w5(32'hb8c0fc75),
	.w6(32'hb7c805ca),
	.w7(32'h37ed8665),
	.w8(32'h37fca12a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae418ca),
	.w1(32'h3b25bf70),
	.w2(32'h3b953d1f),
	.w3(32'h3a54242b),
	.w4(32'h3b372b19),
	.w5(32'h3b56710c),
	.w6(32'hbb2dc7b8),
	.w7(32'hba693cf7),
	.w8(32'hba142402),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09bc71),
	.w1(32'hbb3fa614),
	.w2(32'hbb4ec0e0),
	.w3(32'hb9bf93b6),
	.w4(32'h39d195a5),
	.w5(32'h3aaeeaec),
	.w6(32'hbabf7e28),
	.w7(32'hbaca8be1),
	.w8(32'hb9965768),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b70484),
	.w1(32'hba0b51a7),
	.w2(32'h3884eb5a),
	.w3(32'hb8a9504a),
	.w4(32'hba436449),
	.w5(32'hba0405ce),
	.w6(32'h3a25af64),
	.w7(32'h39e6123f),
	.w8(32'h39bcb15e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8331d0),
	.w1(32'hbb928a43),
	.w2(32'hbbe1bdec),
	.w3(32'h3bd247e3),
	.w4(32'h3bd7fac8),
	.w5(32'h3add1ba8),
	.w6(32'hbabedc49),
	.w7(32'h3b4ccb30),
	.w8(32'hbaf848bd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c897),
	.w1(32'h3b84de5a),
	.w2(32'h3a39ed9d),
	.w3(32'hbb15efef),
	.w4(32'hb9a6d2cb),
	.w5(32'hbaade624),
	.w6(32'hbbd18245),
	.w7(32'hbbccf209),
	.w8(32'hbbc0ae12),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997da1),
	.w1(32'hbb5d63bb),
	.w2(32'hbafe7983),
	.w3(32'hbbd3e1aa),
	.w4(32'hbbfa8cf1),
	.w5(32'hbbeee41f),
	.w6(32'h3aef7d7a),
	.w7(32'hbb235d50),
	.w8(32'hbbca42b0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b135c75),
	.w1(32'h3b61e4c6),
	.w2(32'h3b367f32),
	.w3(32'hbb9659c1),
	.w4(32'hb96fd18a),
	.w5(32'hba9047d8),
	.w6(32'hbb578d7a),
	.w7(32'hbbc3dceb),
	.w8(32'hbbf91a13),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4f6c4),
	.w1(32'h3ca0311a),
	.w2(32'h3c51ac2b),
	.w3(32'h3bde3130),
	.w4(32'h3c000f12),
	.w5(32'h3b318627),
	.w6(32'hbbe7d8cc),
	.w7(32'hbbd87730),
	.w8(32'hbc0985a4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87dbe72),
	.w1(32'hb78b2c9c),
	.w2(32'h383d822a),
	.w3(32'hb86a020a),
	.w4(32'hb849a641),
	.w5(32'h37957fd8),
	.w6(32'h381ce0a2),
	.w7(32'h381f74cc),
	.w8(32'h38878196),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955e210),
	.w1(32'hb8b25386),
	.w2(32'h3902e41b),
	.w3(32'hb819f9ba),
	.w4(32'h37ed7c25),
	.w5(32'h3943567c),
	.w6(32'h39185db8),
	.w7(32'h3954c677),
	.w8(32'h39ae4905),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a08dbe),
	.w1(32'hb7e5bb1d),
	.w2(32'h389491e6),
	.w3(32'hb7f21f75),
	.w4(32'h3721bcef),
	.w5(32'h38df7bac),
	.w6(32'h391b2d0b),
	.w7(32'h3937f126),
	.w8(32'h394bc19a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f998d7),
	.w1(32'h38021c3f),
	.w2(32'h39c2a5d4),
	.w3(32'h39e0aa2f),
	.w4(32'h39e45725),
	.w5(32'h3a2dc755),
	.w6(32'h393e21bf),
	.w7(32'h39c1d8dd),
	.w8(32'h3a17e465),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d421),
	.w1(32'h3a8e6df1),
	.w2(32'h3b5cc86d),
	.w3(32'h3a65d22c),
	.w4(32'h3a9eab10),
	.w5(32'h3b1983dd),
	.w6(32'h3abef9d1),
	.w7(32'h3a28fcf2),
	.w8(32'hb98e5865),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1a47),
	.w1(32'h3a243d85),
	.w2(32'h3a03ed09),
	.w3(32'h3abec89a),
	.w4(32'h39bf97c8),
	.w5(32'hb8a217f5),
	.w6(32'h3a4cd6b2),
	.w7(32'h3a424de9),
	.w8(32'h390e2bb3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33f02e),
	.w1(32'hbc2339c5),
	.w2(32'hbc028be0),
	.w3(32'h398e59a6),
	.w4(32'hba3505e3),
	.w5(32'hb997120d),
	.w6(32'h37d9419a),
	.w7(32'h3b5550ea),
	.w8(32'hbacf9e52),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8119e6),
	.w1(32'hbb882505),
	.w2(32'hbb2e69cc),
	.w3(32'hb989d468),
	.w4(32'hba8579e3),
	.w5(32'hb943a1c8),
	.w6(32'h3b175de7),
	.w7(32'h3aedc193),
	.w8(32'h3b1f1019),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5e67),
	.w1(32'h3be8c9cb),
	.w2(32'hb906331c),
	.w3(32'h3b4003d0),
	.w4(32'h3c6b58c2),
	.w5(32'h3c6ccd30),
	.w6(32'hbc4b09bc),
	.w7(32'hbc449124),
	.w8(32'hbc5f3ddf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc8913),
	.w1(32'hb908e103),
	.w2(32'h3aec60a1),
	.w3(32'hbba07262),
	.w4(32'hbb5d96e7),
	.w5(32'hbb2c2602),
	.w6(32'hbc00cebd),
	.w7(32'hbbb968d7),
	.w8(32'hbbb1a0bb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82dcbe),
	.w1(32'hbb95835c),
	.w2(32'hbb43e4e0),
	.w3(32'h3a25290f),
	.w4(32'hb9f2b10d),
	.w5(32'hbb0277fb),
	.w6(32'h3a65ddf7),
	.w7(32'h39dcb103),
	.w8(32'hbaab2301),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa810dd),
	.w1(32'hbb19693f),
	.w2(32'hba807c94),
	.w3(32'h3ae9d369),
	.w4(32'h3a10dc58),
	.w5(32'h3ac754d9),
	.w6(32'h3b2c1ed1),
	.w7(32'h3b233565),
	.w8(32'h3af37a8f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baca988),
	.w1(32'h3bf0136c),
	.w2(32'h3c0ed89a),
	.w3(32'h3a4aa41c),
	.w4(32'h3ad716ce),
	.w5(32'h3b2656c6),
	.w6(32'hbac81610),
	.w7(32'hbac08668),
	.w8(32'h3b88eb9b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46fe21),
	.w1(32'hbb4497df),
	.w2(32'hbb4f30e6),
	.w3(32'hbb35a0b3),
	.w4(32'hbc1b20bc),
	.w5(32'hbc3a7732),
	.w6(32'h3bc547e2),
	.w7(32'hbad963c8),
	.w8(32'hbbc1e9f7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0285),
	.w1(32'hb7f4c23e),
	.w2(32'hbb827a98),
	.w3(32'h3b0a7ef2),
	.w4(32'h39b7858d),
	.w5(32'hbb2d9945),
	.w6(32'h3a2ded9b),
	.w7(32'hbb350e69),
	.w8(32'hbbb09784),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf299c),
	.w1(32'hbc159b63),
	.w2(32'hbba11863),
	.w3(32'h3aa38b2c),
	.w4(32'hbac74c41),
	.w5(32'h3a877f5a),
	.w6(32'h3bbb2dbb),
	.w7(32'h3b8ab8e7),
	.w8(32'h3b99a7c6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828a5f),
	.w1(32'h39c88893),
	.w2(32'h3a769db8),
	.w3(32'hb93c8a3c),
	.w4(32'h39ac86e9),
	.w5(32'h3a21a9f0),
	.w6(32'hb797eb2f),
	.w7(32'h3a2e8b91),
	.w8(32'h39f0e015),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa211d0),
	.w1(32'h3b0fabdf),
	.w2(32'h39ddcbcf),
	.w3(32'h3aa45441),
	.w4(32'h3b2ee245),
	.w5(32'h3adea904),
	.w6(32'hb9a3537a),
	.w7(32'h39f176b6),
	.w8(32'h395d39d0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af4f30),
	.w1(32'hb89e64ee),
	.w2(32'h378d252d),
	.w3(32'hbad71589),
	.w4(32'hbab924cc),
	.w5(32'hb9a64c60),
	.w6(32'hba9f5391),
	.w7(32'hbace5425),
	.w8(32'h3abd559a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0982d),
	.w1(32'h39efee69),
	.w2(32'hbab5f1f9),
	.w3(32'h3b30c648),
	.w4(32'h3793ee58),
	.w5(32'hba866a25),
	.w6(32'h3a74c248),
	.w7(32'h3b1170f2),
	.w8(32'hbb03c311),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b048),
	.w1(32'h3b93f67c),
	.w2(32'hbaf6f2d4),
	.w3(32'h3b97a087),
	.w4(32'h3bed5828),
	.w5(32'h3b397409),
	.w6(32'hbb9aa9ce),
	.w7(32'hbb8b571f),
	.w8(32'hbb845adf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a67778),
	.w1(32'hbb9e38c9),
	.w2(32'hbb5ca4cd),
	.w3(32'h395e8d7d),
	.w4(32'hbb41a50c),
	.w5(32'hbb37f904),
	.w6(32'hbb1d0826),
	.w7(32'hbacdaa10),
	.w8(32'hba57e6de),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f27a6),
	.w1(32'hbb463fbe),
	.w2(32'hba72ccc9),
	.w3(32'hbac5da82),
	.w4(32'hbb67380e),
	.w5(32'hbb0b3968),
	.w6(32'hba4e595b),
	.w7(32'hb9c2deca),
	.w8(32'hba94a463),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc254f6c),
	.w1(32'hbc3e9e60),
	.w2(32'hbbe62b36),
	.w3(32'hbb4397ca),
	.w4(32'hbb1cdb34),
	.w5(32'hbbdb8ae8),
	.w6(32'h375d6e4b),
	.w7(32'h3ba19f4b),
	.w8(32'hba249b51),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bee72),
	.w1(32'h3bd6668b),
	.w2(32'h3c006d0a),
	.w3(32'hbb9d9a3d),
	.w4(32'hbb8fce6d),
	.w5(32'hb912a9cd),
	.w6(32'hbc4d962a),
	.w7(32'hbc2ac508),
	.w8(32'hbb828960),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088cf5),
	.w1(32'h3a1f06e6),
	.w2(32'h3af46017),
	.w3(32'h3b327380),
	.w4(32'h3a25e99f),
	.w5(32'h39d604d1),
	.w6(32'h3afc63b2),
	.w7(32'h3af821dd),
	.w8(32'h3a23f7c9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393de738),
	.w1(32'hbadfb381),
	.w2(32'hb9bf53a4),
	.w3(32'h3b4eae89),
	.w4(32'h3a55f5d7),
	.w5(32'h3ab7bc5c),
	.w6(32'h3b9d32d6),
	.w7(32'h3b96d51b),
	.w8(32'h3b822f55),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade8d07),
	.w1(32'hbb0b66ae),
	.w2(32'h3ab95913),
	.w3(32'h3aa5d801),
	.w4(32'h3a743bd5),
	.w5(32'hb9860618),
	.w6(32'hba67813c),
	.w7(32'hbb16f3b4),
	.w8(32'hbaab2125),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57fdd9),
	.w1(32'hbb406f5f),
	.w2(32'hbb43e05f),
	.w3(32'hbb6723c0),
	.w4(32'hbaa33782),
	.w5(32'hbb5a4a2c),
	.w6(32'hbb1279f9),
	.w7(32'hb997ff25),
	.w8(32'hbae9d062),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f8a96),
	.w1(32'h3b47f92d),
	.w2(32'h3b31d54a),
	.w3(32'hbb305287),
	.w4(32'hbb4f0214),
	.w5(32'hbb1d0649),
	.w6(32'hb9181631),
	.w7(32'hbb167fa7),
	.w8(32'hbb6cf501),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c29bf),
	.w1(32'hba7be1ac),
	.w2(32'hbb8bab63),
	.w3(32'h3a7e9cdb),
	.w4(32'hb9950ece),
	.w5(32'hbaf91825),
	.w6(32'hba6b0ae0),
	.w7(32'hbb4b84cc),
	.w8(32'hbbf26e2f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule