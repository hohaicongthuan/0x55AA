module layer_10_featuremap_422(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d320fc),
	.w1(32'hb736c58e),
	.w2(32'hb7580f2e),
	.w3(32'h38277f9c),
	.w4(32'h3709ab9a),
	.w5(32'hb694e761),
	.w6(32'h3884aa22),
	.w7(32'h38187129),
	.w8(32'h3720d64d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950e34b),
	.w1(32'h39e5993b),
	.w2(32'hb916ff76),
	.w3(32'h3ae00e8b),
	.w4(32'hbaac619d),
	.w5(32'hbb257f88),
	.w6(32'h392f1108),
	.w7(32'hbb2e1557),
	.w8(32'hbb12d234),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372aa4e7),
	.w1(32'h37113d38),
	.w2(32'h375a72f6),
	.w3(32'h36da82a3),
	.w4(32'h361ec20b),
	.w5(32'h37376444),
	.w6(32'h36e6a205),
	.w7(32'h36ee6114),
	.w8(32'h37588388),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcb5b0),
	.w1(32'h3a621572),
	.w2(32'h39365db1),
	.w3(32'h39286a5b),
	.w4(32'hb7d75ece),
	.w5(32'h39fa38de),
	.w6(32'h399ecc49),
	.w7(32'h399b15c1),
	.w8(32'h3a0a900b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397977cd),
	.w1(32'h399332c0),
	.w2(32'h38e46d60),
	.w3(32'h398ed701),
	.w4(32'h399ecd6a),
	.w5(32'h39358c04),
	.w6(32'h39890b83),
	.w7(32'h399d2c5c),
	.w8(32'h398711bb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ff89bd),
	.w1(32'hb82b1420),
	.w2(32'hb799820a),
	.w3(32'hb7bd92ce),
	.w4(32'hb7db5d8d),
	.w5(32'hb6baf7d2),
	.w6(32'hb7407784),
	.w7(32'h3731e5e1),
	.w8(32'h382aa423),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2463f5),
	.w1(32'h39e0dd26),
	.w2(32'hbaa23efc),
	.w3(32'h3b593129),
	.w4(32'hb95e910f),
	.w5(32'hbb0c50be),
	.w6(32'h361cddb0),
	.w7(32'hb9dc575a),
	.w8(32'hbb822369),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058a40),
	.w1(32'hbb915ff5),
	.w2(32'hbab3234e),
	.w3(32'hbc80f7cd),
	.w4(32'hbb978d69),
	.w5(32'hbb0a94cb),
	.w6(32'hbc261c0a),
	.w7(32'hbc0171ac),
	.w8(32'h3b527927),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddf90f),
	.w1(32'hb9c7ace1),
	.w2(32'hb9d1afed),
	.w3(32'hb9960f99),
	.w4(32'h39befdc3),
	.w5(32'h37d9f9e6),
	.w6(32'hba91f3f8),
	.w7(32'hb99057c7),
	.w8(32'hb9e71fae),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36b2ce),
	.w1(32'hb9e52c8f),
	.w2(32'hbb23991a),
	.w3(32'hbb673e8b),
	.w4(32'hb9bf9d9d),
	.w5(32'hbb9611b1),
	.w6(32'hbb8cfc82),
	.w7(32'h39c3846c),
	.w8(32'hbbbdfc79),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d5964),
	.w1(32'h3aa555c5),
	.w2(32'h3a185bdd),
	.w3(32'h39924766),
	.w4(32'h39dc19ad),
	.w5(32'hb9fb089c),
	.w6(32'h396b08b4),
	.w7(32'h398e7bfd),
	.w8(32'hb98fa2d2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21292a),
	.w1(32'h3af60fff),
	.w2(32'hb92d45aa),
	.w3(32'h3bc2ea8c),
	.w4(32'h3b68b426),
	.w5(32'h3b34f6d8),
	.w6(32'h3b204b68),
	.w7(32'h3bbcd047),
	.w8(32'h3b0498f3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb051a2),
	.w1(32'h3a5b1453),
	.w2(32'h3acb652f),
	.w3(32'hbbf51d27),
	.w4(32'hb9255d6e),
	.w5(32'h3a2a3340),
	.w6(32'hbb7a2d4f),
	.w7(32'h3b47a29a),
	.w8(32'hb93f7f6c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae65bdc),
	.w1(32'h3b08ac53),
	.w2(32'hb9b6db3d),
	.w3(32'hba3a63aa),
	.w4(32'hb9f091eb),
	.w5(32'hbaececf7),
	.w6(32'hb9cbe690),
	.w7(32'hb99fc04d),
	.w8(32'hba7f18fd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7edce4),
	.w1(32'hba060423),
	.w2(32'hbb047df3),
	.w3(32'h3a20b659),
	.w4(32'hba10f9ae),
	.w5(32'hbb01b393),
	.w6(32'h3a49c0b9),
	.w7(32'hb9c4e5fb),
	.w8(32'hbaf39325),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c4b58),
	.w1(32'h3af481ec),
	.w2(32'h3b13099e),
	.w3(32'hbb68b41e),
	.w4(32'hbb1c4639),
	.w5(32'hb78d2e54),
	.w6(32'hbbdd9925),
	.w7(32'hbba44945),
	.w8(32'hbb40860e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ddf053),
	.w1(32'h389f8ad1),
	.w2(32'h39ff60b4),
	.w3(32'hb974631a),
	.w4(32'h38e9e4ba),
	.w5(32'h395b4255),
	.w6(32'hba1c4460),
	.w7(32'hb947b7b0),
	.w8(32'h38d1aede),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84d66f),
	.w1(32'hbac6d774),
	.w2(32'h3a44e463),
	.w3(32'hbc42ddcb),
	.w4(32'hbb0016a6),
	.w5(32'h3a06a40b),
	.w6(32'hbbd1545f),
	.w7(32'hbb3b3555),
	.w8(32'hba8f1ce9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2976a8),
	.w1(32'h3987cd39),
	.w2(32'h3adf5365),
	.w3(32'hbbe9457d),
	.w4(32'hbaf9be93),
	.w5(32'h3aa431c9),
	.w6(32'hbb80bfb0),
	.w7(32'hb7fe1c39),
	.w8(32'h3a41e0d5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8801099),
	.w1(32'h38474320),
	.w2(32'hb7899541),
	.w3(32'h37b30e88),
	.w4(32'h38290ee4),
	.w5(32'hb6c2f0b5),
	.w6(32'h37db78ea),
	.w7(32'h37a05a3d),
	.w8(32'h38325e16),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60c55ea),
	.w1(32'hb914694f),
	.w2(32'hb8887ff0),
	.w3(32'hb848ed54),
	.w4(32'hb9765e2d),
	.w5(32'hb887fe75),
	.w6(32'hb6e24a47),
	.w7(32'hb8705c33),
	.w8(32'h385ace94),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a77ace),
	.w1(32'h39ddc01a),
	.w2(32'h37b7567a),
	.w3(32'h3a063126),
	.w4(32'h39b387a6),
	.w5(32'hb94c26d2),
	.w6(32'h3ad2cdc3),
	.w7(32'h3a979464),
	.w8(32'h39ed4b9a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac12921),
	.w1(32'hbba2a675),
	.w2(32'hbb7c48ad),
	.w3(32'hbbe08a16),
	.w4(32'hbb346f12),
	.w5(32'h3a04e93a),
	.w6(32'hbc015019),
	.w7(32'h3a8a000b),
	.w8(32'hbc02db8d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd54b2),
	.w1(32'h39b7d076),
	.w2(32'hbb170894),
	.w3(32'h3892cca1),
	.w4(32'h39de24e1),
	.w5(32'hbb68399b),
	.w6(32'h399878a2),
	.w7(32'hb7b6588b),
	.w8(32'hbb8816fd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903e35d),
	.w1(32'h3a69f19e),
	.w2(32'hb9cca474),
	.w3(32'hb9a43dc1),
	.w4(32'h3912545f),
	.w5(32'hbb691a79),
	.w6(32'h3aa6ff47),
	.w7(32'hbb6670f1),
	.w8(32'hbb9ea730),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6b011),
	.w1(32'h3a247444),
	.w2(32'h39f5cba6),
	.w3(32'hb9e92b82),
	.w4(32'h393f9201),
	.w5(32'h3774646c),
	.w6(32'hba25c2b0),
	.w7(32'hb7b5c192),
	.w8(32'hb9987819),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af9339),
	.w1(32'h38b22ee5),
	.w2(32'h3939ecf9),
	.w3(32'h39020dca),
	.w4(32'h3892bf3b),
	.w5(32'h3938d09c),
	.w6(32'h390f83e7),
	.w7(32'h38a10ed1),
	.w8(32'h39842883),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28174e),
	.w1(32'h3b027841),
	.w2(32'h39efc465),
	.w3(32'h3aa0340a),
	.w4(32'h3b4fd3dc),
	.w5(32'hbabf48ed),
	.w6(32'h3b5fd548),
	.w7(32'h3bbe29a4),
	.w8(32'h3a7029bb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a481848),
	.w1(32'h3a258cc5),
	.w2(32'h3a20105a),
	.w3(32'h3b11b6c3),
	.w4(32'h3b063112),
	.w5(32'h3aa6c644),
	.w6(32'h3b7cb535),
	.w7(32'h3b3a786b),
	.w8(32'h3b5a51b6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa939a),
	.w1(32'h3b34878f),
	.w2(32'hbad33c19),
	.w3(32'h3ab8303e),
	.w4(32'h38a30039),
	.w5(32'hbbccd4b7),
	.w6(32'h3b8e891e),
	.w7(32'h3a839b4e),
	.w8(32'hbbab0589),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d29970),
	.w1(32'h387bdd46),
	.w2(32'h38e2a183),
	.w3(32'hb6f9c397),
	.w4(32'h3843af7b),
	.w5(32'h38d4c609),
	.w6(32'h3735d484),
	.w7(32'h3874317d),
	.w8(32'h38da533b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386658da),
	.w1(32'h39632c3f),
	.w2(32'h39a0127b),
	.w3(32'h380d92fa),
	.w4(32'h3985b53b),
	.w5(32'h399cb216),
	.w6(32'h3814ff74),
	.w7(32'h398e3989),
	.w8(32'h39a91f4d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37ba1),
	.w1(32'h3aee9425),
	.w2(32'h395a0354),
	.w3(32'h39f48041),
	.w4(32'h3aa75ee5),
	.w5(32'hb93059f1),
	.w6(32'hb93f0083),
	.w7(32'h39d16c23),
	.w8(32'hba947002),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1da43),
	.w1(32'hba8bde6f),
	.w2(32'hba6c2dcf),
	.w3(32'hba247f16),
	.w4(32'hba687056),
	.w5(32'hbab610cc),
	.w6(32'hba512fe4),
	.w7(32'hbb1732dd),
	.w8(32'hbb0d6641),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3eb62),
	.w1(32'h388b27f8),
	.w2(32'h3985758f),
	.w3(32'h385fbf97),
	.w4(32'h35bee776),
	.w5(32'h39ce4282),
	.w6(32'hb8fb2f61),
	.w7(32'h37e35a82),
	.w8(32'h3605775c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389aed18),
	.w1(32'h3a0013fe),
	.w2(32'h39d30878),
	.w3(32'hbb036f0f),
	.w4(32'hb6baab6e),
	.w5(32'h3a20d85e),
	.w6(32'hba16f663),
	.w7(32'h3a1d0a4b),
	.w8(32'hb98ec17a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b23aa),
	.w1(32'h3b03118d),
	.w2(32'h39807e57),
	.w3(32'h395dc9e5),
	.w4(32'hbbb075f3),
	.w5(32'h3a6baaa4),
	.w6(32'hbbdc5acd),
	.w7(32'hbb76f04c),
	.w8(32'h3b32972e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4221),
	.w1(32'hb9709179),
	.w2(32'hbb508b7e),
	.w3(32'h3bcce20d),
	.w4(32'h3b2f4207),
	.w5(32'hbb0c91ad),
	.w6(32'h3b21b85a),
	.w7(32'h3aeb35d5),
	.w8(32'hbae2dead),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48a119),
	.w1(32'h3aef3a6f),
	.w2(32'hbbd69e63),
	.w3(32'h3c1f9502),
	.w4(32'h3b76a60e),
	.w5(32'hbbfc1104),
	.w6(32'h3c09cebf),
	.w7(32'h3b667f02),
	.w8(32'hbb9163de),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a684cc),
	.w1(32'h3abd429f),
	.w2(32'h398655e3),
	.w3(32'hb9a18d0f),
	.w4(32'h3931cdab),
	.w5(32'h39851163),
	.w6(32'hba70b2ec),
	.w7(32'hb7422648),
	.w8(32'h3a58b91d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba215843),
	.w1(32'hb97327f3),
	.w2(32'hb9cfe813),
	.w3(32'hba063eb0),
	.w4(32'hb9877a0f),
	.w5(32'hba0cb578),
	.w6(32'hb9a60e01),
	.w7(32'hb8c2eead),
	.w8(32'hb9ce7181),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b691c),
	.w1(32'hb9ae9b61),
	.w2(32'h3910883c),
	.w3(32'h380334f0),
	.w4(32'hb8f35f48),
	.w5(32'h39890cc5),
	.w6(32'h3975deba),
	.w7(32'h38de5d63),
	.w8(32'h39d74afb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e57e4),
	.w1(32'h3a372d0b),
	.w2(32'h3a4432d0),
	.w3(32'h3ae90ece),
	.w4(32'h3a907492),
	.w5(32'h39a066aa),
	.w6(32'h3985cc71),
	.w7(32'h39816a4e),
	.w8(32'hb9ec8075),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1605e),
	.w1(32'h3af6b8c9),
	.w2(32'hbad198ca),
	.w3(32'hbb9321f6),
	.w4(32'hbab38238),
	.w5(32'hbae3ca88),
	.w6(32'hbb8e4e96),
	.w7(32'h3a881faa),
	.w8(32'hbaf3be70),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9936e),
	.w1(32'hb8e0497b),
	.w2(32'hbb37b6c7),
	.w3(32'hb702b888),
	.w4(32'hb9a25571),
	.w5(32'hbba0faf0),
	.w6(32'h3a29bca7),
	.w7(32'hba8d26ec),
	.w8(32'hbba3d9aa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8195ed),
	.w1(32'h39ca0b8f),
	.w2(32'hbb1f0ef4),
	.w3(32'hbb010195),
	.w4(32'h38eebfcb),
	.w5(32'hbb89d185),
	.w6(32'hbafc492f),
	.w7(32'hbb1a7e88),
	.w8(32'hbba797fd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a0b0),
	.w1(32'hbb5d4ee2),
	.w2(32'hbbb8e9b8),
	.w3(32'hbb204e28),
	.w4(32'hbb0db99a),
	.w5(32'hbb95ead0),
	.w6(32'hbba3ddcc),
	.w7(32'hbb555229),
	.w8(32'hbba75f8b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68ecbe),
	.w1(32'hb9a878e9),
	.w2(32'hb819ea62),
	.w3(32'hbc828e4d),
	.w4(32'hbbad3685),
	.w5(32'h3a6d10a6),
	.w6(32'hbc51955b),
	.w7(32'hbb2c1141),
	.w8(32'hba5a706f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1952b4),
	.w1(32'h38ee82cb),
	.w2(32'hba24a88c),
	.w3(32'h3a5de247),
	.w4(32'h39ec48f6),
	.w5(32'hb8172391),
	.w6(32'h3a3950e8),
	.w7(32'h39db61d2),
	.w8(32'h38e72c5e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29de0b),
	.w1(32'hbaa748b7),
	.w2(32'hbac6a799),
	.w3(32'hbac0713e),
	.w4(32'hba578dff),
	.w5(32'hba9a5c82),
	.w6(32'hbab5cea4),
	.w7(32'hbaebd22e),
	.w8(32'hbafe128b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93bc35),
	.w1(32'h3a56c38a),
	.w2(32'hb939f253),
	.w3(32'h3ac5b6d0),
	.w4(32'h3a9743d6),
	.w5(32'h3a0f6eca),
	.w6(32'h3aa00df4),
	.w7(32'h3a9db0b9),
	.w8(32'h3877aa0c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bedbd),
	.w1(32'hb9759d69),
	.w2(32'hbaa4efd9),
	.w3(32'hbb71973e),
	.w4(32'hba52ee31),
	.w5(32'hbaa52a32),
	.w6(32'hba8389dc),
	.w7(32'hba820721),
	.w8(32'hbb6a2d10),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba175456),
	.w1(32'hba323a79),
	.w2(32'hba10c7c8),
	.w3(32'hba57aef4),
	.w4(32'hb9d6f4f5),
	.w5(32'hba29e3fd),
	.w6(32'hba6b3db8),
	.w7(32'hba3accd5),
	.w8(32'hba7294d6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa18f5b),
	.w1(32'hbad09426),
	.w2(32'hbae062d2),
	.w3(32'hbbdb725c),
	.w4(32'hbafa0d7d),
	.w5(32'h3b050f9b),
	.w6(32'hbb95e93c),
	.w7(32'hb8d3ad9c),
	.w8(32'hb9c28655),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca548b),
	.w1(32'hb9c4d407),
	.w2(32'hb9a92938),
	.w3(32'h38ce8a89),
	.w4(32'h3a6ada5a),
	.w5(32'hb9dbbf45),
	.w6(32'h39920e27),
	.w7(32'hb91bd5b9),
	.w8(32'hb7663667),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d7dc5),
	.w1(32'h3907740a),
	.w2(32'hb6ee953b),
	.w3(32'h38b97567),
	.w4(32'hb8ba0552),
	.w5(32'hb91043b1),
	.w6(32'h37efa9d7),
	.w7(32'hb8d4807f),
	.w8(32'hb9028fcc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7145e80),
	.w1(32'hb75e12db),
	.w2(32'h379e0139),
	.w3(32'h376ba333),
	.w4(32'hb7ccaa47),
	.w5(32'hb7832301),
	.w6(32'h37fc9d55),
	.w7(32'h36abdf02),
	.w8(32'h372aac1f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b2a7d),
	.w1(32'hb87b2029),
	.w2(32'hb8984fbb),
	.w3(32'h39e1f83a),
	.w4(32'h387fbdff),
	.w5(32'hb9d31c1d),
	.w6(32'h3a2c6745),
	.w7(32'h387003ce),
	.w8(32'hb9f313b1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d8230),
	.w1(32'h3a420bf6),
	.w2(32'h3a761b20),
	.w3(32'h3a4a6bfa),
	.w4(32'h3a2ee398),
	.w5(32'h3a13649b),
	.w6(32'h3a3ed6c4),
	.w7(32'h3a23c081),
	.w8(32'h39daf78b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad1b49),
	.w1(32'h39cbb894),
	.w2(32'h3915ff1a),
	.w3(32'h39cd476e),
	.w4(32'h38839c8b),
	.w5(32'hb9869d5d),
	.w6(32'h3a35842a),
	.w7(32'h3897d19e),
	.w8(32'hb9b2ae92),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96a921),
	.w1(32'h3999109b),
	.w2(32'h3a008ee3),
	.w3(32'hbb85a0f2),
	.w4(32'hb9944130),
	.w5(32'h3a7a0fc6),
	.w6(32'hbaa544f3),
	.w7(32'h3aac8af6),
	.w8(32'h394225de),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5642),
	.w1(32'hbaa68975),
	.w2(32'h3ae22119),
	.w3(32'hbbbebc6e),
	.w4(32'hba93b9d0),
	.w5(32'h39383dd5),
	.w6(32'hbb2631bf),
	.w7(32'hba650730),
	.w8(32'hbb138cb9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896b91b),
	.w1(32'h3662f858),
	.w2(32'h37ebb8be),
	.w3(32'hb723bdf9),
	.w4(32'h38c2226c),
	.w5(32'h3938f9ea),
	.w6(32'h380e4ae5),
	.w7(32'h3893a4d1),
	.w8(32'h39343f03),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7518df7),
	.w1(32'hb65730ca),
	.w2(32'h37e5f326),
	.w3(32'hb79115ba),
	.w4(32'hb7377989),
	.w5(32'h3788f592),
	.w6(32'hb6f9ff1d),
	.w7(32'hb6bf2b8d),
	.w8(32'h377d8d9a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e9a57),
	.w1(32'h3971814d),
	.w2(32'h399c78f1),
	.w3(32'h38da91bf),
	.w4(32'hb84bdb47),
	.w5(32'h366374a6),
	.w6(32'h39380408),
	.w7(32'h389d9e67),
	.w8(32'h3981901f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358a7352),
	.w1(32'h37a37a85),
	.w2(32'h3879c6c3),
	.w3(32'h37c2cff0),
	.w4(32'h37f15569),
	.w5(32'h38ab600a),
	.w6(32'h3852e562),
	.w7(32'h383209bc),
	.w8(32'h38f8a8a8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6bee9),
	.w1(32'h3ae81636),
	.w2(32'h3ba6445e),
	.w3(32'h3af35d00),
	.w4(32'h3a487088),
	.w5(32'h3b640232),
	.w6(32'hbb9810f8),
	.w7(32'h3b30858e),
	.w8(32'h3b02b59a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa99556),
	.w1(32'h3a8bf466),
	.w2(32'hbaa4c0f8),
	.w3(32'h3a29db17),
	.w4(32'h3aaabb64),
	.w5(32'hbb80128f),
	.w6(32'hbb6888e6),
	.w7(32'hbbb60626),
	.w8(32'hbbefa7a7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada16d4),
	.w1(32'h3a323330),
	.w2(32'h38cc0432),
	.w3(32'h3ad513e3),
	.w4(32'h3b494c73),
	.w5(32'h3b092bd8),
	.w6(32'h3b2c04ce),
	.w7(32'h39b80860),
	.w8(32'hbb48ac8a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd72a4),
	.w1(32'h3b43ebe6),
	.w2(32'hbb61adb6),
	.w3(32'h3b8b3018),
	.w4(32'h3bc270db),
	.w5(32'hbc4785e7),
	.w6(32'h3ba4a0a6),
	.w7(32'h3bc084b9),
	.w8(32'hbc85ed64),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f850b),
	.w1(32'h3b3f0441),
	.w2(32'h3bb726be),
	.w3(32'h3b83ff7a),
	.w4(32'h3b295d59),
	.w5(32'hbba22447),
	.w6(32'h3b0506a7),
	.w7(32'hbb76f53f),
	.w8(32'hbbc1f35e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47bb62),
	.w1(32'hbb66742c),
	.w2(32'hbbbbc587),
	.w3(32'hbbb99347),
	.w4(32'hbb59a3dd),
	.w5(32'hbbff30fc),
	.w6(32'hbbeaab93),
	.w7(32'hbbadabec),
	.w8(32'hbc095fe5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092503),
	.w1(32'hbbd58c87),
	.w2(32'hbbaccc24),
	.w3(32'hbbf23bc6),
	.w4(32'hbb59606a),
	.w5(32'hbbfeddeb),
	.w6(32'hbb65c952),
	.w7(32'hbab3860f),
	.w8(32'hbbc8d2e1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbb0a),
	.w1(32'hbb5e5604),
	.w2(32'hbba81a56),
	.w3(32'hbc2ad6bb),
	.w4(32'h3a95df2b),
	.w5(32'h3b4c4661),
	.w6(32'hbc4d3780),
	.w7(32'hbae17bb0),
	.w8(32'hbac57fae),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ea9d),
	.w1(32'hbbff6a69),
	.w2(32'hbc07e51c),
	.w3(32'hba268410),
	.w4(32'hbc03672e),
	.w5(32'hbbddf752),
	.w6(32'hbb20eb16),
	.w7(32'h3a9a9f6d),
	.w8(32'h3b88acf8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1deb55),
	.w1(32'hbbc0ec3a),
	.w2(32'hbbe3919a),
	.w3(32'hbc44512a),
	.w4(32'hbb954d72),
	.w5(32'hbb7748a8),
	.w6(32'hbb531da5),
	.w7(32'hb994722c),
	.w8(32'hbb4ea316),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc02f6),
	.w1(32'hbc35a3dd),
	.w2(32'hbbaf13ff),
	.w3(32'hbc2b2d76),
	.w4(32'hbc2b13dd),
	.w5(32'h3a375d95),
	.w6(32'hbc6e3120),
	.w7(32'hbb51b098),
	.w8(32'h3af863e6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc3f6),
	.w1(32'hbb85de9f),
	.w2(32'hbacad4b6),
	.w3(32'h3847058f),
	.w4(32'hbbe733a7),
	.w5(32'hbc028a24),
	.w6(32'hbb100cc9),
	.w7(32'hbb1cace0),
	.w8(32'hbac51c3b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c795f),
	.w1(32'hbade1290),
	.w2(32'hbada297b),
	.w3(32'hbbe84657),
	.w4(32'hb8eb1388),
	.w5(32'h3a98dbfd),
	.w6(32'hbb1466d2),
	.w7(32'h3b5ecf5a),
	.w8(32'hbacb0015),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba957f60),
	.w1(32'hbb8d3abe),
	.w2(32'hbaf003bd),
	.w3(32'h3b7cb56f),
	.w4(32'hbbe393f6),
	.w5(32'hbb891ce4),
	.w6(32'hbb11c17b),
	.w7(32'hbb928fa8),
	.w8(32'hbbc3d2bb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3641),
	.w1(32'h3afdbb8d),
	.w2(32'hbbe82356),
	.w3(32'hba414fdc),
	.w4(32'h3c2d1430),
	.w5(32'h3bc807b3),
	.w6(32'hb8873bc3),
	.w7(32'h3c8f6c75),
	.w8(32'h3c5de198),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef1281),
	.w1(32'hbb0bf7f8),
	.w2(32'h392733ea),
	.w3(32'h3be17c39),
	.w4(32'h39aa3f61),
	.w5(32'h3b96fd08),
	.w6(32'h3c320f95),
	.w7(32'h3b7bf976),
	.w8(32'h3bd44c72),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aee4c),
	.w1(32'h3bb5df39),
	.w2(32'h3af02a5c),
	.w3(32'h3b079630),
	.w4(32'h3b7b7ea3),
	.w5(32'h3bae287d),
	.w6(32'h3c00306f),
	.w7(32'hbac51533),
	.w8(32'h38d1e622),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13948c),
	.w1(32'h3aaa5443),
	.w2(32'hb97bcb85),
	.w3(32'h3b6a42c1),
	.w4(32'h3ab7cb0e),
	.w5(32'hba6067a6),
	.w6(32'h3a16989a),
	.w7(32'hbbc19204),
	.w8(32'hbaae0819),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab757b0),
	.w1(32'hbb1ebd0c),
	.w2(32'hba81bcff),
	.w3(32'hbc022368),
	.w4(32'hbb64fffc),
	.w5(32'hbb59a707),
	.w6(32'hbb1728ce),
	.w7(32'hbb0e1b4b),
	.w8(32'hbb50d1c5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133f4b),
	.w1(32'hb940110f),
	.w2(32'h3c10d588),
	.w3(32'hbba7626b),
	.w4(32'hbb70f647),
	.w5(32'h3c212f04),
	.w6(32'hbb3160e3),
	.w7(32'hbbbf1a16),
	.w8(32'h3bb84a4e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979db84),
	.w1(32'h3b4a5e22),
	.w2(32'h395d33aa),
	.w3(32'h3b95cafd),
	.w4(32'h3abfe706),
	.w5(32'hbbca15d7),
	.w6(32'h3b20f78d),
	.w7(32'hbb27b8fd),
	.w8(32'hbba4d914),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e043),
	.w1(32'h3935e811),
	.w2(32'h3b409830),
	.w3(32'hbbc52811),
	.w4(32'h3b5712fe),
	.w5(32'h3a960a3e),
	.w6(32'hbbca64a6),
	.w7(32'h3a2437ae),
	.w8(32'hbaddf2ba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c00ff),
	.w1(32'h3a2b1e0a),
	.w2(32'hbc097605),
	.w3(32'hbba5bf56),
	.w4(32'hbb57f22b),
	.w5(32'hbb6c0847),
	.w6(32'hbb4c86e9),
	.w7(32'hbb8383ae),
	.w8(32'hbbf17487),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5cf95),
	.w1(32'hbb6e190e),
	.w2(32'hbb8b490d),
	.w3(32'hbad74bdd),
	.w4(32'hbc0cf155),
	.w5(32'hbad71a0c),
	.w6(32'hbbf99ec3),
	.w7(32'hbbf25a63),
	.w8(32'hbaf14df2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabc325),
	.w1(32'hbae4ce04),
	.w2(32'hbbd0607d),
	.w3(32'h3c16db83),
	.w4(32'hb9c71732),
	.w5(32'hbbf9d820),
	.w6(32'h3b026608),
	.w7(32'h3ace0221),
	.w8(32'hbc12be4b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4100b1),
	.w1(32'hbb0c0179),
	.w2(32'hbb8971f7),
	.w3(32'hbb8c4bac),
	.w4(32'hbb0e9d92),
	.w5(32'h3c0e20b3),
	.w6(32'hbc288007),
	.w7(32'h3a522d2b),
	.w8(32'h3c1c1359),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a283f8c),
	.w1(32'hbab0f25c),
	.w2(32'hbb6b1d2b),
	.w3(32'h3a0b5398),
	.w4(32'h3b2a03cd),
	.w5(32'h3bcf4afe),
	.w6(32'h3c4b6d83),
	.w7(32'h37d53067),
	.w8(32'h38e44e40),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1358),
	.w1(32'h3ba8c99d),
	.w2(32'hb9bd6caf),
	.w3(32'h3b4757f5),
	.w4(32'h3be4c078),
	.w5(32'h3a947116),
	.w6(32'h3b6743de),
	.w7(32'hba515fb8),
	.w8(32'hbad84cee),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a2671),
	.w1(32'hbbbcfdbe),
	.w2(32'hbbda6499),
	.w3(32'h3b20d3ba),
	.w4(32'hba46c3ae),
	.w5(32'hbb321237),
	.w6(32'h3aa744dc),
	.w7(32'hbb7402e7),
	.w8(32'hbb9f3954),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf50f7),
	.w1(32'h3c18009f),
	.w2(32'hb926c3ee),
	.w3(32'hbbd24356),
	.w4(32'h3b45c148),
	.w5(32'hbc25a590),
	.w6(32'hb95a0351),
	.w7(32'h3af2ecde),
	.w8(32'hbc0b6c1d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b731728),
	.w1(32'h3b9d71fb),
	.w2(32'h3c3cee67),
	.w3(32'h3a60c6cd),
	.w4(32'h3c0eb932),
	.w5(32'h3c5c75b7),
	.w6(32'hba82779b),
	.w7(32'h3bf86be7),
	.w8(32'h3bec4381),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012373),
	.w1(32'hbbce2f78),
	.w2(32'hbc71f5f6),
	.w3(32'hbb6000f0),
	.w4(32'hbc4f762e),
	.w5(32'hbc1b2d65),
	.w6(32'h3b031582),
	.w7(32'hbc641140),
	.w8(32'hbc21ed08),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bfd8d),
	.w1(32'h36f0876a),
	.w2(32'hba97b498),
	.w3(32'h3c2eb344),
	.w4(32'h3b9bff87),
	.w5(32'h3b7783e1),
	.w6(32'h3b50a7c5),
	.w7(32'h3bbabec2),
	.w8(32'h3b317308),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6610),
	.w1(32'h3aab3af0),
	.w2(32'hbc4475f8),
	.w3(32'hbc5b14ff),
	.w4(32'hbc814cab),
	.w5(32'hbb4ea3a4),
	.w6(32'hbbbc0d9c),
	.w7(32'hbc269e47),
	.w8(32'hbb86b7e0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f4ae),
	.w1(32'h3b9c1942),
	.w2(32'h3aecb8b5),
	.w3(32'h3c650b31),
	.w4(32'h3c76d74b),
	.w5(32'h3bdabcc8),
	.w6(32'hbb895202),
	.w7(32'h3bb39ad5),
	.w8(32'h3a1d250f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99a41c),
	.w1(32'hbb47ac63),
	.w2(32'hbb84352c),
	.w3(32'hbbcced3d),
	.w4(32'hbb15afdb),
	.w5(32'hbbda768a),
	.w6(32'hbb23cabb),
	.w7(32'hbc149210),
	.w8(32'hbc469cf6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf03876),
	.w1(32'hbb1a94be),
	.w2(32'hbb58cb0b),
	.w3(32'h3bcbae49),
	.w4(32'hbb044998),
	.w5(32'h3b40ee57),
	.w6(32'hbb77d1bb),
	.w7(32'h3a5c1eb5),
	.w8(32'hbbfa01f8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff305),
	.w1(32'hba81197a),
	.w2(32'hbad708ab),
	.w3(32'hb9b6053f),
	.w4(32'hbaab81dc),
	.w5(32'hbb272a62),
	.w6(32'h3b128711),
	.w7(32'hbc0c4ed2),
	.w8(32'hbbf199a4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d96b7),
	.w1(32'h3abe7099),
	.w2(32'hbbc721b3),
	.w3(32'hbcb638dd),
	.w4(32'hbc277852),
	.w5(32'h3b9a0792),
	.w6(32'hbc958b12),
	.w7(32'hbc2b358d),
	.w8(32'hbab0f1d0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20da45),
	.w1(32'hbb2d2f37),
	.w2(32'hbb73d5db),
	.w3(32'h3b548fcb),
	.w4(32'h3980702c),
	.w5(32'hbb52c6ce),
	.w6(32'hbb186e56),
	.w7(32'h3b94ea1f),
	.w8(32'h3b9c712a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435ac3),
	.w1(32'h3b81b1e8),
	.w2(32'h3c2976ba),
	.w3(32'h3a34e2e1),
	.w4(32'h3b39782d),
	.w5(32'h3bb95636),
	.w6(32'h3b8e6932),
	.w7(32'hb64688d2),
	.w8(32'h3b174f12),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19d5ed),
	.w1(32'hbb85afd7),
	.w2(32'hba8c0f34),
	.w3(32'h39b5fe2f),
	.w4(32'h3b0e6068),
	.w5(32'hbaf81af0),
	.w6(32'hbc0f6467),
	.w7(32'h3b879a68),
	.w8(32'h3acb4cea),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84492a),
	.w1(32'h3b14dd07),
	.w2(32'hbaba1844),
	.w3(32'hbbff53a0),
	.w4(32'hbb692d25),
	.w5(32'h3a67df4e),
	.w6(32'hbb8d6664),
	.w7(32'hbb9e6685),
	.w8(32'h3a722dc5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6344ff),
	.w1(32'h3aefeedb),
	.w2(32'hbb05c7c0),
	.w3(32'hbaf0d28e),
	.w4(32'h3ac2638b),
	.w5(32'hbbc3a05e),
	.w6(32'h3b36ae8b),
	.w7(32'hb8d39c7a),
	.w8(32'hbbf74c67),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5f8ae),
	.w1(32'h3b919313),
	.w2(32'h3badd934),
	.w3(32'h3be295e4),
	.w4(32'hbb154fa7),
	.w5(32'hbc13cab6),
	.w6(32'h3ac18e61),
	.w7(32'h3b910554),
	.w8(32'h3ba85662),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884fc4),
	.w1(32'hbb0a7eca),
	.w2(32'h3ba1d645),
	.w3(32'h3b917220),
	.w4(32'hb9b9c131),
	.w5(32'h3b28f2fe),
	.w6(32'h3b81c532),
	.w7(32'hbafeef93),
	.w8(32'hba569310),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ad9a8),
	.w1(32'h3bb8f7ac),
	.w2(32'h3c116a13),
	.w3(32'h38f58946),
	.w4(32'h3baa47bc),
	.w5(32'h3c2a9f98),
	.w6(32'h3b224557),
	.w7(32'h3b91b9a9),
	.w8(32'h3b314bb1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31fc7c),
	.w1(32'hb8c7e843),
	.w2(32'h39f352de),
	.w3(32'hbbe88493),
	.w4(32'hbb664a63),
	.w5(32'h3bb3493c),
	.w6(32'hbaf4b997),
	.w7(32'h3bb555d4),
	.w8(32'hbb1cfc00),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc5db),
	.w1(32'h3bda2fee),
	.w2(32'hb9ba08e4),
	.w3(32'h39b66c17),
	.w4(32'hba2c5d08),
	.w5(32'hbbcfc7db),
	.w6(32'hbb83b6fe),
	.w7(32'hbad64eba),
	.w8(32'hbb5d4811),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b689b58),
	.w1(32'hbb876f5b),
	.w2(32'hbbf3062a),
	.w3(32'h3b6bb7b8),
	.w4(32'hbb941f1e),
	.w5(32'hbb6eb0b0),
	.w6(32'h3c1ea725),
	.w7(32'hba90971d),
	.w8(32'hba5693c5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad304a9),
	.w1(32'h3bb67a1e),
	.w2(32'h3b0c74af),
	.w3(32'h39f1d95f),
	.w4(32'hba917c29),
	.w5(32'hbb8b205e),
	.w6(32'h3b0a0d91),
	.w7(32'h3b6d3032),
	.w8(32'h3ada18ce),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8e48e),
	.w1(32'h3b651924),
	.w2(32'hbab4b8ff),
	.w3(32'h3b459802),
	.w4(32'hbb451d55),
	.w5(32'h3b3144ff),
	.w6(32'h3b94ea33),
	.w7(32'hbb162112),
	.w8(32'h3b235958),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe18b5),
	.w1(32'hbb3ac624),
	.w2(32'hbba2a573),
	.w3(32'h3b03a3cf),
	.w4(32'hbb115ddd),
	.w5(32'hba78f9ec),
	.w6(32'h3b3ac610),
	.w7(32'hbb5e68eb),
	.w8(32'hbbcea8d8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9c90),
	.w1(32'hb9e3675e),
	.w2(32'hba66c0de),
	.w3(32'hbbfeb614),
	.w4(32'hbb86070d),
	.w5(32'hbbbb1efa),
	.w6(32'hbba71427),
	.w7(32'hbbf1ec3a),
	.w8(32'hbc0dc111),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4590f),
	.w1(32'hbba7b661),
	.w2(32'hbb9c7e4e),
	.w3(32'hbbd45391),
	.w4(32'hbb45d59a),
	.w5(32'hbad70976),
	.w6(32'hbba7ea15),
	.w7(32'hbb31f6f9),
	.w8(32'hbb97a267),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977afa),
	.w1(32'h3bdf77d9),
	.w2(32'hbb5c0d13),
	.w3(32'hb902d05a),
	.w4(32'h3a86bbe5),
	.w5(32'h3c0745d9),
	.w6(32'hbba5d8bb),
	.w7(32'h3a2c5cbb),
	.w8(32'hbbc99c55),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe48cb),
	.w1(32'hb9ed851c),
	.w2(32'h3b87a5a5),
	.w3(32'h3c2e986c),
	.w4(32'h3ad580df),
	.w5(32'hba833a1f),
	.w6(32'hbb83ee23),
	.w7(32'hbb3f1a15),
	.w8(32'hbbdcc167),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7832),
	.w1(32'hbb8fe895),
	.w2(32'hbbaa9c4c),
	.w3(32'h3b083799),
	.w4(32'h3b7a8342),
	.w5(32'h3bc91cb3),
	.w6(32'h3a89f30d),
	.w7(32'hbb90337c),
	.w8(32'hb7a8a40c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf142),
	.w1(32'hbbb06731),
	.w2(32'hbbab966f),
	.w3(32'h3baeb37d),
	.w4(32'hbc046f07),
	.w5(32'hbb716de3),
	.w6(32'h3b9c9582),
	.w7(32'hbb171a11),
	.w8(32'hba9e6854),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba165f5a),
	.w1(32'hbb92ec2a),
	.w2(32'hbb1d160e),
	.w3(32'hbb111466),
	.w4(32'hbb7f8004),
	.w5(32'h3af55356),
	.w6(32'h3a154cd0),
	.w7(32'h3b205ac0),
	.w8(32'h3ac5bc8e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae90903),
	.w1(32'hbb2fa970),
	.w2(32'h3ba2f24a),
	.w3(32'hbadbef44),
	.w4(32'hbbadf07c),
	.w5(32'hbaee3f87),
	.w6(32'h3b717cb4),
	.w7(32'hbbbcb749),
	.w8(32'hbb24a923),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c63c1),
	.w1(32'hb8dd007e),
	.w2(32'hba9776cf),
	.w3(32'hbc2cf689),
	.w4(32'hbbc674fd),
	.w5(32'hbb947b32),
	.w6(32'hbc1e7ef0),
	.w7(32'hbbd37b46),
	.w8(32'hbb07637a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7db97e),
	.w1(32'hbb977964),
	.w2(32'hbbeb63f7),
	.w3(32'hbb55051e),
	.w4(32'hbbdda3d1),
	.w5(32'hbaa84970),
	.w6(32'hbaaa2e70),
	.w7(32'hbacb621d),
	.w8(32'h3aeecc3b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643ff6),
	.w1(32'hbb304b5c),
	.w2(32'hbb01b739),
	.w3(32'h3b92eacb),
	.w4(32'hbb2d959e),
	.w5(32'h374b6e36),
	.w6(32'h3bbe37d7),
	.w7(32'hbaed1fe4),
	.w8(32'hb8eeb0fb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab006b6),
	.w1(32'hbb01dcf6),
	.w2(32'hbb8a2811),
	.w3(32'hbb3e994b),
	.w4(32'hbb3d1a32),
	.w5(32'hbba5f129),
	.w6(32'hbb086c83),
	.w7(32'hbb5075b9),
	.w8(32'hbbee5c98),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1141b),
	.w1(32'h3b9a162a),
	.w2(32'hb94b167e),
	.w3(32'hbbae6ae5),
	.w4(32'hbb11b7b0),
	.w5(32'hbbc44ea6),
	.w6(32'hbc044102),
	.w7(32'h3ae2bf85),
	.w8(32'hbbe2c468),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827cb9),
	.w1(32'hbb37cbfc),
	.w2(32'hbbbfb24c),
	.w3(32'hbb22a617),
	.w4(32'hba0f0224),
	.w5(32'hbb1d69c6),
	.w6(32'hbb8ec09f),
	.w7(32'hbb9f3165),
	.w8(32'hbb7c4a02),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7539),
	.w1(32'h3aebd8a0),
	.w2(32'hbb35be3c),
	.w3(32'h3c097356),
	.w4(32'hbae4deb0),
	.w5(32'h3c0b54b4),
	.w6(32'h3bb64ff7),
	.w7(32'hbb9376c6),
	.w8(32'hb95e72f4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad632e6),
	.w1(32'hbbab1a1e),
	.w2(32'hbbb65c35),
	.w3(32'hbc1ac9f3),
	.w4(32'h3b1409a3),
	.w5(32'h3b468a34),
	.w6(32'hbb9ddb73),
	.w7(32'h39c3900a),
	.w8(32'hbb2091de),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba052e6),
	.w1(32'h3931c152),
	.w2(32'hb93b4301),
	.w3(32'h3953dd40),
	.w4(32'h3b97af6a),
	.w5(32'h3aa85070),
	.w6(32'h3b33497c),
	.w7(32'h3ad9d6f9),
	.w8(32'h3a6ec005),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb8b51),
	.w1(32'hbba16fdb),
	.w2(32'hbb122d3c),
	.w3(32'hba8e6e8c),
	.w4(32'hb9d6ba3b),
	.w5(32'h38279453),
	.w6(32'h3abf06ba),
	.w7(32'hbb34b583),
	.w8(32'hbc0fbbfe),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8327be),
	.w1(32'h3bef3288),
	.w2(32'hbacad8d1),
	.w3(32'hbc0ac334),
	.w4(32'h3b4f1978),
	.w5(32'h3ba442d2),
	.w6(32'hbc26c24d),
	.w7(32'h3b28f6bd),
	.w8(32'hbabb637d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08fb8f),
	.w1(32'h3a80201b),
	.w2(32'h3b346d8b),
	.w3(32'hbb880678),
	.w4(32'hbb73846b),
	.w5(32'hbb76c3ef),
	.w6(32'hbb84dd28),
	.w7(32'hbbb447be),
	.w8(32'hbba79cb4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd7aa8),
	.w1(32'hbc3957f2),
	.w2(32'hbb947f01),
	.w3(32'hbbae7629),
	.w4(32'hbb47465b),
	.w5(32'h3c0960c8),
	.w6(32'hbb9bbe79),
	.w7(32'hb9d6635b),
	.w8(32'h3b2c4b0d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b7de),
	.w1(32'hb8965871),
	.w2(32'h3bc5cc56),
	.w3(32'h3b1e8ee0),
	.w4(32'hbb144ecb),
	.w5(32'h3b6160c5),
	.w6(32'hba767034),
	.w7(32'hbb75e640),
	.w8(32'hbb89f7a1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f252a),
	.w1(32'h39891da2),
	.w2(32'hbaeb8e8e),
	.w3(32'h3b926874),
	.w4(32'h3b3cc668),
	.w5(32'hbc31b44a),
	.w6(32'h3aa53214),
	.w7(32'hbbdfc33e),
	.w8(32'hbc4ad32a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fda27),
	.w1(32'hbb338fe3),
	.w2(32'h3ac388f7),
	.w3(32'hb71295ec),
	.w4(32'hbb36f862),
	.w5(32'hba94a311),
	.w6(32'hb9154342),
	.w7(32'hbb94f6a5),
	.w8(32'hbb4b634b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9637eb),
	.w1(32'hbb99ad13),
	.w2(32'h3a1678a5),
	.w3(32'hb9252115),
	.w4(32'hbad38607),
	.w5(32'h3b4de451),
	.w6(32'h3b81b696),
	.w7(32'h3b13fcf9),
	.w8(32'h3b6835f1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808078),
	.w1(32'hbb3252b5),
	.w2(32'h39ca7c06),
	.w3(32'hbb1034b8),
	.w4(32'hbb0682a4),
	.w5(32'h38745acb),
	.w6(32'hba832a97),
	.w7(32'hba289f4e),
	.w8(32'hb9595d00),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b7e60),
	.w1(32'hbb0c571c),
	.w2(32'hbc192508),
	.w3(32'hb8fa1b35),
	.w4(32'h39b03151),
	.w5(32'hbad0d899),
	.w6(32'hbb1e48a5),
	.w7(32'h3b951b76),
	.w8(32'h3b74eaad),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6c7b),
	.w1(32'hb90d4e82),
	.w2(32'h3abd768d),
	.w3(32'h3956e953),
	.w4(32'hb90ae6e0),
	.w5(32'h3bcf5bf6),
	.w6(32'h3a8de9bf),
	.w7(32'hbb86b3c5),
	.w8(32'hb9f61c91),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bbb6a),
	.w1(32'h3b7e8414),
	.w2(32'h3bacd2cb),
	.w3(32'hbc44dcb2),
	.w4(32'hbbef3b19),
	.w5(32'hbb9e17c3),
	.w6(32'hbbc2818d),
	.w7(32'hbb6ac9af),
	.w8(32'hbbbbe55b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928310c),
	.w1(32'h3ae64e86),
	.w2(32'h3b344aea),
	.w3(32'hbb920195),
	.w4(32'h3b74c899),
	.w5(32'h3c05ab3a),
	.w6(32'hbbc60743),
	.w7(32'hbbb9e7e6),
	.w8(32'h3b18338e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0ce5),
	.w1(32'hba4bb369),
	.w2(32'h3b9c60be),
	.w3(32'hbb4ea7d5),
	.w4(32'hbafaf839),
	.w5(32'hb9519299),
	.w6(32'hbb03e571),
	.w7(32'hbb824baa),
	.w8(32'hbc3c4c1f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9669df),
	.w1(32'hbae99078),
	.w2(32'hbaa986da),
	.w3(32'hbb19ce06),
	.w4(32'hbbc55b20),
	.w5(32'hbb140e32),
	.w6(32'h3a8ff6fa),
	.w7(32'hbbf0ab1b),
	.w8(32'hbbb399b9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba650f86),
	.w1(32'hbb53161d),
	.w2(32'hbbb87312),
	.w3(32'hbb4c9d70),
	.w4(32'hb7900da9),
	.w5(32'hbb167e63),
	.w6(32'hbc11e45d),
	.w7(32'h3ad24861),
	.w8(32'hbb807ca1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074642),
	.w1(32'hba4fafc1),
	.w2(32'h3bbb94d1),
	.w3(32'h3b7e41b6),
	.w4(32'hba692976),
	.w5(32'hbc6513c7),
	.w6(32'h3c2f824b),
	.w7(32'hba8cb12b),
	.w8(32'hbbf6c435),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9229aa),
	.w1(32'hbbc3cccf),
	.w2(32'hbc496bcc),
	.w3(32'hbb18d7a6),
	.w4(32'hbc069dab),
	.w5(32'hbc22ea7c),
	.w6(32'hbb171ea7),
	.w7(32'hbc08c338),
	.w8(32'hbb853bc7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993d87),
	.w1(32'h3952c167),
	.w2(32'hbbedc9ba),
	.w3(32'h3b324333),
	.w4(32'hbba73c69),
	.w5(32'hbb6b4bfc),
	.w6(32'h3b8ae51a),
	.w7(32'h37b2947d),
	.w8(32'h3bfbfd33),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a10a),
	.w1(32'h39829cc5),
	.w2(32'hbb799de9),
	.w3(32'hbba2f0ef),
	.w4(32'h3ad053d8),
	.w5(32'hbbe1da2c),
	.w6(32'h3c1a32c6),
	.w7(32'h3ba3a4d3),
	.w8(32'hbc08ffb3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2008a),
	.w1(32'hbb820357),
	.w2(32'hbb2726c8),
	.w3(32'h3a7a15e7),
	.w4(32'hbb691fd4),
	.w5(32'hba877b59),
	.w6(32'hbac79779),
	.w7(32'hbb6109b7),
	.w8(32'h3b3e31ff),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f275a),
	.w1(32'hbb94f7ac),
	.w2(32'h3b850d37),
	.w3(32'h39dce9f5),
	.w4(32'hbb44787e),
	.w5(32'h3c248d7e),
	.w6(32'h3934fdc8),
	.w7(32'hb9d4a2d2),
	.w8(32'h3c0d7773),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd85e),
	.w1(32'hbaaffb63),
	.w2(32'hbbcace74),
	.w3(32'h3bbaab56),
	.w4(32'hbbaab6d3),
	.w5(32'h3a2352a8),
	.w6(32'h3a2a2498),
	.w7(32'hbad3fbbf),
	.w8(32'hba0b1745),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a039d),
	.w1(32'hbaa09273),
	.w2(32'h398ab25a),
	.w3(32'h3b2f691b),
	.w4(32'hbb8e58da),
	.w5(32'hbbbb4ded),
	.w6(32'h39aabf8f),
	.w7(32'hbacb370c),
	.w8(32'hbb0e48fd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392486f7),
	.w1(32'h3b935599),
	.w2(32'h3a0cee81),
	.w3(32'hba9b2bed),
	.w4(32'h3b944082),
	.w5(32'h3a9932c9),
	.w6(32'hbb7c6ccc),
	.w7(32'hbac60f98),
	.w8(32'hbb4831cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39266d02),
	.w1(32'h3be74476),
	.w2(32'h39ce117b),
	.w3(32'hb9f2e608),
	.w4(32'h3c14e8c7),
	.w5(32'h3b623f32),
	.w6(32'hb9dc6a5e),
	.w7(32'h3bc0fa7d),
	.w8(32'h3b0b7932),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa6182),
	.w1(32'h3c1f241a),
	.w2(32'h39fa2938),
	.w3(32'h3b439cb9),
	.w4(32'h3bb5df50),
	.w5(32'h3c1a9a02),
	.w6(32'h3c25cf9b),
	.w7(32'hba100024),
	.w8(32'hba2574b2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d9f09),
	.w1(32'h3a3464fd),
	.w2(32'hbb4be1d7),
	.w3(32'h3bd37841),
	.w4(32'h3a87bf7d),
	.w5(32'h3a01a4c7),
	.w6(32'h3bbbbdb9),
	.w7(32'h3c058bbc),
	.w8(32'h3a75db02),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1253e7),
	.w1(32'hbba45867),
	.w2(32'h39631b39),
	.w3(32'h3b4c7158),
	.w4(32'hbbacf836),
	.w5(32'hbb6150a7),
	.w6(32'h3ba28711),
	.w7(32'hbb865455),
	.w8(32'hbba89d11),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26344a),
	.w1(32'hbb11438f),
	.w2(32'hb99aff35),
	.w3(32'hbb1bafe1),
	.w4(32'hba67421d),
	.w5(32'hbb30e7f9),
	.w6(32'hba985c36),
	.w7(32'h3a0fd718),
	.w8(32'hbb2445e0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a4bcc),
	.w1(32'h3bcde314),
	.w2(32'hbaa1bfda),
	.w3(32'hba2b6d1f),
	.w4(32'h3b79efc2),
	.w5(32'hbb750d76),
	.w6(32'h3a3fff49),
	.w7(32'h3be7332d),
	.w8(32'h3b89a1aa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c00d),
	.w1(32'h3a90ce41),
	.w2(32'hbb9dde4a),
	.w3(32'h3b82e422),
	.w4(32'h3b45145a),
	.w5(32'hbbdff753),
	.w6(32'h3b2fdf45),
	.w7(32'h3bc5a1bb),
	.w8(32'hbb12e49f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1539e),
	.w1(32'hbb661ba0),
	.w2(32'hbc1772a1),
	.w3(32'hbb3c06c8),
	.w4(32'hbb270f2f),
	.w5(32'hbb03780d),
	.w6(32'hbc120460),
	.w7(32'hbc5c1ea2),
	.w8(32'hbbfe0121),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e54ae),
	.w1(32'h3a129502),
	.w2(32'h3b6ac5f2),
	.w3(32'hbb0c4a22),
	.w4(32'h3aaeb2db),
	.w5(32'h3bab5184),
	.w6(32'hba7dd0d8),
	.w7(32'hbbb9ccbb),
	.w8(32'hbb8dbfbd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8d20),
	.w1(32'hbb84979b),
	.w2(32'hbb60e700),
	.w3(32'hba3ee6ad),
	.w4(32'hbbcaf8f9),
	.w5(32'hbb875da2),
	.w6(32'h37ad85e8),
	.w7(32'h3a1d0df9),
	.w8(32'hbb697131),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb400667),
	.w1(32'h3bd4fb9b),
	.w2(32'hbb11f4e8),
	.w3(32'h3b78b61b),
	.w4(32'hbaa769b4),
	.w5(32'hbaf5c34a),
	.w6(32'h3b59cbed),
	.w7(32'h3b66106d),
	.w8(32'h3b187ce1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb2118),
	.w1(32'h38c1ab62),
	.w2(32'hbb40eb8c),
	.w3(32'hbb2cb001),
	.w4(32'h3bd29947),
	.w5(32'h3ab5f21d),
	.w6(32'h3b824114),
	.w7(32'h3bc9976d),
	.w8(32'hbbb10f85),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46fe0c),
	.w1(32'hbaad3fde),
	.w2(32'h3ba3b9bf),
	.w3(32'hbb026f51),
	.w4(32'hbabc7267),
	.w5(32'hbb4821bc),
	.w6(32'hbb85a8a7),
	.w7(32'hba0761c2),
	.w8(32'hbb15440a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badbdc6),
	.w1(32'h3befb897),
	.w2(32'h3bc92755),
	.w3(32'hbbf76475),
	.w4(32'h3bea234c),
	.w5(32'h3a544e83),
	.w6(32'hbc1c7c52),
	.w7(32'h3b1d6092),
	.w8(32'hbbaa38df),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d5e9),
	.w1(32'h3ba6e999),
	.w2(32'h3b273956),
	.w3(32'hbac7d391),
	.w4(32'h3bb3b473),
	.w5(32'hb8a22b1f),
	.w6(32'hb5824187),
	.w7(32'h3bbec7bd),
	.w8(32'h379daf34),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af08b8f),
	.w1(32'h3c15ff90),
	.w2(32'h3bfe3d40),
	.w3(32'hbba36e37),
	.w4(32'h3bc05242),
	.w5(32'h3b3362f6),
	.w6(32'hbb25de76),
	.w7(32'h3bbbb4ec),
	.w8(32'hbb348f78),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96f2c2),
	.w1(32'h3b7d4748),
	.w2(32'h3b917300),
	.w3(32'hba7738a1),
	.w4(32'h3b1deae0),
	.w5(32'h3aa7510d),
	.w6(32'hb9cfa8ea),
	.w7(32'h3b4211f7),
	.w8(32'h3b0e2958),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94006d),
	.w1(32'hba8e4945),
	.w2(32'h3a6d226b),
	.w3(32'h3ba29a0a),
	.w4(32'hb9c95fdf),
	.w5(32'hba601857),
	.w6(32'h3a49ac9d),
	.w7(32'hb99f2be4),
	.w8(32'hbb8a907d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6322e0),
	.w1(32'hb9f3db39),
	.w2(32'hbaf78700),
	.w3(32'hbabc7fa1),
	.w4(32'hbad00a4f),
	.w5(32'hbb8dead9),
	.w6(32'h3a1fde02),
	.w7(32'hbaedb748),
	.w8(32'hbbc4d204),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fddfe),
	.w1(32'hbb3f034b),
	.w2(32'hbadf10c4),
	.w3(32'hbc145348),
	.w4(32'hba73caa8),
	.w5(32'h3b21e255),
	.w6(32'hbc0bb7c0),
	.w7(32'hbb04a2e1),
	.w8(32'h3b05ea8d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca40f),
	.w1(32'h3b46fa28),
	.w2(32'h3b1e8dd0),
	.w3(32'h3b1f1d21),
	.w4(32'h3a6cc9b3),
	.w5(32'hbb88cd56),
	.w6(32'h3ba223ff),
	.w7(32'h3b178e83),
	.w8(32'h3b7887bb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb4bd),
	.w1(32'hbbe72cc0),
	.w2(32'hbba7e3e6),
	.w3(32'hbb28e2b1),
	.w4(32'hbb7dc90d),
	.w5(32'hbb990382),
	.w6(32'h3b63eb0b),
	.w7(32'h3bcce7ae),
	.w8(32'hbade9214),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2028d),
	.w1(32'hbba3e87e),
	.w2(32'hbb568711),
	.w3(32'hbbbc8a99),
	.w4(32'hbb132633),
	.w5(32'hbb1302bb),
	.w6(32'hbb81a9f6),
	.w7(32'hbb20376f),
	.w8(32'hbac0446b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84997e),
	.w1(32'hbb9ad952),
	.w2(32'hbc178f68),
	.w3(32'h3b586549),
	.w4(32'hbb0b07ae),
	.w5(32'h3c25583d),
	.w6(32'h3b3d0985),
	.w7(32'h3a7c66d9),
	.w8(32'h3c13f5e8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf94b02),
	.w1(32'h3bb1af16),
	.w2(32'h3b47e40b),
	.w3(32'h3b3885dc),
	.w4(32'hbb93db4f),
	.w5(32'h3b3c2177),
	.w6(32'h3b95a0f0),
	.w7(32'hbbeb68c2),
	.w8(32'h3b9c00a4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee3ee7),
	.w1(32'hbb0f345f),
	.w2(32'hba97fad2),
	.w3(32'h3b583426),
	.w4(32'hbb6cca52),
	.w5(32'h3a7f74eb),
	.w6(32'h3b4effcf),
	.w7(32'hbb184a3a),
	.w8(32'h3a8e926c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc114892),
	.w1(32'hbc4a25bf),
	.w2(32'hba563a0f),
	.w3(32'hbbb27493),
	.w4(32'hbc09e943),
	.w5(32'hbb9a9b37),
	.w6(32'h3afa8e76),
	.w7(32'h3c2ad6dd),
	.w8(32'h3c1ab6aa),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe369e5),
	.w1(32'hbb898ad1),
	.w2(32'hbbf4e553),
	.w3(32'h3ba98b44),
	.w4(32'hbadf119f),
	.w5(32'hbc03b407),
	.w6(32'h3bab65b6),
	.w7(32'h3c0bc122),
	.w8(32'h3c0a787b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad43a),
	.w1(32'hbb97fdbb),
	.w2(32'hbb09d9c9),
	.w3(32'hbb8cd27e),
	.w4(32'h3a324332),
	.w5(32'hba3120b2),
	.w6(32'h3c301a56),
	.w7(32'h3bcc7d60),
	.w8(32'h3b84ee9c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdcef6),
	.w1(32'h3bd6c231),
	.w2(32'h3a537e2b),
	.w3(32'hbb4f326e),
	.w4(32'hbaefc02a),
	.w5(32'hbbcbdba1),
	.w6(32'hba0e0f16),
	.w7(32'hbb27ca16),
	.w8(32'hbc0ebd9d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52d3d),
	.w1(32'hbb8dbba6),
	.w2(32'hbb8af209),
	.w3(32'hbba46bcd),
	.w4(32'h3857fc79),
	.w5(32'h3c14ac15),
	.w6(32'hbc1680c9),
	.w7(32'h3bc3e242),
	.w8(32'h3c006c88),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d0f2a),
	.w1(32'h3b5470b5),
	.w2(32'hba849809),
	.w3(32'h3c1a084d),
	.w4(32'h3bb4e722),
	.w5(32'h3b9a4d8e),
	.w6(32'h3c222734),
	.w7(32'h3c148de0),
	.w8(32'h3c00f596),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ed476),
	.w1(32'h3b405555),
	.w2(32'hba4c6644),
	.w3(32'h3bca1427),
	.w4(32'h3b38664a),
	.w5(32'h3af13783),
	.w6(32'h3ba00ea9),
	.w7(32'h3a08c1c3),
	.w8(32'hb784f403),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3bcd1),
	.w1(32'hbbf474a1),
	.w2(32'hbab65bd9),
	.w3(32'h3b74e727),
	.w4(32'h3ac237e4),
	.w5(32'h3b7c04c2),
	.w6(32'hb9e4dccd),
	.w7(32'hbae8e0a0),
	.w8(32'h3b0e4b7c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae817b),
	.w1(32'hbac683d9),
	.w2(32'hbb60731e),
	.w3(32'hbc028c7a),
	.w4(32'hbba9e021),
	.w5(32'hbc490f4d),
	.w6(32'h39a2c874),
	.w7(32'hba9d31a6),
	.w8(32'hbc04fcad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a67a),
	.w1(32'hba0c0602),
	.w2(32'h3b8e30ef),
	.w3(32'hbc28f2b0),
	.w4(32'hbbc97621),
	.w5(32'hbb5d3c87),
	.w6(32'hbb8f9c5b),
	.w7(32'hbc15eb33),
	.w8(32'hbb5981de),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3af6e),
	.w1(32'h39eb255b),
	.w2(32'h391bdd0d),
	.w3(32'hbbb2dc5a),
	.w4(32'h3b029f1d),
	.w5(32'h3b91445b),
	.w6(32'h3b180c2c),
	.w7(32'h3aa05091),
	.w8(32'h391840b6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976596f),
	.w1(32'h3bd8e4a8),
	.w2(32'h3bb99545),
	.w3(32'h3b0cc291),
	.w4(32'h3b816e7c),
	.w5(32'h3b564750),
	.w6(32'h3ad69e3e),
	.w7(32'hba68871f),
	.w8(32'h3af4c519),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341f70),
	.w1(32'hbc05e256),
	.w2(32'hbbac9d3e),
	.w3(32'h3b28c7f5),
	.w4(32'hbb3d3649),
	.w5(32'hbbeb56f7),
	.w6(32'h3b5a0420),
	.w7(32'hbb4ff8cd),
	.w8(32'hbbc241a0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab60f9),
	.w1(32'hba79bd17),
	.w2(32'hbb85e119),
	.w3(32'hbc16fd44),
	.w4(32'hba069ab8),
	.w5(32'hbbb0f72c),
	.w6(32'hbc224918),
	.w7(32'h3a9eff2b),
	.w8(32'hbb9d360c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6456fb),
	.w1(32'h3bc7d652),
	.w2(32'h3a451d13),
	.w3(32'hbb443b4b),
	.w4(32'h3c196025),
	.w5(32'h3adb5644),
	.w6(32'hba554e54),
	.w7(32'h3bbc4d70),
	.w8(32'h3b64aacd),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa03245),
	.w1(32'h3c848358),
	.w2(32'h3be9b9ba),
	.w3(32'h3b96554e),
	.w4(32'hbb295044),
	.w5(32'hbb937f25),
	.w6(32'h3c04f8bd),
	.w7(32'h3a94ec60),
	.w8(32'hbba09b4d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a8ae4),
	.w1(32'hbb1a506b),
	.w2(32'h3aa9a35d),
	.w3(32'hbb48b2a1),
	.w4(32'hba90555f),
	.w5(32'hbab8ca73),
	.w6(32'h37222bd3),
	.w7(32'hbb820b56),
	.w8(32'h390445d1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed678),
	.w1(32'h3af3680e),
	.w2(32'h3a171ef1),
	.w3(32'h3bbf8b54),
	.w4(32'h3baf07af),
	.w5(32'h3b51b65c),
	.w6(32'h3b5346b2),
	.w7(32'h3b4ac39c),
	.w8(32'h3b25a68b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dc264),
	.w1(32'h3b52a0c4),
	.w2(32'h3c03810e),
	.w3(32'h3acbeb3f),
	.w4(32'hba6c5384),
	.w5(32'h3a3dee07),
	.w6(32'h3a6e6393),
	.w7(32'h3abf5126),
	.w8(32'h3ba05ffa),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea799),
	.w1(32'h3bb3bc87),
	.w2(32'h3aca9ac0),
	.w3(32'h3b2623e7),
	.w4(32'h3a60d78e),
	.w5(32'hbb318056),
	.w6(32'h3b0c53a9),
	.w7(32'h3b5327e1),
	.w8(32'hbaa9dadf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac62e9d),
	.w1(32'h3b20d368),
	.w2(32'hba93f634),
	.w3(32'hbb8fd02e),
	.w4(32'hbb1f48d7),
	.w5(32'h3a349c0e),
	.w6(32'hbb1f5f1e),
	.w7(32'hb872f5e4),
	.w8(32'hbb4d6e82),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad85c4),
	.w1(32'h3ab29b7a),
	.w2(32'hba8bbb39),
	.w3(32'hbbd56a9e),
	.w4(32'h3b6a79df),
	.w5(32'h3b0897f7),
	.w6(32'hbc0c4ecf),
	.w7(32'h3b856e56),
	.w8(32'h3abfcc2f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5af4e),
	.w1(32'hbabd3698),
	.w2(32'hbba4cd7c),
	.w3(32'hbb7c6935),
	.w4(32'hba4f2faf),
	.w5(32'hbbabba39),
	.w6(32'hbae16452),
	.w7(32'hbb3fbae1),
	.w8(32'hbbd3f175),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70d1f),
	.w1(32'hbc9e4d6d),
	.w2(32'hbc0872c6),
	.w3(32'hbc126d73),
	.w4(32'hbc6bd76e),
	.w5(32'hbb776be8),
	.w6(32'hbc2a0007),
	.w7(32'hbc7159f1),
	.w8(32'hbc090bbd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d4560),
	.w1(32'h3be1b5e2),
	.w2(32'h3b62b22b),
	.w3(32'hbabf7296),
	.w4(32'h3bc1e28b),
	.w5(32'h3b6522a1),
	.w6(32'hbc3afa06),
	.w7(32'hbaff8be1),
	.w8(32'h37b48670),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd8a8),
	.w1(32'h3b25a86a),
	.w2(32'hbc42c232),
	.w3(32'hbb12e87f),
	.w4(32'h3c170da7),
	.w5(32'hbc2793c2),
	.w6(32'h3a276a6e),
	.w7(32'h3be04972),
	.w8(32'hbc2c9a53),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f02f),
	.w1(32'h39ca5299),
	.w2(32'hb904f260),
	.w3(32'hbbcd9237),
	.w4(32'hbb337ca2),
	.w5(32'hbbad1f6a),
	.w6(32'hbc110f39),
	.w7(32'hbbbee877),
	.w8(32'hbbdf29f5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c9cc3),
	.w1(32'h3ba2e051),
	.w2(32'h3b57c96a),
	.w3(32'h3b29a653),
	.w4(32'h3b037525),
	.w5(32'h3ba4764a),
	.w6(32'h3a49330d),
	.w7(32'h3b92fafe),
	.w8(32'h37994bd6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbcc3),
	.w1(32'hbb734b10),
	.w2(32'hbbccb36e),
	.w3(32'hbb667b11),
	.w4(32'hbbb6b9d6),
	.w5(32'hbba84392),
	.w6(32'hbaef6325),
	.w7(32'hbb8a6a92),
	.w8(32'hba8aaa0a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec86d9),
	.w1(32'h3bbf60da),
	.w2(32'h3bb84c87),
	.w3(32'hbba5af5c),
	.w4(32'h3b8a7cce),
	.w5(32'h3be752a2),
	.w6(32'hbb85b5e6),
	.w7(32'hbac026d7),
	.w8(32'h3a991ff2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d318),
	.w1(32'hba21c901),
	.w2(32'hbae4e77d),
	.w3(32'hbbdbe0e0),
	.w4(32'hbbbfa7ff),
	.w5(32'hbb2dd7f3),
	.w6(32'hbc1784a9),
	.w7(32'hbb578b90),
	.w8(32'hbb9f0a6d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10b2d0),
	.w1(32'h3b695f50),
	.w2(32'h3b308bc3),
	.w3(32'hbc81c8a8),
	.w4(32'h3bdf04e6),
	.w5(32'h3b2b1651),
	.w6(32'hbc17d091),
	.w7(32'h3bd6834c),
	.w8(32'h3b6acf84),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1a099),
	.w1(32'h3aa28465),
	.w2(32'h3b398742),
	.w3(32'hbbcb8179),
	.w4(32'hbbd1d671),
	.w5(32'h373a93df),
	.w6(32'hbc225cd3),
	.w7(32'hbb704b7e),
	.w8(32'hba08c54b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39672b84),
	.w1(32'hbbca140a),
	.w2(32'hbb48c0da),
	.w3(32'hbb34acdd),
	.w4(32'h3b3878a2),
	.w5(32'h3b56547c),
	.w6(32'hb96da572),
	.w7(32'h3aea3491),
	.w8(32'h3a642275),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16f0e1),
	.w1(32'hba8582e1),
	.w2(32'hbb8e5aef),
	.w3(32'h3ac5bb5a),
	.w4(32'hbabef7cd),
	.w5(32'hbbc653c5),
	.w6(32'hbb3d8d76),
	.w7(32'hbbfb5ed1),
	.w8(32'hbb835466),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449b2f),
	.w1(32'h3afec59c),
	.w2(32'h3ae740ec),
	.w3(32'hbb432631),
	.w4(32'hb93043d1),
	.w5(32'h3b87d820),
	.w6(32'h3a86c082),
	.w7(32'hba582160),
	.w8(32'h3b592262),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b283d),
	.w1(32'h3bb56e8d),
	.w2(32'h3babdfe8),
	.w3(32'h3b8cb855),
	.w4(32'h3bcf6a05),
	.w5(32'h3c137bb0),
	.w6(32'h3be25730),
	.w7(32'h3ba7ebce),
	.w8(32'h3c0502a1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c063),
	.w1(32'h3b85a561),
	.w2(32'hbb324b91),
	.w3(32'h3c510575),
	.w4(32'h3bc36b79),
	.w5(32'h3ac37d8e),
	.w6(32'h3c89ff0f),
	.w7(32'h3b92b8e9),
	.w8(32'h3b6b9fc3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac29dbe),
	.w1(32'h3b6c7bfd),
	.w2(32'hba5edfa2),
	.w3(32'h3c2d5a3a),
	.w4(32'h3b792cdb),
	.w5(32'hbb57b9d4),
	.w6(32'h3c5a93e4),
	.w7(32'h3b8b8a1d),
	.w8(32'hbbd8b1f3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3532ab),
	.w1(32'hbac0b486),
	.w2(32'h39148f69),
	.w3(32'hbbaefc5b),
	.w4(32'hbb41f399),
	.w5(32'hbc0a3663),
	.w6(32'hbc2bd84a),
	.w7(32'hbba66f3f),
	.w8(32'hbb82b19d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b98b),
	.w1(32'hbb772a36),
	.w2(32'hb8496b79),
	.w3(32'hbc315708),
	.w4(32'hbb1a17d0),
	.w5(32'hba7d6c27),
	.w6(32'hbc3ef5f0),
	.w7(32'hba2759e0),
	.w8(32'hbb01c313),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964002),
	.w1(32'h3bb10c3c),
	.w2(32'hbb9c6e0c),
	.w3(32'hba9d85d1),
	.w4(32'h3a54cade),
	.w5(32'hbbf8f45b),
	.w6(32'hb941efb7),
	.w7(32'hbb5b6d66),
	.w8(32'hbbfb305f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5eba),
	.w1(32'h3b8d7e36),
	.w2(32'hbbc89521),
	.w3(32'hbc1ac40c),
	.w4(32'h3b7fc1f9),
	.w5(32'hbc0150bb),
	.w6(32'hbbee53f6),
	.w7(32'hbb12d17d),
	.w8(32'hbc415fed),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866d82),
	.w1(32'hbbae4f33),
	.w2(32'hbc285acb),
	.w3(32'hbc7ace2c),
	.w4(32'hbc541388),
	.w5(32'hbba164fc),
	.w6(32'hbc853a9c),
	.w7(32'hbc2b33d7),
	.w8(32'hbbf6be97),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1548f),
	.w1(32'hbb61d2e2),
	.w2(32'hbca59456),
	.w3(32'hbb987f64),
	.w4(32'h3b232995),
	.w5(32'hbc577eda),
	.w6(32'hbc037fa6),
	.w7(32'hba7abad5),
	.w8(32'hbca50ba2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9b0f),
	.w1(32'hbbe703b5),
	.w2(32'hba679568),
	.w3(32'h3a6cabf8),
	.w4(32'hbb8226a4),
	.w5(32'h3b1882c5),
	.w6(32'hbb549f53),
	.w7(32'h39eca7e9),
	.w8(32'h3b8c162a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad607d5),
	.w1(32'h3a31bac3),
	.w2(32'h3ae78c75),
	.w3(32'h3abe1b3a),
	.w4(32'h3a39c304),
	.w5(32'h3b25114d),
	.w6(32'h3b9ca41d),
	.w7(32'h3a4baf83),
	.w8(32'h3b4c76cb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd2bb6),
	.w1(32'hbbe8cce1),
	.w2(32'h38ff2f6b),
	.w3(32'hba29a0a4),
	.w4(32'hbbfcdf2d),
	.w5(32'hba2d8d05),
	.w6(32'h3ab38e12),
	.w7(32'hbbaf9767),
	.w8(32'hba33e4cb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba5a52),
	.w1(32'h3ba07a83),
	.w2(32'h3b455d03),
	.w3(32'h3a5fc70b),
	.w4(32'h3c0089c9),
	.w5(32'h3b2ae1a6),
	.w6(32'hbaae2faf),
	.w7(32'h3bf8b098),
	.w8(32'h3b98fefa),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8461e),
	.w1(32'hbaca5b2c),
	.w2(32'hbaee7afd),
	.w3(32'h3a8d49d1),
	.w4(32'hbb1a33e1),
	.w5(32'hbba9ce01),
	.w6(32'hb9cb8025),
	.w7(32'hbb0a5f21),
	.w8(32'hbb8ab0d3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a894d19),
	.w1(32'h3b031438),
	.w2(32'h3b4ce50f),
	.w3(32'h3a0033a0),
	.w4(32'hbadf4d02),
	.w5(32'hba8133fa),
	.w6(32'h3684e9bf),
	.w7(32'h3aa2a88a),
	.w8(32'h3b06a586),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea75c2),
	.w1(32'hb993be9d),
	.w2(32'hbb15fef9),
	.w3(32'h3b090dce),
	.w4(32'hbb31af4f),
	.w5(32'hbb97e193),
	.w6(32'h3b9bd913),
	.w7(32'h3a39ea00),
	.w8(32'hba8e7c5a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c3d5),
	.w1(32'h3bb8e4a5),
	.w2(32'h3b815207),
	.w3(32'hb8806b8a),
	.w4(32'h3b5c345f),
	.w5(32'h3b2c6f5c),
	.w6(32'hbb611b4c),
	.w7(32'h3b1f5b84),
	.w8(32'hba94dd64),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21083e),
	.w1(32'h3b39614b),
	.w2(32'hbaebf01e),
	.w3(32'h3b92affa),
	.w4(32'h3b819eae),
	.w5(32'h3a4efc0d),
	.w6(32'h3b218382),
	.w7(32'h3b405ae5),
	.w8(32'h39594fce),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38409),
	.w1(32'hbc05a59a),
	.w2(32'hbbc1e0d4),
	.w3(32'hbbf9e2cc),
	.w4(32'hbc2b3642),
	.w5(32'hbbc597fa),
	.w6(32'hbc135dd5),
	.w7(32'hbbe7bbbb),
	.w8(32'hbb860006),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041edd),
	.w1(32'h3a00aa94),
	.w2(32'hbb6f3f69),
	.w3(32'h3c08096a),
	.w4(32'h3a3e494b),
	.w5(32'hb90e72cd),
	.w6(32'h3c5498e5),
	.w7(32'h3a7c3988),
	.w8(32'hbab9852a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93fed7),
	.w1(32'h3b8283b9),
	.w2(32'h3af81838),
	.w3(32'hbb98ac89),
	.w4(32'h3ba250d3),
	.w5(32'h3b0e9a13),
	.w6(32'hbb99f2b4),
	.w7(32'h3b5119fa),
	.w8(32'h3b564819),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a151),
	.w1(32'hbb691a1a),
	.w2(32'hb9ea363e),
	.w3(32'hba975484),
	.w4(32'hbb1ca052),
	.w5(32'h3b9c6599),
	.w6(32'h3ac4f535),
	.w7(32'hb9874da1),
	.w8(32'h3c1c917b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874330),
	.w1(32'h3ab1a9e2),
	.w2(32'hbbaf03cf),
	.w3(32'h3ba2ede6),
	.w4(32'h3bf1f9c3),
	.w5(32'hbb3f8954),
	.w6(32'h3b9a4c92),
	.w7(32'hba28e60a),
	.w8(32'hbbb6e57d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31af2e),
	.w1(32'h3b3e9f94),
	.w2(32'hba92ddb3),
	.w3(32'h39a72263),
	.w4(32'hba8ffcf6),
	.w5(32'hba3a1775),
	.w6(32'hbb8dd130),
	.w7(32'h3a855962),
	.w8(32'h3b8d1d29),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66114d),
	.w1(32'hbc8af2dd),
	.w2(32'hbb1d24ce),
	.w3(32'hb9492a32),
	.w4(32'hbc96296f),
	.w5(32'hbbe2f2f0),
	.w6(32'h3bddd7c5),
	.w7(32'hbc92023a),
	.w8(32'hbbf380d6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e9976),
	.w1(32'h3abe7fc1),
	.w2(32'h3acb17a5),
	.w3(32'hbc916d67),
	.w4(32'h3b2d0c55),
	.w5(32'h3b567c39),
	.w6(32'hbcbf5e67),
	.w7(32'h39e64b59),
	.w8(32'h3b2d1770),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf3f0),
	.w1(32'h3bbd955a),
	.w2(32'h3b253270),
	.w3(32'hbb60c401),
	.w4(32'h3b12fefe),
	.w5(32'h39212e0e),
	.w6(32'hbb5cccdb),
	.w7(32'h3a8940bd),
	.w8(32'h3bbf53ae),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5b30),
	.w1(32'h3b6b9dd3),
	.w2(32'h3b28a50c),
	.w3(32'h3b31a337),
	.w4(32'h3a5d2c78),
	.w5(32'h3b5a3fd8),
	.w6(32'h3b50873c),
	.w7(32'hbb06eb24),
	.w8(32'h3b947e71),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a9803),
	.w1(32'h3c146da1),
	.w2(32'h3bc4584c),
	.w3(32'h3b590883),
	.w4(32'h3ba83a42),
	.w5(32'h3b7213ad),
	.w6(32'h3aa894b8),
	.w7(32'h3b83a71b),
	.w8(32'h3ba23a4d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071a2a),
	.w1(32'hb938f1cd),
	.w2(32'hbb85baa1),
	.w3(32'h3b84d890),
	.w4(32'h3a946a93),
	.w5(32'hbb32d73b),
	.w6(32'h3c1be568),
	.w7(32'hba56669b),
	.w8(32'hba176664),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364730a5),
	.w1(32'h3bab8821),
	.w2(32'hbaa8045c),
	.w3(32'hb925179c),
	.w4(32'h3b7e0d4e),
	.w5(32'hbb241369),
	.w6(32'hbbc2ef66),
	.w7(32'h3ac3f65c),
	.w8(32'hbaca6ab0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a67c),
	.w1(32'h3a10846c),
	.w2(32'h39582a79),
	.w3(32'hb9a04069),
	.w4(32'hb9b2a3be),
	.w5(32'hbab96300),
	.w6(32'h3b8042d2),
	.w7(32'h3b0a12d2),
	.w8(32'hba136adb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4ac2),
	.w1(32'h3bacb7af),
	.w2(32'h3b9b176a),
	.w3(32'h3abc306c),
	.w4(32'h3affeca5),
	.w5(32'h3a2534cc),
	.w6(32'h39338753),
	.w7(32'hbafe0bcc),
	.w8(32'h39ba496a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule