module layer_10_featuremap_25(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aacd2),
	.w1(32'h3b505a09),
	.w2(32'h3b96d00c),
	.w3(32'h3c031a62),
	.w4(32'h3ac31c76),
	.w5(32'h3c81d2cf),
	.w6(32'h3c5bc36d),
	.w7(32'h3a1b021d),
	.w8(32'h3d083417),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3655b2),
	.w1(32'hbc2e35f4),
	.w2(32'hbb30b5fd),
	.w3(32'h3aee8a24),
	.w4(32'hbbbd05ff),
	.w5(32'hbbddd0f0),
	.w6(32'h3ca256c9),
	.w7(32'h3bc951ac),
	.w8(32'h3ba37262),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba950),
	.w1(32'h3bb8b77f),
	.w2(32'h3c82e53f),
	.w3(32'hbc2ed860),
	.w4(32'hba2d0620),
	.w5(32'h3c777348),
	.w6(32'hbba0b5c1),
	.w7(32'hbc0a3e68),
	.w8(32'h3c83384b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8ccfa),
	.w1(32'h3c613e5b),
	.w2(32'hbc1552f8),
	.w3(32'h3cedb2b6),
	.w4(32'h3cb6f766),
	.w5(32'hbbf3467e),
	.w6(32'h3cc98de5),
	.w7(32'h3c2d5e63),
	.w8(32'hba43bccc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaeade),
	.w1(32'hbb430406),
	.w2(32'hbc73f96f),
	.w3(32'hbc91092c),
	.w4(32'hbc7fbb5c),
	.w5(32'hbba737c2),
	.w6(32'hbc11dbbb),
	.w7(32'hbbedd955),
	.w8(32'h3b7509f0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25dd91),
	.w1(32'h3c366aad),
	.w2(32'hbb799afa),
	.w3(32'hbbbf0a77),
	.w4(32'h3b603a1d),
	.w5(32'hbaa05c71),
	.w6(32'hb7d1a59f),
	.w7(32'hbb185d64),
	.w8(32'hbb5313e8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab469cf),
	.w1(32'h3b5d8595),
	.w2(32'hbbb0514a),
	.w3(32'h3b253b9c),
	.w4(32'h3bbd7aef),
	.w5(32'hbb19f81d),
	.w6(32'hbb058bee),
	.w7(32'hba1e5530),
	.w8(32'hbb8c2e78),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb559482),
	.w1(32'h38afe625),
	.w2(32'hbb5b825c),
	.w3(32'hbb095481),
	.w4(32'hbb6a9bcf),
	.w5(32'hbc129809),
	.w6(32'hba224e92),
	.w7(32'h3bcb92bd),
	.w8(32'hbc43000b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9682),
	.w1(32'hbb24b787),
	.w2(32'h3be99185),
	.w3(32'h3bc253de),
	.w4(32'h3b4e5c13),
	.w5(32'h3b311f5e),
	.w6(32'hba29b026),
	.w7(32'h3bb729a2),
	.w8(32'hbc5d5758),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca3e03),
	.w1(32'hbb7ff922),
	.w2(32'hbac07c2d),
	.w3(32'h3b9e9034),
	.w4(32'h38d5bf23),
	.w5(32'hba9328a0),
	.w6(32'hbc2c40aa),
	.w7(32'hbbc53106),
	.w8(32'h3a388a7b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39314fd1),
	.w1(32'h39c543d1),
	.w2(32'h3c1b6f0d),
	.w3(32'hbae5cc23),
	.w4(32'hb942a9f7),
	.w5(32'h3ca1e160),
	.w6(32'h3a0316e2),
	.w7(32'hba3fd965),
	.w8(32'h3c933ae2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab354f),
	.w1(32'h3c777800),
	.w2(32'hb91b118e),
	.w3(32'h3cd66de1),
	.w4(32'h3cb9f147),
	.w5(32'hbafb7aae),
	.w6(32'h3cc8469f),
	.w7(32'h3cb414a6),
	.w8(32'hbb2f7157),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971e475),
	.w1(32'hbb6145b0),
	.w2(32'h39ff62d5),
	.w3(32'h3aefbb8e),
	.w4(32'h3a4da1f3),
	.w5(32'h375e0887),
	.w6(32'hba4ba161),
	.w7(32'h39fb526f),
	.w8(32'h3baf71e2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a662e),
	.w1(32'hbb8eb27a),
	.w2(32'hbbc6d804),
	.w3(32'hba338052),
	.w4(32'hbb453308),
	.w5(32'h3b2ba0c5),
	.w6(32'h3b004205),
	.w7(32'h3af2c667),
	.w8(32'h3be4b3f2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09379d),
	.w1(32'h3b81f0ef),
	.w2(32'hbc0e7ef0),
	.w3(32'hbc2d70c2),
	.w4(32'hbbe91e69),
	.w5(32'hbb4dc446),
	.w6(32'hbb89e7e0),
	.w7(32'hbb700266),
	.w8(32'h3bd86ecb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391dfee2),
	.w1(32'h3b0ac126),
	.w2(32'hb9f7f9de),
	.w3(32'h3a9ac034),
	.w4(32'h3b17857e),
	.w5(32'h39d36c43),
	.w6(32'h3b9123c3),
	.w7(32'h3bdc8fb7),
	.w8(32'h3b56c122),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b0aa),
	.w1(32'h3af2b715),
	.w2(32'hbbbadd39),
	.w3(32'h3a2602f4),
	.w4(32'h3b13b1f2),
	.w5(32'h39b62dc6),
	.w6(32'h3b10d8bc),
	.w7(32'h3a3d8a9f),
	.w8(32'h3bf8951f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dc26e),
	.w1(32'h3bcba85d),
	.w2(32'h3a30fafd),
	.w3(32'h3ab7a1b1),
	.w4(32'h3b572b7a),
	.w5(32'h3a9649dd),
	.w6(32'h3bd0375f),
	.w7(32'h3b519737),
	.w8(32'h3aafa423),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c77c9),
	.w1(32'hbbacf376),
	.w2(32'h3c6592ad),
	.w3(32'hbc0fe991),
	.w4(32'hbc1753f8),
	.w5(32'h3c3c405e),
	.w6(32'hbbbe0930),
	.w7(32'hbb3b634c),
	.w8(32'h3be50698),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86dd40),
	.w1(32'h3c2d701b),
	.w2(32'hbbfacccd),
	.w3(32'h3cc22376),
	.w4(32'h3ca505cd),
	.w5(32'hbb8f9d08),
	.w6(32'h3cbffc3b),
	.w7(32'h3c120520),
	.w8(32'h3b547183),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d326),
	.w1(32'h3aa44ac6),
	.w2(32'hbc00a978),
	.w3(32'hbc5cef77),
	.w4(32'hbbd93b4a),
	.w5(32'hbc83bd09),
	.w6(32'hbb9e05e3),
	.w7(32'hbb90677b),
	.w8(32'hbba681b3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cc980),
	.w1(32'h392e82a2),
	.w2(32'hbbee0236),
	.w3(32'hbca6ff57),
	.w4(32'hbc7f71c3),
	.w5(32'h3a9e020d),
	.w6(32'hbcbadc8f),
	.w7(32'hbcae2b88),
	.w8(32'h39e8a794),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878e70),
	.w1(32'h3b18a3b8),
	.w2(32'hbb79a690),
	.w3(32'h3bf89d9e),
	.w4(32'h3b8acbd2),
	.w5(32'hb979d8c6),
	.w6(32'h3b6ef42f),
	.w7(32'h3aa85bee),
	.w8(32'h3ac19fc3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49cc3f),
	.w1(32'hba109b90),
	.w2(32'h3bb17765),
	.w3(32'hbaa21ca4),
	.w4(32'hbb3e0e0c),
	.w5(32'h3c12f0e4),
	.w6(32'h3b49ad3e),
	.w7(32'hb9e31bdc),
	.w8(32'h36b05607),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a912aac),
	.w1(32'h3b372454),
	.w2(32'h3c35bcae),
	.w3(32'h3c3d91c7),
	.w4(32'h3b857f7c),
	.w5(32'h3cae4e1c),
	.w6(32'h3bec33a8),
	.w7(32'h3ba2470d),
	.w8(32'h3c81b9cf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e16fa),
	.w1(32'h3bf76082),
	.w2(32'h3c922d5e),
	.w3(32'h3cb8239c),
	.w4(32'h3c661660),
	.w5(32'h3c4c20a5),
	.w6(32'h3cec3151),
	.w7(32'h3cd74bc6),
	.w8(32'h3c48afe4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f947b),
	.w1(32'h3c178653),
	.w2(32'h3a3cc252),
	.w3(32'h3cc0fd82),
	.w4(32'h3c94971a),
	.w5(32'hba32aad6),
	.w6(32'h3c6f9023),
	.w7(32'h3c06594e),
	.w8(32'h3a7a3bad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8968046),
	.w1(32'h39860160),
	.w2(32'hb9819efb),
	.w3(32'hbae1a645),
	.w4(32'hbab42574),
	.w5(32'hbb01ed78),
	.w6(32'h399ffe06),
	.w7(32'h3a321c9b),
	.w8(32'hba00e716),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1241e9),
	.w1(32'hbad95188),
	.w2(32'h3b10b1a9),
	.w3(32'hbb2be197),
	.w4(32'hbb67c67b),
	.w5(32'h3b892230),
	.w6(32'hba9a7bc6),
	.w7(32'hbb049008),
	.w8(32'h3bcac7df),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb405b),
	.w1(32'hb9c8da3f),
	.w2(32'hb9af0df5),
	.w3(32'h3b1115a7),
	.w4(32'h39d99e5f),
	.w5(32'hbb84bb2c),
	.w6(32'h3bb59b1d),
	.w7(32'hbaca21b0),
	.w8(32'h3a6124a2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0fcb2),
	.w1(32'hbaf83c11),
	.w2(32'h3b8e381f),
	.w3(32'hbc2c37a4),
	.w4(32'hbbe86ada),
	.w5(32'h3b898c43),
	.w6(32'hbb9fcbfd),
	.w7(32'hbaadc03c),
	.w8(32'h3c100259),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c341),
	.w1(32'h3b8ffc84),
	.w2(32'h3b85e9b2),
	.w3(32'h3bb4011f),
	.w4(32'h3b287a18),
	.w5(32'hba31bd06),
	.w6(32'h3bc9d33f),
	.w7(32'h3bc04d04),
	.w8(32'h3b536379),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8392b3),
	.w1(32'h3c045677),
	.w2(32'hbc1b0e95),
	.w3(32'hbae4105d),
	.w4(32'hba98859a),
	.w5(32'hbc72ac9b),
	.w6(32'h3b904518),
	.w7(32'h3ba987ae),
	.w8(32'hbc0977d5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84dcb1),
	.w1(32'hbc4b41b0),
	.w2(32'h3849cb62),
	.w3(32'hbccf0fc3),
	.w4(32'hbca02ca9),
	.w5(32'hb8229f9d),
	.w6(32'hbc8b6e67),
	.w7(32'hbc381dd4),
	.w8(32'h39d35158),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c6ae3),
	.w1(32'h3bd8db48),
	.w2(32'hbb6961d9),
	.w3(32'h348b0724),
	.w4(32'h3b829463),
	.w5(32'hbaf5ffca),
	.w6(32'hba6193a8),
	.w7(32'h3bacf445),
	.w8(32'hbb79ef20),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f1e39),
	.w1(32'hbb269d35),
	.w2(32'h3ac44b2d),
	.w3(32'h3ac98bd7),
	.w4(32'hb9285c2a),
	.w5(32'h3aa811df),
	.w6(32'hba306915),
	.w7(32'hbb4f7db1),
	.w8(32'h3898c663),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22948d),
	.w1(32'h3bbd79b4),
	.w2(32'hbc2e091c),
	.w3(32'h3ada2f3f),
	.w4(32'h3b4cdde7),
	.w5(32'hbc867314),
	.w6(32'hbae13cf4),
	.w7(32'h3ad0e2fa),
	.w8(32'hbc22075d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e29c6),
	.w1(32'hbc6885ac),
	.w2(32'h3a5a7057),
	.w3(32'hbcd91a7c),
	.w4(32'hbcbb44db),
	.w5(32'h3a9e3eed),
	.w6(32'hbc93a03b),
	.w7(32'hbc61220b),
	.w8(32'h3a305528),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3acdb3),
	.w1(32'h3b078b15),
	.w2(32'h3ad1f208),
	.w3(32'h39218e43),
	.w4(32'h3b29d760),
	.w5(32'h3b215fd3),
	.w6(32'h39ba6ce8),
	.w7(32'h3b05c5c9),
	.w8(32'h3b56fa0d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a194f),
	.w1(32'hbb92e0d1),
	.w2(32'hb9cc99bf),
	.w3(32'hbac0c8e0),
	.w4(32'hbbb85264),
	.w5(32'hba848d2e),
	.w6(32'h3a9f41a4),
	.w7(32'hbbb607fb),
	.w8(32'h3b015e00),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9591bf8),
	.w1(32'h3ae1d3f9),
	.w2(32'h3a666a70),
	.w3(32'hbabf8f3c),
	.w4(32'h3a472f76),
	.w5(32'hba815ef5),
	.w6(32'h39f6d443),
	.w7(32'h3ac195b2),
	.w8(32'hbb3278d4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e892f),
	.w1(32'h3b38c89f),
	.w2(32'hba8349bd),
	.w3(32'h3a159d1e),
	.w4(32'h3b456061),
	.w5(32'hba3ac500),
	.w6(32'h3a371c4c),
	.w7(32'h39ce5f40),
	.w8(32'hb9ce65ce),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8cb8d),
	.w1(32'hbb6bbdf5),
	.w2(32'hbb26615e),
	.w3(32'h3ab9ff21),
	.w4(32'h3a14ca14),
	.w5(32'h3a926236),
	.w6(32'h3abadaa5),
	.w7(32'h3acbcaec),
	.w8(32'hbb6f0133),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c2f0),
	.w1(32'h3a5fe998),
	.w2(32'h3af5ad14),
	.w3(32'h3c0dfefc),
	.w4(32'h3bd32624),
	.w5(32'h3aaa56d8),
	.w6(32'h3b5019d1),
	.w7(32'h3a2993e5),
	.w8(32'hba82ac6b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1101d),
	.w1(32'hbb861dd8),
	.w2(32'h3bca1ca2),
	.w3(32'hbb8f25af),
	.w4(32'hbbb2a8d9),
	.w5(32'h3b49b5f7),
	.w6(32'hbaceb057),
	.w7(32'hbb92805e),
	.w8(32'h3bfd248f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96aed7),
	.w1(32'h3bcf7c47),
	.w2(32'hba80334b),
	.w3(32'hbaa34a2b),
	.w4(32'h3b761763),
	.w5(32'hbaa05f40),
	.w6(32'h3b257157),
	.w7(32'h3bb467c7),
	.w8(32'hb94daa80),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a159603),
	.w1(32'hb930c88e),
	.w2(32'h3b9c74cf),
	.w3(32'h3ae8e6ae),
	.w4(32'h39982f9c),
	.w5(32'h3b255f03),
	.w6(32'h3ab0897e),
	.w7(32'hbabd71b1),
	.w8(32'h3b8df167),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18fa30),
	.w1(32'h3c1af418),
	.w2(32'hbba670c0),
	.w3(32'h3ba7d406),
	.w4(32'h3c05bb65),
	.w5(32'hbaa639a4),
	.w6(32'h3b9e271e),
	.w7(32'h3bb54032),
	.w8(32'hbbe1a88d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38180f),
	.w1(32'hbb81196d),
	.w2(32'h3b0b8ad1),
	.w3(32'h3bdca777),
	.w4(32'h3ad37917),
	.w5(32'h3a4115ac),
	.w6(32'hb95efd14),
	.w7(32'hbba631e8),
	.w8(32'h3bc8f847),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0a6c8),
	.w1(32'hba256b90),
	.w2(32'hba156b7c),
	.w3(32'h3b35fb14),
	.w4(32'h3b638258),
	.w5(32'h39af1358),
	.w6(32'h3b651e58),
	.w7(32'h3ba58a04),
	.w8(32'hbaf21932),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d602),
	.w1(32'hbabcca61),
	.w2(32'h3ba8b9a4),
	.w3(32'hbb1e1644),
	.w4(32'hbaa8e142),
	.w5(32'h3b07d8a1),
	.w6(32'hba84bbed),
	.w7(32'hbb86ce8e),
	.w8(32'hba6097c8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1228bb),
	.w1(32'h3b349d05),
	.w2(32'hba9d47b1),
	.w3(32'hb9ca405a),
	.w4(32'h3a3e6807),
	.w5(32'h3a403863),
	.w6(32'hbb86380b),
	.w7(32'hbb229e1e),
	.w8(32'h3a9344bc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c9784),
	.w1(32'hbaa8c13e),
	.w2(32'h3b669057),
	.w3(32'h39bc2168),
	.w4(32'hbb6805d3),
	.w5(32'h3b0cc33a),
	.w6(32'hbba04db0),
	.w7(32'hbb5eefcd),
	.w8(32'h3ba53614),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ffc7),
	.w1(32'h3c117de6),
	.w2(32'h3baa6441),
	.w3(32'h3ab871e2),
	.w4(32'h3bc06fda),
	.w5(32'h3bee75a4),
	.w6(32'h3bcf6c05),
	.w7(32'h3c2893c4),
	.w8(32'h3b799109),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bce61),
	.w1(32'h3b5ab722),
	.w2(32'h3b32ab88),
	.w3(32'h3b00dc1d),
	.w4(32'h3b040a1f),
	.w5(32'h3ac86195),
	.w6(32'h3b7fb263),
	.w7(32'h3b54674c),
	.w8(32'h3ba66104),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7415aa),
	.w1(32'h3bb14f47),
	.w2(32'hb9f93c6f),
	.w3(32'hbae0cba1),
	.w4(32'hba8c9dd9),
	.w5(32'h3b4f62b7),
	.w6(32'h3b910835),
	.w7(32'h3be7d2f7),
	.w8(32'h3aa36b03),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811a5a),
	.w1(32'h3a8a5dde),
	.w2(32'hbad3b892),
	.w3(32'hbb660d59),
	.w4(32'hba70e4e8),
	.w5(32'hbb848ff8),
	.w6(32'h3a050350),
	.w7(32'h398a8011),
	.w8(32'hbbaabe00),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e2740),
	.w1(32'hbb33c85b),
	.w2(32'hb9c75d14),
	.w3(32'hbbc1fc0c),
	.w4(32'hbbad5c21),
	.w5(32'hb928142a),
	.w6(32'hbb98f686),
	.w7(32'hbb82ad10),
	.w8(32'h39a46352),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aab448),
	.w1(32'h3b7cfc26),
	.w2(32'h3ad44a2c),
	.w3(32'hbaaeaf24),
	.w4(32'h3b424f0d),
	.w5(32'hbabbe735),
	.w6(32'h3a4303a0),
	.w7(32'h3b9331b2),
	.w8(32'h39919312),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68132e),
	.w1(32'h3b81699a),
	.w2(32'h3a4e6b93),
	.w3(32'hba326db9),
	.w4(32'h3b0df31a),
	.w5(32'hba665d96),
	.w6(32'h3ae64487),
	.w7(32'h3b8e1c7a),
	.w8(32'hbab7bba1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20859a),
	.w1(32'hb9f8a93d),
	.w2(32'h3a1bc117),
	.w3(32'h39368723),
	.w4(32'h3af0719a),
	.w5(32'h3a8170e3),
	.w6(32'hbb28e093),
	.w7(32'hba98f1f4),
	.w8(32'h3b467147),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39e992),
	.w1(32'h3b7c47dd),
	.w2(32'hbb111707),
	.w3(32'h3b472da9),
	.w4(32'h3b6d2aee),
	.w5(32'hbb460699),
	.w6(32'h3b3266e0),
	.w7(32'h3b860499),
	.w8(32'hbbba2363),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a19e3),
	.w1(32'hbbab09e3),
	.w2(32'h3b367b82),
	.w3(32'hbb566739),
	.w4(32'hbbb25cb2),
	.w5(32'hbb01dd1c),
	.w6(32'hbb89875c),
	.w7(32'hbba64043),
	.w8(32'h3a24d1f0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaba62b),
	.w1(32'h3adde829),
	.w2(32'h3b71bccc),
	.w3(32'hbb76b0b1),
	.w4(32'hbb87db01),
	.w5(32'hbade0032),
	.w6(32'hbac17af6),
	.w7(32'hbab74fe0),
	.w8(32'h3b8d98b4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae31b78),
	.w1(32'h3b5c71b8),
	.w2(32'h3a28f071),
	.w3(32'h3ade98ca),
	.w4(32'hbaa7672e),
	.w5(32'h39221f3e),
	.w6(32'h3a27e964),
	.w7(32'h3b2e9443),
	.w8(32'h3966f983),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf3910),
	.w1(32'h3a89ee5a),
	.w2(32'h3a8627da),
	.w3(32'h39e2d867),
	.w4(32'h3a050d1c),
	.w5(32'h3a1d29e1),
	.w6(32'h39102568),
	.w7(32'h39c5e8a8),
	.w8(32'h3ad7a9c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e8a0b),
	.w1(32'h3b12e8c3),
	.w2(32'hb9dc8ec5),
	.w3(32'hb78693a4),
	.w4(32'h3acd1997),
	.w5(32'h362d8aff),
	.w6(32'h3ad03b87),
	.w7(32'h3b655d8f),
	.w8(32'h3b06f102),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b340d2),
	.w1(32'hbaae9bc8),
	.w2(32'hbb57e12f),
	.w3(32'hbba41597),
	.w4(32'hbb174755),
	.w5(32'hbadef248),
	.w6(32'hbb8ef27c),
	.w7(32'hbb17cb7b),
	.w8(32'hbb422a2e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b64f1),
	.w1(32'hbb6f35e8),
	.w2(32'hbb3e1d16),
	.w3(32'hbb98642c),
	.w4(32'hbb69ca40),
	.w5(32'hbb845b14),
	.w6(32'hbb8e8861),
	.w7(32'hbb4ea396),
	.w8(32'hbb50447e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6d11),
	.w1(32'hbb3fc381),
	.w2(32'hbaab8d4c),
	.w3(32'hbb40f36d),
	.w4(32'hbb68a924),
	.w5(32'hbad69db9),
	.w6(32'hbadf32b6),
	.w7(32'hbb1095cd),
	.w8(32'hbaa19702),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba70da),
	.w1(32'hbb01c0b7),
	.w2(32'h3aae66e5),
	.w3(32'hbaa18bea),
	.w4(32'hbb3def1d),
	.w5(32'h3b044937),
	.w6(32'hbad38dca),
	.w7(32'hbb80f55a),
	.w8(32'h3ae234d1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fa080),
	.w1(32'h3986b14d),
	.w2(32'hbaf34534),
	.w3(32'hba38af90),
	.w4(32'hba14fe02),
	.w5(32'h38c699c3),
	.w6(32'h3ad9d287),
	.w7(32'hb98dc4cf),
	.w8(32'h3a3f0caf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4e643),
	.w1(32'h3a195019),
	.w2(32'h3b3c18d1),
	.w3(32'hba857513),
	.w4(32'h3a3cf591),
	.w5(32'h3b1af18e),
	.w6(32'hbb29ef85),
	.w7(32'h3a0b1203),
	.w8(32'h3a29f37b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75c490),
	.w1(32'h3b58261c),
	.w2(32'hbbf6c34a),
	.w3(32'h3ba3fc5f),
	.w4(32'h3b9e6ef4),
	.w5(32'hbbb2ca10),
	.w6(32'h3b41c1c1),
	.w7(32'h3ac75c5c),
	.w8(32'hbbea6cbd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20feaa),
	.w1(32'hbbb84f0e),
	.w2(32'h3b8e8c0a),
	.w3(32'h3b101ba0),
	.w4(32'hba34a052),
	.w5(32'h3b904ed7),
	.w6(32'hb9fbaf7c),
	.w7(32'hbb9cca58),
	.w8(32'h3b8dcd43),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818183),
	.w1(32'h3bd07b0e),
	.w2(32'hbafe9a1b),
	.w3(32'h3bb63ab9),
	.w4(32'h3bf6a5d9),
	.w5(32'hbb09c05a),
	.w6(32'h3bb49276),
	.w7(32'h3c099813),
	.w8(32'h3af605b1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9179636),
	.w1(32'h3922b165),
	.w2(32'hba84b91b),
	.w3(32'hb992a8ff),
	.w4(32'hbabf90ac),
	.w5(32'h3b0b6662),
	.w6(32'hbabb0cd6),
	.w7(32'hbaefdf95),
	.w8(32'h3a43d365),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3203a4),
	.w1(32'h391554f6),
	.w2(32'h3a2cd6c9),
	.w3(32'hb86a2e1e),
	.w4(32'h3b028887),
	.w5(32'hb9c45567),
	.w6(32'hb9f4ce87),
	.w7(32'hbb58783e),
	.w8(32'h3acb360a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adff333),
	.w1(32'h3a4af615),
	.w2(32'h39c8d162),
	.w3(32'h3b438265),
	.w4(32'h39d35a90),
	.w5(32'hbafb00ab),
	.w6(32'h3ba5d661),
	.w7(32'h3a83cc48),
	.w8(32'h3a8ae62e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dd2660),
	.w1(32'h3a83f1b6),
	.w2(32'h3a8932de),
	.w3(32'hbab6d639),
	.w4(32'hba58e0bc),
	.w5(32'h39cc631a),
	.w6(32'h3a952a04),
	.w7(32'h3aef2610),
	.w8(32'h3916b2b8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceeaf8),
	.w1(32'h3b184e91),
	.w2(32'hb942c009),
	.w3(32'h3a8ab163),
	.w4(32'h3ad72af4),
	.w5(32'hbb0de619),
	.w6(32'h3aa14dc4),
	.w7(32'h3b0c9607),
	.w8(32'h3a9a19ae),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2be1c),
	.w1(32'h3a1cd584),
	.w2(32'hbbe1da94),
	.w3(32'hbba9a80d),
	.w4(32'hbad05a8f),
	.w5(32'hbb556021),
	.w6(32'h3909a571),
	.w7(32'h3b5920be),
	.w8(32'hbb9ce9ed),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa019),
	.w1(32'hbb43f1b0),
	.w2(32'hbb209a1b),
	.w3(32'hbbb9c0d4),
	.w4(32'hbb5446d0),
	.w5(32'h39f66d3a),
	.w6(32'hbbe877a9),
	.w7(32'hbba6df5c),
	.w8(32'h39fc74b0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9871c),
	.w1(32'hbb0b3e38),
	.w2(32'hbb036595),
	.w3(32'hba474da8),
	.w4(32'hbae9b292),
	.w5(32'hbb0d27a7),
	.w6(32'hba2263c9),
	.w7(32'hbb909f9b),
	.w8(32'hbb091f29),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fec6),
	.w1(32'hba43988d),
	.w2(32'h3bd67c04),
	.w3(32'hb9f86d5e),
	.w4(32'hbb133c38),
	.w5(32'h3b84cd96),
	.w6(32'h3a22740d),
	.w7(32'h389e1784),
	.w8(32'h3b76707b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b451ab4),
	.w1(32'h3af40764),
	.w2(32'h3aa2c17f),
	.w3(32'h3b52a305),
	.w4(32'h3b1dc24f),
	.w5(32'h3a810bca),
	.w6(32'h3a9a2700),
	.w7(32'h3b333b9b),
	.w8(32'h3a852754),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4ec35),
	.w1(32'hba9d38f2),
	.w2(32'hbb66a1f5),
	.w3(32'hbb4515ab),
	.w4(32'hbb003d51),
	.w5(32'hbb3cc7ee),
	.w6(32'hbb1eaa80),
	.w7(32'hbacab1c2),
	.w8(32'hbb318d26),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de9bd),
	.w1(32'hbae7f899),
	.w2(32'h3ab8d2a5),
	.w3(32'hbae04244),
	.w4(32'hbaa53576),
	.w5(32'h3aa39c99),
	.w6(32'hbac3caae),
	.w7(32'hba412b61),
	.w8(32'hba0e7dfd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf28f37),
	.w1(32'hbadc8149),
	.w2(32'hba30d752),
	.w3(32'hbb834828),
	.w4(32'hbb01e4aa),
	.w5(32'h3b1d7ba8),
	.w6(32'hbb87211a),
	.w7(32'hbb2549ca),
	.w8(32'h3ae21f8e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba7de5),
	.w1(32'h3b9a0f40),
	.w2(32'hba92f3ab),
	.w3(32'h3b311c97),
	.w4(32'h3b97d128),
	.w5(32'hbb8bbbe9),
	.w6(32'hba18a807),
	.w7(32'h3b889671),
	.w8(32'hbba676e7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabf7f3),
	.w1(32'hba64a3a5),
	.w2(32'h3bf39376),
	.w3(32'hbbd253bb),
	.w4(32'hbbc4a5e8),
	.w5(32'h3bd43f38),
	.w6(32'hbbd242db),
	.w7(32'hbbc2b5d7),
	.w8(32'h3b9e5615),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11091c),
	.w1(32'h3be42f14),
	.w2(32'hbbf16145),
	.w3(32'h3be865de),
	.w4(32'h3b8e58f9),
	.w5(32'hbc1803db),
	.w6(32'h3b94374a),
	.w7(32'h3b02dc8c),
	.w8(32'hbc0a6557),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18c3dd),
	.w1(32'hbc12e35e),
	.w2(32'hbbbfce83),
	.w3(32'hbc376108),
	.w4(32'hbc2d5813),
	.w5(32'hbb9a81a4),
	.w6(32'hbc13fc84),
	.w7(32'hbc10d8e8),
	.w8(32'hbbce66fd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a49b),
	.w1(32'hbb3e3acb),
	.w2(32'hbbaa69d2),
	.w3(32'hba0be9dc),
	.w4(32'hba8ab264),
	.w5(32'hbb6dacfd),
	.w6(32'hbb2d7999),
	.w7(32'hbb4ea4ed),
	.w8(32'hbb8c1336),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5538e3),
	.w1(32'hbbac9475),
	.w2(32'h39b038b8),
	.w3(32'hbbae8e61),
	.w4(32'hbb8c6f47),
	.w5(32'h3aec672b),
	.w6(32'hbba6489c),
	.w7(32'hbbac6f2f),
	.w8(32'h3b5a7680),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0c11b),
	.w1(32'h3abe300e),
	.w2(32'h3a132bf3),
	.w3(32'h3a4e768a),
	.w4(32'hb94ee0ac),
	.w5(32'h38b92969),
	.w6(32'h3a873ba6),
	.w7(32'hb975e628),
	.w8(32'h3a256047),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed9aa1),
	.w1(32'h385e0e8c),
	.w2(32'h3a48ed4e),
	.w3(32'h3abf5180),
	.w4(32'h3b30476c),
	.w5(32'hba0eb9bc),
	.w6(32'h3a2b5851),
	.w7(32'h3aa5e3e1),
	.w8(32'hba5f1900),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6e5eb),
	.w1(32'h3a49480a),
	.w2(32'h3b9b173d),
	.w3(32'h3b2f3b81),
	.w4(32'h38400f2b),
	.w5(32'h3b87e47c),
	.w6(32'hba07c435),
	.w7(32'hbad2ab44),
	.w8(32'h3b755b0a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58db4c),
	.w1(32'h3c1258b0),
	.w2(32'hbb59b6bc),
	.w3(32'h3b3338ca),
	.w4(32'h3bf5acdd),
	.w5(32'hbb45ef9e),
	.w6(32'h3b8dd896),
	.w7(32'h3b9c4453),
	.w8(32'hbb376e0d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd02f),
	.w1(32'hbb8112af),
	.w2(32'h3a6c9ba7),
	.w3(32'hbbc3d915),
	.w4(32'hbb912585),
	.w5(32'h386178d6),
	.w6(32'hbb7fe31c),
	.w7(32'hbb0b588b),
	.w8(32'hb9d96b5d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad977a4),
	.w1(32'hba80b5f8),
	.w2(32'hbb306514),
	.w3(32'h39c187da),
	.w4(32'h3ae29dcc),
	.w5(32'h3ae18bb4),
	.w6(32'h3ac1ac83),
	.w7(32'hbad54750),
	.w8(32'hba11a17b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeb020),
	.w1(32'hbb1693a2),
	.w2(32'h3a004a7a),
	.w3(32'hb9e3d9d7),
	.w4(32'h3a093975),
	.w5(32'hb9d9732e),
	.w6(32'h392e7968),
	.w7(32'hb7b1ea18),
	.w8(32'h380badd6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace9846),
	.w1(32'hb79d88a2),
	.w2(32'h3aba2101),
	.w3(32'hbb78b0a8),
	.w4(32'h391b074a),
	.w5(32'hba74e07c),
	.w6(32'hbb5bc574),
	.w7(32'hba2b4091),
	.w8(32'hbad7e469),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9331d19),
	.w1(32'h3ae9e01a),
	.w2(32'h3b0fee51),
	.w3(32'hbb31cec9),
	.w4(32'h3a68c532),
	.w5(32'h393ef0a3),
	.w6(32'hbae7d4d2),
	.w7(32'h39f55a4e),
	.w8(32'h3a360882),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47f3be),
	.w1(32'h3ada465c),
	.w2(32'h3a0289e6),
	.w3(32'h3a8cdb7f),
	.w4(32'hb8b2aa92),
	.w5(32'hbaa7f6ee),
	.w6(32'hba4b3b96),
	.w7(32'h3a46e2e8),
	.w8(32'hbae2192f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962df80),
	.w1(32'hbab318ea),
	.w2(32'h3a0f452c),
	.w3(32'hbb01ea77),
	.w4(32'hbb4c8599),
	.w5(32'hba06ed5c),
	.w6(32'hba3cf1c7),
	.w7(32'hbb0a29d4),
	.w8(32'hbacf8ae4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ca330),
	.w1(32'hb91ae62d),
	.w2(32'hbadce11e),
	.w3(32'hba236aee),
	.w4(32'hba933445),
	.w5(32'hba82abce),
	.w6(32'hb9025608),
	.w7(32'hba96ae14),
	.w8(32'h39982b12),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18ea49),
	.w1(32'hba804d88),
	.w2(32'hbb2d23d1),
	.w3(32'hbae36400),
	.w4(32'hba2e072c),
	.w5(32'hbb168db5),
	.w6(32'h3b2af739),
	.w7(32'h3b19ec43),
	.w8(32'hbb08955f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162185),
	.w1(32'hbb51fd30),
	.w2(32'h3ba9ccf1),
	.w3(32'hbaa253b8),
	.w4(32'hbbcf127f),
	.w5(32'h3af2f70d),
	.w6(32'hba0b1eea),
	.w7(32'hbb9590b0),
	.w8(32'h3b837e70),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f271e),
	.w1(32'h3b5055b5),
	.w2(32'h3b1f4f40),
	.w3(32'h3b5ec2fe),
	.w4(32'h3b686979),
	.w5(32'h3a9f7d7e),
	.w6(32'h3bab8f72),
	.w7(32'h3ba660ab),
	.w8(32'hb90cd20c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb026ac0),
	.w1(32'hbb26e923),
	.w2(32'h3a0b56ba),
	.w3(32'hbae0acd6),
	.w4(32'h3a6d4a50),
	.w5(32'h3b0d967c),
	.w6(32'hba1cc4fc),
	.w7(32'hb9372ee1),
	.w8(32'h3ba23424),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11fef0),
	.w1(32'h3a6ae190),
	.w2(32'h3b3716a7),
	.w3(32'h3b283a63),
	.w4(32'h3af2b335),
	.w5(32'h38f45afd),
	.w6(32'h3b2ccc28),
	.w7(32'h3b0e854f),
	.w8(32'h3b62bd4c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8f076),
	.w1(32'h3b70c225),
	.w2(32'h39b38973),
	.w3(32'h3ada4569),
	.w4(32'h3b090e04),
	.w5(32'h3b94e493),
	.w6(32'hba2da60b),
	.w7(32'h3b4dd59f),
	.w8(32'h3b857139),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334b4d),
	.w1(32'h3a6d80ca),
	.w2(32'h3aec9138),
	.w3(32'h3b6b044c),
	.w4(32'h3bd4e4e6),
	.w5(32'h38d5c09b),
	.w6(32'h3bf6fa5d),
	.w7(32'h3b89a8b5),
	.w8(32'h3b3ea2b0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89510),
	.w1(32'h3b662dbe),
	.w2(32'hbb0bb179),
	.w3(32'h3aaaa807),
	.w4(32'hbb55dadd),
	.w5(32'hbb35b229),
	.w6(32'h3ba4a613),
	.w7(32'h3a416bf1),
	.w8(32'hbaf1f75a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33c5da),
	.w1(32'hbb2d8595),
	.w2(32'h3a9afe97),
	.w3(32'hbb7ed5c5),
	.w4(32'hbb4b3359),
	.w5(32'h3b548692),
	.w6(32'hbac6158b),
	.w7(32'hba96c3d8),
	.w8(32'h3b94517c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d41ad8),
	.w1(32'h3b70df76),
	.w2(32'h3a8e8883),
	.w3(32'h3b7d95b1),
	.w4(32'h3b9b9c4e),
	.w5(32'hb76b5618),
	.w6(32'h3b47bf6d),
	.w7(32'h3b684680),
	.w8(32'h3afe9041),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6284c),
	.w1(32'h3aed57a3),
	.w2(32'h3affdb84),
	.w3(32'hb95835ce),
	.w4(32'h3ab4f5e3),
	.w5(32'h3ba301a4),
	.w6(32'h3b69d5e2),
	.w7(32'h3b9107d0),
	.w8(32'h3ba322c4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c94e),
	.w1(32'h3b65397f),
	.w2(32'hbab516d7),
	.w3(32'h3b8ab192),
	.w4(32'h3bd873ce),
	.w5(32'hba8627d1),
	.w6(32'h3b57a84a),
	.w7(32'h3b8eafe8),
	.w8(32'h3a1bc98a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d2a0e),
	.w1(32'h3a4b2049),
	.w2(32'hbb89e869),
	.w3(32'hbb3a84ed),
	.w4(32'h39a56fcd),
	.w5(32'hbbbb1f4c),
	.w6(32'h3ad88609),
	.w7(32'h3a23390a),
	.w8(32'hbb752dbe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15bc69),
	.w1(32'hbb620e71),
	.w2(32'hbaa80420),
	.w3(32'hbbc6cb10),
	.w4(32'hbb7d9523),
	.w5(32'hbb0b1979),
	.w6(32'hbbab4355),
	.w7(32'hbb8eb4e7),
	.w8(32'hbb0fb803),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dfa6c),
	.w1(32'hbb61b688),
	.w2(32'hbaee204d),
	.w3(32'hbb8029e1),
	.w4(32'hbba07e44),
	.w5(32'hbb88cd8a),
	.w6(32'hbb85f832),
	.w7(32'hbb9a9788),
	.w8(32'hbadf9516),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb251af),
	.w1(32'hbb7535f6),
	.w2(32'hba5f4349),
	.w3(32'hbc0dcaa1),
	.w4(32'hbbc55196),
	.w5(32'hbb437021),
	.w6(32'hbbb86b58),
	.w7(32'hbb47334b),
	.w8(32'h395fc494),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b41ea),
	.w1(32'hbb101924),
	.w2(32'h3a420148),
	.w3(32'hbb0f3a0d),
	.w4(32'hbb8f6a13),
	.w5(32'hb9766ee8),
	.w6(32'hbac96a7c),
	.w7(32'hbb96d677),
	.w8(32'h39842861),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1f98),
	.w1(32'hb85c2636),
	.w2(32'h3b06c46d),
	.w3(32'h39f39482),
	.w4(32'h38937538),
	.w5(32'h3b048643),
	.w6(32'h3ab68f89),
	.w7(32'h3a92f16a),
	.w8(32'h3a1ce558),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e22e2),
	.w1(32'h3a9c577f),
	.w2(32'hba30f31b),
	.w3(32'h3a878da2),
	.w4(32'hbaf86d1c),
	.w5(32'hbafd22a2),
	.w6(32'hbaeba242),
	.w7(32'h3ab1c2f8),
	.w8(32'hba980237),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba9d9f),
	.w1(32'hb887cae8),
	.w2(32'hbb45ac42),
	.w3(32'hbb424ab9),
	.w4(32'hba1d9496),
	.w5(32'hbb4b879c),
	.w6(32'hbb176794),
	.w7(32'hba6932b3),
	.w8(32'hbb00e384),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe158),
	.w1(32'hb99fa375),
	.w2(32'h3a08309b),
	.w3(32'hbbd1fa34),
	.w4(32'hbb20ea40),
	.w5(32'hba276e3e),
	.w6(32'hbbbb103f),
	.w7(32'hbb174818),
	.w8(32'h3b6c9e2a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcf6ab),
	.w1(32'h3abccd81),
	.w2(32'h3adcf697),
	.w3(32'hba7124d1),
	.w4(32'hb9ec5125),
	.w5(32'h3a64aa30),
	.w6(32'hb94dacfa),
	.w7(32'hba402887),
	.w8(32'h3b89ded8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b832877),
	.w1(32'h3b816900),
	.w2(32'h3b3fec3f),
	.w3(32'h3afc75ff),
	.w4(32'h3a373f6b),
	.w5(32'h3a2f951d),
	.w6(32'h3b9948c0),
	.w7(32'h3b8e782d),
	.w8(32'h3aeb0e1f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdbe7e),
	.w1(32'h3bdb043b),
	.w2(32'hbaffaedc),
	.w3(32'h3bc970fc),
	.w4(32'h3b36b774),
	.w5(32'hbae55ac3),
	.w6(32'h3b6f49aa),
	.w7(32'h3b46bf0d),
	.w8(32'hbb68cf3f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7872),
	.w1(32'hbb41a382),
	.w2(32'h39dc4fe0),
	.w3(32'hbb9355c0),
	.w4(32'hbb253d0a),
	.w5(32'h3aadb398),
	.w6(32'hbadcd169),
	.w7(32'hbad2d35e),
	.w8(32'h3a0616cd),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965b3be),
	.w1(32'hb8b3867d),
	.w2(32'h3b4043e5),
	.w3(32'hb9bb9f8a),
	.w4(32'h3a337366),
	.w5(32'h38a4d688),
	.w6(32'hbb130b35),
	.w7(32'hbab2996f),
	.w8(32'h3a5835c3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0921bf),
	.w1(32'hbade1e82),
	.w2(32'hbaf73a09),
	.w3(32'hbb954b13),
	.w4(32'hbbb8f867),
	.w5(32'hba67671d),
	.w6(32'hbb841155),
	.w7(32'hbb3925ad),
	.w8(32'hbb53f0e2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390805),
	.w1(32'h3a3f08ca),
	.w2(32'h3b0f0759),
	.w3(32'h3be83654),
	.w4(32'h3b996703),
	.w5(32'hb917cdff),
	.w6(32'h3b3b353c),
	.w7(32'h388d37ae),
	.w8(32'h3b664ae2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944582),
	.w1(32'h3b8dba5a),
	.w2(32'hba553e95),
	.w3(32'h3a818fc8),
	.w4(32'h3b420a02),
	.w5(32'h378eed02),
	.w6(32'h3bcaf02c),
	.w7(32'h3becc802),
	.w8(32'hbabaec5d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a322518),
	.w1(32'h3b19060d),
	.w2(32'h3ba867ee),
	.w3(32'h361f3c66),
	.w4(32'h3a0b36a1),
	.w5(32'h3b83b143),
	.w6(32'h3b01b6dc),
	.w7(32'h3a20ee2b),
	.w8(32'h3ba4ba9b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e3fc),
	.w1(32'h3bd0c004),
	.w2(32'h3a9d6f0f),
	.w3(32'h3b536042),
	.w4(32'h3b3af814),
	.w5(32'hba494b40),
	.w6(32'h3b6ecd58),
	.w7(32'h3b85d68f),
	.w8(32'h3af32118),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7ae07),
	.w1(32'hb96b36b0),
	.w2(32'h39757f08),
	.w3(32'hbbb4522b),
	.w4(32'hbb46106f),
	.w5(32'hba6581f9),
	.w6(32'hbaf567b5),
	.w7(32'h3a82e188),
	.w8(32'hb9e3572b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64aacd),
	.w1(32'hbb5da3d5),
	.w2(32'hbbab0620),
	.w3(32'hbb278cfa),
	.w4(32'hbb60d2e5),
	.w5(32'hbb97691c),
	.w6(32'hb9959038),
	.w7(32'h3a9ac6a6),
	.w8(32'hbb93cf25),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3b8e),
	.w1(32'hbb035d1c),
	.w2(32'h3be550b7),
	.w3(32'hba3625ad),
	.w4(32'hb9d6909a),
	.w5(32'h3b5d92f0),
	.w6(32'hba96aa78),
	.w7(32'hba87c463),
	.w8(32'h3c213857),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0666d4),
	.w1(32'h3bbc4a7a),
	.w2(32'h3b87215f),
	.w3(32'h3b992893),
	.w4(32'h3bcf919c),
	.w5(32'hb9ef0e40),
	.w6(32'h3bf3f0c6),
	.w7(32'h3c1e32a3),
	.w8(32'h39ecb0ee),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054100),
	.w1(32'h3b64b7ff),
	.w2(32'h3a9ae1af),
	.w3(32'h3aa4c349),
	.w4(32'h3b0c3021),
	.w5(32'h3a214090),
	.w6(32'hba11bcc5),
	.w7(32'h396a3a82),
	.w8(32'h3a7a75d5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f1393),
	.w1(32'h3ac8d305),
	.w2(32'hb9777fa2),
	.w3(32'h39b2275a),
	.w4(32'h3a6a2443),
	.w5(32'hba6cba3c),
	.w6(32'h3ac4ec47),
	.w7(32'h3b1f9c03),
	.w8(32'h39aa14ea),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab49c03),
	.w1(32'hb98b72e5),
	.w2(32'h3b110f13),
	.w3(32'hbb43786a),
	.w4(32'hba98b8e9),
	.w5(32'h3b0f6e63),
	.w6(32'hba8856af),
	.w7(32'h3a44100a),
	.w8(32'h3b1ec50f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa02e90),
	.w1(32'h3afda90e),
	.w2(32'h3bcc2954),
	.w3(32'h3a8c93a1),
	.w4(32'h3b367277),
	.w5(32'h3bcccf8c),
	.w6(32'h3b1d7e80),
	.w7(32'h3b932575),
	.w8(32'h3be61d9c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18cab4),
	.w1(32'h3ba74a96),
	.w2(32'h3af52443),
	.w3(32'h3b2f8e18),
	.w4(32'h3ba6f880),
	.w5(32'hbb0b72fc),
	.w6(32'h3b7f5990),
	.w7(32'h3b991cd4),
	.w8(32'hbaf4996c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18c53b),
	.w1(32'h3a5aac5c),
	.w2(32'hba4e92ea),
	.w3(32'hba2966c8),
	.w4(32'hba9b43ca),
	.w5(32'hbab675f5),
	.w6(32'hbadff823),
	.w7(32'hbb4a25ad),
	.w8(32'hba21f06a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f64ed),
	.w1(32'h3a2104e7),
	.w2(32'h3aaac6da),
	.w3(32'hbb1611b7),
	.w4(32'h398bafde),
	.w5(32'hb8d5841f),
	.w6(32'hba67165b),
	.w7(32'h3b159143),
	.w8(32'hba9df85a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1686b9),
	.w1(32'hbb1560a9),
	.w2(32'h3a4eb296),
	.w3(32'h3b51ef29),
	.w4(32'h3a13e664),
	.w5(32'hb8844c20),
	.w6(32'h3af0a121),
	.w7(32'hbb3993be),
	.w8(32'h3adf28fb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ffa04),
	.w1(32'hba7aad90),
	.w2(32'hbb85113a),
	.w3(32'h39b575c3),
	.w4(32'h3a984d29),
	.w5(32'hbbf5d932),
	.w6(32'hba3ef361),
	.w7(32'h3a6ed6c2),
	.w8(32'hbb87ea20),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc044f29),
	.w1(32'hbbd97000),
	.w2(32'h3be7065c),
	.w3(32'hbc5d2a69),
	.w4(32'hbc39f531),
	.w5(32'h3bae87d1),
	.w6(32'hbc1ef822),
	.w7(32'hbc02e79c),
	.w8(32'h3c071393),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dc5a9),
	.w1(32'h3b8bec6d),
	.w2(32'hba81615b),
	.w3(32'hbb423767),
	.w4(32'h3ae6fc99),
	.w5(32'hba48f5af),
	.w6(32'h3b2de41d),
	.w7(32'h3b6bf3ba),
	.w8(32'hbb1558bb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3554e2),
	.w1(32'h374e4928),
	.w2(32'h3a333f3c),
	.w3(32'h3b672625),
	.w4(32'hbabd3571),
	.w5(32'h3ab577cf),
	.w6(32'hbb606b7d),
	.w7(32'hbb56437a),
	.w8(32'hb93c42df),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa62a),
	.w1(32'hb7a8addd),
	.w2(32'hba497cba),
	.w3(32'hbb458dd5),
	.w4(32'hbb86e10b),
	.w5(32'hbb02840b),
	.w6(32'hbb03f4de),
	.w7(32'hba935d87),
	.w8(32'hba148014),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd13e6),
	.w1(32'hba827fb3),
	.w2(32'hbc40daf6),
	.w3(32'hbb41ba10),
	.w4(32'hbb26eacf),
	.w5(32'hbc1c5ce3),
	.w6(32'hbaa46ff9),
	.w7(32'hbad25fe9),
	.w8(32'hbb84ec0b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515e87),
	.w1(32'h3bc0d904),
	.w2(32'h3b7fa8fe),
	.w3(32'h3bcdaece),
	.w4(32'h3c3a11c6),
	.w5(32'hbbbb324c),
	.w6(32'h3ba85282),
	.w7(32'hbb54b8b3),
	.w8(32'h3bc40515),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82a7a5),
	.w1(32'hbb4f9ea4),
	.w2(32'hbc0d9c3e),
	.w3(32'hbc54a3bd),
	.w4(32'hbb6abc32),
	.w5(32'hbc04db69),
	.w6(32'hbc373572),
	.w7(32'hbbf040e1),
	.w8(32'hbbc8ef86),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4aa5),
	.w1(32'hbbf082ea),
	.w2(32'h3bf0f34c),
	.w3(32'hbbaa5a56),
	.w4(32'hbbe4eb3d),
	.w5(32'h3c0c45e8),
	.w6(32'hbb4427ad),
	.w7(32'hbb1bd2a6),
	.w8(32'h3bc325ac),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af053f0),
	.w1(32'hbb9b3c06),
	.w2(32'h3b906fe0),
	.w3(32'h3a68e935),
	.w4(32'hbbef86dc),
	.w5(32'h3af2e26d),
	.w6(32'h3c060163),
	.w7(32'hba21b348),
	.w8(32'hba6a7119),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fbd97),
	.w1(32'hbb2c15bc),
	.w2(32'hbbd8cbb8),
	.w3(32'h3bd01e53),
	.w4(32'hbb47821a),
	.w5(32'hbb56ec75),
	.w6(32'hbb8b24bf),
	.w7(32'h3ba70541),
	.w8(32'hba85966d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a921),
	.w1(32'h39540e31),
	.w2(32'hbc5bd6e4),
	.w3(32'hba845141),
	.w4(32'h3aeb9bcc),
	.w5(32'hbc0697fc),
	.w6(32'h3af4c13b),
	.w7(32'h3bb728ee),
	.w8(32'hbbc81ab1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8def2b),
	.w1(32'hb9beda46),
	.w2(32'hb9a307a5),
	.w3(32'h3c317b2d),
	.w4(32'h3cdf200c),
	.w5(32'hba3328ac),
	.w6(32'h3c304f8c),
	.w7(32'h3cd967b9),
	.w8(32'hbab0e74e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84d191),
	.w1(32'h3aa94329),
	.w2(32'hbbbb6829),
	.w3(32'hbb049d6a),
	.w4(32'h3b492fd1),
	.w5(32'h3a1f1eb5),
	.w6(32'hbb84d2fe),
	.w7(32'hba3ae657),
	.w8(32'hbb48e5aa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda8293),
	.w1(32'h3c0ebe07),
	.w2(32'hbc03d0e7),
	.w3(32'h3c1ef8fa),
	.w4(32'hbb26c68b),
	.w5(32'hbbfdd338),
	.w6(32'hba141c2e),
	.w7(32'hbc875a60),
	.w8(32'hbbbb1818),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb654d6c),
	.w1(32'hbbd2c580),
	.w2(32'hbb6d8e79),
	.w3(32'h388bb1bf),
	.w4(32'hbb91f9d0),
	.w5(32'hbb9f8467),
	.w6(32'h3ae8f6ea),
	.w7(32'hbad4e935),
	.w8(32'h3bb4433c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf99e35),
	.w1(32'h3954a98e),
	.w2(32'hbb533fa3),
	.w3(32'hbbcbaf9e),
	.w4(32'hbac93693),
	.w5(32'h3bb637f0),
	.w6(32'hbc1ab67c),
	.w7(32'hbbb21f3e),
	.w8(32'h3b147d74),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43d6ce),
	.w1(32'h3b6e9f16),
	.w2(32'hbb334346),
	.w3(32'h3b02c4c2),
	.w4(32'h3b8a8a66),
	.w5(32'hbb65cb4f),
	.w6(32'hb8cb99fa),
	.w7(32'hbb234aa5),
	.w8(32'hbc0ac358),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce211),
	.w1(32'h3c26ce55),
	.w2(32'hbb3a9ab3),
	.w3(32'h3b8420df),
	.w4(32'h3c8ad3a3),
	.w5(32'hbbd95826),
	.w6(32'h3bd3b8eb),
	.w7(32'h3c9e343b),
	.w8(32'hbb1393fd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd77fee),
	.w1(32'hbbb21573),
	.w2(32'h3bf20751),
	.w3(32'hbbc95bd4),
	.w4(32'hbbc7c133),
	.w5(32'h3ae0a2f8),
	.w6(32'hbbbace3e),
	.w7(32'hbc4c1e3a),
	.w8(32'h3be15f6c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9304),
	.w1(32'hbad9652f),
	.w2(32'h3b7533d7),
	.w3(32'h3ba3bdf7),
	.w4(32'h3a8dea45),
	.w5(32'hb89ffc33),
	.w6(32'h39f4b5f9),
	.w7(32'h3b2c367f),
	.w8(32'h3ab1d027),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e64c6),
	.w1(32'hbaaffa15),
	.w2(32'hbae371fd),
	.w3(32'hbbbc2b59),
	.w4(32'hbb22a71c),
	.w5(32'hbbf09648),
	.w6(32'hbb87ba48),
	.w7(32'hbb3f8efb),
	.w8(32'hbc21c2f0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23a9ac),
	.w1(32'h3c2d8b1b),
	.w2(32'hbbde5b58),
	.w3(32'hb9e3debe),
	.w4(32'h3b9b0aad),
	.w5(32'hbbb2866e),
	.w6(32'hbb8ac468),
	.w7(32'h3b958f66),
	.w8(32'hba398f8e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0b715),
	.w1(32'h3bfcd7ac),
	.w2(32'h3c2a311c),
	.w3(32'hbbe36fff),
	.w4(32'h3ab1e165),
	.w5(32'hbb47fbb5),
	.w6(32'hbbb7ccd9),
	.w7(32'h3c05335a),
	.w8(32'h3b777dea),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ebc30),
	.w1(32'h3a014277),
	.w2(32'hbb29ef55),
	.w3(32'hbb568806),
	.w4(32'hbbb695b4),
	.w5(32'hbb852404),
	.w6(32'h3b8c060a),
	.w7(32'hbb177d22),
	.w8(32'h3b9d9864),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7270c),
	.w1(32'hbb59c74c),
	.w2(32'h398169d8),
	.w3(32'h3ac61292),
	.w4(32'h3b643f52),
	.w5(32'hbb6ef08a),
	.w6(32'h3ad91f7b),
	.w7(32'hba02e2af),
	.w8(32'hbb87b84e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a679),
	.w1(32'hbbc1a056),
	.w2(32'h3c0ae671),
	.w3(32'hbb9ed1cc),
	.w4(32'hbbc86694),
	.w5(32'h3c493358),
	.w6(32'hbbbda1df),
	.w7(32'hbc08fb5f),
	.w8(32'h3c3c3bf7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c29a),
	.w1(32'hbbc78eb5),
	.w2(32'h3bef4726),
	.w3(32'h3b8ac6c5),
	.w4(32'hbbff1297),
	.w5(32'h3b1a055d),
	.w6(32'hbbadb2aa),
	.w7(32'hbb089dd7),
	.w8(32'h3acde115),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c08016),
	.w1(32'hbb906348),
	.w2(32'hba6d7655),
	.w3(32'hbadd34a4),
	.w4(32'h39f0fbfd),
	.w5(32'hbac3ff17),
	.w6(32'hbb9e06a9),
	.w7(32'h3bdbf9cd),
	.w8(32'hbb058e5f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21e538),
	.w1(32'hbc10369c),
	.w2(32'h3c722406),
	.w3(32'hbc9ce1dc),
	.w4(32'hbb0ddbd8),
	.w5(32'h3bcf816d),
	.w6(32'hbbaae413),
	.w7(32'h3c139666),
	.w8(32'h3b01f668),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d37fa),
	.w1(32'h3c4416b1),
	.w2(32'h3bb9d293),
	.w3(32'h3c44f963),
	.w4(32'h3c22cc83),
	.w5(32'h3c0f25c1),
	.w6(32'hbaffb0fd),
	.w7(32'h3bba5ba9),
	.w8(32'h3b893349),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addb0bf),
	.w1(32'hbc13a4bc),
	.w2(32'hb9fff1ff),
	.w3(32'hbb94cdb3),
	.w4(32'hbbf191d5),
	.w5(32'h3a21a63f),
	.w6(32'hbbdd6d48),
	.w7(32'h39a1c92d),
	.w8(32'h393480c2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fb160),
	.w1(32'hbac95de8),
	.w2(32'hbc1c2521),
	.w3(32'hbbd0cb58),
	.w4(32'h3c5a10a4),
	.w5(32'hbbc23998),
	.w6(32'hbb4acb64),
	.w7(32'hbba0ff2c),
	.w8(32'hbb4948f9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0bf6),
	.w1(32'hb913c408),
	.w2(32'h3bab965d),
	.w3(32'hbc3ea1bb),
	.w4(32'hbc62a80c),
	.w5(32'h3b13d730),
	.w6(32'hbbd2ae86),
	.w7(32'hbb046c48),
	.w8(32'h3b6d3c92),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f4a3d),
	.w1(32'h3c64140a),
	.w2(32'h3c3c87fd),
	.w3(32'h3c866f8b),
	.w4(32'h3cf56e13),
	.w5(32'h3c31e1e9),
	.w6(32'h3c4ff868),
	.w7(32'h3c9d4709),
	.w8(32'h3c23bfb1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29ef8f),
	.w1(32'hbb5ee195),
	.w2(32'hb92c209c),
	.w3(32'hbb496b35),
	.w4(32'hbbc9914b),
	.w5(32'h3a17bc0f),
	.w6(32'hbba0b254),
	.w7(32'hbc0cde70),
	.w8(32'hbbc6837f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3b867),
	.w1(32'hba766a45),
	.w2(32'h3bbfcf6a),
	.w3(32'hba3cd7de),
	.w4(32'h3bb3d1d7),
	.w5(32'h3b079d55),
	.w6(32'hbba698fb),
	.w7(32'h3adf6475),
	.w8(32'hbb15ea95),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05553f),
	.w1(32'hba68a41a),
	.w2(32'h3c794156),
	.w3(32'hbac4b70e),
	.w4(32'h3b3e711b),
	.w5(32'h3cb97218),
	.w6(32'hbb4efde1),
	.w7(32'hbbb5da6e),
	.w8(32'h3c92485f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dfcd5),
	.w1(32'hbbc74ad7),
	.w2(32'hbb8755cb),
	.w3(32'h3cc8962f),
	.w4(32'hbc16bd38),
	.w5(32'hbb66309b),
	.w6(32'h3c9c4fb0),
	.w7(32'hbc974803),
	.w8(32'hbb91039e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89b163),
	.w1(32'hba547fb6),
	.w2(32'hbba37df6),
	.w3(32'hbd059e27),
	.w4(32'hbb668c47),
	.w5(32'h3bb67026),
	.w6(32'hbccb78a3),
	.w7(32'hbc28ae32),
	.w8(32'h3beed411),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb81fa0),
	.w1(32'h3c1cc1ec),
	.w2(32'h3beffa07),
	.w3(32'hbb5aefc3),
	.w4(32'hba4116df),
	.w5(32'h3b84a371),
	.w6(32'h3b4c0e51),
	.w7(32'h3a298708),
	.w8(32'h3aa6c94b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb864516a),
	.w1(32'hbc1e5987),
	.w2(32'h3ab3fa3b),
	.w3(32'hbbcfbfad),
	.w4(32'hbc7898a1),
	.w5(32'h3b12e55b),
	.w6(32'hbc101cc8),
	.w7(32'hbc351e43),
	.w8(32'h3bee1d05),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57c513),
	.w1(32'h3b85cfc8),
	.w2(32'h3b3f6764),
	.w3(32'h3a242fe4),
	.w4(32'h3b847979),
	.w5(32'hbaf7304c),
	.w6(32'h3bbb26cc),
	.w7(32'hbb377e02),
	.w8(32'hbbb141fb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68780a),
	.w1(32'h391ce01c),
	.w2(32'h39b19107),
	.w3(32'h3b46f01b),
	.w4(32'h3b5972fe),
	.w5(32'h3a10c6b8),
	.w6(32'hb9a64f31),
	.w7(32'h3ba46fe9),
	.w8(32'h3b607c3c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df7ad),
	.w1(32'hbb23f93a),
	.w2(32'h3ba0fdd9),
	.w3(32'hbab3ae95),
	.w4(32'hbb09640f),
	.w5(32'h3bc95d40),
	.w6(32'h3b038352),
	.w7(32'h39f67d3f),
	.w8(32'h3b84b146),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb3bd),
	.w1(32'hbb9529db),
	.w2(32'h3b8df800),
	.w3(32'h3b345d68),
	.w4(32'hbb0a5d5b),
	.w5(32'h3b998843),
	.w6(32'h3bbd2e6e),
	.w7(32'h3b553254),
	.w8(32'hbb6e26ee),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c7ab),
	.w1(32'h3b15d18d),
	.w2(32'hba288647),
	.w3(32'hb905da41),
	.w4(32'h389adeed),
	.w5(32'hb7c3896e),
	.w6(32'hbb123543),
	.w7(32'hbbdfb5f9),
	.w8(32'hbab0ee00),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21737),
	.w1(32'hbbae0f82),
	.w2(32'hbc3ab64a),
	.w3(32'hba99204d),
	.w4(32'hbbcfb79a),
	.w5(32'hbbde23d1),
	.w6(32'hbb1afcbf),
	.w7(32'hbbd2f7c2),
	.w8(32'hbc0c3cb1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53605),
	.w1(32'h39a382d1),
	.w2(32'h39874cab),
	.w3(32'h3b0895cc),
	.w4(32'hbbbc1922),
	.w5(32'h398704d6),
	.w6(32'h3b3cf8c3),
	.w7(32'hbb723e86),
	.w8(32'hb9bd8f94),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39641d14),
	.w1(32'h3bce726a),
	.w2(32'h3c45844c),
	.w3(32'hbbd817c7),
	.w4(32'h3c5664e3),
	.w5(32'h3b9cc4df),
	.w6(32'h3b62fbf3),
	.w7(32'h3c86f3df),
	.w8(32'h3c1142ce),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42b68),
	.w1(32'h3c370de0),
	.w2(32'hbc6f7d20),
	.w3(32'h3bb57dc8),
	.w4(32'h3ca1139e),
	.w5(32'hbc3ed753),
	.w6(32'h3b4735ff),
	.w7(32'h3c2f35f6),
	.w8(32'hbc76ab4c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97e005),
	.w1(32'h38a8bf6e),
	.w2(32'hbadfc1e4),
	.w3(32'hba85f838),
	.w4(32'h3b93ea84),
	.w5(32'hbb8892ec),
	.w6(32'hbc0578cc),
	.w7(32'h3b888c6c),
	.w8(32'hbafd6bb7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a68559),
	.w1(32'h37d709e0),
	.w2(32'h3a45b572),
	.w3(32'h3a569451),
	.w4(32'h3b0b370c),
	.w5(32'hba127b67),
	.w6(32'h3b56e1c8),
	.w7(32'h3b23f116),
	.w8(32'h39df66bc),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098db9),
	.w1(32'hbaed7a5e),
	.w2(32'h3b7f0486),
	.w3(32'hbc7cdc28),
	.w4(32'hba7046c8),
	.w5(32'h3aab4c55),
	.w6(32'hbc030e39),
	.w7(32'h3b77ec2a),
	.w8(32'h3bd11301),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0010a5),
	.w1(32'h3bb07b38),
	.w2(32'h3b0e7809),
	.w3(32'h3ad1298f),
	.w4(32'h3b3899d2),
	.w5(32'hba6307c7),
	.w6(32'h3b3bc60f),
	.w7(32'h3ba46250),
	.w8(32'h3ba73b84),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e5f86),
	.w1(32'h392fccfa),
	.w2(32'h3c0bba00),
	.w3(32'h3b7e58d2),
	.w4(32'h3c373736),
	.w5(32'h3bcaad09),
	.w6(32'hbbcaca8f),
	.w7(32'h3c1f4a5d),
	.w8(32'h3bd8f839),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24c30f),
	.w1(32'h3c82a5d7),
	.w2(32'h38943312),
	.w3(32'h3c9d7de3),
	.w4(32'h3caee0eb),
	.w5(32'h37688266),
	.w6(32'h3c16221a),
	.w7(32'h3c5620fb),
	.w8(32'h3a135f30),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995cf3),
	.w1(32'hb9e8fcc0),
	.w2(32'h3bde5b6b),
	.w3(32'hbab607e8),
	.w4(32'hba559a92),
	.w5(32'h3c2792a5),
	.w6(32'hbab98c0d),
	.w7(32'hbafbecab),
	.w8(32'h3c0b22c2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e8b2d),
	.w1(32'hbc1ecc68),
	.w2(32'hbb6a8552),
	.w3(32'hba6a5021),
	.w4(32'hbc760bc2),
	.w5(32'hbad45c6b),
	.w6(32'hb8cf0ff9),
	.w7(32'hbbfeae9b),
	.w8(32'h3a47bd0e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb237),
	.w1(32'hbba8fb7e),
	.w2(32'hbc62b5b3),
	.w3(32'hbaea9795),
	.w4(32'hbba9d04a),
	.w5(32'hbc33129e),
	.w6(32'h3aa019bd),
	.w7(32'hba363ef2),
	.w8(32'hbc9109ee),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba020483),
	.w1(32'h3bc3e3e1),
	.w2(32'h3c7efcb9),
	.w3(32'hbc2c9a24),
	.w4(32'h3c2ac2b4),
	.w5(32'h3c2324bc),
	.w6(32'hba7add74),
	.w7(32'h3b8ca835),
	.w8(32'h3b88fffb),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e7faa),
	.w1(32'hbca0eb29),
	.w2(32'h3c0edc33),
	.w3(32'hbc311749),
	.w4(32'hbd0ae0d1),
	.w5(32'h3ba2d1c7),
	.w6(32'hbbfe44e4),
	.w7(32'hbccb45f6),
	.w8(32'hbb814d15),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d7dd),
	.w1(32'h3bbc34be),
	.w2(32'hbc31058c),
	.w3(32'hbba09439),
	.w4(32'h3b85f450),
	.w5(32'hbc9895ca),
	.w6(32'h3b9a1855),
	.w7(32'hbb562758),
	.w8(32'hbc0d6cb1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb94b),
	.w1(32'h3d08ce34),
	.w2(32'h3b4c7e23),
	.w3(32'h3c582315),
	.w4(32'h3d48f33f),
	.w5(32'h3b1be7e0),
	.w6(32'h3cd1f6eb),
	.w7(32'h3d1f467b),
	.w8(32'h39e2d6dd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd751),
	.w1(32'h3a2c54c2),
	.w2(32'hbb17aad0),
	.w3(32'h3bd4c81a),
	.w4(32'h3b6d1bda),
	.w5(32'hbaafe0fa),
	.w6(32'h3bba0dce),
	.w7(32'h3bbfa60c),
	.w8(32'hba83c9c8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cee92),
	.w1(32'hb8b957f2),
	.w2(32'h3bf0cc7a),
	.w3(32'hbb7cdad6),
	.w4(32'h3b2fd463),
	.w5(32'h3bc76222),
	.w6(32'hba493e5d),
	.w7(32'h3b291535),
	.w8(32'h3bf10a25),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c7934),
	.w1(32'hbba1e0c8),
	.w2(32'hbbcf9d92),
	.w3(32'h3bed0f8a),
	.w4(32'h3a18c86b),
	.w5(32'hbbadf39b),
	.w6(32'h3b939d3e),
	.w7(32'h3b36088e),
	.w8(32'h3be2904c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc238091),
	.w1(32'h39e7e4af),
	.w2(32'h3bba67c4),
	.w3(32'hbbd7183b),
	.w4(32'h3acab7cf),
	.w5(32'h3abe548d),
	.w6(32'h3bdf09f9),
	.w7(32'h3bda6701),
	.w8(32'hbb8a4ea1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c674de1),
	.w1(32'hbacc0780),
	.w2(32'h3b69311d),
	.w3(32'h3b29ff96),
	.w4(32'hbb3ad6a9),
	.w5(32'h3c31919d),
	.w6(32'hbb35c7cb),
	.w7(32'h3c0cf127),
	.w8(32'h3c150ded),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30fe84),
	.w1(32'h3ae7a246),
	.w2(32'h3af027c1),
	.w3(32'h3c93c23c),
	.w4(32'h3b514501),
	.w5(32'h3a153b4f),
	.w6(32'h3c73b954),
	.w7(32'hbb4bd386),
	.w8(32'h3b246e67),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b037e88),
	.w1(32'h3be0c76d),
	.w2(32'h3b7db1b7),
	.w3(32'h3b1a0523),
	.w4(32'h3c0de9a9),
	.w5(32'h3bbb2939),
	.w6(32'h3b93564d),
	.w7(32'h3c4fb782),
	.w8(32'h3b9a5bfe),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ba3c5),
	.w1(32'h39dfed43),
	.w2(32'h3b4de68e),
	.w3(32'h3b38ec00),
	.w4(32'h3b336de4),
	.w5(32'h38fb322b),
	.w6(32'h3b19d58b),
	.w7(32'h3ab6f534),
	.w8(32'hbbb39d0e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f7f31),
	.w1(32'h3c1a3bd9),
	.w2(32'h3bf94fdc),
	.w3(32'hbb1e5a00),
	.w4(32'h3b2b86bf),
	.w5(32'h3acd487e),
	.w6(32'hbb901d6f),
	.w7(32'h3b085f9b),
	.w8(32'hbc0123b0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42240),
	.w1(32'hbbf5962f),
	.w2(32'h3bd58dba),
	.w3(32'hbc922740),
	.w4(32'hbb8f9fd1),
	.w5(32'h3bf1b30c),
	.w6(32'hbc7f9c39),
	.w7(32'h3be87aa3),
	.w8(32'h3b86d8f9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8448e6),
	.w1(32'h3b91754d),
	.w2(32'h3c1556ce),
	.w3(32'hbb57ec65),
	.w4(32'h3c019e48),
	.w5(32'h3bfa6476),
	.w6(32'h3ac0379c),
	.w7(32'h3c478dab),
	.w8(32'hba5d2502),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc884c1),
	.w1(32'hbb268e9d),
	.w2(32'h3c4611fe),
	.w3(32'hbba4eb79),
	.w4(32'h3b3739cf),
	.w5(32'h3c730e3d),
	.w6(32'h3b8dc582),
	.w7(32'hbab61217),
	.w8(32'h3c7856b8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c885),
	.w1(32'hbc3a844c),
	.w2(32'h3b9282a3),
	.w3(32'hbc2934aa),
	.w4(32'hbc2e2e85),
	.w5(32'h3be6a1af),
	.w6(32'hbad56c74),
	.w7(32'h399915b7),
	.w8(32'h3c3f00fa),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05aebf),
	.w1(32'hbc375385),
	.w2(32'h3aa5adca),
	.w3(32'hbbe6c6df),
	.w4(32'hbcbe2588),
	.w5(32'hbb57db34),
	.w6(32'h3a8cf2bb),
	.w7(32'hbc8b66bb),
	.w8(32'h3b7aa952),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44fdf6),
	.w1(32'h3b7259a1),
	.w2(32'hba89af64),
	.w3(32'h3ba1e3e5),
	.w4(32'h3c1f84a9),
	.w5(32'hbb811691),
	.w6(32'h3b599b84),
	.w7(32'h3b30f2eb),
	.w8(32'h3b214505),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad81d0d),
	.w1(32'h3b800bcf),
	.w2(32'h3b8a063a),
	.w3(32'h3a61ed78),
	.w4(32'hb9692ee3),
	.w5(32'h3b1b7311),
	.w6(32'h3c2d5a4c),
	.w7(32'h3bc7f180),
	.w8(32'h3bb8a3ad),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7677),
	.w1(32'h3af21645),
	.w2(32'h3b8bcfd8),
	.w3(32'hbaf098cb),
	.w4(32'h3a2b8a3c),
	.w5(32'h3c0c2912),
	.w6(32'hba8c7a76),
	.w7(32'hbb4deacd),
	.w8(32'h3b10446f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba73ab),
	.w1(32'hbc26cc84),
	.w2(32'h3c2100eb),
	.w3(32'hbbe36f93),
	.w4(32'hbc9255ff),
	.w5(32'h3c6e5d51),
	.w6(32'hbbd98070),
	.w7(32'hbc64bd70),
	.w8(32'h3c27bfdd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bee16),
	.w1(32'h3c63dcc7),
	.w2(32'hbb94e913),
	.w3(32'h3c922f16),
	.w4(32'h3d0580b5),
	.w5(32'hbb421fe7),
	.w6(32'h3c8e4411),
	.w7(32'h3cc4c744),
	.w8(32'hb9c861f2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb709774),
	.w1(32'hba0fdaad),
	.w2(32'h3bd2c1df),
	.w3(32'hbc229684),
	.w4(32'h3b164101),
	.w5(32'h3b915687),
	.w6(32'hbb6dcfd4),
	.w7(32'h3be2a0b8),
	.w8(32'h3b8b7d08),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b591b68),
	.w1(32'h3b5e521e),
	.w2(32'h3bd409ea),
	.w3(32'h3b4c88fd),
	.w4(32'h3c233d6b),
	.w5(32'h3c064583),
	.w6(32'h3b924ba5),
	.w7(32'h3c301a99),
	.w8(32'h3c2bcfec),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ff80),
	.w1(32'hbc821367),
	.w2(32'h3acee761),
	.w3(32'hbbba6587),
	.w4(32'hbc07de30),
	.w5(32'h3a61b69d),
	.w6(32'h3bbfa75a),
	.w7(32'hbc1046d3),
	.w8(32'h3ae5fd5d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692ae3),
	.w1(32'h3b8a205a),
	.w2(32'h3b8486b5),
	.w3(32'h3b54959f),
	.w4(32'h3b4b4b1c),
	.w5(32'h3c2ce5db),
	.w6(32'hbb9f5217),
	.w7(32'h3b2a6f57),
	.w8(32'h3b7ca9e6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e6459),
	.w1(32'hbb79a9cf),
	.w2(32'h3c146ab1),
	.w3(32'h3b8176d9),
	.w4(32'hbbb0ae81),
	.w5(32'h3bbe206d),
	.w6(32'h3b275128),
	.w7(32'hbb88c645),
	.w8(32'h3b6a65d3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27071e),
	.w1(32'h3c11ba1f),
	.w2(32'hbbecb192),
	.w3(32'h3b7d024e),
	.w4(32'h3b038a58),
	.w5(32'hbba14530),
	.w6(32'h39fd91d7),
	.w7(32'hbb5d5e2f),
	.w8(32'hbab8f80f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb19fe),
	.w1(32'h3c2b7698),
	.w2(32'hb926005d),
	.w3(32'h3c923e1f),
	.w4(32'h3c82c476),
	.w5(32'hb904e420),
	.w6(32'h3c5d18e1),
	.w7(32'h3c851c76),
	.w8(32'h3ab45381),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1552dc),
	.w1(32'hbc8f6ad1),
	.w2(32'hb9a387fe),
	.w3(32'hbc0e6192),
	.w4(32'hbca6234a),
	.w5(32'hbb4d3a16),
	.w6(32'hbbbbb54a),
	.w7(32'hbc266eb7),
	.w8(32'h3b1bb576),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a64e5),
	.w1(32'hbbef2a10),
	.w2(32'hba42a1ab),
	.w3(32'hbb16a80a),
	.w4(32'hbc47a925),
	.w5(32'h392f20bc),
	.w6(32'hbbcbbb6a),
	.w7(32'hbc0f7d30),
	.w8(32'h3b2f386b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba66290),
	.w1(32'hba014b21),
	.w2(32'hbb1cf484),
	.w3(32'h3b9a0f33),
	.w4(32'h3a462764),
	.w5(32'h3a5041e7),
	.w6(32'h3be9b20f),
	.w7(32'hbaab87f4),
	.w8(32'h3b9b757a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c61ea4),
	.w1(32'h3bf6d93d),
	.w2(32'hbc5a3035),
	.w3(32'h39a8cfc8),
	.w4(32'h3b391979),
	.w5(32'hbb12e81f),
	.w6(32'h3b5c5b72),
	.w7(32'hbbd92af7),
	.w8(32'hbb3fe0db),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee15d4),
	.w1(32'hbc1bcc77),
	.w2(32'h3abbf458),
	.w3(32'hb90278c3),
	.w4(32'h3b44f005),
	.w5(32'h3bb19a36),
	.w6(32'hb992b579),
	.w7(32'h3c0a8f93),
	.w8(32'h3b8d5f9c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a5fb9),
	.w1(32'h3ba0830a),
	.w2(32'h3b910117),
	.w3(32'h3b0ebb4f),
	.w4(32'h3b6c7598),
	.w5(32'h3c320823),
	.w6(32'h39a19cee),
	.w7(32'hbbe5c273),
	.w8(32'h3c276ef9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1662),
	.w1(32'hbb9064bc),
	.w2(32'hba4d70ab),
	.w3(32'h3b8c1329),
	.w4(32'hbaa3cfd4),
	.w5(32'h3924d6f9),
	.w6(32'h3bd44929),
	.w7(32'h3bed77fd),
	.w8(32'h3b8a2e3d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6b35e),
	.w1(32'h3c1b5ed1),
	.w2(32'h3b1110e2),
	.w3(32'hb84151b8),
	.w4(32'h3bcb0417),
	.w5(32'h3b60a3a2),
	.w6(32'h3ba66430),
	.w7(32'h3bc5c0bb),
	.w8(32'h3b218606),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ee0e4),
	.w1(32'h3b8c030d),
	.w2(32'hbba9b761),
	.w3(32'hb9841c19),
	.w4(32'h3ba8e78e),
	.w5(32'hbbeb6846),
	.w6(32'h3b61baad),
	.w7(32'h3c5a1a0b),
	.w8(32'hbbad70a9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb611325),
	.w1(32'hbbba7952),
	.w2(32'hbb9b6470),
	.w3(32'hbb5b7b10),
	.w4(32'hbba4872f),
	.w5(32'hbbae39aa),
	.w6(32'hbb6296fb),
	.w7(32'hbb93a3b9),
	.w8(32'hbbcad6f5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe77886),
	.w1(32'hba4df2f8),
	.w2(32'h3c228c62),
	.w3(32'hbc067f9d),
	.w4(32'hb9e65b32),
	.w5(32'h3c7c368f),
	.w6(32'hbbf9b3fc),
	.w7(32'h3b073bbe),
	.w8(32'h3cac026f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26915a),
	.w1(32'hbc27c6f6),
	.w2(32'hba6beef9),
	.w3(32'hbae00ec4),
	.w4(32'hbc8aea63),
	.w5(32'h3b2f0f8b),
	.w6(32'hbbca1267),
	.w7(32'hbc767907),
	.w8(32'h3b9dae45),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a2e7a),
	.w1(32'h3bed7993),
	.w2(32'h3c3129d7),
	.w3(32'h3bef2cb9),
	.w4(32'h3c0210b9),
	.w5(32'hba0b714a),
	.w6(32'h3bba2f2b),
	.w7(32'h3a33d138),
	.w8(32'hbab44746),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9918aa),
	.w1(32'hbcc72f43),
	.w2(32'h3bbcecc8),
	.w3(32'hbcfe1f13),
	.w4(32'hbcc1c470),
	.w5(32'h3c07ea08),
	.w6(32'hbc57a2fd),
	.w7(32'hbc2c92ed),
	.w8(32'h3c591c8d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab3d4),
	.w1(32'hbb8b67de),
	.w2(32'h3bb37194),
	.w3(32'hbc38cfe8),
	.w4(32'hbb8fc904),
	.w5(32'h3b71b996),
	.w6(32'hbc434a6e),
	.w7(32'hb9e44bfe),
	.w8(32'h3b35e693),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9260d5),
	.w1(32'h3c88b3bd),
	.w2(32'hbb888d9e),
	.w3(32'h3c1fe5c1),
	.w4(32'h3d1dec5c),
	.w5(32'hbc23d827),
	.w6(32'h3c5b7f50),
	.w7(32'h3ce5978e),
	.w8(32'h3a986708),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule