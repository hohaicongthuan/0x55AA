module layer_8_featuremap_117(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf05de),
	.w1(32'h38576fb1),
	.w2(32'hb859e024),
	.w3(32'hb6c3f5e4),
	.w4(32'hb839944b),
	.w5(32'hb8b5d0bb),
	.w6(32'h38314100),
	.w7(32'hb806bedc),
	.w8(32'hb7d64674),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399147e4),
	.w1(32'h3999e222),
	.w2(32'h3996ef4b),
	.w3(32'h39ca0f18),
	.w4(32'h39a9414c),
	.w5(32'h395f00bb),
	.w6(32'h39ba4b25),
	.w7(32'h39ada858),
	.w8(32'h391b2a0c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399445e7),
	.w1(32'h3997143c),
	.w2(32'h39bb6e6d),
	.w3(32'h39d3a45c),
	.w4(32'h39bd9736),
	.w5(32'h39d7da63),
	.w6(32'h39e79076),
	.w7(32'h39f4cbdc),
	.w8(32'h39d5a5f9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78af593),
	.w1(32'h36297cc4),
	.w2(32'hb71543fb),
	.w3(32'hb81c86dd),
	.w4(32'hb76bdb4e),
	.w5(32'hb83ce73c),
	.w6(32'hb82032e8),
	.w7(32'hb7d8911f),
	.w8(32'hb83e9a0a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d6bd3),
	.w1(32'h38e6313f),
	.w2(32'h38aa0167),
	.w3(32'h390f2621),
	.w4(32'h38d4b21e),
	.w5(32'h37742d23),
	.w6(32'h395c113f),
	.w7(32'h393e38d1),
	.w8(32'h375e053c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383e019d),
	.w1(32'hb908a1ed),
	.w2(32'hb895da88),
	.w3(32'h36efdf9d),
	.w4(32'hb88b477b),
	.w5(32'hb65cc973),
	.w6(32'h38b1f5e8),
	.w7(32'hb79aedcf),
	.w8(32'hb80b7d90),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3755e6ba),
	.w1(32'hb6429192),
	.w2(32'hb79e379d),
	.w3(32'h36d6e82b),
	.w4(32'hb6663953),
	.w5(32'hb4bd3724),
	.w6(32'h374afa5d),
	.w7(32'hb70b81f9),
	.w8(32'hb7ba1ff5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a34a6e),
	.w1(32'h3983c71a),
	.w2(32'h3904058a),
	.w3(32'h39c82071),
	.w4(32'h39852939),
	.w5(32'h38314e7a),
	.w6(32'h396c2fde),
	.w7(32'h392fbfa0),
	.w8(32'hb8b11ffc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfc193),
	.w1(32'h397ca606),
	.w2(32'h38639241),
	.w3(32'h39bcd93c),
	.w4(32'h397d6f91),
	.w5(32'h38889be4),
	.w6(32'h39a48d10),
	.w7(32'h39919cc7),
	.w8(32'h3865bb4f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968cb6f),
	.w1(32'h3937e2c2),
	.w2(32'h399b31d5),
	.w3(32'h3992c43d),
	.w4(32'h395b6c66),
	.w5(32'h39345a28),
	.w6(32'h399f8894),
	.w7(32'h398f07bd),
	.w8(32'h394f8eb6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809f709),
	.w1(32'hb7865969),
	.w2(32'hb8476c1b),
	.w3(32'hb72c4d5c),
	.w4(32'hb8b0b8a4),
	.w5(32'hb85f204a),
	.w6(32'hb7b55c68),
	.w7(32'hb85b40a1),
	.w8(32'hb5eaea0b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920670f),
	.w1(32'h38fb9b3c),
	.w2(32'h388eec9d),
	.w3(32'h38fb8836),
	.w4(32'h38d58b10),
	.w5(32'h38f5f2a7),
	.w6(32'h38daf451),
	.w7(32'h391c0d40),
	.w8(32'h38c86382),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a437bf),
	.w1(32'h39805678),
	.w2(32'h39daa9e9),
	.w3(32'h39c66ef6),
	.w4(32'h3b0ac1f1),
	.w5(32'h3a5dac9f),
	.w6(32'h399ae567),
	.w7(32'h3a50414c),
	.w8(32'h3a64eeba),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c7ff6),
	.w1(32'hba3dce30),
	.w2(32'h3a55263d),
	.w3(32'hb887e86e),
	.w4(32'hb9848cfd),
	.w5(32'hbae3c8cf),
	.w6(32'hb9231077),
	.w7(32'hbb262c9f),
	.w8(32'hbb7d41b5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0534e5),
	.w1(32'hba8bd2f5),
	.w2(32'hba741654),
	.w3(32'hb90b0fc3),
	.w4(32'hb987bfe4),
	.w5(32'hbaa353bd),
	.w6(32'hbb3696ce),
	.w7(32'hbb144290),
	.w8(32'hbb76a3d0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01fb33),
	.w1(32'hbaf31853),
	.w2(32'h3a14277d),
	.w3(32'hbaac5d3c),
	.w4(32'hbb0411d6),
	.w5(32'hbba2f0d0),
	.w6(32'hbb6daffc),
	.w7(32'h3a002962),
	.w8(32'h3b1ee52e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ca0a),
	.w1(32'hbb99568f),
	.w2(32'hbb5fa1de),
	.w3(32'hbb8fd0b9),
	.w4(32'hbad26c14),
	.w5(32'hba86a7a3),
	.w6(32'hbbbe2d42),
	.w7(32'hbbaeb3a2),
	.w8(32'hba962baa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75943a),
	.w1(32'hbb574124),
	.w2(32'hbb51593d),
	.w3(32'h3a1d039e),
	.w4(32'hbb6e8d40),
	.w5(32'hbb0e86e2),
	.w6(32'h3ae26575),
	.w7(32'hb9c523f5),
	.w8(32'h3b0aa54c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc8903),
	.w1(32'hbba489f1),
	.w2(32'hbb945eff),
	.w3(32'hbbc32dd5),
	.w4(32'h3adec14b),
	.w5(32'hbb1270f7),
	.w6(32'hba802c59),
	.w7(32'hbba596bc),
	.w8(32'h3b7e95d7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f7972),
	.w1(32'h3a3dba05),
	.w2(32'hbbb252cb),
	.w3(32'h38bad3ad),
	.w4(32'h3a8adfaf),
	.w5(32'hbaea1ad7),
	.w6(32'h3c041bb5),
	.w7(32'hbb1164db),
	.w8(32'hbad0247a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44befc),
	.w1(32'hbb5acd88),
	.w2(32'hbacf5733),
	.w3(32'hbb867464),
	.w4(32'hba645ea5),
	.w5(32'h3b82cb43),
	.w6(32'h3bbcad39),
	.w7(32'hbb9017e6),
	.w8(32'hbb5f6a32),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac65548),
	.w1(32'h3aac7ab2),
	.w2(32'h3c0bcc91),
	.w3(32'h3b63938c),
	.w4(32'hbafa2649),
	.w5(32'h3aacfadb),
	.w6(32'h3b6516b4),
	.w7(32'hbbde4745),
	.w8(32'hbb848cf9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba2a24),
	.w1(32'h397fba2b),
	.w2(32'h3a623606),
	.w3(32'h3a392184),
	.w4(32'h3a97c8de),
	.w5(32'hb9ad50f4),
	.w6(32'hbbc1d092),
	.w7(32'h3b7830a4),
	.w8(32'h3b2b94fc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831c4c),
	.w1(32'h3bff13ab),
	.w2(32'h3b4e6d11),
	.w3(32'h3ae6e895),
	.w4(32'h3a2d369e),
	.w5(32'h3905b758),
	.w6(32'h3ba7aa0f),
	.w7(32'h3a746ff8),
	.w8(32'h399b274e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d181ea),
	.w1(32'h3a482dc4),
	.w2(32'h3a82b674),
	.w3(32'h3a763a9f),
	.w4(32'hbab9ee1b),
	.w5(32'hbb170a96),
	.w6(32'h3a46a7a8),
	.w7(32'hba505035),
	.w8(32'hbb835dc6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b7cd0),
	.w1(32'hb9b0236d),
	.w2(32'hbb54a316),
	.w3(32'hba239d02),
	.w4(32'hbb3429b7),
	.w5(32'hbb6b5ab1),
	.w6(32'hbaf20e7c),
	.w7(32'h3b399f47),
	.w8(32'hbb16c342),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba249b5d),
	.w1(32'hba1a8f76),
	.w2(32'hb9d05c9c),
	.w3(32'hba456917),
	.w4(32'h3b09d2ee),
	.w5(32'h3b25bb65),
	.w6(32'h3bb04207),
	.w7(32'h3c11f0b3),
	.w8(32'h3b843f63),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38e14d),
	.w1(32'h388cdac8),
	.w2(32'h3af42aa3),
	.w3(32'h3b98776d),
	.w4(32'hbb8db011),
	.w5(32'hbc215d7a),
	.w6(32'h3bf2496a),
	.w7(32'h3c3e8280),
	.w8(32'h3bb87a88),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c141b),
	.w1(32'h3b3dfa0f),
	.w2(32'h396810f5),
	.w3(32'hbc19b4dd),
	.w4(32'hbb38e5ab),
	.w5(32'hbbc079eb),
	.w6(32'h3b119e4b),
	.w7(32'hbb27eb2a),
	.w8(32'hba243eed),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a80a3),
	.w1(32'h3b484bcd),
	.w2(32'h3a1d215a),
	.w3(32'h392b2666),
	.w4(32'hbbd9e993),
	.w5(32'hbbb8cb1f),
	.w6(32'h3bd6c9cf),
	.w7(32'hbc0745b9),
	.w8(32'hbc92a10b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa9768),
	.w1(32'hbbafe87b),
	.w2(32'hbabb58b7),
	.w3(32'hbac1cebf),
	.w4(32'hba71f685),
	.w5(32'hbb001970),
	.w6(32'hbc80e526),
	.w7(32'hbb93d177),
	.w8(32'hbba44deb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5790c),
	.w1(32'hbae6cbe6),
	.w2(32'h3bbf1fc6),
	.w3(32'hba9a2442),
	.w4(32'h3bec5543),
	.w5(32'h3b1212a3),
	.w6(32'hbb8c8634),
	.w7(32'hbb4d3261),
	.w8(32'hbb325b6f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898374),
	.w1(32'h3bba7578),
	.w2(32'hbc25373d),
	.w3(32'h3b03642a),
	.w4(32'hbb9a3dc2),
	.w5(32'hba66f12b),
	.w6(32'hba8c4771),
	.w7(32'hbba8f70d),
	.w8(32'hbabd8e63),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25e091),
	.w1(32'hbc48e548),
	.w2(32'hba5f33bc),
	.w3(32'hbb00c1fb),
	.w4(32'hbb14a094),
	.w5(32'hbb106fcb),
	.w6(32'hba3c3f7d),
	.w7(32'hbb2dc5b2),
	.w8(32'hbbeb576a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d4bb),
	.w1(32'hbbebd8a6),
	.w2(32'hbab6f92f),
	.w3(32'hbb86ccef),
	.w4(32'h3ad6f6b9),
	.w5(32'h3b26f6aa),
	.w6(32'hbb802260),
	.w7(32'hb93f7a2f),
	.w8(32'hb9d4fc51),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0424bf),
	.w1(32'hbaf7fe64),
	.w2(32'hbbbcb3d4),
	.w3(32'h3aa2df5a),
	.w4(32'h3ac20a8a),
	.w5(32'h3ad6b0be),
	.w6(32'h3a5887f1),
	.w7(32'h39e401c5),
	.w8(32'hba8ee1a1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280314),
	.w1(32'hbaf00ad3),
	.w2(32'hbb6d8c35),
	.w3(32'hb9a0cc51),
	.w4(32'h3c44dc0e),
	.w5(32'h3c84f305),
	.w6(32'hbbc16e6c),
	.w7(32'hba95d0e5),
	.w8(32'h3ba73f64),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3573),
	.w1(32'h3a081390),
	.w2(32'h3baaedbf),
	.w3(32'h3c54cd96),
	.w4(32'hb9c81727),
	.w5(32'hb94503ae),
	.w6(32'h3c17ee81),
	.w7(32'h3aabecb0),
	.w8(32'hbaa925fa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc2b93),
	.w1(32'h39699d78),
	.w2(32'hba8bd78e),
	.w3(32'hba024cba),
	.w4(32'h3b67f474),
	.w5(32'h3a34dc07),
	.w6(32'hbb1c81be),
	.w7(32'h3ad43bfe),
	.w8(32'h3b822716),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7c5a),
	.w1(32'hbb85c975),
	.w2(32'h3b3660db),
	.w3(32'hbb7c3709),
	.w4(32'hbb277541),
	.w5(32'hbb3f8a66),
	.w6(32'h3c1095fe),
	.w7(32'h3c205139),
	.w8(32'h3bc0d2ff),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b433a99),
	.w1(32'h3bb31139),
	.w2(32'hbae373ea),
	.w3(32'hbac1d37a),
	.w4(32'hbb3a06fa),
	.w5(32'hbbf40797),
	.w6(32'h3bca9692),
	.w7(32'h3b9dba02),
	.w8(32'h3b30b34a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b28c1),
	.w1(32'hbbd75584),
	.w2(32'hbb951fa8),
	.w3(32'hbbd5e03d),
	.w4(32'hbb5b8ce0),
	.w5(32'hbb8bffe7),
	.w6(32'hbb9af902),
	.w7(32'h3aed9ba1),
	.w8(32'h3b056eb8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b781d),
	.w1(32'h3b45e02b),
	.w2(32'hbb65d9f2),
	.w3(32'hbbdf9ee4),
	.w4(32'hb9f9ce4e),
	.w5(32'h3bb28855),
	.w6(32'h3abe89a5),
	.w7(32'hbc5cfa3a),
	.w8(32'hbc22244f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ab37),
	.w1(32'hbc2855f3),
	.w2(32'hb88ff596),
	.w3(32'hba40455c),
	.w4(32'h3a9b1c2c),
	.w5(32'h39350247),
	.w6(32'hbb8e6092),
	.w7(32'h3a03ea7d),
	.w8(32'h395db623),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5937eb),
	.w1(32'hba60e8ab),
	.w2(32'h3b9ef9bc),
	.w3(32'hb9af3161),
	.w4(32'h3a5f5c17),
	.w5(32'hbb0e12fa),
	.w6(32'hb8837c6c),
	.w7(32'h3a927289),
	.w8(32'hbaeb6024),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27b3c8),
	.w1(32'h3ab45c49),
	.w2(32'hbb240acf),
	.w3(32'h386f50fd),
	.w4(32'hba8731bb),
	.w5(32'hba48a1e0),
	.w6(32'hbb888d72),
	.w7(32'h3b22fe10),
	.w8(32'h3b9ad239),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4439dc),
	.w1(32'h3bb327ef),
	.w2(32'h3bbf5871),
	.w3(32'hbbdee712),
	.w4(32'hb9e534e1),
	.w5(32'hbb90a59b),
	.w6(32'hbae2d2a3),
	.w7(32'hbb4ff810),
	.w8(32'hbb6a808d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d15f0),
	.w1(32'h3972e235),
	.w2(32'h3b85f210),
	.w3(32'hbb405835),
	.w4(32'h3bb579ad),
	.w5(32'hbaa6d630),
	.w6(32'h3b1496b1),
	.w7(32'h3b7b6c1b),
	.w8(32'h3b0fc46c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94199aa),
	.w1(32'hbb33148f),
	.w2(32'h3b1dd056),
	.w3(32'hba357f0e),
	.w4(32'hba8ffa86),
	.w5(32'hbb8d50e2),
	.w6(32'hbb7dfeec),
	.w7(32'h3c113d37),
	.w8(32'h3bf717f9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac781c),
	.w1(32'h3bb5fdf8),
	.w2(32'h3c25c6ac),
	.w3(32'hbb903e7e),
	.w4(32'h3937b62f),
	.w5(32'hbb85ea82),
	.w6(32'h3b1bf4ac),
	.w7(32'h3bed4aaa),
	.w8(32'h3bc5df1c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c51a),
	.w1(32'h3c2df441),
	.w2(32'hbbebe08a),
	.w3(32'h39635bd3),
	.w4(32'hbbfe0d32),
	.w5(32'hbb9a7f2f),
	.w6(32'h3be761cf),
	.w7(32'h39e3ffa8),
	.w8(32'hba824c1a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea3790),
	.w1(32'hbc20fbe1),
	.w2(32'hb90b20fd),
	.w3(32'hbbd59688),
	.w4(32'hbb857a43),
	.w5(32'hba1b81c9),
	.w6(32'hbbd5625a),
	.w7(32'hbbc88e6b),
	.w8(32'hbbc0fafa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a873573),
	.w1(32'h3b118315),
	.w2(32'h3b1c992d),
	.w3(32'hbba1c91b),
	.w4(32'h3af4c295),
	.w5(32'hbab2701f),
	.w6(32'hbb4bb87b),
	.w7(32'hb95b918a),
	.w8(32'hbabfe240),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9777103),
	.w1(32'h39aca45d),
	.w2(32'h3ac7fc99),
	.w3(32'h3aa73082),
	.w4(32'h3abed04a),
	.w5(32'h398998b1),
	.w6(32'h3b930112),
	.w7(32'hb80b0ff2),
	.w8(32'hba860c71),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1cad5),
	.w1(32'hb8d84a0d),
	.w2(32'hbbb335bd),
	.w3(32'h39ccd567),
	.w4(32'h3bd77337),
	.w5(32'hbb786bc7),
	.w6(32'hba88d020),
	.w7(32'h3c18015d),
	.w8(32'h3b7c5b80),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8e18c),
	.w1(32'h3bb0ab6e),
	.w2(32'h3ba9fa28),
	.w3(32'hbb90882f),
	.w4(32'h3aaff6bd),
	.w5(32'hbada91bc),
	.w6(32'h3b57df35),
	.w7(32'h3c2c16a5),
	.w8(32'h3c36193d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb62f0),
	.w1(32'h3b92e165),
	.w2(32'h3ac18516),
	.w3(32'hbaec60ec),
	.w4(32'hbb407c56),
	.w5(32'hbb2d9a37),
	.w6(32'h3b314377),
	.w7(32'hba262b6d),
	.w8(32'hbafd7ebd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32e565),
	.w1(32'hba4f0452),
	.w2(32'hbc1ee531),
	.w3(32'hbb10b301),
	.w4(32'hbbb40a43),
	.w5(32'hbbb86688),
	.w6(32'hbaa7c3f2),
	.w7(32'h3ac14019),
	.w8(32'h3b1c6d01),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2f796),
	.w1(32'hbc269b7a),
	.w2(32'h39c5e091),
	.w3(32'hbbb11120),
	.w4(32'h3a92e6da),
	.w5(32'h371e6825),
	.w6(32'hbba46022),
	.w7(32'h3a058803),
	.w8(32'hb999c879),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7367d1),
	.w1(32'hba5a8b44),
	.w2(32'hbbe3bb08),
	.w3(32'h395f6f61),
	.w4(32'h3b412471),
	.w5(32'h3c07aa00),
	.w6(32'hba1adef3),
	.w7(32'h3c2bbabe),
	.w8(32'h3c8716cd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994e50a),
	.w1(32'hbbae5fc7),
	.w2(32'hbb789345),
	.w3(32'h3b62681b),
	.w4(32'hbb776575),
	.w5(32'hbb082838),
	.w6(32'h3c802228),
	.w7(32'hbbb962f1),
	.w8(32'hbbc403b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ac1d),
	.w1(32'hbc3722aa),
	.w2(32'hbadb320b),
	.w3(32'hbbe87288),
	.w4(32'hbad9fe14),
	.w5(32'h3a23ff35),
	.w6(32'hbbfb08c3),
	.w7(32'hbb560372),
	.w8(32'hbb25cbdc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12eb66),
	.w1(32'hba859c7e),
	.w2(32'h3bcade01),
	.w3(32'hb6879ee1),
	.w4(32'hbbb01986),
	.w5(32'hbbac79af),
	.w6(32'h3b1e1a8a),
	.w7(32'h3ac4fdd8),
	.w8(32'hbbdfee48),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a0e4d),
	.w1(32'hbb915440),
	.w2(32'h39b353db),
	.w3(32'hbb48b320),
	.w4(32'h3a42be0e),
	.w5(32'hbb61e267),
	.w6(32'hbb899f5e),
	.w7(32'h3a6db9c4),
	.w8(32'h39ef1641),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991d32f),
	.w1(32'h395a64c7),
	.w2(32'h3beda8c8),
	.w3(32'hbb639df8),
	.w4(32'h3a9ddc8b),
	.w5(32'h3ac74b4b),
	.w6(32'h3b17ecbd),
	.w7(32'hbaf199ee),
	.w8(32'hbb4aaec8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5421bb),
	.w1(32'h3c317240),
	.w2(32'hbaf2c7e0),
	.w3(32'h3ad1ece5),
	.w4(32'hbafd9331),
	.w5(32'hbb03dd2c),
	.w6(32'h3b9ed1b4),
	.w7(32'hbb43a5c6),
	.w8(32'hbb4847be),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078b66),
	.w1(32'hbb3af533),
	.w2(32'hbbb71df4),
	.w3(32'hbad64fd9),
	.w4(32'h3b4e115e),
	.w5(32'h3a17a9a4),
	.w6(32'hbb4b5822),
	.w7(32'hb893b6a8),
	.w8(32'h3b1a83c6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0eea2),
	.w1(32'hb9bbbbdc),
	.w2(32'hbc29ac9a),
	.w3(32'hbb51412d),
	.w4(32'h3c31aa89),
	.w5(32'h3c19bf04),
	.w6(32'h3bde3928),
	.w7(32'hbb27e310),
	.w8(32'hbb9d84eb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d1f6),
	.w1(32'hbbdc1b4f),
	.w2(32'hbc01d667),
	.w3(32'h3b55f00b),
	.w4(32'hbadf3826),
	.w5(32'hbbf47997),
	.w6(32'hbb59117c),
	.w7(32'h3b86e3f6),
	.w8(32'h3bd41cb4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef06ce),
	.w1(32'hba6f089c),
	.w2(32'hbba05a07),
	.w3(32'hbbf665be),
	.w4(32'hbb61e088),
	.w5(32'hbb06ef17),
	.w6(32'h3a6555b1),
	.w7(32'hbb1f2010),
	.w8(32'hbb02ffd7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42e7ea),
	.w1(32'hbbd25c1c),
	.w2(32'hbb542d39),
	.w3(32'hbb0e936b),
	.w4(32'h3a5b7f43),
	.w5(32'hba18ade7),
	.w6(32'hbb094e65),
	.w7(32'hbb8cebe4),
	.w8(32'hbc0b419d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30f10),
	.w1(32'h3ba1f6e1),
	.w2(32'h3ba40353),
	.w3(32'h3b4f6792),
	.w4(32'h3b2fb33c),
	.w5(32'h3a69af08),
	.w6(32'hbb709855),
	.w7(32'h3be600fc),
	.w8(32'h3ad05b3b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b092),
	.w1(32'hbbcb681f),
	.w2(32'h3ad1fe47),
	.w3(32'hba961009),
	.w4(32'h3bcc3fa6),
	.w5(32'h3b90870a),
	.w6(32'hbb348c6f),
	.w7(32'hbb6827fd),
	.w8(32'hbba0c024),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f545),
	.w1(32'h3b9fad11),
	.w2(32'hbc13e702),
	.w3(32'h3b9c3b10),
	.w4(32'h3bbb3a07),
	.w5(32'h3a6efd36),
	.w6(32'hba0747f2),
	.w7(32'hb7eb9958),
	.w8(32'h3bcc9360),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe644a),
	.w1(32'hbb1ac295),
	.w2(32'h3c0fb75d),
	.w3(32'h3b533f88),
	.w4(32'hbb53c3f5),
	.w5(32'hba0ebe83),
	.w6(32'h3b4d5e93),
	.w7(32'h3b82bdb4),
	.w8(32'hbb140ffd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12a788),
	.w1(32'h3b6b66b5),
	.w2(32'hb9f80715),
	.w3(32'h3ba3d592),
	.w4(32'hb95e38b2),
	.w5(32'hba4e50f7),
	.w6(32'h3a0043d9),
	.w7(32'h3a570e96),
	.w8(32'hba93a00a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab07c0b),
	.w1(32'hbb62c92e),
	.w2(32'h3b8e9548),
	.w3(32'hbb1ffe15),
	.w4(32'h3b4f9905),
	.w5(32'hba193ed1),
	.w6(32'hbb3d008b),
	.w7(32'hbb950752),
	.w8(32'h3c535731),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ce262),
	.w1(32'h3ad46e56),
	.w2(32'h3a698039),
	.w3(32'h39bfe276),
	.w4(32'h3a518900),
	.w5(32'h3828b44e),
	.w6(32'h3bf89dc7),
	.w7(32'h3b680af0),
	.w8(32'h3ac60ba2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89eac2),
	.w1(32'hbad0c860),
	.w2(32'h3b8f291c),
	.w3(32'h395cf801),
	.w4(32'h3a9922f4),
	.w5(32'h3bbe2f89),
	.w6(32'hbbd15e62),
	.w7(32'h3b3b274b),
	.w8(32'h371baa73),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b9ed6),
	.w1(32'hbae9026c),
	.w2(32'hbafd0826),
	.w3(32'h3ae4e217),
	.w4(32'h3b38f8b1),
	.w5(32'hbbb09403),
	.w6(32'hbb0bbbfe),
	.w7(32'hbc01c014),
	.w8(32'hbc41cb53),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1faa18),
	.w1(32'hbbe17f49),
	.w2(32'h3b3e1b01),
	.w3(32'hbc0771b1),
	.w4(32'hbbdf56b0),
	.w5(32'hbb947c1a),
	.w6(32'h3b70c0d7),
	.w7(32'hbb869922),
	.w8(32'h3ba6006d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9db8),
	.w1(32'h3c151ece),
	.w2(32'h39386524),
	.w3(32'h3c0d473c),
	.w4(32'hb97063d5),
	.w5(32'hbc2f5f54),
	.w6(32'hbac9c19e),
	.w7(32'hbc59d949),
	.w8(32'hbc1cf342),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bf3bb),
	.w1(32'hbc1a1a97),
	.w2(32'h3a20d630),
	.w3(32'hbb163ed6),
	.w4(32'hbbf4829f),
	.w5(32'hbafbc1a1),
	.w6(32'hbc28a43c),
	.w7(32'hbba1ceb8),
	.w8(32'hbc68bc9f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf34e01),
	.w1(32'hbbe242c9),
	.w2(32'hbca85f47),
	.w3(32'hbb384a8c),
	.w4(32'hbc76e4a5),
	.w5(32'hbb9bfdf5),
	.w6(32'hb9cd9c18),
	.w7(32'hbbd579ac),
	.w8(32'h3cb52730),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6db15),
	.w1(32'h3c7cfb89),
	.w2(32'hbca030f6),
	.w3(32'h3c5aa3ac),
	.w4(32'h3bd251c7),
	.w5(32'h3b7be82a),
	.w6(32'hbca3a332),
	.w7(32'h3c3d90b7),
	.w8(32'hbc04aae3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096338),
	.w1(32'hbbfe5f9b),
	.w2(32'hbb6f6ed6),
	.w3(32'h3c4dd336),
	.w4(32'hbaaf5df3),
	.w5(32'hbae75dbc),
	.w6(32'hbc0cf9df),
	.w7(32'hbc3a9e7c),
	.w8(32'hbcf70644),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f3a6c),
	.w1(32'h3752369f),
	.w2(32'hbbeb71a2),
	.w3(32'hbbbb1584),
	.w4(32'hba7ea3e1),
	.w5(32'h39cab4df),
	.w6(32'hbad901ea),
	.w7(32'hbc835b5f),
	.w8(32'hbb73ed8e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c138906),
	.w1(32'h3bc814ce),
	.w2(32'h3cb0e1d7),
	.w3(32'hbb8d414f),
	.w4(32'h3c6e7abc),
	.w5(32'hbaba3ec6),
	.w6(32'hbc5faf19),
	.w7(32'h3c066a47),
	.w8(32'h3b15af91),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c322320),
	.w1(32'hbba9f04e),
	.w2(32'hbb9e185a),
	.w3(32'hbae63fba),
	.w4(32'h3b13727a),
	.w5(32'h3b60a07c),
	.w6(32'hbbce064e),
	.w7(32'h3a51e230),
	.w8(32'h3bd6e5bd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ffb93),
	.w1(32'hbadfe784),
	.w2(32'hbd243e68),
	.w3(32'hbb409e90),
	.w4(32'hbc7f38f4),
	.w5(32'h3b309467),
	.w6(32'hbbf8c753),
	.w7(32'h3d528654),
	.w8(32'hbcfa9d7b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfeea38),
	.w1(32'h3d00bc03),
	.w2(32'h397084b9),
	.w3(32'h3bab3069),
	.w4(32'h3c3c5291),
	.w5(32'hbcbfd039),
	.w6(32'hbd5c9dea),
	.w7(32'h3c2254da),
	.w8(32'h3cae1382),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19256a),
	.w1(32'hbca81f32),
	.w2(32'hbc396638),
	.w3(32'h3bfaa106),
	.w4(32'hbc1ebf0c),
	.w5(32'h3b86610a),
	.w6(32'hbbe9f5d6),
	.w7(32'h3c04901c),
	.w8(32'h3cc6ef6a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e2ac6),
	.w1(32'hba2cd82b),
	.w2(32'hbb8d8a17),
	.w3(32'h3c267d72),
	.w4(32'h3a48688e),
	.w5(32'h3b7e483e),
	.w6(32'hbca163cd),
	.w7(32'hbc05e326),
	.w8(32'hbcb956f4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59cb8),
	.w1(32'h3b46616c),
	.w2(32'h3b831920),
	.w3(32'h3bf18934),
	.w4(32'h3c082517),
	.w5(32'hbc2d96d8),
	.w6(32'hbc71ae86),
	.w7(32'hbd34a1f6),
	.w8(32'h3d893fcd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4999e6),
	.w1(32'h3c37a47b),
	.w2(32'h3aa03fd6),
	.w3(32'hbbf0db97),
	.w4(32'h3a1002de),
	.w5(32'hba8ec5ca),
	.w6(32'h3b324c8d),
	.w7(32'hba07af9f),
	.w8(32'hbb5ca199),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33caa5),
	.w1(32'h39e897f5),
	.w2(32'hbb38a5f6),
	.w3(32'h3aae2001),
	.w4(32'hbc4dfc01),
	.w5(32'h3c672314),
	.w6(32'hbaf30c8b),
	.w7(32'hbd043c54),
	.w8(32'h3b5e0fab),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd024990),
	.w1(32'h3b262f40),
	.w2(32'h3be82d61),
	.w3(32'hbba8744a),
	.w4(32'h3c5c7c7c),
	.w5(32'hbc96faa8),
	.w6(32'h3b0634b9),
	.w7(32'h386c749a),
	.w8(32'h3d0d69ff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd717),
	.w1(32'h3ad14930),
	.w2(32'hbba1dcb1),
	.w3(32'h37b6dd3f),
	.w4(32'h3bb49e79),
	.w5(32'hbc3e2915),
	.w6(32'h3bec0b89),
	.w7(32'h3bad0a84),
	.w8(32'hbbead977),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd591a),
	.w1(32'h3c8f3ba1),
	.w2(32'h3b98d62c),
	.w3(32'h3be81007),
	.w4(32'h3bea95ce),
	.w5(32'h3bfe6f88),
	.w6(32'hbce1bc7a),
	.w7(32'hb9390b43),
	.w8(32'hbb17c606),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6eaa6),
	.w1(32'h3b7f553e),
	.w2(32'h3c15a85d),
	.w3(32'h3be4f9ad),
	.w4(32'hbb847bad),
	.w5(32'hbb0b5da4),
	.w6(32'h3bbb3bbd),
	.w7(32'hbc37a4ba),
	.w8(32'hbc007d25),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62a409),
	.w1(32'h3c32146d),
	.w2(32'h3b2143f0),
	.w3(32'hbc49db31),
	.w4(32'h3b81d58d),
	.w5(32'h3b309b64),
	.w6(32'h3c1f41c0),
	.w7(32'hbb4ed1dd),
	.w8(32'hbc08a290),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f650),
	.w1(32'hbc065ffb),
	.w2(32'hbb604eec),
	.w3(32'h3bbdd84c),
	.w4(32'h3bc94f16),
	.w5(32'h3bc24742),
	.w6(32'hbc88a7bb),
	.w7(32'h3ae1d850),
	.w8(32'hbb97ede6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42de5b),
	.w1(32'h3b40e2fe),
	.w2(32'hbc39a523),
	.w3(32'h3c40c2e8),
	.w4(32'hbc2c53fd),
	.w5(32'hbba49c96),
	.w6(32'hbc338e47),
	.w7(32'hbc9d8507),
	.w8(32'hbcd4eaa5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe35a),
	.w1(32'hbbf6972d),
	.w2(32'h3a7addca),
	.w3(32'hb941ee81),
	.w4(32'h3bb6096e),
	.w5(32'hbbdc7c52),
	.w6(32'hbc1b5e01),
	.w7(32'h3b0d21d3),
	.w8(32'h3b222316),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151a6b),
	.w1(32'h3b095352),
	.w2(32'h378e765c),
	.w3(32'hbc3c42d4),
	.w4(32'hbb854af2),
	.w5(32'hbc418047),
	.w6(32'h3c4838a5),
	.w7(32'hbc52a4ad),
	.w8(32'h3c172874),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0675fb),
	.w1(32'h3c420e45),
	.w2(32'hbbcaf405),
	.w3(32'hbc56209a),
	.w4(32'h3c3c2406),
	.w5(32'hbc7028d9),
	.w6(32'hbc56d01c),
	.w7(32'h3cebbaee),
	.w8(32'h3d16774e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dc41f),
	.w1(32'hbc6eb3f5),
	.w2(32'h3ca1aa32),
	.w3(32'h3c447ff3),
	.w4(32'hb979e3e9),
	.w5(32'h3cc80d95),
	.w6(32'hbcaf1193),
	.w7(32'hbd122e04),
	.w8(32'hbd276786),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a4d1),
	.w1(32'hbcc3e183),
	.w2(32'h3b6d336f),
	.w3(32'hbb9a4dd1),
	.w4(32'h3af4920f),
	.w5(32'hbb504eb3),
	.w6(32'h3d2a1fb6),
	.w7(32'hbb6301bd),
	.w8(32'h3c3e54fa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad28727),
	.w1(32'h3a1c0af9),
	.w2(32'h3ba90dbe),
	.w3(32'hb94c899f),
	.w4(32'hbb8b3ebc),
	.w5(32'hbbc5f0c4),
	.w6(32'h3b45ea24),
	.w7(32'hbc1e50e1),
	.w8(32'hbbea664d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894bc68),
	.w1(32'hbb20f5bc),
	.w2(32'h3cadd7bf),
	.w3(32'hbc28a34b),
	.w4(32'h3b92eaca),
	.w5(32'h3b6b76ec),
	.w6(32'h3b030e8a),
	.w7(32'hbd08e131),
	.w8(32'h3be27ad7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab706b1),
	.w1(32'hbc50e800),
	.w2(32'hba2773d1),
	.w3(32'hbcfd883f),
	.w4(32'h3bcd9d45),
	.w5(32'hb98f25e5),
	.w6(32'h3cbade5f),
	.w7(32'h3c989bd4),
	.w8(32'hbcbd4044),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9506b0),
	.w1(32'hbaf0071f),
	.w2(32'h3ac1917d),
	.w3(32'hbaa2fb06),
	.w4(32'h3b81b0ce),
	.w5(32'h3c0f2541),
	.w6(32'h3c644970),
	.w7(32'hb90a5a9d),
	.w8(32'h3c600615),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4032ee),
	.w1(32'hbb43d051),
	.w2(32'hbc76b036),
	.w3(32'h3b82a833),
	.w4(32'h3c964e54),
	.w5(32'hbcca42e6),
	.w6(32'hbc056f24),
	.w7(32'hbc73dbba),
	.w8(32'h3d669821),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97f065),
	.w1(32'hbc9e3a4d),
	.w2(32'hbb935dbf),
	.w3(32'hbc87f0e2),
	.w4(32'hbc82b1e6),
	.w5(32'hbcaac335),
	.w6(32'hbc8149c4),
	.w7(32'hbbd9b0d6),
	.w8(32'hbb16a727),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71b2b1),
	.w1(32'hbcd2c14f),
	.w2(32'hbc82a609),
	.w3(32'hbc787413),
	.w4(32'hbac37416),
	.w5(32'h3b63f8d8),
	.w6(32'hbc6fa5e3),
	.w7(32'h3ccb76a7),
	.w8(32'h3c24d9ab),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f31ea),
	.w1(32'h3c3bbc0a),
	.w2(32'hbc8857eb),
	.w3(32'h3aa7e578),
	.w4(32'h3c167982),
	.w5(32'h3b215305),
	.w6(32'hbcd32615),
	.w7(32'h3c66f1f7),
	.w8(32'hbbe9ebc4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bdeda),
	.w1(32'hba287701),
	.w2(32'hbb3baace),
	.w3(32'h3c589d0d),
	.w4(32'hbc0ec9c2),
	.w5(32'hbbcae902),
	.w6(32'hbb35434a),
	.w7(32'h3b0b3b55),
	.w8(32'h3be294dd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4f03b),
	.w1(32'h3b9e45fb),
	.w2(32'h3b1bf8e9),
	.w3(32'hba8ce835),
	.w4(32'h39df0b1b),
	.w5(32'hbb35a876),
	.w6(32'hbc53acb8),
	.w7(32'hba75e0a4),
	.w8(32'h3c2aeca9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c10bc),
	.w1(32'hba44d57f),
	.w2(32'hba94d714),
	.w3(32'hba8ed29a),
	.w4(32'hbc218751),
	.w5(32'hbc23585e),
	.w6(32'h3b15e569),
	.w7(32'h3b7a68af),
	.w8(32'hbba355a1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dff4b),
	.w1(32'hbc272792),
	.w2(32'hbb7c59df),
	.w3(32'hbc19e22b),
	.w4(32'hbc456812),
	.w5(32'hbbf3f52d),
	.w6(32'hbc5869f2),
	.w7(32'hbc00ae23),
	.w8(32'hbb8a291c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc013cc4),
	.w1(32'hbbbe5ac2),
	.w2(32'hbc216a9e),
	.w3(32'hbbbd1a23),
	.w4(32'hba7dab67),
	.w5(32'h3b4e8e08),
	.w6(32'hbc90311b),
	.w7(32'h3c2bce33),
	.w8(32'h3c3a5e2b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae498),
	.w1(32'h3b3e1313),
	.w2(32'h3c0ce6fe),
	.w3(32'h3ba02950),
	.w4(32'hbc83ed7c),
	.w5(32'h3c4cdf90),
	.w6(32'hbb8bd7cf),
	.w7(32'h3c3c9300),
	.w8(32'hb9a67fe4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba275a2),
	.w1(32'h39ae42cd),
	.w2(32'h3b657412),
	.w3(32'hbb85805c),
	.w4(32'h3a8c087e),
	.w5(32'hbb6f740a),
	.w6(32'h3c50e367),
	.w7(32'hbb2baafd),
	.w8(32'h3c161ac1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba997dfd),
	.w1(32'hba33dacc),
	.w2(32'hbb793aa9),
	.w3(32'h38bb19f6),
	.w4(32'hbc8cc79f),
	.w5(32'h3cfe4923),
	.w6(32'h39d78367),
	.w7(32'h3d16e8e2),
	.w8(32'hbde7822b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d12de88),
	.w1(32'hbbc7320e),
	.w2(32'h3b5e20fa),
	.w3(32'h3c02bdab),
	.w4(32'hbc07c39c),
	.w5(32'h3b8cfc6d),
	.w6(32'hbbfc314d),
	.w7(32'h3bec5648),
	.w8(32'hbc586157),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ac9bf),
	.w1(32'h3bb0840a),
	.w2(32'hb94f7ad0),
	.w3(32'h3bfeab0c),
	.w4(32'hbaa7e4a1),
	.w5(32'h3b1f8705),
	.w6(32'hbb80291f),
	.w7(32'h3b6955c8),
	.w8(32'hbae8797f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e226),
	.w1(32'hbb5616d5),
	.w2(32'h3abafeee),
	.w3(32'h3b9a0dbe),
	.w4(32'h3aa8fdf2),
	.w5(32'h3b4cc450),
	.w6(32'h3b06ad33),
	.w7(32'h3bce9816),
	.w8(32'hbc1f04e0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3d4b6),
	.w1(32'hbb538ad1),
	.w2(32'hbb4ba2a4),
	.w3(32'hbbc50e01),
	.w4(32'h3c026704),
	.w5(32'h3c294c03),
	.w6(32'hbc1a108b),
	.w7(32'hbbd2ada9),
	.w8(32'h3bd21dee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule