module layer_8_featuremap_27(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9659582),
	.w1(32'hbc30b51b),
	.w2(32'h3bbfabe2),
	.w3(32'h3c8f18da),
	.w4(32'h3b5e2407),
	.w5(32'h3b20d236),
	.w6(32'h3c1deb9a),
	.w7(32'h3bf5015b),
	.w8(32'h3bd20439),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85966e),
	.w1(32'h3b0d0be0),
	.w2(32'h3b4bad6d),
	.w3(32'h3b92fab5),
	.w4(32'h39f70571),
	.w5(32'h3b0e3b31),
	.w6(32'h3b1d372d),
	.w7(32'hbad9b7cf),
	.w8(32'h3adf2a7e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d334c),
	.w1(32'hbb3d3fc1),
	.w2(32'hb7d3a900),
	.w3(32'h3b9e3beb),
	.w4(32'hb9dfe09c),
	.w5(32'h3b4ea169),
	.w6(32'h3b91ff5a),
	.w7(32'hbb61f668),
	.w8(32'h3c195fba),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8a70d),
	.w1(32'hbc533cb7),
	.w2(32'h3c9c6b43),
	.w3(32'hbc3d0ffc),
	.w4(32'hbced056e),
	.w5(32'h3a3bf4cd),
	.w6(32'h3cc91b63),
	.w7(32'h3c8bdd37),
	.w8(32'h3c9f2164),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51dd00),
	.w1(32'h3b65223c),
	.w2(32'h3b93a5c5),
	.w3(32'h3c32f299),
	.w4(32'h3af7a911),
	.w5(32'h3afa067d),
	.w6(32'h3c756561),
	.w7(32'h3b547c4b),
	.w8(32'h3b9fd521),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1af8be),
	.w1(32'hbc5dcae2),
	.w2(32'hbcc3898f),
	.w3(32'h3d4063e5),
	.w4(32'hbc1b360c),
	.w5(32'h3a2de576),
	.w6(32'h3d2a5206),
	.w7(32'hbc2da0b3),
	.w8(32'hbbeeec8b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06fc53),
	.w1(32'hbb195e65),
	.w2(32'hb95eb60b),
	.w3(32'h3bf55d05),
	.w4(32'h3c0c4ab1),
	.w5(32'h3bd4bffc),
	.w6(32'hba396802),
	.w7(32'h3a0d4239),
	.w8(32'hbb889eed),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93a765),
	.w1(32'hbc1ce7b2),
	.w2(32'hbbad3f07),
	.w3(32'h3be612e3),
	.w4(32'hbbaebcbc),
	.w5(32'hbbeb33aa),
	.w6(32'h3c352a37),
	.w7(32'hbb4ba7f8),
	.w8(32'h3c1b1368),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16ee66),
	.w1(32'h3b6b1f4c),
	.w2(32'h3b801b72),
	.w3(32'h3c45f8ab),
	.w4(32'h3c26dcef),
	.w5(32'h3c2418a8),
	.w6(32'h3bbb1859),
	.w7(32'h3b41974e),
	.w8(32'h3c6e884c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bf95e),
	.w1(32'h3b9a3487),
	.w2(32'h3d045122),
	.w3(32'h3c8ff145),
	.w4(32'h3bdefd6c),
	.w5(32'hbb87b566),
	.w6(32'h3d3b0213),
	.w7(32'h3c619ac4),
	.w8(32'h3bad8da6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db0767),
	.w1(32'hbc2fd042),
	.w2(32'hbb272ba2),
	.w3(32'h3bbd9834),
	.w4(32'hbbfb93ea),
	.w5(32'hbb354738),
	.w6(32'h3c62b6fa),
	.w7(32'h3b1d4dfe),
	.w8(32'hbb3f5ecd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caaa2f4),
	.w1(32'h3a9a6544),
	.w2(32'h3b04941b),
	.w3(32'h3cd8fb9f),
	.w4(32'h3c17483f),
	.w5(32'h3bfb6bcd),
	.w6(32'h3cc5dbfe),
	.w7(32'h3b5e73de),
	.w8(32'h3bdb5c04),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c769481),
	.w1(32'hbb5385e3),
	.w2(32'h3b00a5e2),
	.w3(32'h3c3a8af3),
	.w4(32'hbad79a29),
	.w5(32'h398b4947),
	.w6(32'h3c8c1dfa),
	.w7(32'hbb08a24f),
	.w8(32'h3b7a1c9c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61f310),
	.w1(32'hbb8ab546),
	.w2(32'hbabdfad3),
	.w3(32'h3cb9da21),
	.w4(32'h3c807a61),
	.w5(32'h3c7d4503),
	.w6(32'h3a97f655),
	.w7(32'hbab87b2e),
	.w8(32'hba78f3a9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868fea),
	.w1(32'hbbcd6400),
	.w2(32'hbb4a79a7),
	.w3(32'h3c548393),
	.w4(32'h3c2103b0),
	.w5(32'h3bdf3a0c),
	.w6(32'hba05b4be),
	.w7(32'hb9e04ffb),
	.w8(32'h38948814),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa53a),
	.w1(32'h3b1708dc),
	.w2(32'h3b57da85),
	.w3(32'hbb2a047c),
	.w4(32'hbb1dbc29),
	.w5(32'hbb9f59ac),
	.w6(32'h3b0d7501),
	.w7(32'h3b0741fc),
	.w8(32'h3c8feccb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c463533),
	.w1(32'h3d28e989),
	.w2(32'h3c6dad65),
	.w3(32'h3c0a0b84),
	.w4(32'h3b50b6af),
	.w5(32'h3c89757f),
	.w6(32'hbba26b7d),
	.w7(32'hbb16a4d8),
	.w8(32'hbbca89a4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd18ce4),
	.w1(32'h3bd1d6f0),
	.w2(32'h3c1d5093),
	.w3(32'h3c0bed15),
	.w4(32'h3be1fca1),
	.w5(32'h3c66e32e),
	.w6(32'h3c70b5ef),
	.w7(32'h3b9434dd),
	.w8(32'h3bda56d9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c959ce7),
	.w1(32'hbd2b417c),
	.w2(32'hbcba7cd6),
	.w3(32'h3d67af3a),
	.w4(32'hbc13af09),
	.w5(32'hbcb5d6c1),
	.w6(32'h3d2b6f28),
	.w7(32'h3bb43b25),
	.w8(32'h3afa7350),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4c36d3),
	.w1(32'h3d3e0acb),
	.w2(32'h3cd0255e),
	.w3(32'h3d35f842),
	.w4(32'hbc41f16a),
	.w5(32'h3baa59af),
	.w6(32'h3d45caf3),
	.w7(32'h3bf3be52),
	.w8(32'h3cb4822e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdbc09),
	.w1(32'hbc807479),
	.w2(32'hbc3c69fe),
	.w3(32'h3a6c7d4d),
	.w4(32'hbc900d79),
	.w5(32'hbc850704),
	.w6(32'h3c61c179),
	.w7(32'hbbfb291b),
	.w8(32'hbc174ac9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22bce9),
	.w1(32'hbbc19844),
	.w2(32'h3a47be06),
	.w3(32'h3bb45212),
	.w4(32'hbadff87e),
	.w5(32'h3b484b46),
	.w6(32'h3bdd3304),
	.w7(32'hbb635926),
	.w8(32'h3c7e2c8d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2445a),
	.w1(32'hbc12a924),
	.w2(32'hbb924b16),
	.w3(32'h3b32c6d4),
	.w4(32'h3b5c3398),
	.w5(32'hbaf735d7),
	.w6(32'h3c8cb934),
	.w7(32'h3d0a2671),
	.w8(32'h3c4012ec),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04c19c),
	.w1(32'hbb09f8d7),
	.w2(32'h3bb49a8f),
	.w3(32'h3c0773f7),
	.w4(32'hbbfd2e1b),
	.w5(32'hbba5e5fa),
	.w6(32'h3bfe619f),
	.w7(32'h38da07aa),
	.w8(32'hbb0a1f65),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592ba2),
	.w1(32'hbbcdb1fa),
	.w2(32'hbb775cc6),
	.w3(32'hbc0e997c),
	.w4(32'hbb9037c7),
	.w5(32'hbb4e445e),
	.w6(32'hbb4268db),
	.w7(32'hbb32ef1c),
	.w8(32'h3c424561),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cddfcea),
	.w1(32'hba09cd1a),
	.w2(32'h3b8fac8a),
	.w3(32'h3cacbdbf),
	.w4(32'hbab1169d),
	.w5(32'hbb7755a6),
	.w6(32'h3d0f9db3),
	.w7(32'h3c9e2870),
	.w8(32'h3c309c0b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75fa8d),
	.w1(32'h3b5cdb62),
	.w2(32'h3bf34eb7),
	.w3(32'hbbb71e17),
	.w4(32'hbb2937c9),
	.w5(32'h3a551c19),
	.w6(32'h3b99a108),
	.w7(32'h3c5f3745),
	.w8(32'hb9c2e085),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6a56d4),
	.w1(32'hbdacd634),
	.w2(32'hbdad00b3),
	.w3(32'h3d6cc5de),
	.w4(32'hbd47a136),
	.w5(32'hbd6ed742),
	.w6(32'h3d8e3a64),
	.w7(32'hbcada3dc),
	.w8(32'h3ca54089),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb3fca),
	.w1(32'h3b483485),
	.w2(32'h3c45f615),
	.w3(32'h3c3e968d),
	.w4(32'hbc64ed65),
	.w5(32'hbca9ddc9),
	.w6(32'h3d1e2985),
	.w7(32'h3c70c9ea),
	.w8(32'h3b74bb2a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba11aac),
	.w1(32'hba3e7288),
	.w2(32'h3a777d23),
	.w3(32'h3bb7ed18),
	.w4(32'hb8215280),
	.w5(32'h3a8410e6),
	.w6(32'h3b6d7c7d),
	.w7(32'hbac04376),
	.w8(32'hbbc616e3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7911d),
	.w1(32'h3d04408a),
	.w2(32'h3a53d7c0),
	.w3(32'hbbcc5c97),
	.w4(32'h3c0bfce4),
	.w5(32'hbc719e78),
	.w6(32'hbc18ff6d),
	.w7(32'hbadac935),
	.w8(32'h3ba45de0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0385d),
	.w1(32'hbcc02e6d),
	.w2(32'hbbdf745e),
	.w3(32'h3b6d8790),
	.w4(32'hbc19e2a8),
	.w5(32'hbb9bacf7),
	.w6(32'h3cc05c22),
	.w7(32'h3ba97d2f),
	.w8(32'h3c336ddf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a17d3),
	.w1(32'hbc018372),
	.w2(32'hbc122669),
	.w3(32'h3c4ca067),
	.w4(32'h3d04cd02),
	.w5(32'h3c2a490c),
	.w6(32'hbb36ac3f),
	.w7(32'h3c314d4b),
	.w8(32'hbc8205c0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd69f72),
	.w1(32'h3b8640f5),
	.w2(32'hbb5a1a15),
	.w3(32'hbcb1643c),
	.w4(32'hbcc6794d),
	.w5(32'hbc824519),
	.w6(32'h3c3aa1d0),
	.w7(32'hbb8a7b7c),
	.w8(32'h3976986b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c088e),
	.w1(32'h3ad02237),
	.w2(32'h3c4c7dda),
	.w3(32'h3d07012a),
	.w4(32'h3be79f1e),
	.w5(32'h3c9a4942),
	.w6(32'h3cab2972),
	.w7(32'h3b6ce771),
	.w8(32'h3c5126dd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976a50),
	.w1(32'hbc803324),
	.w2(32'hbc3c221d),
	.w3(32'h3c23e571),
	.w4(32'hbaf9a8ba),
	.w5(32'hbc3b1cdc),
	.w6(32'h3b7c96ca),
	.w7(32'hbb843c18),
	.w8(32'hbb3dc5ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8953fc),
	.w1(32'h3c2b5681),
	.w2(32'hbc0237ba),
	.w3(32'hbbb4c692),
	.w4(32'hbb661e3c),
	.w5(32'h3b932e41),
	.w6(32'h39457324),
	.w7(32'hbbafa865),
	.w8(32'hbb59f3ca),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95c45f),
	.w1(32'hba9c22c8),
	.w2(32'h3a7cc950),
	.w3(32'h3b2849e4),
	.w4(32'h3b083db1),
	.w5(32'h3aaf2e40),
	.w6(32'h392df1f9),
	.w7(32'hbb051776),
	.w8(32'hbb99d9f8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc548981),
	.w1(32'hbc87566d),
	.w2(32'hbc27b5b8),
	.w3(32'h3cd9918a),
	.w4(32'h3cb359d0),
	.w5(32'h3c820d77),
	.w6(32'hbb8b0d87),
	.w7(32'hba41636c),
	.w8(32'hba8a7040),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3960e),
	.w1(32'hbba25719),
	.w2(32'hbb8601d4),
	.w3(32'hbbbdb3fa),
	.w4(32'hbb757f5c),
	.w5(32'hbb0ac68e),
	.w6(32'h3b83b211),
	.w7(32'h3b76e610),
	.w8(32'h3b967e1a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dada00a),
	.w1(32'hbcd4d3cd),
	.w2(32'hbcc83015),
	.w3(32'h3dba1757),
	.w4(32'hbc15f23a),
	.w5(32'hbce77582),
	.w6(32'h3df40c10),
	.w7(32'h3c9af290),
	.w8(32'hbb55cbcf),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48d9a),
	.w1(32'hbc27e3b1),
	.w2(32'hbba74233),
	.w3(32'h3b71b291),
	.w4(32'hbc217e4c),
	.w5(32'hbbfc209a),
	.w6(32'h3b39e0bb),
	.w7(32'hba9513b6),
	.w8(32'hbbc600a4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8321d),
	.w1(32'h3b38e006),
	.w2(32'h3c9a93f1),
	.w3(32'h3b644786),
	.w4(32'hba6b862e),
	.w5(32'h3ccdd01a),
	.w6(32'h3c5b13b3),
	.w7(32'h3c9a8d28),
	.w8(32'hbbcd23da),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62c450),
	.w1(32'hbc261e8a),
	.w2(32'hbb82b1a5),
	.w3(32'h3c7414ad),
	.w4(32'hbb896ed1),
	.w5(32'hbc08dafd),
	.w6(32'h3cab0677),
	.w7(32'h3a5fdcfb),
	.w8(32'hbbfd75ab),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd449f7),
	.w1(32'hbcbc2385),
	.w2(32'hbbf43bac),
	.w3(32'h3ca1e871),
	.w4(32'hbc03c806),
	.w5(32'hbb6d62d1),
	.w6(32'h3c82a609),
	.w7(32'h3b791b08),
	.w8(32'h3c8d4af9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e3f40),
	.w1(32'hbc6f4b6f),
	.w2(32'hbbe498cd),
	.w3(32'h3c21fce9),
	.w4(32'hbc9154f4),
	.w5(32'hbc58d9b2),
	.w6(32'h3b319298),
	.w7(32'hbbfec188),
	.w8(32'hbc379684),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7539e6),
	.w1(32'hbc382853),
	.w2(32'hbbc15af4),
	.w3(32'hbc20027e),
	.w4(32'h3c884bb9),
	.w5(32'hbc67e20d),
	.w6(32'hbc6d764e),
	.w7(32'hbbd31d1d),
	.w8(32'h3c7012ac),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc656b0),
	.w1(32'hbbf7e609),
	.w2(32'hbcec97ab),
	.w3(32'h3c25d295),
	.w4(32'h3bcc7f57),
	.w5(32'hbb2f7999),
	.w6(32'h3caf8f44),
	.w7(32'hbc0b0c32),
	.w8(32'h39c02e7c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86d2a0),
	.w1(32'h3a9e4e82),
	.w2(32'hbc7a1e53),
	.w3(32'h3c14610d),
	.w4(32'hbc0a1458),
	.w5(32'hbc3d3eed),
	.w6(32'h3c0aa1c3),
	.w7(32'hbc67a3fa),
	.w8(32'h3ac71c5c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c050125),
	.w1(32'hbc5910e8),
	.w2(32'h3c1e9d65),
	.w3(32'h3c3791bd),
	.w4(32'hbbe177e0),
	.w5(32'hbb8242f9),
	.w6(32'h3c485215),
	.w7(32'h3bacbe65),
	.w8(32'h3bc229d9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5a3c4),
	.w1(32'h39c36016),
	.w2(32'hbbbfbbd2),
	.w3(32'h3c438f30),
	.w4(32'hbc5100bc),
	.w5(32'hbc7342d5),
	.w6(32'h3cce506d),
	.w7(32'hba74bb1c),
	.w8(32'hbc718ade),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5db6a9),
	.w1(32'hbc9fc177),
	.w2(32'hbc26c6de),
	.w3(32'h3d8655e5),
	.w4(32'hbbbdba83),
	.w5(32'hbcaf8e6d),
	.w6(32'h3d8c7a24),
	.w7(32'h3c74a0be),
	.w8(32'h3cdd0c09),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5e48a4),
	.w1(32'hbbd8735d),
	.w2(32'h3cd79703),
	.w3(32'h3d2cc853),
	.w4(32'hb9492d25),
	.w5(32'h3d15d35e),
	.w6(32'h3c733df9),
	.w7(32'h3c2e7ff4),
	.w8(32'h3c1fba89),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63ff6b),
	.w1(32'h3b7d0fa6),
	.w2(32'h3cad5978),
	.w3(32'h3cac2e1e),
	.w4(32'hba1faf6f),
	.w5(32'h3b34e40b),
	.w6(32'h3c4738fd),
	.w7(32'h3c89539e),
	.w8(32'h3cb28474),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5032e),
	.w1(32'hbb97ec49),
	.w2(32'hbbca2a52),
	.w3(32'hbbe1c281),
	.w4(32'h3c80f305),
	.w5(32'h3c1047f4),
	.w6(32'hbc8d3799),
	.w7(32'h3c030c8e),
	.w8(32'hba3f7fb7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1216d6),
	.w1(32'h3c874814),
	.w2(32'h3c76c9b3),
	.w3(32'h3d2ae4a2),
	.w4(32'h3cfdd1fb),
	.w5(32'h3c954ac8),
	.w6(32'h3cd8c3f4),
	.w7(32'h3c6a9d8d),
	.w8(32'h3c153334),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56a0df),
	.w1(32'h3cbbb81d),
	.w2(32'hbbcbce6f),
	.w3(32'h3c769c36),
	.w4(32'h3ca8b801),
	.w5(32'hbaeafcc7),
	.w6(32'h3c0de9b9),
	.w7(32'hbb853f78),
	.w8(32'h3a962151),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d344),
	.w1(32'h3c5888d1),
	.w2(32'hbc6d2b55),
	.w3(32'h3cd19408),
	.w4(32'hbb9b7917),
	.w5(32'h3b25d3db),
	.w6(32'h3d043b9a),
	.w7(32'hbbf8e4ed),
	.w8(32'hbbebc003),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac47af),
	.w1(32'hbbac9079),
	.w2(32'hbc6a9254),
	.w3(32'h3b2457e7),
	.w4(32'hbb2b666b),
	.w5(32'hbc18be12),
	.w6(32'h3ba6ab39),
	.w7(32'hbb8a50d5),
	.w8(32'h3bbf6725),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda6463),
	.w1(32'hbc922126),
	.w2(32'h3c5131ce),
	.w3(32'h3ca3ad52),
	.w4(32'hbb3e98ab),
	.w5(32'h3c061d8d),
	.w6(32'h3cb2c5c2),
	.w7(32'h3ce07e41),
	.w8(32'hbb75de32),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c480371),
	.w1(32'h3c05ea32),
	.w2(32'hbcb8040d),
	.w3(32'hbb8e3cad),
	.w4(32'hbc8dcaa6),
	.w5(32'hbb977e99),
	.w6(32'hbb39a86e),
	.w7(32'hbcdd7831),
	.w8(32'h3c321ac3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6978f7),
	.w1(32'h3c23d2c2),
	.w2(32'h3b13a6a0),
	.w3(32'h3b7cf6b6),
	.w4(32'h3a573b7e),
	.w5(32'h3b879c34),
	.w6(32'hbbbbdf46),
	.w7(32'h3b0480ee),
	.w8(32'hbb472821),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d655520),
	.w1(32'hbc729c77),
	.w2(32'hbccc46fb),
	.w3(32'h3d74bb44),
	.w4(32'hbc89c667),
	.w5(32'hbd265018),
	.w6(32'h3d60f7da),
	.w7(32'hbbf77e8c),
	.w8(32'hbce30be2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9614ce0),
	.w1(32'hbd0b0a1b),
	.w2(32'hbbeaec33),
	.w3(32'h3a4e36d0),
	.w4(32'h3c08a02c),
	.w5(32'hbc95aab0),
	.w6(32'h3addd1bc),
	.w7(32'hbbbfb9bd),
	.w8(32'hbbad1bae),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe511),
	.w1(32'hbb8cb97d),
	.w2(32'hbbd7563f),
	.w3(32'hbb7a0aab),
	.w4(32'h39f536d8),
	.w5(32'hbbc9cb37),
	.w6(32'h3a0f99e7),
	.w7(32'hbbac2bb9),
	.w8(32'hbad096ac),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2b4d3),
	.w1(32'hbbb52231),
	.w2(32'hbb799c22),
	.w3(32'h3bd25977),
	.w4(32'hba264243),
	.w5(32'hbb6ec76f),
	.w6(32'h3c288af4),
	.w7(32'h3bac0251),
	.w8(32'h39eb5813),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbb2a6),
	.w1(32'h3b3c0a09),
	.w2(32'hbad6c88c),
	.w3(32'h3c9bef25),
	.w4(32'hbaf1fb43),
	.w5(32'hbb6990b2),
	.w6(32'h3cd9ac6f),
	.w7(32'h3b840353),
	.w8(32'h3c18930b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3d507a),
	.w1(32'h3b8eb786),
	.w2(32'hbbbf6aed),
	.w3(32'h3d20f23c),
	.w4(32'hbafa2d58),
	.w5(32'hbced80ae),
	.w6(32'h3ce91181),
	.w7(32'h3bc0cf0b),
	.w8(32'hbbc6571a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefd82f),
	.w1(32'hbbde2668),
	.w2(32'h3a9fb678),
	.w3(32'h39010841),
	.w4(32'hbb9cf0f4),
	.w5(32'hbb8eb8f9),
	.w6(32'hba53855b),
	.w7(32'h3ae63225),
	.w8(32'hbc316655),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb79be),
	.w1(32'hbd03ceb7),
	.w2(32'hbc750b0f),
	.w3(32'h3cdcd336),
	.w4(32'h399d71e5),
	.w5(32'hbc060a8b),
	.w6(32'h3d189b0d),
	.w7(32'h3bd8cd15),
	.w8(32'h3bda396d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38001792),
	.w1(32'hbaef702f),
	.w2(32'h3ab5ca1f),
	.w3(32'hba4e51ee),
	.w4(32'hbb241815),
	.w5(32'hbb1e83e3),
	.w6(32'h3af2587e),
	.w7(32'h3adb473d),
	.w8(32'h3a1276e7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7263c),
	.w1(32'hbb63912a),
	.w2(32'h3c1e0350),
	.w3(32'h3c98dfed),
	.w4(32'hbba9ff38),
	.w5(32'hb9b8d213),
	.w6(32'h3ca30be4),
	.w7(32'h3b3630f9),
	.w8(32'h3bb4f733),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b90c4),
	.w1(32'h3a85308c),
	.w2(32'h3c04f103),
	.w3(32'hbab3a72f),
	.w4(32'h3a72c0d9),
	.w5(32'h3af4df3f),
	.w6(32'h3bdeb7ab),
	.w7(32'h3c182ef0),
	.w8(32'h3cab680c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceea5e2),
	.w1(32'h3d052a75),
	.w2(32'h3ccd008f),
	.w3(32'h3c60908a),
	.w4(32'h3bf37972),
	.w5(32'h3c9e92bc),
	.w6(32'h3bf36ecb),
	.w7(32'hbaa54ea0),
	.w8(32'h3c9c6047),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7732d),
	.w1(32'h3b8da462),
	.w2(32'h3c038244),
	.w3(32'h3a9064f3),
	.w4(32'hba5f5a52),
	.w5(32'h3b88d7c1),
	.w6(32'h3bef17c4),
	.w7(32'h3bcc91ad),
	.w8(32'hbaac2ab2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73c7c1),
	.w1(32'hbaa3af76),
	.w2(32'h3b2e15ce),
	.w3(32'h3c2974e0),
	.w4(32'hbb7deb3b),
	.w5(32'h3a079f6c),
	.w6(32'h3c604215),
	.w7(32'h3bba857e),
	.w8(32'h3beae29b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b843173),
	.w1(32'h3a9acd0a),
	.w2(32'h3b3a3257),
	.w3(32'h3ad3b0d6),
	.w4(32'hba5659c0),
	.w5(32'h3a360fd6),
	.w6(32'h3b84d4ec),
	.w7(32'h3b7e4cf3),
	.w8(32'hbc61218c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd877d),
	.w1(32'hbc901ba7),
	.w2(32'hbc9002b8),
	.w3(32'h3cdacb18),
	.w4(32'hba4d4f03),
	.w5(32'hbc7f25d5),
	.w6(32'h3d0ed469),
	.w7(32'h3bfad1c1),
	.w8(32'hbc5f5c17),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23aac7),
	.w1(32'hbc0893f9),
	.w2(32'hbc0b3dd2),
	.w3(32'h3c344f58),
	.w4(32'hba9d0cb2),
	.w5(32'hbc4091b1),
	.w6(32'h3bd1d3b3),
	.w7(32'h3bb7dbd1),
	.w8(32'hbbd1c87e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716e7d),
	.w1(32'h3b4abcf6),
	.w2(32'h3b8dd8a4),
	.w3(32'hbb8aaea4),
	.w4(32'h3b52391c),
	.w5(32'h3b99a2f2),
	.w6(32'h3c114681),
	.w7(32'h3b40b741),
	.w8(32'h3cbef45a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdecce8),
	.w1(32'h3c714f3c),
	.w2(32'hbc016ad9),
	.w3(32'h3c20438e),
	.w4(32'h3b82c21d),
	.w5(32'h3c0bdb11),
	.w6(32'hba3c1593),
	.w7(32'hbbf190ce),
	.w8(32'h3ae5e855),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63653b),
	.w1(32'hbbc5354b),
	.w2(32'hbc0f985c),
	.w3(32'h3c433e82),
	.w4(32'hbc3f535a),
	.w5(32'hbbb8cdda),
	.w6(32'h3c950c9f),
	.w7(32'h3bb37e97),
	.w8(32'h3b1a53f1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d138c22),
	.w1(32'hbcab4fc9),
	.w2(32'hbc07fe64),
	.w3(32'h3d151ab4),
	.w4(32'hbc3a2c89),
	.w5(32'hbc357cbc),
	.w6(32'h3d496cfd),
	.w7(32'h3c1d2570),
	.w8(32'hbbb73ff1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd71ebb),
	.w1(32'h3c33bbdd),
	.w2(32'hbb363b1d),
	.w3(32'h3dcf6117),
	.w4(32'h3b9d97d3),
	.w5(32'hbce86490),
	.w6(32'h3dc7b89e),
	.w7(32'h3c95d792),
	.w8(32'h3b914f18),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4d398c),
	.w1(32'hbcbf4a2d),
	.w2(32'hbc4c6e75),
	.w3(32'h3d6412e6),
	.w4(32'hbc93c6fa),
	.w5(32'hbcbeb301),
	.w6(32'h3d7ac792),
	.w7(32'hba6e77d6),
	.w8(32'hbbc3d5dc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33d4d9),
	.w1(32'h3a03b60a),
	.w2(32'h3aa85ce6),
	.w3(32'h3c48d9dc),
	.w4(32'hbb906fe7),
	.w5(32'hbbb6b7c9),
	.w6(32'h3c558134),
	.w7(32'h3c6bbf35),
	.w8(32'h3b04e83f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc909a2d),
	.w1(32'h3b1c1e13),
	.w2(32'hbcb68735),
	.w3(32'hbc1013ac),
	.w4(32'hbc1686f9),
	.w5(32'hbc7f821c),
	.w6(32'hbc5dea08),
	.w7(32'hbca5c7ec),
	.w8(32'hbb8a3524),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9970aa),
	.w1(32'hbc12657d),
	.w2(32'hbc3c9011),
	.w3(32'h3bc5921d),
	.w4(32'h3b8bcc5e),
	.w5(32'hbc2b53e2),
	.w6(32'hba59c72f),
	.w7(32'hba8163bb),
	.w8(32'h3be95f4d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40ca7a),
	.w1(32'hbcce5bd7),
	.w2(32'h3bdce3ce),
	.w3(32'hbb7ac247),
	.w4(32'hbc9ad576),
	.w5(32'hbb9aebae),
	.w6(32'hbaba8f25),
	.w7(32'h3c59d1f2),
	.w8(32'hbbcc3076),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f6ed2),
	.w1(32'h3b0d11d1),
	.w2(32'hbca24ca5),
	.w3(32'hbc0bd2df),
	.w4(32'hbbe9af03),
	.w5(32'hbc520947),
	.w6(32'hbc420d0d),
	.w7(32'hbc8a3f80),
	.w8(32'hbb3abcdf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c220298),
	.w1(32'h3bd797eb),
	.w2(32'hbc7c1523),
	.w3(32'h3c8c76de),
	.w4(32'hbbdfa749),
	.w5(32'hbc8a5c61),
	.w6(32'h3c5cdefe),
	.w7(32'hbc57f83d),
	.w8(32'h3bbd9647),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7392ea),
	.w1(32'hbb8b0ad8),
	.w2(32'hba60cfc5),
	.w3(32'h3ae6dcc6),
	.w4(32'hbc3c1503),
	.w5(32'hbbac183a),
	.w6(32'hb9c04488),
	.w7(32'h3ba0f00f),
	.w8(32'hbb908ea9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf9c15a),
	.w1(32'h3d157598),
	.w2(32'hbc17d550),
	.w3(32'h3ccd363a),
	.w4(32'h3d1149bc),
	.w5(32'h3c85f21b),
	.w6(32'h3d7cce93),
	.w7(32'hbcb6a06e),
	.w8(32'h3b0c23d5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c632d07),
	.w1(32'hbbced947),
	.w2(32'hbac9d165),
	.w3(32'h3c72332a),
	.w4(32'hbb40c986),
	.w5(32'hbb3fc15f),
	.w6(32'h3c961743),
	.w7(32'h3ac556b1),
	.w8(32'h3bc94e8e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd7fb),
	.w1(32'hbb87c0f3),
	.w2(32'hbc3ab7f1),
	.w3(32'h3bb78508),
	.w4(32'hbad9c2fc),
	.w5(32'hbafdbdd0),
	.w6(32'hbb473d87),
	.w7(32'h3a17d519),
	.w8(32'h3c2bdbaa),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ffca8),
	.w1(32'hbcccdc44),
	.w2(32'hbc9ff523),
	.w3(32'h3cd0765f),
	.w4(32'hbcb2bff4),
	.w5(32'hbce4d820),
	.w6(32'h3c36529a),
	.w7(32'hbbb065bb),
	.w8(32'hbc1ad91a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d526970),
	.w1(32'h3c3ed70c),
	.w2(32'hbccb8320),
	.w3(32'h3ce70594),
	.w4(32'hbbaf0c75),
	.w5(32'hbcb93bfa),
	.w6(32'h3cb6a3ba),
	.w7(32'hbbc92ddf),
	.w8(32'h3b5d79d0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825ac7),
	.w1(32'h3bb2d1dd),
	.w2(32'hbaee5224),
	.w3(32'h3c3a6cc7),
	.w4(32'h3d0f0027),
	.w5(32'hb91b5459),
	.w6(32'hbc9c267b),
	.w7(32'hbb6422c3),
	.w8(32'hbc4423d9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cf3bf),
	.w1(32'hbb1e75f8),
	.w2(32'hb8934316),
	.w3(32'hbb82e0db),
	.w4(32'h3bf5aef2),
	.w5(32'h3b370a7b),
	.w6(32'h3ba7229c),
	.w7(32'h3c310232),
	.w8(32'hbb852412),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2fd48),
	.w1(32'hbbcf2f64),
	.w2(32'hbb50b20c),
	.w3(32'h3ac19130),
	.w4(32'h3b7a7728),
	.w5(32'hbb5bb81a),
	.w6(32'h3aca6da2),
	.w7(32'h3b78f84a),
	.w8(32'h3bdbccbe),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbba202),
	.w1(32'hbcc4d071),
	.w2(32'h3aa56d58),
	.w3(32'h3c0c24f5),
	.w4(32'hbc37eadd),
	.w5(32'h39a29ae7),
	.w6(32'hbace9f69),
	.w7(32'h3c329a11),
	.w8(32'hba2139cb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986ce4),
	.w1(32'h39bb0703),
	.w2(32'hbb0fe2e1),
	.w3(32'h3ad4d831),
	.w4(32'h39b2e1d2),
	.w5(32'hbb0e0af3),
	.w6(32'h3b2623b6),
	.w7(32'h3b05c2b0),
	.w8(32'hbb46b044),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c442242),
	.w1(32'hbb60291e),
	.w2(32'hbb2ad401),
	.w3(32'h3c1ab758),
	.w4(32'h3b8f4ab2),
	.w5(32'hbb84e360),
	.w6(32'h3bad6d61),
	.w7(32'h3ba965c8),
	.w8(32'h3b5eaad1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4619ff),
	.w1(32'hbc1fb6dd),
	.w2(32'h3b9d61ef),
	.w3(32'h3c827aca),
	.w4(32'hbc8d2d53),
	.w5(32'h39e9a76a),
	.w6(32'h3ca32a4d),
	.w7(32'h3c034017),
	.w8(32'h3b3693fe),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcf8e8),
	.w1(32'h39dcdcae),
	.w2(32'hbb3ee54d),
	.w3(32'h3b0ca3c3),
	.w4(32'hbbcedd40),
	.w5(32'hbb189d9e),
	.w6(32'h3ac7bd9b),
	.w7(32'hbc1748d0),
	.w8(32'h3b5b0100),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca041d),
	.w1(32'hbc858387),
	.w2(32'hbbf37826),
	.w3(32'h3c852264),
	.w4(32'hbb37d8f2),
	.w5(32'hbb43d941),
	.w6(32'h3c6679aa),
	.w7(32'hbb28eb50),
	.w8(32'h3bd53422),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b754ce),
	.w1(32'hba84884a),
	.w2(32'h39208601),
	.w3(32'hbacf57d7),
	.w4(32'hbb1843ba),
	.w5(32'h39c32cdc),
	.w6(32'hbb888c84),
	.w7(32'hba853c52),
	.w8(32'h3afee248),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c4225),
	.w1(32'hbba867cf),
	.w2(32'h3bcbe51c),
	.w3(32'h3c2b8b98),
	.w4(32'hbc0705d3),
	.w5(32'h3b23b9cf),
	.w6(32'h3c4fa4a4),
	.w7(32'hbbbb716b),
	.w8(32'h3bab49ca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5fc3b),
	.w1(32'hb9834af4),
	.w2(32'h3b5357c5),
	.w3(32'h3baf40c7),
	.w4(32'hba8755bf),
	.w5(32'h3aac49d2),
	.w6(32'h3bc97ea0),
	.w7(32'h38e9dbf3),
	.w8(32'h3b272055),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e89a95),
	.w1(32'h3b679202),
	.w2(32'h3b1e8857),
	.w3(32'h39fc4ff3),
	.w4(32'h3b119543),
	.w5(32'h3aa2c71c),
	.w6(32'hb98d8194),
	.w7(32'h3a68d679),
	.w8(32'h39bd1630),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d034b56),
	.w1(32'h3a9728fe),
	.w2(32'h3a00e78f),
	.w3(32'h3cd44016),
	.w4(32'hbc301b8e),
	.w5(32'hbbfb8daf),
	.w6(32'h3cf46fcf),
	.w7(32'hbb06c199),
	.w8(32'h3a8b1d09),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b4d11),
	.w1(32'h3a8a9bb7),
	.w2(32'h3b4e78b7),
	.w3(32'h3d0d2d95),
	.w4(32'hbb7205ed),
	.w5(32'h3a85b77c),
	.w6(32'h3d1ff3e7),
	.w7(32'hbac88768),
	.w8(32'h3bff3b8c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2d73),
	.w1(32'hbbd50955),
	.w2(32'h3c1e4892),
	.w3(32'h3b54c198),
	.w4(32'hbc03571d),
	.w5(32'h3bee0fef),
	.w6(32'h3b578e5f),
	.w7(32'hbbb882b4),
	.w8(32'h3bf06314),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4068d4),
	.w1(32'h3a1a0916),
	.w2(32'h3a472726),
	.w3(32'hbb0bd8c0),
	.w4(32'h3a90ea0b),
	.w5(32'h3a88c387),
	.w6(32'hbb42a22b),
	.w7(32'h3a72dc58),
	.w8(32'h3a2f22da),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b19df),
	.w1(32'h3aa475b2),
	.w2(32'h38c51390),
	.w3(32'hba03c8de),
	.w4(32'h3b875ed2),
	.w5(32'h3af023e1),
	.w6(32'hb9b4e742),
	.w7(32'h3b956774),
	.w8(32'h3aac3489),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf10659),
	.w1(32'hbae98609),
	.w2(32'hba948c6e),
	.w3(32'hb8fa0080),
	.w4(32'hba0a1676),
	.w5(32'hba3bffa9),
	.w6(32'hba2eac29),
	.w7(32'hba683103),
	.w8(32'h3a9d62ba),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7dad6),
	.w1(32'hbb0f513e),
	.w2(32'h3b861cb2),
	.w3(32'h3c8a69a8),
	.w4(32'hbbd67d02),
	.w5(32'h384b214a),
	.w6(32'h3c878912),
	.w7(32'h398b8215),
	.w8(32'hb93c2f50),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91775b),
	.w1(32'hbc3feb2a),
	.w2(32'hbc32120c),
	.w3(32'h3caffb11),
	.w4(32'hbb277ea4),
	.w5(32'hbbc21f97),
	.w6(32'h3ccc8f45),
	.w7(32'hbba0851c),
	.w8(32'hbbaddb47),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8987cf),
	.w1(32'h3b54d084),
	.w2(32'hbb160e14),
	.w3(32'hbb042013),
	.w4(32'h3ab919a3),
	.w5(32'hbb86b779),
	.w6(32'h383c678d),
	.w7(32'hbb38df2b),
	.w8(32'h3b86e0c1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b534dd4),
	.w1(32'hbb1b9ad1),
	.w2(32'h3b162a6f),
	.w3(32'h3bbd4fae),
	.w4(32'h3af54977),
	.w5(32'h3b6236d7),
	.w6(32'h3b6bda3e),
	.w7(32'h3b2d766e),
	.w8(32'hbb24d4ff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c525465),
	.w1(32'h3c0ca744),
	.w2(32'h3bd9cd09),
	.w3(32'h3c1dac6a),
	.w4(32'hbb83b4f2),
	.w5(32'hbb432fa0),
	.w6(32'h3c8f9fcc),
	.w7(32'h3c031ef1),
	.w8(32'h3c10e791),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0100e),
	.w1(32'h3bf71ada),
	.w2(32'h3a78c843),
	.w3(32'hb972dedd),
	.w4(32'h3b9cf859),
	.w5(32'h3ac187f9),
	.w6(32'h3b8dfb88),
	.w7(32'h3baeea8e),
	.w8(32'h3c10f19c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae656b6),
	.w1(32'hba3c374a),
	.w2(32'h3abd782c),
	.w3(32'h3b73904e),
	.w4(32'h3a921d12),
	.w5(32'h3b5ddad3),
	.w6(32'hb9ec3b04),
	.w7(32'h3b57541f),
	.w8(32'h39ad5fda),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb877e97b),
	.w1(32'hbb1207b0),
	.w2(32'hbb67673c),
	.w3(32'hb998df12),
	.w4(32'hbb79fc6e),
	.w5(32'hbb97ab28),
	.w6(32'hba7fc6d3),
	.w7(32'hbb4dea9d),
	.w8(32'hba7505e4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dc88a),
	.w1(32'hbb4d259c),
	.w2(32'hba7a5c5d),
	.w3(32'hba9144f7),
	.w4(32'h389f07bb),
	.w5(32'h3acba7f0),
	.w6(32'hbb263f45),
	.w7(32'h3a56731d),
	.w8(32'hb8214e11),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec648),
	.w1(32'hbae0569f),
	.w2(32'h3b548dbc),
	.w3(32'h3bee4e8c),
	.w4(32'h3a033895),
	.w5(32'h3a78f339),
	.w6(32'h3ba6c553),
	.w7(32'hba6d7a95),
	.w8(32'hb7bae6e7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b798d05),
	.w1(32'hbb4bc8f8),
	.w2(32'hba876e9d),
	.w3(32'h3ba58ca8),
	.w4(32'hbb236385),
	.w5(32'h3a5c569d),
	.w6(32'h3bb4fa85),
	.w7(32'h399cdb21),
	.w8(32'h3be95bb9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3610c3),
	.w1(32'hbc2d2c30),
	.w2(32'hbc4b5cbb),
	.w3(32'h3b9e7a3e),
	.w4(32'hbba9321d),
	.w5(32'hbbc89003),
	.w6(32'h3b5e91ac),
	.w7(32'hbb2fe9e8),
	.w8(32'hbbe1e5bc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule