module layer_8_featuremap_69(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39887113),
	.w1(32'h3a846a4f),
	.w2(32'h3b8c2172),
	.w3(32'hb8edf0d7),
	.w4(32'hb9995d69),
	.w5(32'h3be19130),
	.w6(32'h3bd52c70),
	.w7(32'h3b841766),
	.w8(32'h3c1aa188),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7f8e),
	.w1(32'h3b83bc25),
	.w2(32'h3a999adb),
	.w3(32'hbbee815b),
	.w4(32'h3b22eb7e),
	.w5(32'h399ad540),
	.w6(32'hbb5f441c),
	.w7(32'h3a8d2094),
	.w8(32'hbb36f314),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b2cc9),
	.w1(32'h3bc640be),
	.w2(32'h3bcaf0f1),
	.w3(32'hbc23d6a6),
	.w4(32'h3ba12a2a),
	.w5(32'h3bd21e40),
	.w6(32'hbc5e9dcb),
	.w7(32'hbb26f6f3),
	.w8(32'hbad2ce57),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c609c),
	.w1(32'hbbcbe852),
	.w2(32'hbc2c1764),
	.w3(32'hbc2faf58),
	.w4(32'hbc12aa9f),
	.w5(32'hbc2404ac),
	.w6(32'hbc24bbf3),
	.w7(32'hbbf95ac4),
	.w8(32'hbbcfe92b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c6dd8),
	.w1(32'hbc04d432),
	.w2(32'hbbe5f91e),
	.w3(32'hbbdec495),
	.w4(32'hbb361f05),
	.w5(32'hbb6cb658),
	.w6(32'h3b419aaa),
	.w7(32'h3b441d8d),
	.w8(32'h3bb519db),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f1acb),
	.w1(32'hbbb493fa),
	.w2(32'hbbba0f9a),
	.w3(32'hbc1da672),
	.w4(32'hba9e0938),
	.w5(32'hbbba46db),
	.w6(32'hbbe48dee),
	.w7(32'h3bad7dbe),
	.w8(32'hbb5ca994),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14da50),
	.w1(32'h38b616ca),
	.w2(32'hba49c3bc),
	.w3(32'hba5a7931),
	.w4(32'hba2c0930),
	.w5(32'hbaa353aa),
	.w6(32'hb9beb6c9),
	.w7(32'hbab34709),
	.w8(32'hbae7ff8a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e80d7),
	.w1(32'hb96f70ab),
	.w2(32'hbb55f444),
	.w3(32'hbcb72636),
	.w4(32'hbc1f44f9),
	.w5(32'hbbcace46),
	.w6(32'hbc104ca9),
	.w7(32'h3af8bf85),
	.w8(32'h39e081da),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0f73),
	.w1(32'h3bbf2965),
	.w2(32'h3be16cdc),
	.w3(32'hbbaef66b),
	.w4(32'h3ad6305c),
	.w5(32'h3b1ab87f),
	.w6(32'h3b53fc3d),
	.w7(32'h3b869516),
	.w8(32'h3b73ad6e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb74ab8),
	.w1(32'h3c3a1b18),
	.w2(32'h3c7bd2ea),
	.w3(32'hbc3644e6),
	.w4(32'h3aa5a27b),
	.w5(32'h3c0bacdd),
	.w6(32'hbb1a424c),
	.w7(32'h3b962065),
	.w8(32'h3a78eb10),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f1b4),
	.w1(32'hbc246f4a),
	.w2(32'hbc1eae49),
	.w3(32'hbc14dcff),
	.w4(32'hbbf18892),
	.w5(32'hbba2dbf0),
	.w6(32'hbac25e1a),
	.w7(32'hba5cd339),
	.w8(32'h39b7fc94),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb8c97),
	.w1(32'hba6800d2),
	.w2(32'hbba229c4),
	.w3(32'hbbe42459),
	.w4(32'hbb8f344e),
	.w5(32'hbbbc8966),
	.w6(32'hbbb4e9b5),
	.w7(32'hbbb8fc9c),
	.w8(32'hbba51758),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54be9b),
	.w1(32'h3b7666ec),
	.w2(32'h3a78f741),
	.w3(32'hbc64cef5),
	.w4(32'h39e54356),
	.w5(32'hbb352ce6),
	.w6(32'hbc0eb015),
	.w7(32'h3b0d691a),
	.w8(32'h3bbc69d5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9b29d),
	.w1(32'h3b0e31be),
	.w2(32'h3b927707),
	.w3(32'h3bbc256f),
	.w4(32'h3b009c1b),
	.w5(32'h3b471fa1),
	.w6(32'h3b914503),
	.w7(32'h3bbaa130),
	.w8(32'h3b75c56d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d97b0),
	.w1(32'h3ae734b9),
	.w2(32'h3b1d921e),
	.w3(32'h3b3425c0),
	.w4(32'h3ae5f317),
	.w5(32'h3aca58dc),
	.w6(32'h3b1cfa23),
	.w7(32'h3b4f8072),
	.w8(32'hb7e9880e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64164e),
	.w1(32'h394abb70),
	.w2(32'h3851c102),
	.w3(32'hba8c020f),
	.w4(32'hba347b9a),
	.w5(32'hba53e7d0),
	.w6(32'hb8dc9431),
	.w7(32'hb9ae4231),
	.w8(32'hbaf6c4a5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d1a0),
	.w1(32'hbbd3091d),
	.w2(32'h3a9f2f10),
	.w3(32'hbbbde8f8),
	.w4(32'hbb984c61),
	.w5(32'hba2886a2),
	.w6(32'hbb10ea13),
	.w7(32'hbb705563),
	.w8(32'h3a54699a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc470e1b),
	.w1(32'h3b286f56),
	.w2(32'h3bee79f2),
	.w3(32'hbc7ea869),
	.w4(32'hbb291e85),
	.w5(32'h3ac78f7b),
	.w6(32'hbc41b0f7),
	.w7(32'hbb053206),
	.w8(32'hbb93c577),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3f656d),
	.w1(32'hbcf0260d),
	.w2(32'hbcb605da),
	.w3(32'hbd1f6c00),
	.w4(32'hbce5e044),
	.w5(32'hbb4457fb),
	.w6(32'hbd0dedda),
	.w7(32'hbc69b9be),
	.w8(32'hb79fec0c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc55382),
	.w1(32'hbb596ac0),
	.w2(32'hbc29edf3),
	.w3(32'hbc85d25f),
	.w4(32'h3ae749f4),
	.w5(32'hbb5cdaac),
	.w6(32'hba4e4e1c),
	.w7(32'h3c0d78de),
	.w8(32'hbc44b1dd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15be2c),
	.w1(32'hbc1f6051),
	.w2(32'hbc28a861),
	.w3(32'hbb29bb6a),
	.w4(32'hbc3ae856),
	.w5(32'hbc85319e),
	.w6(32'hb8b3f9f4),
	.w7(32'hbbace806),
	.w8(32'hbc06a57a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e7548),
	.w1(32'h3c6fe83c),
	.w2(32'h3c377d0d),
	.w3(32'hbb189801),
	.w4(32'h3c49e7e1),
	.w5(32'h3c5ecd46),
	.w6(32'hbb9855a2),
	.w7(32'h3c19eac9),
	.w8(32'h3bd25b86),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd0c3),
	.w1(32'h3ae877be),
	.w2(32'h3c9f18cd),
	.w3(32'h3c2d9d6c),
	.w4(32'h3bf004cf),
	.w5(32'h3d0e8b07),
	.w6(32'h3cede43f),
	.w7(32'h3cf5e571),
	.w8(32'h3d53ca73),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1319e1),
	.w1(32'h3c0717fb),
	.w2(32'h3c020ab2),
	.w3(32'h3b87aa9b),
	.w4(32'h3c0ee2d4),
	.w5(32'h3bb626ae),
	.w6(32'h3bf51ba2),
	.w7(32'h3c0e749f),
	.w8(32'h3aa09089),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f571),
	.w1(32'hbb55be31),
	.w2(32'hbb96e065),
	.w3(32'hbbd83e78),
	.w4(32'hbbbbad30),
	.w5(32'hbb8086d3),
	.w6(32'hbbcf3729),
	.w7(32'hbbc329d4),
	.w8(32'hbb87c736),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57cff8),
	.w1(32'hbc4af834),
	.w2(32'hbc3e0511),
	.w3(32'hbb9a6c7a),
	.w4(32'hbc173736),
	.w5(32'hbba79c83),
	.w6(32'h3c2c9e46),
	.w7(32'h3b8fff40),
	.w8(32'h3aec91e3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35be74f7),
	.w1(32'hbac1ef10),
	.w2(32'hbb17d16c),
	.w3(32'h3a29e6c9),
	.w4(32'hba26e257),
	.w5(32'hba3f857b),
	.w6(32'h39ec63ed),
	.w7(32'hbabc8985),
	.w8(32'hbaf35385),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd68f2fd),
	.w1(32'hbc7bf75f),
	.w2(32'hbc363852),
	.w3(32'hbdb3e459),
	.w4(32'hbdb6ac51),
	.w5(32'hbdc36b82),
	.w6(32'h3c81074a),
	.w7(32'hba40cc55),
	.w8(32'h3c468bd6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d8b24),
	.w1(32'hbc276a28),
	.w2(32'hbb892b28),
	.w3(32'hbc6ad18e),
	.w4(32'hbc36a1b1),
	.w5(32'hbbb1171b),
	.w6(32'h3a2a1f2c),
	.w7(32'h3b8665be),
	.w8(32'h3abafd16),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9fad9),
	.w1(32'hba91c515),
	.w2(32'hb8beb658),
	.w3(32'hbb9c8533),
	.w4(32'hba2d151a),
	.w5(32'h39d8ba83),
	.w6(32'hbb95a230),
	.w7(32'hb9e88312),
	.w8(32'hbb6c373d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5399d9),
	.w1(32'hbb55afc6),
	.w2(32'hbaea0517),
	.w3(32'h3968ff43),
	.w4(32'h39db3d1f),
	.w5(32'hba85fd5d),
	.w6(32'hbbbe8fed),
	.w7(32'hba9e3d11),
	.w8(32'h3b302020),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214edd),
	.w1(32'hbb5a3973),
	.w2(32'hbbf3fbce),
	.w3(32'hbbe546f6),
	.w4(32'hbb87060a),
	.w5(32'hbbe8979c),
	.w6(32'hbb9bc4b8),
	.w7(32'hbb425ca5),
	.w8(32'hbc001ba8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70ed3a),
	.w1(32'hbaac4d09),
	.w2(32'hbaae608b),
	.w3(32'hba52fd84),
	.w4(32'hba5d6a52),
	.w5(32'hbae5a1a7),
	.w6(32'hbaac3a32),
	.w7(32'hbb23378f),
	.w8(32'hba1c7636),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3986dc),
	.w1(32'h3814dc0c),
	.w2(32'hba342fa0),
	.w3(32'hbb0afa83),
	.w4(32'hbaec2cf0),
	.w5(32'hb9cda8ab),
	.w6(32'hba7ebe73),
	.w7(32'hba4d0168),
	.w8(32'h3bbeb74a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41fb65),
	.w1(32'h3c7ea1ac),
	.w2(32'h3c30573d),
	.w3(32'h3ae6f2c1),
	.w4(32'h3c7433cf),
	.w5(32'h3b9d80a8),
	.w6(32'hbb6468f5),
	.w7(32'h3c6499cd),
	.w8(32'hbb5f6719),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4a01),
	.w1(32'hbc1e70bf),
	.w2(32'hbb286ff1),
	.w3(32'hbc695915),
	.w4(32'hbc37eb37),
	.w5(32'hbb60face),
	.w6(32'hbbf301be),
	.w7(32'hbbcfbf5b),
	.w8(32'hbc0e02b5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817d61),
	.w1(32'hbb6f82f0),
	.w2(32'hbb3483b9),
	.w3(32'hbbb08d28),
	.w4(32'hbb9e894c),
	.w5(32'hbb22c2fa),
	.w6(32'hbb892a13),
	.w7(32'hbb7539fb),
	.w8(32'hbaaaeccb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe66d3d),
	.w1(32'hbab296d8),
	.w2(32'h39d038b1),
	.w3(32'hbbb476e0),
	.w4(32'hbb15a88a),
	.w5(32'hba6ca208),
	.w6(32'hbb1ca674),
	.w7(32'hb9ec299a),
	.w8(32'h3bb1c3dd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971e7f),
	.w1(32'h3b4dd788),
	.w2(32'h3b77f013),
	.w3(32'h3b9c7bb9),
	.w4(32'h3b6966c6),
	.w5(32'h3b0b66f0),
	.w6(32'h3b89c273),
	.w7(32'h3bb930ad),
	.w8(32'hbabc3611),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0520a6),
	.w1(32'h3a74df5a),
	.w2(32'hb9b9a779),
	.w3(32'hbae00720),
	.w4(32'hbb3b6b4e),
	.w5(32'hbb16d772),
	.w6(32'h3af88e89),
	.w7(32'hbb01f64f),
	.w8(32'h3a70a90a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd67d850),
	.w1(32'hbcc5ed74),
	.w2(32'hbd0905fa),
	.w3(32'hbd73285b),
	.w4(32'hbccd769a),
	.w5(32'hbd036838),
	.w6(32'hbd4a090c),
	.w7(32'hbca9cce3),
	.w8(32'hbd0ff90f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc512af7),
	.w1(32'hbb00c183),
	.w2(32'hbb4a4e7c),
	.w3(32'hbc614603),
	.w4(32'hbb81fe09),
	.w5(32'hb8e55c29),
	.w6(32'hbc2746f3),
	.w7(32'hbaed59a1),
	.w8(32'h3b67ab28),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eb74d),
	.w1(32'hbbf586c0),
	.w2(32'h3b51b4e4),
	.w3(32'h3b3c6a65),
	.w4(32'hbb09fda5),
	.w5(32'hbb3b1c87),
	.w6(32'hbb96f00c),
	.w7(32'h3c81cd90),
	.w8(32'hbb608b0a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc311706),
	.w1(32'hbb31b1d3),
	.w2(32'hbbc27c72),
	.w3(32'hbc179d62),
	.w4(32'hbb74f973),
	.w5(32'hba97bf4b),
	.w6(32'hbbb240da),
	.w7(32'h3a2664cd),
	.w8(32'hbb80c35b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb323b4),
	.w1(32'hbc9bce04),
	.w2(32'hbc226051),
	.w3(32'hbc8dd631),
	.w4(32'hbc71ccd7),
	.w5(32'hbb40be40),
	.w6(32'hbbb6886d),
	.w7(32'h3bf98b2b),
	.w8(32'h3baac861),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d43b9),
	.w1(32'h3b75662b),
	.w2(32'h3bd228cd),
	.w3(32'hbc4ff41d),
	.w4(32'h3bbe877a),
	.w5(32'h3b8c4e11),
	.w6(32'hbc473962),
	.w7(32'h3b0dafd1),
	.w8(32'h3c61f782),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb595050),
	.w1(32'hbc01ff54),
	.w2(32'hbbec3924),
	.w3(32'hbcc3163a),
	.w4(32'hba7cf539),
	.w5(32'h3afc00cd),
	.w6(32'hbc220f36),
	.w7(32'hbc63718e),
	.w8(32'hbb8ce6dd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02146b),
	.w1(32'h3bef0105),
	.w2(32'hbc3f2b11),
	.w3(32'hbae1ff0c),
	.w4(32'hbb542436),
	.w5(32'hbbc06070),
	.w6(32'h3cb76499),
	.w7(32'hbbf0a958),
	.w8(32'h3c914d3b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2035f7),
	.w1(32'hbb99427c),
	.w2(32'hbbce441e),
	.w3(32'h3ac069a9),
	.w4(32'h3ae86403),
	.w5(32'hbbd0608a),
	.w6(32'hbb82bc1a),
	.w7(32'h3b4441e5),
	.w8(32'hbba2f378),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74c608),
	.w1(32'hbb8b7c03),
	.w2(32'hbbd37f73),
	.w3(32'hbc374c32),
	.w4(32'hbb269173),
	.w5(32'hbbb4fcf5),
	.w6(32'hbbe6b0bf),
	.w7(32'hbb531558),
	.w8(32'hbb7c21f9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06a202),
	.w1(32'h39b0e635),
	.w2(32'hbaaedf2c),
	.w3(32'hbc1efd7e),
	.w4(32'h38bfa3af),
	.w5(32'hbb0b482e),
	.w6(32'hbbe84b12),
	.w7(32'h3ab0c451),
	.w8(32'hbc029454),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5c77b0),
	.w1(32'hbd06613c),
	.w2(32'hbceba737),
	.w3(32'hbd81cb79),
	.w4(32'hbd3ab561),
	.w5(32'hbcba3caa),
	.w6(32'hbce63aed),
	.w7(32'hbbc3be02),
	.w8(32'h3c01e675),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6beae7),
	.w1(32'h3c997386),
	.w2(32'hbc2a0490),
	.w3(32'hbbfcf4fb),
	.w4(32'h3c160d49),
	.w5(32'hbb76f17f),
	.w6(32'h3c892147),
	.w7(32'hba23dcd4),
	.w8(32'hbac634ca),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566d90),
	.w1(32'hbc87b2ec),
	.w2(32'hbb9a1cc5),
	.w3(32'hbc87b6aa),
	.w4(32'hbc843a3e),
	.w5(32'hbbb40195),
	.w6(32'hbc57284c),
	.w7(32'hbc2ad815),
	.w8(32'hbbb53934),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9434f8),
	.w1(32'h3bd72878),
	.w2(32'h3acc1992),
	.w3(32'h3a97ae61),
	.w4(32'h3aa39929),
	.w5(32'h3a53e69f),
	.w6(32'hbb713a2b),
	.w7(32'h3ba209d4),
	.w8(32'hbb83f6fc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5e103),
	.w1(32'h3d231d8f),
	.w2(32'h3c57254a),
	.w3(32'hbbb5fcfe),
	.w4(32'h3bb9b7a4),
	.w5(32'h3c2a738a),
	.w6(32'h3c2ab389),
	.w7(32'h3bc4a142),
	.w8(32'hbbc31ec3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cb4f8),
	.w1(32'h3bd23775),
	.w2(32'h3c044113),
	.w3(32'hbca18903),
	.w4(32'h3bd19823),
	.w5(32'hbc9f155b),
	.w6(32'hbca9a67a),
	.w7(32'hbad58056),
	.w8(32'hba56ee96),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16aaf9),
	.w1(32'h3c25aeb2),
	.w2(32'h3b3c91bb),
	.w3(32'hbcca3b72),
	.w4(32'hbc0c1bec),
	.w5(32'hbbf9a4ee),
	.w6(32'hbc592ed4),
	.w7(32'hbb63ebe4),
	.w8(32'h3bab1239),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034939),
	.w1(32'hbb0dac64),
	.w2(32'h3ba23666),
	.w3(32'h3a2a447f),
	.w4(32'h3b400a61),
	.w5(32'h3c28c688),
	.w6(32'h3c540466),
	.w7(32'h3c990046),
	.w8(32'h3b84d7ed),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff70c4),
	.w1(32'hbc8bcfc3),
	.w2(32'hbc98a6dd),
	.w3(32'hbcca561f),
	.w4(32'hbc9384f2),
	.w5(32'hbca292b0),
	.w6(32'hbc60340f),
	.w7(32'hbc694757),
	.w8(32'hbc3eff16),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba196c2),
	.w1(32'hbcb3905a),
	.w2(32'h3bef9bde),
	.w3(32'hbc381d8e),
	.w4(32'h3bc7cc7a),
	.w5(32'h3c2b8ed2),
	.w6(32'hbabad653),
	.w7(32'h39bdf750),
	.w8(32'hbb8ba4be),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784489),
	.w1(32'h3cc13427),
	.w2(32'h3b90ee60),
	.w3(32'hba9fd960),
	.w4(32'h3bfdf597),
	.w5(32'hbbcf17cb),
	.w6(32'h3c2dadda),
	.w7(32'h3a45da13),
	.w8(32'hbc3203ce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd44fb7f),
	.w1(32'hbce77503),
	.w2(32'hbce4baff),
	.w3(32'hbd43a948),
	.w4(32'hbcca27fb),
	.w5(32'hbc811733),
	.w6(32'hbd0b86bf),
	.w7(32'hbc34d8b6),
	.w8(32'hbcc4be52),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30d753),
	.w1(32'hba8f15fb),
	.w2(32'h3c8594c0),
	.w3(32'hbbf16886),
	.w4(32'hbc8caf0b),
	.w5(32'h3aa5f9d3),
	.w6(32'hbc6c7f88),
	.w7(32'h3bc99d05),
	.w8(32'hbba27288),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65c121),
	.w1(32'h3a8a7ad6),
	.w2(32'h3bea6305),
	.w3(32'h394c9e10),
	.w4(32'h39ffc3fd),
	.w5(32'h3bb7b9f2),
	.w6(32'h3b4350de),
	.w7(32'h3c0098d6),
	.w8(32'h3aa4359d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043678),
	.w1(32'h3b9a5e81),
	.w2(32'h3bb8c203),
	.w3(32'hbbae81dc),
	.w4(32'h3ba36756),
	.w5(32'h3c27c96c),
	.w6(32'h3a27b4d1),
	.w7(32'h3c16f2c2),
	.w8(32'h3bb366c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9da5a9),
	.w1(32'hbbdfe97f),
	.w2(32'hbc1e2069),
	.w3(32'hbc7d5635),
	.w4(32'hba91242b),
	.w5(32'hbb0a1cb2),
	.w6(32'hbc44adc8),
	.w7(32'hb90655b7),
	.w8(32'hbc042acd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88a45a),
	.w1(32'h3c00f8e1),
	.w2(32'hbc5a3083),
	.w3(32'hbc6246d7),
	.w4(32'h3a55a239),
	.w5(32'hbbc0e7b3),
	.w6(32'h3b2b2d8a),
	.w7(32'h3ac51c03),
	.w8(32'h3a3147db),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f46b9),
	.w1(32'h394b0742),
	.w2(32'h3b80f194),
	.w3(32'hbb24daff),
	.w4(32'h3a49e866),
	.w5(32'h3b1e5aab),
	.w6(32'h39ba3936),
	.w7(32'h3b15ae4d),
	.w8(32'hbca4edd7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4c4e8d),
	.w1(32'hbc82b3b1),
	.w2(32'h3a5c2e7d),
	.w3(32'hbd0e140a),
	.w4(32'hbca02436),
	.w5(32'h3bb4d7d3),
	.w6(32'hbb7a0824),
	.w7(32'h3c5befb3),
	.w8(32'h3c17a507),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25a4ac),
	.w1(32'hbad31a1f),
	.w2(32'hba4a6e4f),
	.w3(32'hba6a49f6),
	.w4(32'hbaa9a197),
	.w5(32'h3b10ed5e),
	.w6(32'h3a994034),
	.w7(32'h3b15661b),
	.w8(32'hbb3f40f7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e857c),
	.w1(32'h3b608f2f),
	.w2(32'hbb825814),
	.w3(32'hbc9976b3),
	.w4(32'hbb601eca),
	.w5(32'hbc06e69f),
	.w6(32'hbbee7f51),
	.w7(32'hbb0860a9),
	.w8(32'hbc548903),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25856e),
	.w1(32'hbaeb89ea),
	.w2(32'h3a1bf7a0),
	.w3(32'hbb623f95),
	.w4(32'hba718abd),
	.w5(32'h3b6c6381),
	.w6(32'h3848e785),
	.w7(32'h3acb1261),
	.w8(32'h3c6d57a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa5592),
	.w1(32'h3cdfa077),
	.w2(32'hbba545df),
	.w3(32'hbcc719ad),
	.w4(32'hbcdd420c),
	.w5(32'hbb61a3b1),
	.w6(32'hbca6ea1f),
	.w7(32'hbc82d572),
	.w8(32'hbc6b8002),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0ac8),
	.w1(32'hba690f93),
	.w2(32'h3b954828),
	.w3(32'hbbceca96),
	.w4(32'hbb516225),
	.w5(32'h3bcc0a21),
	.w6(32'h3ac803f9),
	.w7(32'h3bb8f142),
	.w8(32'hbb4c3ba9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc377da4),
	.w1(32'hbbf04c0f),
	.w2(32'hbbf1494b),
	.w3(32'hbc248ecd),
	.w4(32'hbbf4763d),
	.w5(32'hbbb52742),
	.w6(32'h3c009a38),
	.w7(32'h3be6b8d6),
	.w8(32'h3a2f564c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40759e),
	.w1(32'h3af3dc5f),
	.w2(32'h3b49a250),
	.w3(32'hba921a6c),
	.w4(32'hb99f81a0),
	.w5(32'h3aeaf7d9),
	.w6(32'h3b6ecfd4),
	.w7(32'h3b29bc25),
	.w8(32'hbcca9b88),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd47f95c),
	.w1(32'hbbdf0d6b),
	.w2(32'h3b586500),
	.w3(32'hbd08638d),
	.w4(32'hbb580635),
	.w5(32'h3c80c019),
	.w6(32'h39a2d996),
	.w7(32'h3c951958),
	.w8(32'hbc58eaf2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d818a),
	.w1(32'h3c2ec2be),
	.w2(32'h3ca3a593),
	.w3(32'hbc75097e),
	.w4(32'h3c22f985),
	.w5(32'h3cd6ed0e),
	.w6(32'hba06fd8b),
	.w7(32'h3c2cdb53),
	.w8(32'hbac00667),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb6f76),
	.w1(32'h3b78fc8e),
	.w2(32'h392e25ef),
	.w3(32'hbbf025e9),
	.w4(32'hbb1103d6),
	.w5(32'hba1de7f7),
	.w6(32'hba5d4aa5),
	.w7(32'hbb1cd4c3),
	.w8(32'hbaadc6f9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d4a52),
	.w1(32'h3b8edae9),
	.w2(32'hbc0e032c),
	.w3(32'hbc19a77f),
	.w4(32'h3c130a9f),
	.w5(32'hbb6f8f7f),
	.w6(32'hbbd646e8),
	.w7(32'hbbf8eeb4),
	.w8(32'hbb5dc015),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca330a7),
	.w1(32'hbb8dae53),
	.w2(32'hba9c3cb0),
	.w3(32'hbc33fe4d),
	.w4(32'hbb6fa288),
	.w5(32'hbb4a19c4),
	.w6(32'hbc45e080),
	.w7(32'hbb4f129f),
	.w8(32'hbbcbd6db),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3687e),
	.w1(32'hba4e9f85),
	.w2(32'hbc160bbf),
	.w3(32'hbcb056d7),
	.w4(32'h3825b5b1),
	.w5(32'hbbf75d4d),
	.w6(32'hbb9ff1ce),
	.w7(32'hb8ad2bd4),
	.w8(32'hbc5a06ba),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08c9c8),
	.w1(32'h3b0ef8d4),
	.w2(32'hbd64a3e4),
	.w3(32'hbd4cba93),
	.w4(32'hbd27e405),
	.w5(32'hbd581735),
	.w6(32'hbd439f65),
	.w7(32'hbc4a8dfa),
	.w8(32'hbd41a6fd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0dc0df),
	.w1(32'hbc8cd5bc),
	.w2(32'hbc9a1e7b),
	.w3(32'hbcce380d),
	.w4(32'hbc79c3a3),
	.w5(32'hbc0bc157),
	.w6(32'hbb6e13e2),
	.w7(32'h3bb4b224),
	.w8(32'hba764413),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83c18c),
	.w1(32'hbc8317ae),
	.w2(32'hbc647130),
	.w3(32'hbc38a0ec),
	.w4(32'hbc8f27fa),
	.w5(32'hbc76170f),
	.w6(32'h3c8caa64),
	.w7(32'h3ba31ee7),
	.w8(32'h3c5cc899),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122585),
	.w1(32'hbc24aa2c),
	.w2(32'hbc261cb1),
	.w3(32'h3c82e710),
	.w4(32'h3aae508d),
	.w5(32'hbbe0aca7),
	.w6(32'h3c10b95a),
	.w7(32'h3b12e7f5),
	.w8(32'hbbabe1b9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b030a4),
	.w1(32'hbb5b3197),
	.w2(32'h3be435c8),
	.w3(32'hbae8af0d),
	.w4(32'h3a351c16),
	.w5(32'h3c2d2553),
	.w6(32'hbb963b44),
	.w7(32'h3b59c4c7),
	.w8(32'hbc1aa33e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b704d67),
	.w1(32'h3b5d6362),
	.w2(32'hbc73683f),
	.w3(32'hbc1145d7),
	.w4(32'hbc0f461b),
	.w5(32'hbbb6fa61),
	.w6(32'hbbb27a8c),
	.w7(32'hbacbf625),
	.w8(32'h3c53ddc6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8b49e),
	.w1(32'hbc4b5435),
	.w2(32'hbc422461),
	.w3(32'h3c60666f),
	.w4(32'hbb809ac3),
	.w5(32'hbc622560),
	.w6(32'h3c67f31f),
	.w7(32'h3b74dc7d),
	.w8(32'h3c049f99),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0a63),
	.w1(32'hbc78d5b7),
	.w2(32'hbc935c04),
	.w3(32'h39183ce8),
	.w4(32'hbbf9e068),
	.w5(32'hbc866485),
	.w6(32'hb9a1a047),
	.w7(32'hba9c588d),
	.w8(32'hba9aea10),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae92300),
	.w1(32'hbbc93daf),
	.w2(32'h39db7d01),
	.w3(32'h3a94c3c9),
	.w4(32'hbae74cdf),
	.w5(32'h3b3ac26a),
	.w6(32'h3a17445d),
	.w7(32'h3a8d85e0),
	.w8(32'hbcf85d63),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd184004),
	.w1(32'h3c577c08),
	.w2(32'hbb6dd677),
	.w3(32'hbd3c8ad5),
	.w4(32'hbc69de34),
	.w5(32'hbc9ba9f3),
	.w6(32'hbd01ae7e),
	.w7(32'hbc9715eb),
	.w8(32'hbbf696fc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40fb6e),
	.w1(32'hb9c44ec9),
	.w2(32'hbb067c0c),
	.w3(32'hbc2b0ee6),
	.w4(32'hba7d5e25),
	.w5(32'hba526287),
	.w6(32'hbba7ff4b),
	.w7(32'h3b4195bd),
	.w8(32'hbc98d317),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1455c9),
	.w1(32'h3d0b6107),
	.w2(32'hbb289c24),
	.w3(32'h3c609704),
	.w4(32'h3b0f2138),
	.w5(32'hbc49d103),
	.w6(32'hbc478bc6),
	.w7(32'hbc1bdc35),
	.w8(32'h3bd2f842),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096ae0),
	.w1(32'hbbe59260),
	.w2(32'hbb97070e),
	.w3(32'h3adad323),
	.w4(32'hbbc7288c),
	.w5(32'h39eedcdc),
	.w6(32'h3c2c85b0),
	.w7(32'h3bde3e61),
	.w8(32'hbc6a75c9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4e1c54),
	.w1(32'hbb9fc0a7),
	.w2(32'hbc13b747),
	.w3(32'hbd2df7a2),
	.w4(32'hbb907beb),
	.w5(32'hbc935241),
	.w6(32'h3c5db751),
	.w7(32'h3c338afa),
	.w8(32'hbc43d67b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fdb49),
	.w1(32'h3c47e4e2),
	.w2(32'hbc2a1b8f),
	.w3(32'hbaebfb9f),
	.w4(32'hbc9e0e8a),
	.w5(32'hbb800a24),
	.w6(32'h3bdc94d9),
	.w7(32'h3be14f86),
	.w8(32'hbcb07482),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7bc9e),
	.w1(32'h3bf045a8),
	.w2(32'h3c7d809e),
	.w3(32'hbc7cc485),
	.w4(32'h3c006950),
	.w5(32'h3cbe8158),
	.w6(32'h3bd0de27),
	.w7(32'h3c852db0),
	.w8(32'hbb3f86ff),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99bc90),
	.w1(32'h3b27dd1a),
	.w2(32'h3bb8e124),
	.w3(32'h388baa0d),
	.w4(32'h3bb1f49e),
	.w5(32'h3bc629b5),
	.w6(32'h3b3043c7),
	.w7(32'h3b894e21),
	.w8(32'hbbb0800e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb070b),
	.w1(32'hbc2d94d6),
	.w2(32'hbbb4e68f),
	.w3(32'hbc75a04b),
	.w4(32'hbb6d1a32),
	.w5(32'h3a20c8f2),
	.w6(32'hbb8777db),
	.w7(32'hbc072c32),
	.w8(32'hbbb16410),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3294b1),
	.w1(32'hbbf1261a),
	.w2(32'hbbc97626),
	.w3(32'hbc1af8a6),
	.w4(32'hbbf03bdb),
	.w5(32'hbb8608fe),
	.w6(32'hbbd6167f),
	.w7(32'hbbb82d36),
	.w8(32'hbcd05faa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd027382),
	.w1(32'h3c8c8543),
	.w2(32'h3cb17d78),
	.w3(32'hbcb28710),
	.w4(32'h3c4da22b),
	.w5(32'h3ce867c5),
	.w6(32'h3b91ca76),
	.w7(32'h3c7312e4),
	.w8(32'h3b6bdd60),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066718),
	.w1(32'h3b945186),
	.w2(32'h3a9d391a),
	.w3(32'hbc43f6d3),
	.w4(32'h3bdbdea6),
	.w5(32'h3b2129d2),
	.w6(32'hbc155acb),
	.w7(32'h3b802bbf),
	.w8(32'h3b07d751),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ce70c),
	.w1(32'h3b7da7db),
	.w2(32'hbb0a8930),
	.w3(32'h3b98882f),
	.w4(32'h3be3a9d2),
	.w5(32'hbb1d17aa),
	.w6(32'hb980f413),
	.w7(32'h3b88ee4d),
	.w8(32'h3ac3c4f9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc431b6c),
	.w1(32'hbc48b09f),
	.w2(32'hbc4b6ba8),
	.w3(32'hbb8f113b),
	.w4(32'hbc3575fd),
	.w5(32'hbbfff85b),
	.w6(32'h3b9b7f44),
	.w7(32'hba26d3dd),
	.w8(32'hbb0a135f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eed80),
	.w1(32'h3be6ab13),
	.w2(32'h3becefb6),
	.w3(32'h3c51f773),
	.w4(32'h3c6533ff),
	.w5(32'h39fac74f),
	.w6(32'h3b872e10),
	.w7(32'h3c25445c),
	.w8(32'h3bdd39ef),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a5fc),
	.w1(32'h3bfe9c4e),
	.w2(32'hbb7e2ebf),
	.w3(32'hbbb27bc0),
	.w4(32'hba84f2e3),
	.w5(32'hbc113418),
	.w6(32'h399ef392),
	.w7(32'h3b73f7a0),
	.w8(32'h3b8c1fa6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c2006),
	.w1(32'h3b59ca33),
	.w2(32'hbbaf7cd0),
	.w3(32'h3b15b373),
	.w4(32'hba1dcd85),
	.w5(32'hbc104253),
	.w6(32'h3b15e51e),
	.w7(32'h3b4b664b),
	.w8(32'hbb57bbad),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5561ed),
	.w1(32'hbba180e5),
	.w2(32'h3b56d55a),
	.w3(32'hbb96c800),
	.w4(32'hbb2cc66b),
	.w5(32'hbb0eddf7),
	.w6(32'h395a521d),
	.w7(32'h3b37bd0a),
	.w8(32'hbc36730b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0105f),
	.w1(32'hb9cdaab3),
	.w2(32'h3b6d4bc4),
	.w3(32'hbc233856),
	.w4(32'h3b0de481),
	.w5(32'hbc53a593),
	.w6(32'hbc5f3b35),
	.w7(32'h3c195a08),
	.w8(32'hb9dfc653),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e51ab),
	.w1(32'h3c07d5ba),
	.w2(32'h3a628455),
	.w3(32'hbc5d09d8),
	.w4(32'h3bde8c0c),
	.w5(32'h3ba6f74f),
	.w6(32'hbc100bce),
	.w7(32'h3c7e2f0c),
	.w8(32'hbcc2dd4d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73511f),
	.w1(32'h3ca844be),
	.w2(32'h3cffdad9),
	.w3(32'hb94fb423),
	.w4(32'h3d148b3e),
	.w5(32'h3d3fd223),
	.w6(32'hbca17a53),
	.w7(32'h3c8f5a5f),
	.w8(32'h3c60f83e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f8d60),
	.w1(32'hbb3815cb),
	.w2(32'hbbecca24),
	.w3(32'h3aa7e3d2),
	.w4(32'hbbc38a7d),
	.w5(32'hbc3990be),
	.w6(32'h3b67dcbd),
	.w7(32'hbb1f1f4f),
	.w8(32'h3b8a0df4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dfe23),
	.w1(32'hbb37c799),
	.w2(32'hbbc1e536),
	.w3(32'h3a1567fa),
	.w4(32'hbbe7b5e8),
	.w5(32'hbc0601e0),
	.w6(32'h3b32181a),
	.w7(32'hbb7c514f),
	.w8(32'h3c02bbbc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a854188),
	.w1(32'hbbf14dcc),
	.w2(32'hbc7f6e79),
	.w3(32'hbb7c2d7c),
	.w4(32'hbc6f9297),
	.w5(32'hbc8f7acc),
	.w6(32'h3b8c2321),
	.w7(32'hbb784087),
	.w8(32'hbbc29079),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc204cd8),
	.w1(32'h3b4e6f9f),
	.w2(32'h3b850c23),
	.w3(32'hbbc93b66),
	.w4(32'hbc2e6d02),
	.w5(32'h3a11b093),
	.w6(32'hbc02a787),
	.w7(32'h3c2429ab),
	.w8(32'hbca4d8cc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd19f49),
	.w1(32'hbb959c50),
	.w2(32'h3c336f80),
	.w3(32'hbc8749cd),
	.w4(32'h3bf7193d),
	.w5(32'h3c91decf),
	.w6(32'hbca52bcf),
	.w7(32'h3b6108d5),
	.w8(32'hbc2beb3b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf4dd1),
	.w1(32'hbb8ef41d),
	.w2(32'h3aac2638),
	.w3(32'hbb7243e5),
	.w4(32'hbb9f6a9f),
	.w5(32'hbbed07e8),
	.w6(32'hbbfa4a47),
	.w7(32'h3b69a4e6),
	.w8(32'hbabda6f8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06856e),
	.w1(32'h3c44bb83),
	.w2(32'h3b098dfd),
	.w3(32'h3b6c321e),
	.w4(32'h3bc007bc),
	.w5(32'h3b82f4b1),
	.w6(32'h3bee4f67),
	.w7(32'h3b5d5f7b),
	.w8(32'hbb277f61),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc138b8d),
	.w1(32'hba3bcb16),
	.w2(32'h3b62e003),
	.w3(32'hbc8c7a3d),
	.w4(32'hbc815e19),
	.w5(32'hbca11a5c),
	.w6(32'hbb1d6d97),
	.w7(32'hbabff6c7),
	.w8(32'hbc2f81af),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9a97e),
	.w1(32'hbbc91d3f),
	.w2(32'h3a85aed6),
	.w3(32'hbb3dc360),
	.w4(32'hbb0e3ca4),
	.w5(32'h3a862ee7),
	.w6(32'h3bb50236),
	.w7(32'h3bed473b),
	.w8(32'h3c5e747d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed3ab),
	.w1(32'hba33e906),
	.w2(32'hbbaffbd5),
	.w3(32'h3b78adac),
	.w4(32'hbb6313d5),
	.w5(32'hbb9989e2),
	.w6(32'h3b9da171),
	.w7(32'h38858d01),
	.w8(32'hbbe5f992),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf79a4),
	.w1(32'hbb7cf421),
	.w2(32'h3bfdea9f),
	.w3(32'hbab2400b),
	.w4(32'h3b6ca71e),
	.w5(32'h3c04b69c),
	.w6(32'hbc753dc4),
	.w7(32'h3b0cfaa7),
	.w8(32'h3b761724),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1638d),
	.w1(32'hbb263f04),
	.w2(32'h3be94a49),
	.w3(32'hbb869e24),
	.w4(32'h3bb75926),
	.w5(32'h3b8c8812),
	.w6(32'hbc02cfd0),
	.w7(32'h3b3aeba8),
	.w8(32'hbb9cac52),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb8c74),
	.w1(32'h3b8db9de),
	.w2(32'hbb6ff2fb),
	.w3(32'h3b837bdc),
	.w4(32'hba87c87a),
	.w5(32'hbb855b04),
	.w6(32'hbb3656af),
	.w7(32'hbb18de2a),
	.w8(32'h3c063bc9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00eada),
	.w1(32'h3b7a1ef1),
	.w2(32'hbb88386b),
	.w3(32'hbbec95e2),
	.w4(32'hbb510be6),
	.w5(32'hbbc0ef3c),
	.w6(32'h3a28fd01),
	.w7(32'hba8ed029),
	.w8(32'h3b38a7c7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09ed27),
	.w1(32'h3b96525c),
	.w2(32'h3bbe51e8),
	.w3(32'h3c16b947),
	.w4(32'h3b2c3749),
	.w5(32'h3c22f97e),
	.w6(32'hbc03d921),
	.w7(32'hbb9add19),
	.w8(32'h3c060b43),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule