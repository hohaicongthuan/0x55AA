module layer_10_featuremap_237(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a097a67),
	.w1(32'hbaccdde8),
	.w2(32'hbaace08b),
	.w3(32'hb9ab52cb),
	.w4(32'h39b87cac),
	.w5(32'h38c2c8d1),
	.w6(32'hb744adf6),
	.w7(32'hba0fedaa),
	.w8(32'hb9cd7e46),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fa1b4),
	.w1(32'h3a262492),
	.w2(32'h3a15a9db),
	.w3(32'h3a872383),
	.w4(32'h3af2ff8a),
	.w5(32'hba2a1b6d),
	.w6(32'hba1241dd),
	.w7(32'hba2b903f),
	.w8(32'hbaeaa533),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8213b2),
	.w1(32'h3942cf3a),
	.w2(32'h3a92be3a),
	.w3(32'hba8fff0f),
	.w4(32'hb9cdc0be),
	.w5(32'h3a80d2ae),
	.w6(32'hba16abf4),
	.w7(32'hbae7a820),
	.w8(32'h3a9fb9f7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a529307),
	.w1(32'h39b20d6b),
	.w2(32'h39a48054),
	.w3(32'h3a658c3e),
	.w4(32'h3a222938),
	.w5(32'hba8fc8f2),
	.w6(32'h39c9861c),
	.w7(32'h37d4840d),
	.w8(32'hba86226c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb1890),
	.w1(32'hb9f86221),
	.w2(32'h39a0d0c7),
	.w3(32'hba79ef8d),
	.w4(32'hba32592d),
	.w5(32'h3a61e35c),
	.w6(32'hbab16ded),
	.w7(32'h39dd46fb),
	.w8(32'h3a0b5117),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008230),
	.w1(32'h37a1c2da),
	.w2(32'h38e088df),
	.w3(32'h3a8e0c54),
	.w4(32'h3aa8e3d7),
	.w5(32'h3ab86807),
	.w6(32'h384d8867),
	.w7(32'hb8e7a99f),
	.w8(32'h3a981ba5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88179bc),
	.w1(32'hba170c1c),
	.w2(32'hb989eefe),
	.w3(32'h37bef7e4),
	.w4(32'h39d13f95),
	.w5(32'h3ac79d06),
	.w6(32'h39a783ad),
	.w7(32'h3a44d597),
	.w8(32'h3b2164de),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2102b),
	.w1(32'hbb472a3b),
	.w2(32'hba9ba890),
	.w3(32'hb8c45128),
	.w4(32'h39ec409d),
	.w5(32'hba369f88),
	.w6(32'hba15b533),
	.w7(32'hba09fd43),
	.w8(32'hbaf1f431),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1397c4),
	.w1(32'hba102633),
	.w2(32'hb99ff473),
	.w3(32'h3a8dd3fc),
	.w4(32'h3b0b7342),
	.w5(32'h3a6e5b72),
	.w6(32'h39bad88e),
	.w7(32'h3a1b47b7),
	.w8(32'h3a23b046),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2332dd),
	.w1(32'h3aaa4121),
	.w2(32'h39860c93),
	.w3(32'hba52a3ed),
	.w4(32'h3b0977ba),
	.w5(32'h3b04c0d8),
	.w6(32'hbbb5a251),
	.w7(32'hbb98a997),
	.w8(32'hbb56b5b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d15b42),
	.w1(32'hb9d2dc3f),
	.w2(32'h38b4f357),
	.w3(32'h3a1a5673),
	.w4(32'h3a19783e),
	.w5(32'hb96c694f),
	.w6(32'hb7634620),
	.w7(32'hb8abdb59),
	.w8(32'hb9c39feb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cee9d),
	.w1(32'hba2864f0),
	.w2(32'hba84d2e1),
	.w3(32'hbb0f9246),
	.w4(32'hbabe84ac),
	.w5(32'hbbb04c4e),
	.w6(32'hb9c441b2),
	.w7(32'hbac1a0f8),
	.w8(32'hbb69b177),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc2286),
	.w1(32'h38c62006),
	.w2(32'h3890ee0d),
	.w3(32'hbb326330),
	.w4(32'hb9eef69b),
	.w5(32'h39f91a16),
	.w6(32'hbb444bb4),
	.w7(32'hbb826267),
	.w8(32'hbb20ec30),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76a820),
	.w1(32'hbac5ceb7),
	.w2(32'hba85978f),
	.w3(32'hbac8f93b),
	.w4(32'hba98deed),
	.w5(32'hbaeeeb20),
	.w6(32'hbaececdb),
	.w7(32'hbab89028),
	.w8(32'hba6947e2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad26346),
	.w1(32'h3a51ca96),
	.w2(32'h39984aa8),
	.w3(32'h3ab2fd26),
	.w4(32'h3b18a648),
	.w5(32'h3a453137),
	.w6(32'hbb20b1b5),
	.w7(32'hbab416f2),
	.w8(32'hbb0f6305),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1087d),
	.w1(32'hba4321fa),
	.w2(32'hba93390d),
	.w3(32'hba844c36),
	.w4(32'h3ad30fd5),
	.w5(32'h3b1c6ae1),
	.w6(32'hbb96536c),
	.w7(32'hbb5ae868),
	.w8(32'hbb19501a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61ae4f),
	.w1(32'h3a3243b1),
	.w2(32'h39bb3f77),
	.w3(32'h3ab299e5),
	.w4(32'h3ae98ace),
	.w5(32'hbab0cbf2),
	.w6(32'h3aa30460),
	.w7(32'h3a4e4185),
	.w8(32'hbaf5ec76),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa1cc),
	.w1(32'hbb848eb2),
	.w2(32'hbb368394),
	.w3(32'hbb5779f8),
	.w4(32'hbb4965d3),
	.w5(32'hbc02c5d3),
	.w6(32'hbb8fab5e),
	.w7(32'hbb62a7b6),
	.w8(32'hbc188f13),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae53f1b),
	.w1(32'hbadcafd7),
	.w2(32'hbaf1dd84),
	.w3(32'hbb7403a8),
	.w4(32'hbb6323c1),
	.w5(32'hbb18d375),
	.w6(32'hbb3495db),
	.w7(32'hbb1ab920),
	.w8(32'hbb3c1cad),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7677f),
	.w1(32'hb9b01e9a),
	.w2(32'hbabdf607),
	.w3(32'hba312203),
	.w4(32'hb9b650d4),
	.w5(32'h3a1e8bc7),
	.w6(32'hbb06f9ac),
	.w7(32'hba696e1c),
	.w8(32'h399636f3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a930f0d),
	.w1(32'h3a3266c5),
	.w2(32'h3899c4ca),
	.w3(32'h3a3657b7),
	.w4(32'h3a92f826),
	.w5(32'h3b4e7879),
	.w6(32'hb9a4b49d),
	.w7(32'h39f01b7b),
	.w8(32'h3b58e878),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aa8a7),
	.w1(32'h3b1d30d3),
	.w2(32'h3af769b4),
	.w3(32'h3b7e2909),
	.w4(32'h3b7a15ce),
	.w5(32'hb9219e2d),
	.w6(32'h3b334d6d),
	.w7(32'h3b4bb579),
	.w8(32'hb996a926),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac548ba),
	.w1(32'h3b915cd0),
	.w2(32'hbb194e75),
	.w3(32'h3acfedad),
	.w4(32'hbb30e9c8),
	.w5(32'hbc18616c),
	.w6(32'hbc17824b),
	.w7(32'hbc32fa3f),
	.w8(32'hbc90e270),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3fb61),
	.w1(32'h3a94dcc8),
	.w2(32'hbad8e452),
	.w3(32'hbace287c),
	.w4(32'h3a4dc442),
	.w5(32'h39f7befd),
	.w6(32'hbbc6d4e4),
	.w7(32'hbbb7dc33),
	.w8(32'hbbd79c8b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8957fb),
	.w1(32'h3a602435),
	.w2(32'hba71db59),
	.w3(32'hbaaae6e9),
	.w4(32'h3b394c2b),
	.w5(32'h3b98c72f),
	.w6(32'hbbf13303),
	.w7(32'hbc088e7d),
	.w8(32'hbb4b56d8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a6151),
	.w1(32'h39959040),
	.w2(32'hb9abd1db),
	.w3(32'h3a487d57),
	.w4(32'h3a1820b1),
	.w5(32'hb88cb341),
	.w6(32'h3a9b82ab),
	.w7(32'h3a9cfe04),
	.w8(32'hba8bc802),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac580ab),
	.w1(32'hbaa39b1a),
	.w2(32'hbad9081f),
	.w3(32'hb8b6f686),
	.w4(32'hb999f3d2),
	.w5(32'hb9b526c4),
	.w6(32'hba35995f),
	.w7(32'hba5b3caf),
	.w8(32'hba216635),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0624b0),
	.w1(32'hba3adfb5),
	.w2(32'hba51217f),
	.w3(32'h39bf4282),
	.w4(32'h3a4c7c96),
	.w5(32'hb8358cea),
	.w6(32'hb8ff5bf4),
	.w7(32'hba983543),
	.w8(32'hbaaf90e1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984702a),
	.w1(32'hb9866efb),
	.w2(32'hba2a522a),
	.w3(32'h3ac28ac4),
	.w4(32'h3a7692f6),
	.w5(32'hbabde7e5),
	.w6(32'hb9dfd1ff),
	.w7(32'h3a68832b),
	.w8(32'hba902055),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd2366),
	.w1(32'h3ae7724d),
	.w2(32'h3a626ebc),
	.w3(32'hb87d8971),
	.w4(32'h3b1d50b2),
	.w5(32'hbab96945),
	.w6(32'hbb4c6205),
	.w7(32'hbb13bb05),
	.w8(32'hbb894ff5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440bdd),
	.w1(32'hbb1f169a),
	.w2(32'hbaf6407e),
	.w3(32'hbb86436e),
	.w4(32'hbb2016a7),
	.w5(32'hb90a1ed1),
	.w6(32'hb87d1f45),
	.w7(32'h39a35c23),
	.w8(32'hba4e2a42),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b72417),
	.w1(32'hba31739e),
	.w2(32'h38e2673a),
	.w3(32'hb7997aa2),
	.w4(32'h395da39b),
	.w5(32'hb98ce486),
	.w6(32'hba49b36e),
	.w7(32'hbb27fd40),
	.w8(32'h3a0883b3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9a145),
	.w1(32'h39fd4f33),
	.w2(32'hbb043d1b),
	.w3(32'hbaaa4471),
	.w4(32'hb9f44528),
	.w5(32'hbb0282ad),
	.w6(32'h3a51b9f1),
	.w7(32'hbad6e3d6),
	.w8(32'hbb929086),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5f4e),
	.w1(32'hbaaeb7b0),
	.w2(32'hb9f8998d),
	.w3(32'hbac6f380),
	.w4(32'hb9aec314),
	.w5(32'hba14ba51),
	.w6(32'hbb54c54d),
	.w7(32'hbb0e6a7b),
	.w8(32'hbad13fe1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9402f),
	.w1(32'hb9b0783f),
	.w2(32'hba92df94),
	.w3(32'hba368f2b),
	.w4(32'hba77fefb),
	.w5(32'hbb033bf5),
	.w6(32'hbadb1a1a),
	.w7(32'hba56f132),
	.w8(32'hbad2e744),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6df90),
	.w1(32'hba9d84b2),
	.w2(32'hba7e3fb9),
	.w3(32'hbb0096a2),
	.w4(32'hbab447a6),
	.w5(32'hba4b5558),
	.w6(32'hbaedd4db),
	.w7(32'hbaba4c89),
	.w8(32'h39dd4d3d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e44a5),
	.w1(32'hba3e59c6),
	.w2(32'hbb662760),
	.w3(32'h3ad2e9e1),
	.w4(32'hb9c3fedb),
	.w5(32'hbb04b405),
	.w6(32'h3b3f508e),
	.w7(32'h3b0e5e48),
	.w8(32'hbb4a38e6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87704d),
	.w1(32'h3ac82433),
	.w2(32'hba8b246f),
	.w3(32'h3b2fd3f8),
	.w4(32'h3aa9162e),
	.w5(32'hbb13dfa3),
	.w6(32'hbb9c27df),
	.w7(32'hbbb539be),
	.w8(32'hbbbbdb71),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0808bd),
	.w1(32'h395d37ce),
	.w2(32'hbb49e89d),
	.w3(32'h397b9119),
	.w4(32'hb95ccefe),
	.w5(32'hba3385c0),
	.w6(32'hbab2d564),
	.w7(32'hbb32c39a),
	.w8(32'hbb29f038),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0da8),
	.w1(32'h3a148834),
	.w2(32'h3a9d5604),
	.w3(32'h3b0cda5a),
	.w4(32'h3b2cedb0),
	.w5(32'hb9bafb34),
	.w6(32'hba8ae617),
	.w7(32'h3aa25bb2),
	.w8(32'hba68f35c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba430c37),
	.w1(32'hba99ea25),
	.w2(32'h3844ecfe),
	.w3(32'hb7d3fc99),
	.w4(32'hba8054f0),
	.w5(32'h3af14f0f),
	.w6(32'hb7cd99c9),
	.w7(32'hba166df6),
	.w8(32'h3b05db28),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17195),
	.w1(32'h3a701dbb),
	.w2(32'h3a97edb0),
	.w3(32'h3abca16f),
	.w4(32'h3b058191),
	.w5(32'hbab33a29),
	.w6(32'h3abdcf13),
	.w7(32'h3ade1a9b),
	.w8(32'hbab2d344),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e6347),
	.w1(32'hbb1dd20e),
	.w2(32'hbb4aec23),
	.w3(32'hbb015094),
	.w4(32'hbb0ccbce),
	.w5(32'hbb21724f),
	.w6(32'hbb411b6f),
	.w7(32'hbae6dc2b),
	.w8(32'hbba3c0d3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff27f3),
	.w1(32'hbaa104ba),
	.w2(32'hbae2c379),
	.w3(32'hbb46db13),
	.w4(32'hba47a6ea),
	.w5(32'h39c24066),
	.w6(32'hbc0537e5),
	.w7(32'hbbdc2867),
	.w8(32'hbb40ae63),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae94b19),
	.w1(32'h3a9d809b),
	.w2(32'hbae6f654),
	.w3(32'h39f2d348),
	.w4(32'h3ac9c69f),
	.w5(32'h3b3ba1ad),
	.w6(32'hbb8b786b),
	.w7(32'hbb5d3893),
	.w8(32'hbb0b18da),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7e197),
	.w1(32'h3b5b77d1),
	.w2(32'h3a766b23),
	.w3(32'h36a75999),
	.w4(32'h3b79cf91),
	.w5(32'h3ae839ca),
	.w6(32'hbb844fe4),
	.w7(32'hbb2465ad),
	.w8(32'hbbae1b73),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802ef94),
	.w1(32'h3a3254fa),
	.w2(32'hbb1d915c),
	.w3(32'hba2332f7),
	.w4(32'h3b247db9),
	.w5(32'h3b2c10fb),
	.w6(32'hbb99759d),
	.w7(32'hbb882c3f),
	.w8(32'hbb1c3dfd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffcd6f),
	.w1(32'hbb087500),
	.w2(32'hbb28cfcd),
	.w3(32'h399a79f4),
	.w4(32'hba8825de),
	.w5(32'hbc3bf3b8),
	.w6(32'hbb0fc4c5),
	.w7(32'hbb4eba2c),
	.w8(32'hbc25f9f8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb790982),
	.w1(32'hbb6d1c8f),
	.w2(32'hbb4b3671),
	.w3(32'hbb4a8f36),
	.w4(32'hbb22a98c),
	.w5(32'h3b25e010),
	.w6(32'hbb3b01a7),
	.w7(32'hbb584524),
	.w8(32'h3b27d270),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedab25),
	.w1(32'h3a7ec6c8),
	.w2(32'h3aba2dd8),
	.w3(32'h3b196907),
	.w4(32'h3b38a046),
	.w5(32'hba622fee),
	.w6(32'h3ad303ce),
	.w7(32'h3b092963),
	.w8(32'hbaee923a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62d69),
	.w1(32'h38744ef9),
	.w2(32'h3a185c01),
	.w3(32'hba2e9cef),
	.w4(32'hb72045b6),
	.w5(32'h3a6813ae),
	.w6(32'hba977ede),
	.w7(32'hb97c6e21),
	.w8(32'hb9a5c70d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ccb89),
	.w1(32'h39c0f0c5),
	.w2(32'h3a134d97),
	.w3(32'h39ca9050),
	.w4(32'hb97bdad5),
	.w5(32'hbb0f04a0),
	.w6(32'hbb718d44),
	.w7(32'hbb313f30),
	.w8(32'hbb848de5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c26d),
	.w1(32'hbb0bf963),
	.w2(32'hb9de19ed),
	.w3(32'hbb16e106),
	.w4(32'hba3cd191),
	.w5(32'hb7a3052e),
	.w6(32'hbb009d04),
	.w7(32'hba47ea2d),
	.w8(32'hba9abf89),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f0cb),
	.w1(32'hb93539dd),
	.w2(32'hbaeca266),
	.w3(32'hbb047036),
	.w4(32'hbb2391d2),
	.w5(32'hbb82d8cc),
	.w6(32'hbb52226c),
	.w7(32'hbb5a2757),
	.w8(32'hbb92a63b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc0270),
	.w1(32'hba9972ee),
	.w2(32'hbacb21de),
	.w3(32'hb943fe14),
	.w4(32'hb985c765),
	.w5(32'hbb3bf639),
	.w6(32'hbaa39cfa),
	.w7(32'hbac867b0),
	.w8(32'hbb2eea89),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8899051),
	.w1(32'hb95b15a1),
	.w2(32'hb980fd69),
	.w3(32'hbacd97ab),
	.w4(32'hba1681e9),
	.w5(32'h39f991d8),
	.w6(32'hbb177a3d),
	.w7(32'hbb0412a1),
	.w8(32'hb8e72a84),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f468a3),
	.w1(32'h38d66c57),
	.w2(32'hb9841315),
	.w3(32'h397b77a8),
	.w4(32'hb8948fa3),
	.w5(32'h37cd8246),
	.w6(32'hba909efe),
	.w7(32'hba120e17),
	.w8(32'h399e1002),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38305f04),
	.w1(32'hb8a1a202),
	.w2(32'hba1529f5),
	.w3(32'h3a42fdb4),
	.w4(32'hb9fe261d),
	.w5(32'h3b0e3787),
	.w6(32'hb7390483),
	.w7(32'hba95b4f5),
	.w8(32'h3ad81259),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba508c),
	.w1(32'h3a1d8f51),
	.w2(32'h3a725e5a),
	.w3(32'h3afe9fa1),
	.w4(32'h3b21dd33),
	.w5(32'h3a7acec2),
	.w6(32'h3a97cc98),
	.w7(32'h3adb829b),
	.w8(32'h3a159f6c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba9152),
	.w1(32'h39212495),
	.w2(32'h3a02fbea),
	.w3(32'h3af1e904),
	.w4(32'h3a943cb0),
	.w5(32'hbab37de3),
	.w6(32'h3aa0b469),
	.w7(32'h3ab4968f),
	.w8(32'hba9e18d9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2011b),
	.w1(32'hbac4ebfb),
	.w2(32'hbb1f782e),
	.w3(32'hbab7feb8),
	.w4(32'hba997669),
	.w5(32'hba671497),
	.w6(32'hbb0023a8),
	.w7(32'hbb236465),
	.w8(32'hba12e319),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1e5e),
	.w1(32'h3a5ab646),
	.w2(32'hb9d2d0e3),
	.w3(32'h39fbf608),
	.w4(32'hb97fab53),
	.w5(32'hbb27b726),
	.w6(32'hb847d3e4),
	.w7(32'hb98ae666),
	.w8(32'hbb93f7bd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89bd41),
	.w1(32'hbaddaeb3),
	.w2(32'hba76a77b),
	.w3(32'hbad02398),
	.w4(32'hb9457446),
	.w5(32'hba4969c8),
	.w6(32'h392d6482),
	.w7(32'h3a77416f),
	.w8(32'hba944ac4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34094f),
	.w1(32'hb979ffc7),
	.w2(32'hb9c30965),
	.w3(32'hb925eb59),
	.w4(32'hba33692a),
	.w5(32'hb9139bbb),
	.w6(32'hbafb447d),
	.w7(32'hbac30a7c),
	.w8(32'h3601e436),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9daa040),
	.w1(32'hb9212bc1),
	.w2(32'hba46ab2b),
	.w3(32'hb9e94779),
	.w4(32'h38bccbbd),
	.w5(32'hba944bf0),
	.w6(32'hbaa2437a),
	.w7(32'hb9baffea),
	.w8(32'hbb23230f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee298f),
	.w1(32'hbb0c683b),
	.w2(32'hba9823d0),
	.w3(32'hbaf0bfa7),
	.w4(32'hbaa7bfc6),
	.w5(32'h3a923c73),
	.w6(32'hba55969f),
	.w7(32'hba99936d),
	.w8(32'h3ada6e02),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92711f),
	.w1(32'h3a2e52fd),
	.w2(32'h3a8e0ad8),
	.w3(32'hbaa4d45a),
	.w4(32'hba9e08f3),
	.w5(32'hbb4803b1),
	.w6(32'hba5ed90b),
	.w7(32'hbaae3c88),
	.w8(32'hbb6550ca),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab502da),
	.w1(32'hbaa715e7),
	.w2(32'hbb5374f6),
	.w3(32'hba9da5bf),
	.w4(32'h3b264350),
	.w5(32'h3aa0bef3),
	.w6(32'hbbc75fc3),
	.w7(32'hbbb652f9),
	.w8(32'hbba6cd48),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dbc4c),
	.w1(32'h398c2377),
	.w2(32'hbb977a2f),
	.w3(32'h3a9d183b),
	.w4(32'hba1d2ae5),
	.w5(32'hbbbd2005),
	.w6(32'hbbc40bca),
	.w7(32'hbbc7926a),
	.w8(32'hbc2045f5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad138),
	.w1(32'h3b5521a8),
	.w2(32'hbabeac5e),
	.w3(32'hba966296),
	.w4(32'h3b4dde35),
	.w5(32'h3b2b0103),
	.w6(32'hbc1394fd),
	.w7(32'hbc020206),
	.w8(32'hbbda3521),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810867),
	.w1(32'hbb0a2564),
	.w2(32'hbb07c646),
	.w3(32'hba90a7e1),
	.w4(32'hbae9ab82),
	.w5(32'h3a3a4a28),
	.w6(32'hba042f8d),
	.w7(32'hba7c89d7),
	.w8(32'h3a7d05ec),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb688bcf9),
	.w1(32'hb964de52),
	.w2(32'h3a7613b9),
	.w3(32'hba0bf2d9),
	.w4(32'h3a06bef8),
	.w5(32'hbac867ce),
	.w6(32'h3968a0c6),
	.w7(32'h3a854f94),
	.w8(32'h39df0356),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9ff5f),
	.w1(32'h39c02ed0),
	.w2(32'hb8d4425f),
	.w3(32'hba0c0747),
	.w4(32'hb8c43dad),
	.w5(32'h3864db22),
	.w6(32'h3aa53b45),
	.w7(32'hba04fc94),
	.w8(32'hb9df2733),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8c797),
	.w1(32'hbb1a76fb),
	.w2(32'hbada68ca),
	.w3(32'h39fa71e1),
	.w4(32'hb937d787),
	.w5(32'hbabbb1cf),
	.w6(32'hba97f82c),
	.w7(32'hb9d7cd62),
	.w8(32'hbae64858),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0183f2),
	.w1(32'hba7cb6ec),
	.w2(32'hb9e4c02e),
	.w3(32'hb962b2ea),
	.w4(32'h38c3ad3f),
	.w5(32'hbb437bde),
	.w6(32'hb937a22a),
	.w7(32'hba17eb67),
	.w8(32'hbb50f9c0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab3bd),
	.w1(32'hbb2e59d6),
	.w2(32'hbb7b0b27),
	.w3(32'hbb8488c7),
	.w4(32'hbb9a9892),
	.w5(32'hbb8109db),
	.w6(32'hbb7c0331),
	.w7(32'hbb8aa650),
	.w8(32'hbaf2f3a5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28766a),
	.w1(32'hbb099e19),
	.w2(32'hbb0680f9),
	.w3(32'hba377b9e),
	.w4(32'hbab3e445),
	.w5(32'hbb674339),
	.w6(32'hbb5032b7),
	.w7(32'hbb9c2c21),
	.w8(32'hbbb321b2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45dd19),
	.w1(32'h38aa1b73),
	.w2(32'h3ad17111),
	.w3(32'hbaea7698),
	.w4(32'h3926ae53),
	.w5(32'h3b341916),
	.w6(32'hbba32886),
	.w7(32'hbb68e411),
	.w8(32'hbac1d263),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09fa0f),
	.w1(32'hb910630c),
	.w2(32'h3aa235d4),
	.w3(32'hbac39743),
	.w4(32'hba9f9375),
	.w5(32'hba561c17),
	.w6(32'hbb6082a5),
	.w7(32'hbb1bf6be),
	.w8(32'hbb149a5c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f68d9),
	.w1(32'hba3517d0),
	.w2(32'hbaa964d7),
	.w3(32'hba554ca0),
	.w4(32'h3a9b393a),
	.w5(32'h3ab8b1ef),
	.w6(32'hbab1fb8e),
	.w7(32'hbaf2b5e6),
	.w8(32'hba5421ba),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d646f),
	.w1(32'hbaf37176),
	.w2(32'hbaea5140),
	.w3(32'h3a1d04f3),
	.w4(32'h3aa12e1c),
	.w5(32'hbaa39819),
	.w6(32'hbb607c78),
	.w7(32'hbad2c66b),
	.w8(32'hbb40a10e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e177),
	.w1(32'hbb25bca9),
	.w2(32'hbaf98335),
	.w3(32'hbb317baf),
	.w4(32'hbb2414ac),
	.w5(32'hbb2f1968),
	.w6(32'hbb3e96fa),
	.w7(32'hbac1420d),
	.w8(32'hbb1d8c07),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba796508),
	.w1(32'h393f25b4),
	.w2(32'hba3af85d),
	.w3(32'h39518309),
	.w4(32'hba0e33bd),
	.w5(32'hba402eb8),
	.w6(32'h3a20b6d1),
	.w7(32'hba89933d),
	.w8(32'hba9fff8c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c81eb),
	.w1(32'hb8b4c479),
	.w2(32'hba493167),
	.w3(32'h39866926),
	.w4(32'hb98e8802),
	.w5(32'hb98ae675),
	.w6(32'h3a29346a),
	.w7(32'h3893036b),
	.w8(32'hba12fba0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a59c97),
	.w1(32'hba0f25c1),
	.w2(32'hba68c0b7),
	.w3(32'hba0c1e5e),
	.w4(32'hba828e46),
	.w5(32'hb8ad1ba3),
	.w6(32'h3a8d9837),
	.w7(32'hba0fc83a),
	.w8(32'hba1e15be),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf2602),
	.w1(32'hbaa5e26b),
	.w2(32'h39652189),
	.w3(32'h3521c5c8),
	.w4(32'hb92c580d),
	.w5(32'hb9070394),
	.w6(32'hb86c4b56),
	.w7(32'h3a1057b3),
	.w8(32'h3a9a5447),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc3dac),
	.w1(32'h3b329ff6),
	.w2(32'hbabed5f3),
	.w3(32'hba864abc),
	.w4(32'h3a0b14cc),
	.w5(32'hba2fc0dc),
	.w6(32'hbb385b71),
	.w7(32'hbb8d0747),
	.w8(32'hbb75fe19),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995fc60),
	.w1(32'hb9a8ce04),
	.w2(32'hba9770ff),
	.w3(32'h3917d829),
	.w4(32'h393cdda2),
	.w5(32'h3a39cdc3),
	.w6(32'hba1292e8),
	.w7(32'h3a01298d),
	.w8(32'hb8efb038),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5b1b),
	.w1(32'hb9b27142),
	.w2(32'hbadfeb70),
	.w3(32'hb9ae392e),
	.w4(32'h3ac19f58),
	.w5(32'hb85d4d19),
	.w6(32'hbb320a61),
	.w7(32'hbb04475e),
	.w8(32'hbb4e315e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ad05e),
	.w1(32'hba87ada3),
	.w2(32'hbb46b2a9),
	.w3(32'hbb36c5e5),
	.w4(32'hbb40f99d),
	.w5(32'hbb8c595b),
	.w6(32'hbc1644bd),
	.w7(32'hbbae36e1),
	.w8(32'hbbfb40e4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf27a1),
	.w1(32'h3ac31845),
	.w2(32'h3a9cc7f9),
	.w3(32'h3ac9d36e),
	.w4(32'h3acccb1d),
	.w5(32'hba84a7b6),
	.w6(32'h3a2cc523),
	.w7(32'h3795de8f),
	.w8(32'hbb4a4801),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf52ee),
	.w1(32'h3a983253),
	.w2(32'h3b0a3765),
	.w3(32'hba2bc9af),
	.w4(32'hba9685d5),
	.w5(32'hba9c4960),
	.w6(32'hbb3b46e5),
	.w7(32'hbb69e569),
	.w8(32'hbba22aa3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cdb90),
	.w1(32'hb9a6ff33),
	.w2(32'hba731ae3),
	.w3(32'hba6f6faa),
	.w4(32'h39da1e75),
	.w5(32'h3a82173d),
	.w6(32'hbb05f597),
	.w7(32'hbb08c96a),
	.w8(32'hba73ee58),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d90e9),
	.w1(32'h3ad6763c),
	.w2(32'hba380b73),
	.w3(32'h3a516a70),
	.w4(32'hba03bbd6),
	.w5(32'hba76389c),
	.w6(32'hbba60a1f),
	.w7(32'hbbbda08e),
	.w8(32'hbba8e02f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9dae8),
	.w1(32'hba408f7c),
	.w2(32'hbacf7757),
	.w3(32'h3984b63c),
	.w4(32'h39a7f8ce),
	.w5(32'hbaaf5812),
	.w6(32'hbb34c730),
	.w7(32'hbb16ebe1),
	.w8(32'hbb97a90f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ccb06),
	.w1(32'h393221b6),
	.w2(32'hb90f9539),
	.w3(32'h3935d376),
	.w4(32'h3a523da8),
	.w5(32'h3b22e251),
	.w6(32'hbbb1c68e),
	.w7(32'hbbb3996d),
	.w8(32'hb836c6f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab14380),
	.w1(32'h3b08fcf1),
	.w2(32'h3b03a18b),
	.w3(32'h3ab73879),
	.w4(32'h3a29295a),
	.w5(32'h3afe0a1a),
	.w6(32'h3a39b99e),
	.w7(32'h3ae264d4),
	.w8(32'h3afc415a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67e3c),
	.w1(32'h3ad2169d),
	.w2(32'hbabf926d),
	.w3(32'h371f3bd6),
	.w4(32'h39ae4e6c),
	.w5(32'hbaa45fea),
	.w6(32'hbaf839cc),
	.w7(32'hbb70bf0d),
	.w8(32'hbb90dcac),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21c35f),
	.w1(32'hba1e84d8),
	.w2(32'hbb048a2c),
	.w3(32'hba678884),
	.w4(32'hbb091aa3),
	.w5(32'hb74e7229),
	.w6(32'hba91dd9c),
	.w7(32'hbb777e45),
	.w8(32'hbb390cea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fbb72),
	.w1(32'hb9af086d),
	.w2(32'hbad58b89),
	.w3(32'hba60898f),
	.w4(32'hb9000863),
	.w5(32'hbbbc9066),
	.w6(32'hbb3911b3),
	.w7(32'hbacdc788),
	.w8(32'hbb894ba0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf3ce3),
	.w1(32'h3bb08771),
	.w2(32'hba868ab8),
	.w3(32'h3ba5bf62),
	.w4(32'h3b2c79ed),
	.w5(32'hbb5725be),
	.w6(32'hbb3b4b44),
	.w7(32'hbbad1f1b),
	.w8(32'hbc18d56e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986f1d3),
	.w1(32'h3b17fda7),
	.w2(32'h3a397409),
	.w3(32'hba891b4f),
	.w4(32'h3a7c487a),
	.w5(32'h3b2438a7),
	.w6(32'hbbd6b2bb),
	.w7(32'hbb8fb530),
	.w8(32'hbb3bf8ac),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad58d6),
	.w1(32'hbaac7112),
	.w2(32'hbb6de878),
	.w3(32'hbb08fd3a),
	.w4(32'hbb3aa3a3),
	.w5(32'hbb944e37),
	.w6(32'hbb507519),
	.w7(32'hbb6d4a23),
	.w8(32'hbb9ab5af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f7365),
	.w1(32'h3a0b072b),
	.w2(32'h39b548f3),
	.w3(32'h39e10d0f),
	.w4(32'h3a97857b),
	.w5(32'hbafcc90c),
	.w6(32'h3a028260),
	.w7(32'h3a9a412e),
	.w8(32'hbae684bb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d6b2),
	.w1(32'hbb4e25c0),
	.w2(32'hbbcbc582),
	.w3(32'hbb62c5f1),
	.w4(32'hbb9a6a6e),
	.w5(32'hbbfc18ee),
	.w6(32'hbb4d9648),
	.w7(32'hbbd6b580),
	.w8(32'hbba6b3f8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390745ad),
	.w1(32'h3a95d509),
	.w2(32'h3ab7cd91),
	.w3(32'hba1c7b66),
	.w4(32'hb9f187a0),
	.w5(32'h3a3e190b),
	.w6(32'hbabece36),
	.w7(32'hbadc4acb),
	.w8(32'hba9c66e6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc601a),
	.w1(32'hbaa5dfe7),
	.w2(32'h3aee4ef4),
	.w3(32'h39c23902),
	.w4(32'hb8f9a819),
	.w5(32'h3a64e81d),
	.w6(32'h3b048d6f),
	.w7(32'hb9598918),
	.w8(32'h3a9f03b8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e456fb),
	.w1(32'hbac5755a),
	.w2(32'hba199f80),
	.w3(32'h39b8f5a8),
	.w4(32'h39e59619),
	.w5(32'hba6e1a6f),
	.w6(32'hbac1a341),
	.w7(32'hba1dfeeb),
	.w8(32'hba50b2bf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855d36),
	.w1(32'h3a81e966),
	.w2(32'h395f9c85),
	.w3(32'hba81c269),
	.w4(32'hba1d26e2),
	.w5(32'h3ae3f787),
	.w6(32'hbae2d978),
	.w7(32'hbb3d93ff),
	.w8(32'hbb1b5830),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76cc21),
	.w1(32'h3ab31115),
	.w2(32'h3a6e0163),
	.w3(32'hb8d28390),
	.w4(32'h3b1bbcc1),
	.w5(32'h3ac9067d),
	.w6(32'hbb5150d4),
	.w7(32'hbac9ed44),
	.w8(32'hba042c5f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a803c34),
	.w1(32'hbacb27c1),
	.w2(32'hbb45c634),
	.w3(32'hb90fe96a),
	.w4(32'hbb061047),
	.w5(32'h3a2a2924),
	.w6(32'hba58161e),
	.w7(32'hbb43a834),
	.w8(32'hbb84f33c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9841477),
	.w1(32'h39e26282),
	.w2(32'hba11afb3),
	.w3(32'h3a82904c),
	.w4(32'h3a44306d),
	.w5(32'hba65fd68),
	.w6(32'hbaa66847),
	.w7(32'hba7933e2),
	.w8(32'hbb2dd559),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1029c),
	.w1(32'h3a215502),
	.w2(32'h3a29256b),
	.w3(32'hb9c25a95),
	.w4(32'hba15cc39),
	.w5(32'hb8836464),
	.w6(32'hbb1c1763),
	.w7(32'hbabfa216),
	.w8(32'hbb0fad02),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eb6f7),
	.w1(32'h3b011e74),
	.w2(32'hb9e81250),
	.w3(32'hb98d1a4b),
	.w4(32'h391ef61c),
	.w5(32'h388c432b),
	.w6(32'hbb3ea250),
	.w7(32'hbabf9764),
	.w8(32'hbb9a3b8c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a257f93),
	.w1(32'hbae4c6ba),
	.w2(32'hbaced86b),
	.w3(32'hb9b8e87f),
	.w4(32'h3ab0f4d0),
	.w5(32'h3b25b2c4),
	.w6(32'hbb78de67),
	.w7(32'hbb390d67),
	.w8(32'hbac3ab11),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cbd0c),
	.w1(32'hbaa2abf7),
	.w2(32'hba1131d9),
	.w3(32'h3a770494),
	.w4(32'h3a37d8b3),
	.w5(32'h3a9ff3fb),
	.w6(32'hb9eebc34),
	.w7(32'h39a85d49),
	.w8(32'h3ad99d6a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b154),
	.w1(32'h3b2b9ed3),
	.w2(32'h3af9e670),
	.w3(32'h3abb4f75),
	.w4(32'h3a5d9369),
	.w5(32'hba8d2c81),
	.w6(32'h3a963120),
	.w7(32'h3a392efa),
	.w8(32'hbab233d9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba410ca7),
	.w1(32'hb9a74771),
	.w2(32'hbadf4da0),
	.w3(32'hbac65488),
	.w4(32'hba000ac6),
	.w5(32'hb87a1148),
	.w6(32'hba3dd884),
	.w7(32'hbae55ab1),
	.w8(32'hba917638),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f61f1),
	.w1(32'hba8255e7),
	.w2(32'hba6e1c06),
	.w3(32'hba4741fd),
	.w4(32'hb936a6c1),
	.w5(32'hbb146e12),
	.w6(32'hba83cbf8),
	.w7(32'hb9c304ee),
	.w8(32'hbb1976f9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2ef8e),
	.w1(32'h3af0a4b0),
	.w2(32'hba325359),
	.w3(32'hba679974),
	.w4(32'hbaeeb501),
	.w5(32'h3b4c1445),
	.w6(32'hb9a2980e),
	.w7(32'hbb8704e1),
	.w8(32'hbb26668c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90e24d),
	.w1(32'h3ad4fd12),
	.w2(32'h3a36d05f),
	.w3(32'h3a22d9df),
	.w4(32'h3ac93599),
	.w5(32'h3a2418e9),
	.w6(32'hbaa2ccbc),
	.w7(32'h3abb3e22),
	.w8(32'h394e51bd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997eb69),
	.w1(32'hba4d176d),
	.w2(32'hbac09de9),
	.w3(32'h391fd0da),
	.w4(32'h3838b75e),
	.w5(32'hbadba0e5),
	.w6(32'hba4f4959),
	.w7(32'hba68187b),
	.w8(32'hbae6ae04),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add239a),
	.w1(32'h3b293f6f),
	.w2(32'h3aa07e89),
	.w3(32'hba122bcb),
	.w4(32'hba911ec6),
	.w5(32'hba3d005c),
	.w6(32'hbaf84092),
	.w7(32'hbb6875b2),
	.w8(32'hbb4eb870),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d72f4e),
	.w1(32'hba59f5c2),
	.w2(32'h39c4e084),
	.w3(32'hba4b2e2f),
	.w4(32'hbadb509c),
	.w5(32'hbad5d3af),
	.w6(32'hba704dde),
	.w7(32'h3a15439e),
	.w8(32'hba8f4d14),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c6c9a),
	.w1(32'h3a149fb8),
	.w2(32'hb9bb9e15),
	.w3(32'hbb0adccc),
	.w4(32'hba506bd8),
	.w5(32'h3989d376),
	.w6(32'hbad542d7),
	.w7(32'hbaa4e0e5),
	.w8(32'hbac754d0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba065340),
	.w1(32'hb801a931),
	.w2(32'h398f907e),
	.w3(32'h3a7926d5),
	.w4(32'hb9c5328f),
	.w5(32'h3acca9de),
	.w6(32'hb91a5e40),
	.w7(32'hb98e8a8f),
	.w8(32'h3aa28b9d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf40b),
	.w1(32'hb9a446c8),
	.w2(32'hbaa51ac3),
	.w3(32'h3a8d606f),
	.w4(32'hba6ecd38),
	.w5(32'h3aeccb31),
	.w6(32'h3978b068),
	.w7(32'hbaca1d06),
	.w8(32'h3ad1a210),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9003e),
	.w1(32'h3922a665),
	.w2(32'hba6ef5d7),
	.w3(32'hb74118d0),
	.w4(32'hb6259b5e),
	.w5(32'h38b7ec3a),
	.w6(32'hbb01ad8a),
	.w7(32'hbb063980),
	.w8(32'hbb1e5505),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf14ab),
	.w1(32'h3a8197f1),
	.w2(32'h3b0ce99a),
	.w3(32'hb9a4f9bd),
	.w4(32'h3ac283e4),
	.w5(32'h3900971b),
	.w6(32'hbb56a72e),
	.w7(32'hbadba72c),
	.w8(32'hba7d2872),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976a840),
	.w1(32'hb71e206a),
	.w2(32'hb96e8599),
	.w3(32'hba0d2a7a),
	.w4(32'hbaa91409),
	.w5(32'hbabbe0c2),
	.w6(32'hb9e90448),
	.w7(32'h3843ab80),
	.w8(32'hb7488566),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92514a1),
	.w1(32'hba200f8a),
	.w2(32'hbac94972),
	.w3(32'h3a529c4f),
	.w4(32'hb9058d2a),
	.w5(32'hbaf38abc),
	.w6(32'hbadcad86),
	.w7(32'hba212f27),
	.w8(32'hba9b1ff5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b03b86),
	.w1(32'hb907d1a3),
	.w2(32'hbac969b7),
	.w3(32'hba7ca1f2),
	.w4(32'hbaa1dbb7),
	.w5(32'hba1dc59a),
	.w6(32'h3985f8e8),
	.w7(32'hbad32111),
	.w8(32'hb88f0b1a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01964b),
	.w1(32'hba42a856),
	.w2(32'hba98eada),
	.w3(32'hbaa22c47),
	.w4(32'h3a185fd8),
	.w5(32'hb9e2dd7f),
	.w6(32'hbb0329c8),
	.w7(32'hba4ebb37),
	.w8(32'hbae7622c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccb500),
	.w1(32'h3a86588b),
	.w2(32'h3a6bb6a4),
	.w3(32'hbb03a9f1),
	.w4(32'h398d9d8c),
	.w5(32'h3ab7be38),
	.w6(32'hbb34a208),
	.w7(32'hba4a2923),
	.w8(32'h3a5737e2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d4090),
	.w1(32'hb921cd8c),
	.w2(32'hbb013fe4),
	.w3(32'hbacd6011),
	.w4(32'hbb4be0f0),
	.w5(32'hbb8dd7f3),
	.w6(32'hbb65e656),
	.w7(32'hbb98c69b),
	.w8(32'hbba2eddd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf70c4),
	.w1(32'h3acd92cf),
	.w2(32'hb9be12c7),
	.w3(32'h3a25465e),
	.w4(32'h3b04a5b9),
	.w5(32'h3ae705b5),
	.w6(32'hba851dbc),
	.w7(32'hbb10f99a),
	.w8(32'hbafa25e4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfd0db),
	.w1(32'h39458fa7),
	.w2(32'h39c30068),
	.w3(32'hba0b736b),
	.w4(32'hba4e9a22),
	.w5(32'hba8adb95),
	.w6(32'hbb40bf05),
	.w7(32'hbb4e0101),
	.w8(32'hbb35eccd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ae99e),
	.w1(32'hba78a70c),
	.w2(32'hbb2846ce),
	.w3(32'hbad3cb51),
	.w4(32'hbb3cd893),
	.w5(32'hbb76402c),
	.w6(32'hbb56e884),
	.w7(32'hbb525d66),
	.w8(32'hbb462b64),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33edb5),
	.w1(32'h3a4680d3),
	.w2(32'hbae69112),
	.w3(32'hba02144f),
	.w4(32'hb9818545),
	.w5(32'h3a1f17f6),
	.w6(32'hbb252683),
	.w7(32'hbb670f1f),
	.w8(32'hbae08ddd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b2877),
	.w1(32'h39fb344c),
	.w2(32'hbae3643b),
	.w3(32'hb9fbc6da),
	.w4(32'hb9bc62a1),
	.w5(32'hbb1f25ff),
	.w6(32'hbb378b86),
	.w7(32'hbaf60047),
	.w8(32'hbb95c46e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba064089),
	.w1(32'h3a25ed90),
	.w2(32'hb88e4f3b),
	.w3(32'hbb046261),
	.w4(32'hbb4db912),
	.w5(32'hb8b6596a),
	.w6(32'hbb0d8e24),
	.w7(32'hbb299b1d),
	.w8(32'hbaa721ba),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac14866),
	.w1(32'h3a3fd145),
	.w2(32'h3a9c8cc1),
	.w3(32'h39232949),
	.w4(32'h3b2b8d24),
	.w5(32'hba0b7667),
	.w6(32'hbb46b37d),
	.w7(32'hbacb1901),
	.w8(32'hbb5b70b6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee5eaa),
	.w1(32'hbac08928),
	.w2(32'hbb3e3467),
	.w3(32'hbb0762c9),
	.w4(32'hbb6419fb),
	.w5(32'hbb6e877f),
	.w6(32'hba596325),
	.w7(32'hbb58228c),
	.w8(32'hbb7c845a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39d474),
	.w1(32'hba8b0008),
	.w2(32'hba77e746),
	.w3(32'hba762257),
	.w4(32'hba79e6f4),
	.w5(32'hba2789b4),
	.w6(32'hbaab92cd),
	.w7(32'hbab082bc),
	.w8(32'hba0295b3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad4b27),
	.w1(32'hbabf08a8),
	.w2(32'hba66b0a7),
	.w3(32'h384d298c),
	.w4(32'hbac0a151),
	.w5(32'hb912e77d),
	.w6(32'hbab92c0c),
	.w7(32'hba2dd08c),
	.w8(32'hb9d94f5c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38043e),
	.w1(32'h3a525774),
	.w2(32'hb97f8cb1),
	.w3(32'hba48117b),
	.w4(32'h3950aa11),
	.w5(32'h3b4e5b25),
	.w6(32'hbacc47b0),
	.w7(32'hbabda1a4),
	.w8(32'h3b099aee),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a51f),
	.w1(32'h3b24b160),
	.w2(32'h39bf6519),
	.w3(32'h3b8a4fc9),
	.w4(32'h3ba5dbbc),
	.w5(32'hb8399486),
	.w6(32'h3afc8fb0),
	.w7(32'h3a649c76),
	.w8(32'hbb3aae26),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9911dea),
	.w1(32'h3abef736),
	.w2(32'h3ad06ab1),
	.w3(32'hba976615),
	.w4(32'hb9f764e3),
	.w5(32'h3aa6ebb5),
	.w6(32'hbb61636b),
	.w7(32'hbb7aa980),
	.w8(32'hbaae4900),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a106808),
	.w1(32'hb8ed49cd),
	.w2(32'hba2aef83),
	.w3(32'h3a151b3c),
	.w4(32'hb98a7be5),
	.w5(32'h3a37e139),
	.w6(32'h3a5ebfbd),
	.w7(32'hb7ab6111),
	.w8(32'h3a81df5c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc4b62),
	.w1(32'h3b42ad24),
	.w2(32'h3ac491ef),
	.w3(32'hb9ed1099),
	.w4(32'h3a876aed),
	.w5(32'h39984bac),
	.w6(32'hbb0e7b17),
	.w7(32'hbaf9ddf6),
	.w8(32'hbb4cf7ac),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960f7a9),
	.w1(32'h39a10412),
	.w2(32'hb9815de6),
	.w3(32'hbac5c897),
	.w4(32'h39e25181),
	.w5(32'h3924c065),
	.w6(32'hbb3ddb12),
	.w7(32'hbb49d913),
	.w8(32'hbac791ab),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb92b7),
	.w1(32'hbb147b87),
	.w2(32'hbb2aa105),
	.w3(32'hbb436f06),
	.w4(32'hbb0ffc2c),
	.w5(32'hbb1099a1),
	.w6(32'hbb10c22c),
	.w7(32'hbb6ab494),
	.w8(32'hbb391b02),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15e7db),
	.w1(32'h3ab6fc0d),
	.w2(32'h3a7826dc),
	.w3(32'h3b2a203c),
	.w4(32'h3b0b4960),
	.w5(32'h3a829405),
	.w6(32'hbaddb0fb),
	.w7(32'h3a56b72b),
	.w8(32'hbb104ae1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9768870),
	.w1(32'hba70c63e),
	.w2(32'hbac4ad6f),
	.w3(32'hba6368d3),
	.w4(32'hbb083e67),
	.w5(32'hbb013035),
	.w6(32'hba86df0b),
	.w7(32'hbb387e1c),
	.w8(32'hba95dba4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a7482),
	.w1(32'h3a2b7a88),
	.w2(32'hb9be5fee),
	.w3(32'h39d3a0e3),
	.w4(32'hba010162),
	.w5(32'h3a7387d5),
	.w6(32'h3ac5add2),
	.w7(32'h38b95e95),
	.w8(32'hb8a53c21),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3e8a9),
	.w1(32'h39c2c310),
	.w2(32'h39f0c47b),
	.w3(32'h3a9e8348),
	.w4(32'h3b00c115),
	.w5(32'hba2e59ff),
	.w6(32'hbb1d8594),
	.w7(32'hba411396),
	.w8(32'hbaefcfeb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad36fda),
	.w1(32'hba6a7b60),
	.w2(32'hbaf6d6ec),
	.w3(32'hba16a999),
	.w4(32'hbac6118f),
	.w5(32'hbad2f5a4),
	.w6(32'hbb49d15d),
	.w7(32'hbb4b5660),
	.w8(32'hbb12076e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b04e1),
	.w1(32'hba1e65ae),
	.w2(32'h37b117d8),
	.w3(32'h3a53346b),
	.w4(32'h3ac89ec2),
	.w5(32'hb9e0c1e8),
	.w6(32'hb9f7e6cc),
	.w7(32'h3ab65966),
	.w8(32'hbb0b5fca),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30acea),
	.w1(32'hba936548),
	.w2(32'hba88b910),
	.w3(32'hbaa26cbd),
	.w4(32'hba5e527c),
	.w5(32'hba338693),
	.w6(32'hbabd9de0),
	.w7(32'hbb436276),
	.w8(32'hba30ab4d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39926283),
	.w1(32'h39f0fc52),
	.w2(32'h37ef3423),
	.w3(32'hb9caef39),
	.w4(32'h39ae7859),
	.w5(32'h3b1571fb),
	.w6(32'hb98592c5),
	.w7(32'h3a21d73c),
	.w8(32'h3991c1f9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bf18f),
	.w1(32'h3a628405),
	.w2(32'h3afd3978),
	.w3(32'h3ab57d8e),
	.w4(32'h39da51d5),
	.w5(32'hbae86aac),
	.w6(32'hbb224d4f),
	.w7(32'hbaf60369),
	.w8(32'hbb50fec4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc4779),
	.w1(32'h398cd37a),
	.w2(32'h3908b68b),
	.w3(32'hba651bcd),
	.w4(32'hba6f5bdb),
	.w5(32'h396bfbeb),
	.w6(32'h3956f23a),
	.w7(32'hba005d0b),
	.w8(32'hb94f79d5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5058e),
	.w1(32'h3a2c0a04),
	.w2(32'hba102203),
	.w3(32'h3a314afb),
	.w4(32'h3a490303),
	.w5(32'h3b14f25b),
	.w6(32'hbaa74e6e),
	.w7(32'hbab6d121),
	.w8(32'h39767288),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38559468),
	.w1(32'h398a42ff),
	.w2(32'h38941e08),
	.w3(32'h38b756f1),
	.w4(32'h3963c8dc),
	.w5(32'h3a01a373),
	.w6(32'h3a30e7be),
	.w7(32'h3a47bb5c),
	.w8(32'hbb0bb599),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cc448),
	.w1(32'h3ae860b9),
	.w2(32'h3a1dd538),
	.w3(32'hba8f55fc),
	.w4(32'hb9e8ec45),
	.w5(32'hbb01cbd9),
	.w6(32'hba96a9c3),
	.w7(32'h3723f61d),
	.w8(32'hb8bb6b27),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0c8da),
	.w1(32'h3b161ee9),
	.w2(32'hb984838e),
	.w3(32'h3aa67bb2),
	.w4(32'hba2408a3),
	.w5(32'hba964175),
	.w6(32'h3b0e38c3),
	.w7(32'hb6d14686),
	.w8(32'hbac88a46),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13afb0),
	.w1(32'h39cf11ee),
	.w2(32'h3a030147),
	.w3(32'hba705482),
	.w4(32'hbabb90fa),
	.w5(32'h3b26ef66),
	.w6(32'hba0751ed),
	.w7(32'h381ca807),
	.w8(32'h3b527f51),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb05a39),
	.w1(32'h3b0705b8),
	.w2(32'h3a4f9ea2),
	.w3(32'h3b413bc3),
	.w4(32'h3b7aac3c),
	.w5(32'hb90949a9),
	.w6(32'h3a0314d3),
	.w7(32'h3a1fea5f),
	.w8(32'hbb027bb4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194d0d),
	.w1(32'h3a3c2f26),
	.w2(32'hba87d3ac),
	.w3(32'h3a89e5d1),
	.w4(32'h3b11f828),
	.w5(32'hbaf6c666),
	.w6(32'hbb8a4a28),
	.w7(32'hbb633eb7),
	.w8(32'hbb9fedbe),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7457a),
	.w1(32'hba39eb88),
	.w2(32'hbaeb6a85),
	.w3(32'h391fe634),
	.w4(32'hbaab822d),
	.w5(32'hb9e5ee87),
	.w6(32'h3901c73d),
	.w7(32'hba20f3bb),
	.w8(32'hb8b3ca01),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144ad5),
	.w1(32'h3af26bb1),
	.w2(32'hba36902e),
	.w3(32'hb96e14a7),
	.w4(32'h3a84ba72),
	.w5(32'hbab7dd97),
	.w6(32'hbb22c75a),
	.w7(32'hbb668c2d),
	.w8(32'hbb7edb1f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f462),
	.w1(32'hbb5c8845),
	.w2(32'hbb00403f),
	.w3(32'hbb50d87d),
	.w4(32'hbb43b133),
	.w5(32'h3ab5750e),
	.w6(32'hbb17ed80),
	.w7(32'hbae3803d),
	.w8(32'hb9176321),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeef74),
	.w1(32'h3ad41a9b),
	.w2(32'h3a869d11),
	.w3(32'hb946bc36),
	.w4(32'h38df52e7),
	.w5(32'hbb04d733),
	.w6(32'hbb80f61d),
	.w7(32'hbb910df1),
	.w8(32'hbba2442e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab95b96),
	.w1(32'hba9ef7cd),
	.w2(32'hbb41b297),
	.w3(32'hba6fffd1),
	.w4(32'hbabf2247),
	.w5(32'hb9f1d649),
	.w6(32'hbb99810a),
	.w7(32'hbbc45da0),
	.w8(32'hbaee0398),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52778),
	.w1(32'h3a976c56),
	.w2(32'h38e21a8c),
	.w3(32'hb91b200e),
	.w4(32'hbaba09e7),
	.w5(32'hbb133a90),
	.w6(32'hba649a87),
	.w7(32'hbb226c0e),
	.w8(32'hbb08c6b3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff02e4),
	.w1(32'h3b024de7),
	.w2(32'h3b05c9de),
	.w3(32'hba5e5f19),
	.w4(32'hbaa59ddd),
	.w5(32'hbaf3fe4f),
	.w6(32'hb9caf2f2),
	.w7(32'h39e5d6eb),
	.w8(32'hbb01b886),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45610a),
	.w1(32'hba09a029),
	.w2(32'hbadfc386),
	.w3(32'hbb1c01f0),
	.w4(32'hbb5b9c28),
	.w5(32'hb9a5eb49),
	.w6(32'hbb145607),
	.w7(32'hbb60c711),
	.w8(32'hba824a7d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c24a),
	.w1(32'h3b1d1a38),
	.w2(32'h3a8c6572),
	.w3(32'h3a9e1a02),
	.w4(32'h3937d05b),
	.w5(32'h3ae6da80),
	.w6(32'h3ae077ba),
	.w7(32'h3a5cc5f5),
	.w8(32'h3a77de63),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b01da),
	.w1(32'hbae84219),
	.w2(32'h3ae9d390),
	.w3(32'hba6cea79),
	.w4(32'h3b0873fb),
	.w5(32'hbaaf6cf6),
	.w6(32'hbaeefe4f),
	.w7(32'h3b1e7834),
	.w8(32'hbb07933d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf648e),
	.w1(32'hba5fc789),
	.w2(32'hba9d10b8),
	.w3(32'hbb2ef69f),
	.w4(32'h394b971f),
	.w5(32'hb7c5de0d),
	.w6(32'hb60dee75),
	.w7(32'hbaa7332e),
	.w8(32'hba89f375),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd7550),
	.w1(32'h3a2c09c2),
	.w2(32'hba2ad000),
	.w3(32'hbae21b65),
	.w4(32'h393200c1),
	.w5(32'hbafb4ba2),
	.w6(32'hbaff105e),
	.w7(32'hbaf2232a),
	.w8(32'hbb340d01),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999f7e0),
	.w1(32'hbad0a87d),
	.w2(32'hba0043fa),
	.w3(32'hb9bb2d65),
	.w4(32'hb92f0ad2),
	.w5(32'h3a95ea46),
	.w6(32'hbaee21fc),
	.w7(32'hba2f378c),
	.w8(32'h3a3a8ad5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62a7a2),
	.w1(32'h3a4fa00f),
	.w2(32'h39ef9877),
	.w3(32'h3a2b4af0),
	.w4(32'hb90ae066),
	.w5(32'h3a1ee18a),
	.w6(32'hba1a41d5),
	.w7(32'hb9d3ff67),
	.w8(32'h3a5761f5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109ed2),
	.w1(32'hb9285030),
	.w2(32'hbae7ebe6),
	.w3(32'h3af999c1),
	.w4(32'h3addd528),
	.w5(32'hba38045e),
	.w6(32'hbaaba41d),
	.w7(32'hba8a991f),
	.w8(32'hba3aa7ee),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47018),
	.w1(32'h3a292fe4),
	.w2(32'hb9dc143c),
	.w3(32'h3a8e313d),
	.w4(32'h3a9fcf82),
	.w5(32'hb9c95cd9),
	.w6(32'hbb28663f),
	.w7(32'hbb8cbc42),
	.w8(32'hbb87b07b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900869d),
	.w1(32'hbaa97851),
	.w2(32'h399482e4),
	.w3(32'hb98760a0),
	.w4(32'h39875c3d),
	.w5(32'h3a1b805a),
	.w6(32'hba8c8d14),
	.w7(32'h3a05fbd3),
	.w8(32'h3aa286f7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab81c63),
	.w1(32'h3b25707e),
	.w2(32'h3a877d16),
	.w3(32'h3aa1b683),
	.w4(32'hb9ba393d),
	.w5(32'hb9ec5f76),
	.w6(32'h3abe90d4),
	.w7(32'h39c98b5b),
	.w8(32'hbad27e53),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac30a6b),
	.w1(32'h3bccad0e),
	.w2(32'h3ba32194),
	.w3(32'hbad1698c),
	.w4(32'h3b735342),
	.w5(32'h3a260b06),
	.w6(32'hbb709a2d),
	.w7(32'hba4d9065),
	.w8(32'hbb2f0f99),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2251c8),
	.w1(32'h3aa62870),
	.w2(32'hba9d82f3),
	.w3(32'h3a688b88),
	.w4(32'h39ba007c),
	.w5(32'hba8f60a8),
	.w6(32'hbb8c34a4),
	.w7(32'hbb58fee8),
	.w8(32'hbba78d0b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3f1c8),
	.w1(32'hbaaface7),
	.w2(32'hbaf29c87),
	.w3(32'hb79b2c93),
	.w4(32'hba7cfe59),
	.w5(32'h392bd352),
	.w6(32'h3796da38),
	.w7(32'hbb070534),
	.w8(32'h394729a7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54a86c),
	.w1(32'h3a560569),
	.w2(32'h3a1136ef),
	.w3(32'h390cd031),
	.w4(32'h3a31e3ba),
	.w5(32'hb92a9e04),
	.w6(32'hb9f6d8a9),
	.w7(32'h39a6070a),
	.w8(32'h3a3696e8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a630e37),
	.w1(32'hba09fdbd),
	.w2(32'h3950ea22),
	.w3(32'h3998c2ff),
	.w4(32'hb7befd1b),
	.w5(32'h3a883579),
	.w6(32'h39dcf4b6),
	.w7(32'h3944a388),
	.w8(32'h3ad3990a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafd38c),
	.w1(32'h39abe07a),
	.w2(32'h39905284),
	.w3(32'h3a724ebf),
	.w4(32'h3a263eee),
	.w5(32'h3a1faa45),
	.w6(32'h3a11b4f5),
	.w7(32'hb9b9e520),
	.w8(32'hba1be19d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c966a),
	.w1(32'h3a467d84),
	.w2(32'hba164410),
	.w3(32'hb93fbd62),
	.w4(32'h39fae515),
	.w5(32'hb94d8c89),
	.w6(32'hbab6eb03),
	.w7(32'hba288cf5),
	.w8(32'hbaf32a9c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb4545),
	.w1(32'hb911159d),
	.w2(32'hbb2de9d6),
	.w3(32'h3ab0a54a),
	.w4(32'h39d078b4),
	.w5(32'hbb1ff918),
	.w6(32'hbb0cc33f),
	.w7(32'hbb4d8e1e),
	.w8(32'hbb64546b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947e97),
	.w1(32'h3b68e28e),
	.w2(32'h3adb776c),
	.w3(32'h39a72232),
	.w4(32'h39f0dcb3),
	.w5(32'h3bb620be),
	.w6(32'hba09b0b9),
	.w7(32'hbae72535),
	.w8(32'h3acc3415),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af836f9),
	.w1(32'hba829d5a),
	.w2(32'hba79207b),
	.w3(32'h39f59f54),
	.w4(32'hb8ff054d),
	.w5(32'h3b196d9d),
	.w6(32'hb9964ebe),
	.w7(32'hba9551b7),
	.w8(32'h3a815e94),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8631a),
	.w1(32'h3b3a6fbf),
	.w2(32'h3aedc0ea),
	.w3(32'h3a809228),
	.w4(32'h3a7f4fda),
	.w5(32'h3a7f5438),
	.w6(32'hbb19e5e6),
	.w7(32'hbb011685),
	.w8(32'hbb14b299),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2432ad),
	.w1(32'h3aae32e8),
	.w2(32'h391ccd6e),
	.w3(32'h385fc648),
	.w4(32'hbad21152),
	.w5(32'hb81902d7),
	.w6(32'h3ae7faa3),
	.w7(32'hbaafe015),
	.w8(32'hbac52564),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900bb6f),
	.w1(32'hb9c07d79),
	.w2(32'h396a4ad7),
	.w3(32'h3a17e3a2),
	.w4(32'hb940148f),
	.w5(32'h3a2ac2d9),
	.w6(32'h3ab0f2f0),
	.w7(32'h3a9932be),
	.w8(32'h395c5ee9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b5720),
	.w1(32'h3a0fca82),
	.w2(32'hba31b624),
	.w3(32'hb982cefe),
	.w4(32'hba1b7fe7),
	.w5(32'hb8da71a6),
	.w6(32'h3a114b8b),
	.w7(32'hb8be516c),
	.w8(32'hb9dde014),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0bb19),
	.w1(32'h399354a1),
	.w2(32'h37ea6f54),
	.w3(32'hb9b36e40),
	.w4(32'hb9a6f393),
	.w5(32'hb8c284b6),
	.w6(32'hba9f4e0a),
	.w7(32'hb9802fe5),
	.w8(32'hbab08a1f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905d62c),
	.w1(32'h3a9c17d2),
	.w2(32'hb9e8333e),
	.w3(32'h3a0c435d),
	.w4(32'hb84389f0),
	.w5(32'hba53f47b),
	.w6(32'hbb7bf266),
	.w7(32'hbb70264e),
	.w8(32'hbb2be4e8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af39976),
	.w1(32'h3a988577),
	.w2(32'hba2c553e),
	.w3(32'hbaa57495),
	.w4(32'hb9bbdc10),
	.w5(32'hba99132c),
	.w6(32'hbb53088d),
	.w7(32'hbae886b2),
	.w8(32'hbb821043),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a671cbc),
	.w1(32'h3a7986a2),
	.w2(32'h39c6ddbb),
	.w3(32'hba370bb1),
	.w4(32'h3a284693),
	.w5(32'h3ad04d8d),
	.w6(32'hbb83fb0a),
	.w7(32'hbb3a8620),
	.w8(32'hbb3d8da6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a29d65),
	.w1(32'hb8fd49a2),
	.w2(32'h3981cd38),
	.w3(32'h3a0dc7e3),
	.w4(32'h399ed931),
	.w5(32'hbb6795b6),
	.w6(32'h3a60af74),
	.w7(32'h395882d4),
	.w8(32'hbb33610f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5eeb4),
	.w1(32'hba9c40e1),
	.w2(32'hbb9a71ec),
	.w3(32'hba8c0add),
	.w4(32'hba26bd55),
	.w5(32'h37e40988),
	.w6(32'hbaf25b88),
	.w7(32'hbba25b3f),
	.w8(32'hbba0e258),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8839ae),
	.w1(32'hb9ce6685),
	.w2(32'hba052966),
	.w3(32'hbb11a073),
	.w4(32'hba6b0c2f),
	.w5(32'hb825f1a8),
	.w6(32'hbb77fe8a),
	.w7(32'hbb1358e4),
	.w8(32'h392c680e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae971d7),
	.w1(32'h3b319c75),
	.w2(32'h3b0cba08),
	.w3(32'hbaf97eef),
	.w4(32'hba03fa80),
	.w5(32'h3b044d17),
	.w6(32'hbb3b368c),
	.w7(32'hbb4dba8c),
	.w8(32'hbb715466),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dcb55),
	.w1(32'hba10b87f),
	.w2(32'hba4bdad8),
	.w3(32'hba86a0f1),
	.w4(32'hba40796f),
	.w5(32'h3a5cc2f7),
	.w6(32'hba69f652),
	.w7(32'hba6bd562),
	.w8(32'h3a8fbf1e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae85d74),
	.w1(32'hb8f349d5),
	.w2(32'h39ff9fb2),
	.w3(32'hb910e9aa),
	.w4(32'hb9f1712a),
	.w5(32'hbb0a5308),
	.w6(32'h398a8ec1),
	.w7(32'h3a0db136),
	.w8(32'hba482244),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17bc10),
	.w1(32'hbaf95436),
	.w2(32'hbb316470),
	.w3(32'hbb439038),
	.w4(32'hbb15d4d2),
	.w5(32'h3b0d6014),
	.w6(32'hbbc13113),
	.w7(32'hbbe430c2),
	.w8(32'hbb2b33e5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f2937),
	.w1(32'h3b221abb),
	.w2(32'hbb203516),
	.w3(32'h3ab8d476),
	.w4(32'h3b660311),
	.w5(32'hbaa527e7),
	.w6(32'hbbac4df3),
	.w7(32'hbbc2f94a),
	.w8(32'hbbdc95eb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebee9f),
	.w1(32'hbac379ad),
	.w2(32'hbb29f405),
	.w3(32'hbad213b9),
	.w4(32'h3a9572b3),
	.w5(32'h3a98ad0c),
	.w6(32'hbba67384),
	.w7(32'hbbb90fd3),
	.w8(32'hbb379fae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f12312),
	.w1(32'hbb07a5a4),
	.w2(32'hba9de161),
	.w3(32'hba013904),
	.w4(32'hbb2e677f),
	.w5(32'hbab01baf),
	.w6(32'hba0d36e5),
	.w7(32'hba4a9c3c),
	.w8(32'hba81e35c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab9780),
	.w1(32'h3a8198f1),
	.w2(32'h3a7a3a8a),
	.w3(32'hb9a2f095),
	.w4(32'hb8f55670),
	.w5(32'h382099f7),
	.w6(32'hb92558fc),
	.w7(32'h39bc18e9),
	.w8(32'hb9c81312),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9861ca1),
	.w1(32'h38a409ad),
	.w2(32'h389e1271),
	.w3(32'hb7977c75),
	.w4(32'hba66946f),
	.w5(32'h3ac7bd3d),
	.w6(32'hb9de5201),
	.w7(32'hb9f57f52),
	.w8(32'h3a60c5ad),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364bff66),
	.w1(32'hb9e8d51a),
	.w2(32'h3abe8200),
	.w3(32'h3aa69951),
	.w4(32'h3a9cb682),
	.w5(32'hbaf998e6),
	.w6(32'h391f0159),
	.w7(32'h3b0a9144),
	.w8(32'h3a3dd3d6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c062a),
	.w1(32'h393cdfe5),
	.w2(32'hbb19cedb),
	.w3(32'hbb4c6e3b),
	.w4(32'hb8b250e6),
	.w5(32'h398eaa90),
	.w6(32'hbb8bc519),
	.w7(32'hbb1f7a3a),
	.w8(32'hbafdf6d9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9fe12),
	.w1(32'hbb27259e),
	.w2(32'hbb2c75dd),
	.w3(32'hba3cfdab),
	.w4(32'hba90c511),
	.w5(32'hbbaaa672),
	.w6(32'hbb06e0f5),
	.w7(32'hbb292d35),
	.w8(32'hbb80c617),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb782),
	.w1(32'hbb05f06d),
	.w2(32'hbb172f7b),
	.w3(32'hba3bfb69),
	.w4(32'hba055e93),
	.w5(32'hb9b80c8f),
	.w6(32'hbb86f7e2),
	.w7(32'hba1c624b),
	.w8(32'hbaac05bb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab026fb),
	.w1(32'h39580799),
	.w2(32'hbaf14ad4),
	.w3(32'h3ab011db),
	.w4(32'h3abfc4d1),
	.w5(32'h3aa33d02),
	.w6(32'hba4ffe05),
	.w7(32'hb9e057e4),
	.w8(32'hbb0fb365),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bf07f),
	.w1(32'h3a81c102),
	.w2(32'h3a0954e1),
	.w3(32'h3aa7390b),
	.w4(32'h3a0286f7),
	.w5(32'hba507758),
	.w6(32'h3a297307),
	.w7(32'h3933a26c),
	.w8(32'h3ab7e9ff),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8667c6),
	.w1(32'h3b4d81de),
	.w2(32'h3aedbacf),
	.w3(32'hb8b26be8),
	.w4(32'hba82715a),
	.w5(32'hba8042e2),
	.w6(32'h3bb2e734),
	.w7(32'h3b1d072f),
	.w8(32'hb994d924),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b92b7),
	.w1(32'hba28798b),
	.w2(32'hbad837cf),
	.w3(32'hba1c845a),
	.w4(32'h39d5cb4a),
	.w5(32'h3a57f02c),
	.w6(32'h39e890ac),
	.w7(32'h38e7d5eb),
	.w8(32'h3a14028b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8159a90),
	.w1(32'hba517c17),
	.w2(32'h3a3683d8),
	.w3(32'hb9e00ca9),
	.w4(32'hb8a75676),
	.w5(32'h3aba154e),
	.w6(32'hb8834c45),
	.w7(32'h3a857e42),
	.w8(32'h3a8d9df7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3e57),
	.w1(32'hbb390334),
	.w2(32'hbba2971c),
	.w3(32'hbb8e4cb0),
	.w4(32'hbb222cd3),
	.w5(32'hbbc09839),
	.w6(32'hbb827ecf),
	.w7(32'hbbf95a43),
	.w8(32'hbbd0f556),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b6755),
	.w1(32'h3ac9d2d2),
	.w2(32'h3c3088cb),
	.w3(32'hbb162a16),
	.w4(32'h3c35edba),
	.w5(32'hbbb0f8b2),
	.w6(32'hbc3e97ac),
	.w7(32'h3c8b636d),
	.w8(32'hbb81fa76),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f48e),
	.w1(32'hbb59196c),
	.w2(32'hbbb60d0a),
	.w3(32'hb9bb64bb),
	.w4(32'hbb9096d6),
	.w5(32'hbacb6be7),
	.w6(32'h3aed5c37),
	.w7(32'hbc35f04d),
	.w8(32'hba9190d0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab533fb),
	.w1(32'h3b545c5a),
	.w2(32'h3c54a4a2),
	.w3(32'hbbc5b0e0),
	.w4(32'hbb46baa4),
	.w5(32'h39ab548e),
	.w6(32'hbae18f8c),
	.w7(32'h3c167454),
	.w8(32'hb99e2d06),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5975cd),
	.w1(32'hbab26ff5),
	.w2(32'hba309bd5),
	.w3(32'hba8f3f7c),
	.w4(32'hb6c196ab),
	.w5(32'hbb9025bd),
	.w6(32'hbb006857),
	.w7(32'h3b609dd5),
	.w8(32'hbab96705),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff367c),
	.w1(32'h394b0f5a),
	.w2(32'h3bb4ea68),
	.w3(32'h3a867b31),
	.w4(32'h3c28ad6c),
	.w5(32'hbb9c4dd6),
	.w6(32'hbbe963ef),
	.w7(32'h3c0e28e9),
	.w8(32'h3b2f945c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a369856),
	.w1(32'hbb84cf61),
	.w2(32'hbc328418),
	.w3(32'hbbc06cc5),
	.w4(32'hbc3091fb),
	.w5(32'hbb9fac1f),
	.w6(32'h3bbd1d86),
	.w7(32'hbc0d4e83),
	.w8(32'hbc10b6ea),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb7b0),
	.w1(32'hbb8c0043),
	.w2(32'h3c00729c),
	.w3(32'hbb804440),
	.w4(32'h3bc94622),
	.w5(32'hbbe1dcad),
	.w6(32'hbbed61ad),
	.w7(32'h3ba78ecf),
	.w8(32'hbbcf8f45),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4b30e),
	.w1(32'hbb964265),
	.w2(32'hba4966b7),
	.w3(32'hbc0dc48a),
	.w4(32'hbb09b376),
	.w5(32'h3972f771),
	.w6(32'h3b0953d8),
	.w7(32'h3b3b7c9b),
	.w8(32'hb8f0410c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97caf4),
	.w1(32'hb99906da),
	.w2(32'hbafdaa90),
	.w3(32'hba4a5391),
	.w4(32'hbac6451a),
	.w5(32'h3ba7bbc7),
	.w6(32'h3abd53bf),
	.w7(32'hba575f13),
	.w8(32'h3b2b4828),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8855f2),
	.w1(32'hbb4a41a2),
	.w2(32'hbb948905),
	.w3(32'hbb1703d0),
	.w4(32'hba8d331c),
	.w5(32'h3b42424a),
	.w6(32'hbb8a63c8),
	.w7(32'hbb985494),
	.w8(32'h3ab79e69),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a336678),
	.w1(32'h39eb89ba),
	.w2(32'hbb2475c6),
	.w3(32'h3b1ce4ef),
	.w4(32'h392caae5),
	.w5(32'hba890c66),
	.w6(32'h3a16a245),
	.w7(32'hbb8cb01f),
	.w8(32'h3b45242a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6444ae),
	.w1(32'hb95ac9c1),
	.w2(32'h3acb9808),
	.w3(32'h3b113fde),
	.w4(32'hbb3d0196),
	.w5(32'hb9028aa5),
	.w6(32'h3bb69645),
	.w7(32'h3abd0240),
	.w8(32'hbbbc3e20),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebd7c9),
	.w1(32'hba84f868),
	.w2(32'hba0c34cc),
	.w3(32'hbb57f646),
	.w4(32'hbb11cd5f),
	.w5(32'h3b56b396),
	.w6(32'hbc3ba957),
	.w7(32'h3b4b5c50),
	.w8(32'h3a242248),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1720dc),
	.w1(32'h3b964f2b),
	.w2(32'hbad3afa2),
	.w3(32'h3aec0ea4),
	.w4(32'hbacb1549),
	.w5(32'hbab806d1),
	.w6(32'h3be2b1d3),
	.w7(32'hbbabb774),
	.w8(32'h3b1ea796),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb4cc),
	.w1(32'hbad8435a),
	.w2(32'hbb279d27),
	.w3(32'hb9fa7bae),
	.w4(32'hbb075f9a),
	.w5(32'hb9c4571f),
	.w6(32'h3bdc5eea),
	.w7(32'hbb7cbe34),
	.w8(32'hbafb620f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b2c9b),
	.w1(32'h3b701f14),
	.w2(32'h3c82812f),
	.w3(32'h3a17a399),
	.w4(32'h3b4c7db0),
	.w5(32'hba84afba),
	.w6(32'hbbc879bd),
	.w7(32'h3bffce5f),
	.w8(32'hbba7e22e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc3c8f),
	.w1(32'hbb745247),
	.w2(32'h3bb76235),
	.w3(32'hbbafa2b3),
	.w4(32'hba376820),
	.w5(32'hbbcf581b),
	.w6(32'hbc505e73),
	.w7(32'h3c07ceb3),
	.w8(32'hbbf8ae1b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc4af),
	.w1(32'hbb345f60),
	.w2(32'hbaa5bd05),
	.w3(32'hbbad11b3),
	.w4(32'hba7ccad1),
	.w5(32'h3b91bcc9),
	.w6(32'hbbce6b18),
	.w7(32'hbad979f5),
	.w8(32'h3b205781),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c0ad),
	.w1(32'hbadb647d),
	.w2(32'hbbf03223),
	.w3(32'hbb067fc9),
	.w4(32'h3b2b4c89),
	.w5(32'h3a79a945),
	.w6(32'h3c25dce7),
	.w7(32'h3b2a26e7),
	.w8(32'hbb3b1081),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185b8b),
	.w1(32'hbb931376),
	.w2(32'hbbe12a8b),
	.w3(32'hbb9706f9),
	.w4(32'hbb4dcec5),
	.w5(32'hbb03504d),
	.w6(32'hbc15f201),
	.w7(32'hbc209485),
	.w8(32'h3ac40982),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852981),
	.w1(32'hbb43bb6f),
	.w2(32'hbbc07afa),
	.w3(32'hbb3eccc0),
	.w4(32'h3807faa8),
	.w5(32'h3b4f0b38),
	.w6(32'h3afc280d),
	.w7(32'hba0c3dcd),
	.w8(32'h3ae2d69b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42e644),
	.w1(32'h3c3ef068),
	.w2(32'h3c11eddb),
	.w3(32'hba74bc5d),
	.w4(32'h3c535796),
	.w5(32'hba3608b2),
	.w6(32'hbc289303),
	.w7(32'h3c6de04e),
	.w8(32'hbb091eb6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ef22a),
	.w1(32'hbb14688d),
	.w2(32'h3b265ee6),
	.w3(32'hba707666),
	.w4(32'h3a8aac01),
	.w5(32'hbbc85dfb),
	.w6(32'hbb260c1c),
	.w7(32'h3b060edf),
	.w8(32'hbb9ab80d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850313),
	.w1(32'hbb81eca4),
	.w2(32'h3bb2d444),
	.w3(32'hbb790dc9),
	.w4(32'hbab5d100),
	.w5(32'hbad21060),
	.w6(32'hbaef1480),
	.w7(32'h3b2c5018),
	.w8(32'h3b2b7800),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99617df),
	.w1(32'h3b214219),
	.w2(32'h3ba6b385),
	.w3(32'hba17cd05),
	.w4(32'h3bb36419),
	.w5(32'hbb5a6167),
	.w6(32'hb9d8b920),
	.w7(32'h3af83dcc),
	.w8(32'hbba471bc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb234d91),
	.w1(32'hb9cb9ae2),
	.w2(32'h3ba9501b),
	.w3(32'hbbb7bf8b),
	.w4(32'hbb5d0dbf),
	.w5(32'h3c4b05f1),
	.w6(32'hbb20295e),
	.w7(32'hba0bee11),
	.w8(32'h3baa983b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c9238),
	.w1(32'hbb303864),
	.w2(32'hbba220b1),
	.w3(32'h3c66ed59),
	.w4(32'hb87948ca),
	.w5(32'h38900bb8),
	.w6(32'h3c00af61),
	.w7(32'h3b689065),
	.w8(32'hba34958c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a9d7f),
	.w1(32'h3b558ce1),
	.w2(32'hbb10ed4a),
	.w3(32'hbabdffba),
	.w4(32'hba127991),
	.w5(32'hba3df603),
	.w6(32'h3b0bab8c),
	.w7(32'hbb4b5667),
	.w8(32'hb97bb99a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b439b39),
	.w1(32'h3b9539ba),
	.w2(32'h3b9e1f60),
	.w3(32'h3bbd7832),
	.w4(32'h3b367b6b),
	.w5(32'hbaa3bcdf),
	.w6(32'h3ba4f386),
	.w7(32'h3b1c07ad),
	.w8(32'hbb3497be),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule