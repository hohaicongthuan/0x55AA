module layer_10_featuremap_103(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f011d),
	.w1(32'hb80e4af5),
	.w2(32'hb81204f5),
	.w3(32'h37ad9599),
	.w4(32'hb81c9940),
	.w5(32'hb8112db7),
	.w6(32'h37e75467),
	.w7(32'hb7c0e588),
	.w8(32'hb78648ff),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a317b),
	.w1(32'hba80952a),
	.w2(32'hba9813bd),
	.w3(32'hbb1d2be3),
	.w4(32'hbb5214af),
	.w5(32'hbb4a66eb),
	.w6(32'hbadabb45),
	.w7(32'hbb3d20e0),
	.w8(32'hbb5dc49f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb558d3e6),
	.w1(32'hb5d30910),
	.w2(32'h35d4bb4f),
	.w3(32'h35ff8094),
	.w4(32'h348afb3f),
	.w5(32'h363fedd1),
	.w6(32'hb63c2a8f),
	.w7(32'h35caebc8),
	.w8(32'h36036a4f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5b972),
	.w1(32'h3ad329e7),
	.w2(32'h3a9b2018),
	.w3(32'h384b2ed0),
	.w4(32'h3a7f0a04),
	.w5(32'hb67ec768),
	.w6(32'h3943ddd9),
	.w7(32'h3a393ecc),
	.w8(32'hb98a50b7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c1eaf8),
	.w1(32'hb89f0c6c),
	.w2(32'h37c5dec9),
	.w3(32'hb912908d),
	.w4(32'hb901c531),
	.w5(32'h373c70d6),
	.w6(32'hb91add29),
	.w7(32'hb92bda7c),
	.w8(32'hb7c39913),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366859bf),
	.w1(32'h3735d5a3),
	.w2(32'h37727c53),
	.w3(32'hb72ebaa2),
	.w4(32'h3690d9b5),
	.w5(32'h3668e476),
	.w6(32'hb7a736c5),
	.w7(32'hb7027d91),
	.w8(32'hb61a8eb6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b929a3d),
	.w1(32'h3b8083c5),
	.w2(32'hbbea5213),
	.w3(32'h3c16a344),
	.w4(32'h3b922688),
	.w5(32'hbb468b1c),
	.w6(32'h3b9c7113),
	.w7(32'h3bda6292),
	.w8(32'hba8c25cb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171767),
	.w1(32'h3a855a95),
	.w2(32'hbbb8cc61),
	.w3(32'h397d05d7),
	.w4(32'hba2d8dda),
	.w5(32'h3ba2519b),
	.w6(32'hbbf8532b),
	.w7(32'hbc38071e),
	.w8(32'hbb53e8a6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39525d48),
	.w1(32'hba7fcbd3),
	.w2(32'hba30a1a2),
	.w3(32'hba130cab),
	.w4(32'hbaab3af9),
	.w5(32'hba8560ab),
	.w6(32'hba4876ed),
	.w7(32'hbabe4c9a),
	.w8(32'hba8e7db9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf9704),
	.w1(32'h3ad0c4fc),
	.w2(32'hbba7f31a),
	.w3(32'h3be1a6ca),
	.w4(32'h3b88975d),
	.w5(32'hbb8c227c),
	.w6(32'h3bd329da),
	.w7(32'h3b8802e6),
	.w8(32'hbb0510ce),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393be004),
	.w1(32'h398b7edd),
	.w2(32'h3836db5a),
	.w3(32'h3a014a74),
	.w4(32'h39b466c4),
	.w5(32'h3936b362),
	.w6(32'h395f2fdb),
	.w7(32'h38af0e8f),
	.w8(32'hb8ebe47e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897a5a),
	.w1(32'h3c059fd9),
	.w2(32'hbc33a9ec),
	.w3(32'h3bf8505c),
	.w4(32'h3c3a9d20),
	.w5(32'hbbd3a604),
	.w6(32'h3ae5b808),
	.w7(32'h3be1cf22),
	.w8(32'hbb93e132),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0133ce),
	.w1(32'h3b8281d4),
	.w2(32'hbb2df0df),
	.w3(32'h3bc99d83),
	.w4(32'h3baa7735),
	.w5(32'hb9c5d9f1),
	.w6(32'h3bb77925),
	.w7(32'h3b984ec4),
	.w8(32'hb9c5ff4e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d5e70),
	.w1(32'hb9d35593),
	.w2(32'hbb649de9),
	.w3(32'h3b526ac4),
	.w4(32'hbb021b6e),
	.w5(32'hbb077afc),
	.w6(32'h3acec0d3),
	.w7(32'hbb06020e),
	.w8(32'hbb0abd3a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bf373),
	.w1(32'h3a3d475e),
	.w2(32'h39739ce6),
	.w3(32'h390aeb9d),
	.w4(32'hb9480675),
	.w5(32'hbaf036c3),
	.w6(32'h38485423),
	.w7(32'hba2dde13),
	.w8(32'hbb1de0ac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08a865),
	.w1(32'hbb812eb5),
	.w2(32'hbbb25e83),
	.w3(32'h3b3a34f9),
	.w4(32'hbba3642b),
	.w5(32'hbbcd089b),
	.w6(32'hbb62a426),
	.w7(32'hbbde5ad2),
	.w8(32'hbb8e67ae),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9127feb),
	.w1(32'hb80472db),
	.w2(32'hb85d0e60),
	.w3(32'h389410ab),
	.w4(32'hb7e46ebd),
	.w5(32'hb9963c80),
	.w6(32'h3a1d0f0f),
	.w7(32'h397cc184),
	.w8(32'hb98c31a2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36258e),
	.w1(32'h3b470c06),
	.w2(32'hbbb58898),
	.w3(32'h3bbd31ed),
	.w4(32'h3b04caee),
	.w5(32'hbb201ec7),
	.w6(32'hbaf06a8e),
	.w7(32'hba5f3670),
	.w8(32'hbb35f535),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c979),
	.w1(32'h3accd2fe),
	.w2(32'hbafe9c74),
	.w3(32'h3b892204),
	.w4(32'h3b35fa84),
	.w5(32'hb922ee3f),
	.w6(32'h3b03e1d3),
	.w7(32'h3ad776f3),
	.w8(32'hb944b5e3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9b113),
	.w1(32'h39a68f8e),
	.w2(32'h388435ef),
	.w3(32'h38ecd48c),
	.w4(32'h399c9ef2),
	.w5(32'h382ecd26),
	.w6(32'h387f63e2),
	.w7(32'h38803775),
	.w8(32'hb857b541),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b2b50),
	.w1(32'h39f7219b),
	.w2(32'h392b396c),
	.w3(32'h38c9b692),
	.w4(32'h39091dcb),
	.w5(32'h39019069),
	.w6(32'h38d568e7),
	.w7(32'h3697bf3f),
	.w8(32'hb73b3f75),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6797ec),
	.w1(32'h3aaabe85),
	.w2(32'h3a9c693f),
	.w3(32'hbac03636),
	.w4(32'h39fae5d1),
	.w5(32'h39c34228),
	.w6(32'hba325bbe),
	.w7(32'h39f045e4),
	.w8(32'h39be7656),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad99ce),
	.w1(32'hba07c0d0),
	.w2(32'hbc69b5b6),
	.w3(32'h3b2cf746),
	.w4(32'hbaab1fb3),
	.w5(32'hbc44f53a),
	.w6(32'h3bad12f8),
	.w7(32'h3937fae2),
	.w8(32'hbc40fae7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b409e0f),
	.w1(32'h3ad01db6),
	.w2(32'hba967512),
	.w3(32'h3b56a0b9),
	.w4(32'h3b13efda),
	.w5(32'hbaa98260),
	.w6(32'h3b474164),
	.w7(32'h3b27934a),
	.w8(32'hba34fb97),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bc009),
	.w1(32'h3bc01499),
	.w2(32'h3badfab1),
	.w3(32'hbb9654eb),
	.w4(32'hbb2773f4),
	.w5(32'hbae00813),
	.w6(32'hbab06ced),
	.w7(32'hbae11ec4),
	.w8(32'hbb89e089),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9365b32),
	.w1(32'hba92bb54),
	.w2(32'hbaa66174),
	.w3(32'h39f185e0),
	.w4(32'hba0a87d6),
	.w5(32'hba5cdcb8),
	.w6(32'h391ecd55),
	.w7(32'hb9e5322f),
	.w8(32'hba88c83c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e19c67),
	.w1(32'h3835ee24),
	.w2(32'h38a8b049),
	.w3(32'hb8d5dd02),
	.w4(32'h3818f623),
	.w5(32'h38b42592),
	.w6(32'hb8ba7878),
	.w7(32'hb7096907),
	.w8(32'h37c851ea),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18db39),
	.w1(32'hbb821484),
	.w2(32'h3b318650),
	.w3(32'hbc33eb9f),
	.w4(32'hbbc2c42c),
	.w5(32'hbb77f671),
	.w6(32'h3ac9a93a),
	.w7(32'h3b3e15cc),
	.w8(32'h3bb5bed1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd7b0c),
	.w1(32'h39d14061),
	.w2(32'h38922151),
	.w3(32'hb9bf4103),
	.w4(32'h3866426b),
	.w5(32'h387e5904),
	.w6(32'hba49c071),
	.w7(32'hb9ecd420),
	.w8(32'hba072adb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38305a08),
	.w1(32'hbb34d9fb),
	.w2(32'h3b7a52ba),
	.w3(32'hbb656bfe),
	.w4(32'hbc0562d9),
	.w5(32'hbba1f31a),
	.w6(32'h3b7e91be),
	.w7(32'hbb1e27ed),
	.w8(32'hba605897),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8558af5),
	.w1(32'hb76b356d),
	.w2(32'hb7f35747),
	.w3(32'hb80ce04d),
	.w4(32'hb708280a),
	.w5(32'hb7dc9406),
	.w6(32'hb7643736),
	.w7(32'hb6c593a4),
	.w8(32'hb810e177),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39368ab8),
	.w1(32'h39623ab3),
	.w2(32'h385f5128),
	.w3(32'h3965ea70),
	.w4(32'h390a136d),
	.w5(32'hb90eb61b),
	.w6(32'h3987b7b5),
	.w7(32'h3841f1e4),
	.w8(32'hb968b57f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b652e76),
	.w1(32'h3acd7a6b),
	.w2(32'hbacd69cc),
	.w3(32'h3b5b099f),
	.w4(32'h3b142659),
	.w5(32'hba940277),
	.w6(32'h3ac6e9ea),
	.w7(32'h3a8e1648),
	.w8(32'hba9c0731),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921d330),
	.w1(32'h3a375ef7),
	.w2(32'h39870d69),
	.w3(32'hba9e2e87),
	.w4(32'hbabb2c2f),
	.w5(32'hbaf22bcb),
	.w6(32'h389d5103),
	.w7(32'hba7a2928),
	.w8(32'hbb0fca78),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac313b1),
	.w1(32'h3a8ad3cb),
	.w2(32'hb988fc73),
	.w3(32'h3a613c75),
	.w4(32'h3a3356b7),
	.w5(32'hba9e07b8),
	.w6(32'h38fd77bc),
	.w7(32'h399a791a),
	.w8(32'h396775e8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a0ed9),
	.w1(32'h3b869fc0),
	.w2(32'hbaeb9747),
	.w3(32'h3b2dea58),
	.w4(32'h3a888c55),
	.w5(32'hba88b12c),
	.w6(32'h39e27af1),
	.w7(32'h396c669a),
	.w8(32'hbb382430),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c9fa3),
	.w1(32'h3c7d67d4),
	.w2(32'hbc86d3df),
	.w3(32'hbc26ce10),
	.w4(32'h3bebf483),
	.w5(32'hbc2a43cc),
	.w6(32'hbbc56292),
	.w7(32'hbb8b3dc4),
	.w8(32'hbcadce0f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0902c2),
	.w1(32'h3bc3b501),
	.w2(32'h3b97b86b),
	.w3(32'hbba24f37),
	.w4(32'h3b5c0749),
	.w5(32'hbb27fa90),
	.w6(32'hba5e0af2),
	.w7(32'h3ba3e1c0),
	.w8(32'hba2ae537),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba94f1e),
	.w1(32'hbbf775d2),
	.w2(32'hba3564b6),
	.w3(32'hbb2157ec),
	.w4(32'hbb9f3814),
	.w5(32'hbb1088d8),
	.w6(32'h3b454f85),
	.w7(32'h3b769e3e),
	.w8(32'h3bbc8205),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0129c4),
	.w1(32'h3b0a3155),
	.w2(32'h3ae61d60),
	.w3(32'hbac4e441),
	.w4(32'h3a7df439),
	.w5(32'h39a450e1),
	.w6(32'hba1507ae),
	.w7(32'h3ab427de),
	.w8(32'h39f42294),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a1940),
	.w1(32'h39806d06),
	.w2(32'h39154aed),
	.w3(32'h395d635b),
	.w4(32'h394dd291),
	.w5(32'h3937fde8),
	.w6(32'h39303721),
	.w7(32'h392a1858),
	.w8(32'h3834916c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70a59b6),
	.w1(32'h39539695),
	.w2(32'h398d923b),
	.w3(32'hb9865e80),
	.w4(32'h38af5310),
	.w5(32'h3936ee73),
	.w6(32'hb9721761),
	.w7(32'h388e3fea),
	.w8(32'h39314491),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d492c2),
	.w1(32'h3afac52b),
	.w2(32'hbab86980),
	.w3(32'h3a2482e9),
	.w4(32'h3aac7b3f),
	.w5(32'hbac84304),
	.w6(32'h3a12d8b6),
	.w7(32'h3a9845f3),
	.w8(32'hbae1e87b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbef332),
	.w1(32'hbac82070),
	.w2(32'hbb9533f4),
	.w3(32'h3b567864),
	.w4(32'h3a3c6f90),
	.w5(32'hba9df27b),
	.w6(32'h3b79cdcb),
	.w7(32'h3a346478),
	.w8(32'hba7c09f1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e11b),
	.w1(32'h3aec95b3),
	.w2(32'h36c96a85),
	.w3(32'hbaafb2ef),
	.w4(32'hb754d8c4),
	.w5(32'hbb31490e),
	.w6(32'h3b27d20a),
	.w7(32'h3af287e9),
	.w8(32'hbb0f6266),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888d02),
	.w1(32'h3b93e72e),
	.w2(32'hba14c6f5),
	.w3(32'h3a2a3b51),
	.w4(32'h39e35504),
	.w5(32'hbb088809),
	.w6(32'h3b4b0969),
	.w7(32'h3a6febe4),
	.w8(32'hbb816c17),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f24f4a),
	.w1(32'hba43f140),
	.w2(32'hbb08a01e),
	.w3(32'hba53602c),
	.w4(32'hbac05634),
	.w5(32'hbb525940),
	.w6(32'h3921c12f),
	.w7(32'h39a51739),
	.w8(32'h3a3de07c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c4ac1),
	.w1(32'h3b92b473),
	.w2(32'hbc1b091e),
	.w3(32'h3c1dee0a),
	.w4(32'h3bbfcfea),
	.w5(32'hbb78a970),
	.w6(32'h3bc28f45),
	.w7(32'h3b3c538f),
	.w8(32'hbba755b8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925b035),
	.w1(32'h38fa65f3),
	.w2(32'h394f05ed),
	.w3(32'hb971ef79),
	.w4(32'hb88af337),
	.w5(32'h399020a6),
	.w6(32'hb94c4641),
	.w7(32'hb865d860),
	.w8(32'h399049e7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3f0e6),
	.w1(32'hba2d5109),
	.w2(32'hb94dc3eb),
	.w3(32'hba633dd7),
	.w4(32'hba1c3405),
	.w5(32'h388880d1),
	.w6(32'hba1d24e8),
	.w7(32'hb938e4a0),
	.w8(32'h39a00fcd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9704641),
	.w1(32'hb9e2e6ef),
	.w2(32'h38133e94),
	.w3(32'hba3a46ef),
	.w4(32'hba42f730),
	.w5(32'hb857f4fc),
	.w6(32'hba21410a),
	.w7(32'hba3485d8),
	.w8(32'hb9268c41),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da4ede),
	.w1(32'hba72f136),
	.w2(32'h3a98204a),
	.w3(32'hba497390),
	.w4(32'hb7870fbd),
	.w5(32'h39430806),
	.w6(32'h3afcba4a),
	.w7(32'h3accc74d),
	.w8(32'hb9bd0acf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b18918),
	.w1(32'h39c6bbd5),
	.w2(32'hba2f066f),
	.w3(32'hba466f7f),
	.w4(32'hb9ec3f3f),
	.w5(32'hb9654654),
	.w6(32'hba47de53),
	.w7(32'hba26e165),
	.w8(32'hba6fe5bd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ee4b),
	.w1(32'h3a90f67d),
	.w2(32'hbbff90d5),
	.w3(32'h3c248b64),
	.w4(32'h3bda0057),
	.w5(32'hbb499a9b),
	.w6(32'h3b9d3d09),
	.w7(32'h3ae0d422),
	.w8(32'hbb50e958),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a16785),
	.w1(32'h39b13b3f),
	.w2(32'hbaae20c7),
	.w3(32'hba85d997),
	.w4(32'hba48b8ef),
	.w5(32'hba926320),
	.w6(32'hb90aed4d),
	.w7(32'hb956a312),
	.w8(32'hb9c3c366),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbe968),
	.w1(32'hb961bd65),
	.w2(32'hb9545290),
	.w3(32'h3885c358),
	.w4(32'hb91244f1),
	.w5(32'hb989ff89),
	.w6(32'h395de23f),
	.w7(32'hb90f7896),
	.w8(32'hb9cf81a6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807a0bb),
	.w1(32'hb668062a),
	.w2(32'hb7d3ceed),
	.w3(32'hb7d3da91),
	.w4(32'hb73ba9af),
	.w5(32'hb845b776),
	.w6(32'hb85ae989),
	.w7(32'hb813caf2),
	.w8(32'hb8821546),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1019f),
	.w1(32'hb988ed1a),
	.w2(32'h394c775f),
	.w3(32'hb7bc1175),
	.w4(32'hb9d97979),
	.w5(32'hb976eede),
	.w6(32'h39c8f1a5),
	.w7(32'hb7a6f331),
	.w8(32'h37e5fe83),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f44c3),
	.w1(32'h3a3493aa),
	.w2(32'h37fd7027),
	.w3(32'hb88c8944),
	.w4(32'h39eb71c5),
	.w5(32'hb991ec0f),
	.w6(32'h38015008),
	.w7(32'h3a0a6e40),
	.w8(32'hb8408a0e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5f025),
	.w1(32'h39740e28),
	.w2(32'hb9b28d58),
	.w3(32'h3a0a2919),
	.w4(32'h38c30239),
	.w5(32'hba9757f9),
	.w6(32'hb958cf5c),
	.w7(32'h3843d1c0),
	.w8(32'hb9acbf10),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4baed8),
	.w1(32'hb822d448),
	.w2(32'hbb016180),
	.w3(32'h3b44b229),
	.w4(32'h3ab3d8a9),
	.w5(32'hbab0b98d),
	.w6(32'h3a96433c),
	.w7(32'hb9c24a39),
	.w8(32'hbb03f416),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa412),
	.w1(32'hbb62aa1a),
	.w2(32'hbb587654),
	.w3(32'hbb6eeabf),
	.w4(32'hbb493c35),
	.w5(32'hbb46521e),
	.w6(32'hbb16ca6a),
	.w7(32'hbb4133ee),
	.w8(32'hbadf7649),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38294228),
	.w1(32'h383a6d62),
	.w2(32'h38a889cd),
	.w3(32'hb78eec63),
	.w4(32'hb785dec1),
	.w5(32'h37ba0c41),
	.w6(32'hb6d6c32a),
	.w7(32'hb82e7f80),
	.w8(32'hb7be9f46),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739a67b),
	.w1(32'h375559b3),
	.w2(32'h38485194),
	.w3(32'hb6cfa7d1),
	.w4(32'h3724cf0f),
	.w5(32'h38102eda),
	.w6(32'hb6812a9a),
	.w7(32'h37aa1fcf),
	.w8(32'h38159aeb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91def2d),
	.w1(32'hb8b9a977),
	.w2(32'hb858cb80),
	.w3(32'hb8f7ab3e),
	.w4(32'hb57cfbd7),
	.w5(32'h38860c8c),
	.w6(32'hb8c678b1),
	.w7(32'h37126d04),
	.w8(32'h3885a1c6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3753675d),
	.w1(32'h3896faff),
	.w2(32'h3873884e),
	.w3(32'h361bc50c),
	.w4(32'h381beb33),
	.w5(32'h382e0438),
	.w6(32'hb7a39744),
	.w7(32'h379daff9),
	.w8(32'h37694127),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c400705),
	.w1(32'hbb0db277),
	.w2(32'hbc356308),
	.w3(32'h3bb15055),
	.w4(32'h3b82d46d),
	.w5(32'hbc31d3c0),
	.w6(32'hbb055dc0),
	.w7(32'hb7a9e5e8),
	.w8(32'h3b3c56c0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8511e8),
	.w1(32'h3c8033e4),
	.w2(32'h3a320afb),
	.w3(32'h3a65c612),
	.w4(32'h3a107a51),
	.w5(32'hbb4f4db4),
	.w6(32'h39b7f25a),
	.w7(32'hbb636b1f),
	.w8(32'hbc45889c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22377d),
	.w1(32'hba227a69),
	.w2(32'hbb8e45a7),
	.w3(32'hba4e2c5b),
	.w4(32'hbb74590a),
	.w5(32'hbbbf8504),
	.w6(32'hb8c6abd4),
	.w7(32'hbb42342b),
	.w8(32'hbba0ef60),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446265),
	.w1(32'h3ba0ccba),
	.w2(32'h3b778743),
	.w3(32'hbbaeacaf),
	.w4(32'hbb6c0fcd),
	.w5(32'hbba7c460),
	.w6(32'hbae2b02b),
	.w7(32'hbb1e3771),
	.w8(32'hbbec60dd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d505c7),
	.w1(32'h38981f1f),
	.w2(32'h37c2e87b),
	.w3(32'h37dfbea1),
	.w4(32'h3866a8a9),
	.w5(32'h37b0f821),
	.w6(32'h368d85f2),
	.w7(32'hb72b8f05),
	.w8(32'hb76db41a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8153e5f),
	.w1(32'h37807f87),
	.w2(32'h3891522f),
	.w3(32'hb86232da),
	.w4(32'hb780771e),
	.w5(32'h38763953),
	.w6(32'hb8a43ab2),
	.w7(32'hb7533257),
	.w8(32'h382e8f65),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7810ea9),
	.w1(32'h38078ab9),
	.w2(32'h38b4662f),
	.w3(32'hb85a03dd),
	.w4(32'h36e1817a),
	.w5(32'h3886afb1),
	.w6(32'hb88385d3),
	.w7(32'h3738eacd),
	.w8(32'h37d004ca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c0a70),
	.w1(32'h3adb63f8),
	.w2(32'hba58fe74),
	.w3(32'h3b017b2f),
	.w4(32'h3aabf37d),
	.w5(32'hb911b5da),
	.w6(32'h3aad1857),
	.w7(32'h39ca5b50),
	.w8(32'hb98d36b6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872b095),
	.w1(32'h38ccfa81),
	.w2(32'h3931e0a7),
	.w3(32'hb92b6174),
	.w4(32'h373f6e2c),
	.w5(32'h3927c475),
	.w6(32'hb9279b99),
	.w7(32'hb732ae46),
	.w8(32'h3903d3ad),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88eb63),
	.w1(32'h3b42ba4f),
	.w2(32'hbb7a4a80),
	.w3(32'h3b637e01),
	.w4(32'h3b963469),
	.w5(32'h39dc9b41),
	.w6(32'h3b609b6e),
	.w7(32'h3b45684e),
	.w8(32'h39867f03),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9bf37),
	.w1(32'h3bccb604),
	.w2(32'hbb816fa3),
	.w3(32'h3b894a1b),
	.w4(32'h3ae6a1b1),
	.w5(32'hbb42c65a),
	.w6(32'hb7def0f0),
	.w7(32'hbb2ae666),
	.w8(32'hbbf1ae8b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963bc0b),
	.w1(32'h3ad53cd0),
	.w2(32'hb7eb84fb),
	.w3(32'hbaa7b1af),
	.w4(32'hbabd5261),
	.w5(32'hbb505c21),
	.w6(32'h3a52d20c),
	.w7(32'h3a1933b1),
	.w8(32'hbadc363a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4874c6),
	.w1(32'h39ad9b35),
	.w2(32'hbb1a48f1),
	.w3(32'h3b11f8e2),
	.w4(32'hb98e6263),
	.w5(32'hbaf33eb6),
	.w6(32'h39ecd63e),
	.w7(32'hbacd7ca7),
	.w8(32'hbb0437ef),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8762d),
	.w1(32'h3b995352),
	.w2(32'hbb434f79),
	.w3(32'h3b5567b6),
	.w4(32'h3b18de57),
	.w5(32'hbb90dfe6),
	.w6(32'h3a9ad371),
	.w7(32'h3acc9a8e),
	.w8(32'h392a5fc3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0df68b),
	.w1(32'hba2736f3),
	.w2(32'hba73fca1),
	.w3(32'hb93fc110),
	.w4(32'hba1c725a),
	.w5(32'hbaf13b22),
	.w6(32'h3b088c69),
	.w7(32'h39f759b9),
	.w8(32'hba89c3c7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7025df),
	.w1(32'h3b0bae09),
	.w2(32'hbb3e09e6),
	.w3(32'h3b561b82),
	.w4(32'h3b4449b7),
	.w5(32'hba259273),
	.w6(32'h3b2f2aa3),
	.w7(32'h3b19c62d),
	.w8(32'hb9c1a61f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d4c2e3),
	.w1(32'h37122c0e),
	.w2(32'h375bc19b),
	.w3(32'hb7847697),
	.w4(32'hb304415c),
	.w5(32'h373145cb),
	.w6(32'hb7a9973a),
	.w7(32'hb71ef203),
	.w8(32'h3791ae52),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f6ba2e),
	.w1(32'hb79f3787),
	.w2(32'hb71a6fa0),
	.w3(32'h37abb121),
	.w4(32'hb811b4d8),
	.w5(32'hb72262f3),
	.w6(32'h37ce9196),
	.w7(32'hb7b974c3),
	.w8(32'hb70ff68c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68c2738),
	.w1(32'h35b26511),
	.w2(32'h366f79d6),
	.w3(32'hb6fa958c),
	.w4(32'hb614ee9b),
	.w5(32'hb562a025),
	.w6(32'hb64a8621),
	.w7(32'hb6ff6f4d),
	.w8(32'hb4cc3d9c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68e8b2),
	.w1(32'hb95a7ed7),
	.w2(32'h39a5e6d7),
	.w3(32'hba56bfc5),
	.w4(32'hb9eb9221),
	.w5(32'h38819e42),
	.w6(32'hb8aa787e),
	.w7(32'h396f1f1f),
	.w8(32'h393d1d4a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfcbd2),
	.w1(32'h398476f6),
	.w2(32'hbb0f4c51),
	.w3(32'hbb4f7c97),
	.w4(32'hba93f057),
	.w5(32'hbba0bf4d),
	.w6(32'hba9e696d),
	.w7(32'hba99ddc6),
	.w8(32'hbb9500f8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a79ebd),
	.w1(32'h3a897543),
	.w2(32'hb8f8088c),
	.w3(32'hb919cab6),
	.w4(32'h3a2b8b40),
	.w5(32'hb9b1cdff),
	.w6(32'hb908ff6f),
	.w7(32'h3a50adf2),
	.w8(32'hb94009f3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9816b),
	.w1(32'h3b602772),
	.w2(32'h3aed1290),
	.w3(32'hbb424d36),
	.w4(32'hba563480),
	.w5(32'hb978a168),
	.w6(32'hbae773e2),
	.w7(32'hbaf25eb1),
	.w8(32'hbb591d57),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e08fb),
	.w1(32'h3b93e7f8),
	.w2(32'hbb65d12b),
	.w3(32'h3be44a8f),
	.w4(32'h3bb74dc1),
	.w5(32'hba882247),
	.w6(32'h3b97e9f1),
	.w7(32'h3b14c46f),
	.w8(32'hbb08e83b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b956),
	.w1(32'hbad842d5),
	.w2(32'h3ac16375),
	.w3(32'hba998123),
	.w4(32'hba63f8fa),
	.w5(32'hba077a5e),
	.w6(32'h3aff90b5),
	.w7(32'h3ba05323),
	.w8(32'h3b9aae05),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11429b),
	.w1(32'h3b0b990a),
	.w2(32'hbc5356c9),
	.w3(32'h3c066445),
	.w4(32'h3b623bc7),
	.w5(32'hbc3c6c7d),
	.w6(32'h3b3ba884),
	.w7(32'h3a982928),
	.w8(32'hbc2a172f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2712f),
	.w1(32'h3afa7e20),
	.w2(32'h3abfb3f8),
	.w3(32'hba9609a9),
	.w4(32'h3af24186),
	.w5(32'h3a636ba2),
	.w6(32'h3a86a0de),
	.w7(32'h3b3651ce),
	.w8(32'h3aa6ec32),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4eb615),
	.w1(32'h3b22b2b4),
	.w2(32'hbbb156b2),
	.w3(32'h3c04ec54),
	.w4(32'h3a0b1e0a),
	.w5(32'hbbcaaaa7),
	.w6(32'h3a534395),
	.w7(32'hbbbcd054),
	.w8(32'hbbeec108),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa85b),
	.w1(32'hba89e93f),
	.w2(32'hba8cf435),
	.w3(32'h3aa618d4),
	.w4(32'hbac097ef),
	.w5(32'hbb9befda),
	.w6(32'h39ccc2f0),
	.w7(32'h3911460b),
	.w8(32'hba9988f9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af971),
	.w1(32'hba9462e1),
	.w2(32'h3b45c4b8),
	.w3(32'hbb4905b8),
	.w4(32'hbb4afbc1),
	.w5(32'hbaf6416d),
	.w6(32'h39c47cd0),
	.w7(32'hb9281c41),
	.w8(32'h3a26eb59),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e6750),
	.w1(32'hba2608cc),
	.w2(32'h39d71e80),
	.w3(32'hb9c947e9),
	.w4(32'hb92e071f),
	.w5(32'h3a0bc3be),
	.w6(32'h391a0685),
	.w7(32'h3999e4df),
	.w8(32'h3a2e28bf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35c32),
	.w1(32'hb7e15fcc),
	.w2(32'hbb8459be),
	.w3(32'h3b82f1ac),
	.w4(32'h3a8c9b79),
	.w5(32'hbb2e4293),
	.w6(32'h3b0fc31b),
	.w7(32'h3a5fab52),
	.w8(32'hbb52442d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8485d),
	.w1(32'h3aa835a1),
	.w2(32'hbbd436ab),
	.w3(32'h3c003cc1),
	.w4(32'h3bedab46),
	.w5(32'hbb66fe82),
	.w6(32'h3bd8dcdf),
	.w7(32'h3bc2a362),
	.w8(32'h3b57c26f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a966ddf),
	.w1(32'h3c86b13a),
	.w2(32'hbacdec5e),
	.w3(32'hbc3a0f0d),
	.w4(32'h3ad38d2c),
	.w5(32'hbbbd69ed),
	.w6(32'hbc24c55a),
	.w7(32'hbb915c78),
	.w8(32'hbc9eb053),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ec080),
	.w1(32'h3c2bed91),
	.w2(32'h3b00e60c),
	.w3(32'hbb65c474),
	.w4(32'h3ba168e5),
	.w5(32'hbb85fd33),
	.w6(32'hbb6c5659),
	.w7(32'h3bc9e410),
	.w8(32'h3a801c7a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24224f),
	.w1(32'h3b5f3bf8),
	.w2(32'h3b271596),
	.w3(32'hbaf02d01),
	.w4(32'hb9366fe2),
	.w5(32'hba897d78),
	.w6(32'h39c9ad1a),
	.w7(32'h39981c5d),
	.w8(32'hbb5791b1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba14389),
	.w1(32'h3b8a5af4),
	.w2(32'hbc33e069),
	.w3(32'h3bc03352),
	.w4(32'h39d0ba08),
	.w5(32'hbbea19da),
	.w6(32'h3af5a3cc),
	.w7(32'h3b27b648),
	.w8(32'hbbc283af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db8290),
	.w1(32'h386cd137),
	.w2(32'h3a195799),
	.w3(32'hba854fe1),
	.w4(32'hb9ace9e0),
	.w5(32'h39d968b7),
	.w6(32'hb8e9b8b0),
	.w7(32'hb99ded92),
	.w8(32'h3a599006),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f0e86),
	.w1(32'h3b5fc2d1),
	.w2(32'hbbde0889),
	.w3(32'hbbd52b25),
	.w4(32'hbacde6fa),
	.w5(32'hbb4577ef),
	.w6(32'hbad3d071),
	.w7(32'hbc2aaa08),
	.w8(32'hbc10607e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81941),
	.w1(32'h3a2e658a),
	.w2(32'hbbb5d725),
	.w3(32'h3b26f638),
	.w4(32'h3b9435d8),
	.w5(32'hbb95c58d),
	.w6(32'h3bb088c2),
	.w7(32'h3bbac76e),
	.w8(32'hbb191195),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931645d),
	.w1(32'h38ce7522),
	.w2(32'h391e5e37),
	.w3(32'hb90c3df7),
	.w4(32'hb6995a8d),
	.w5(32'h389e514b),
	.w6(32'h3831de5f),
	.w7(32'h391ca7a7),
	.w8(32'h399146ed),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7513af),
	.w1(32'h3a749029),
	.w2(32'hb9a1669e),
	.w3(32'h386b8bc0),
	.w4(32'hb9899bce),
	.w5(32'hbaffaaf9),
	.w6(32'hba8b17d8),
	.w7(32'hba7ea7f0),
	.w8(32'hbb1d2c3c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4580),
	.w1(32'hb9a54c86),
	.w2(32'hbb99afe2),
	.w3(32'h3b6b9d27),
	.w4(32'h3b0986d0),
	.w5(32'hbadd976a),
	.w6(32'h3b611ed9),
	.w7(32'h3b2edb76),
	.w8(32'hbab2f6a6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d403f),
	.w1(32'hba43cd0f),
	.w2(32'h3a038bfc),
	.w3(32'hba859914),
	.w4(32'hbac83d33),
	.w5(32'hbae29137),
	.w6(32'h3abc0173),
	.w7(32'h3aa5b3af),
	.w8(32'hbafe8aa1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9393d6),
	.w1(32'hbb93eb69),
	.w2(32'hba9c072c),
	.w3(32'h3a5de7a2),
	.w4(32'hbb386196),
	.w5(32'hbafb4572),
	.w6(32'h3b6bcb16),
	.w7(32'h3a519aac),
	.w8(32'h3af306be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd49c1),
	.w1(32'hba38737a),
	.w2(32'hb9f17ab8),
	.w3(32'hba6169f6),
	.w4(32'hbacb590f),
	.w5(32'hbafd9a9e),
	.w6(32'hba24eb7f),
	.w7(32'hbabf66c0),
	.w8(32'hbabdf203),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c453471),
	.w1(32'h3c3e75b5),
	.w2(32'h3b87cea8),
	.w3(32'hb8824c6d),
	.w4(32'h3b39329f),
	.w5(32'hb9ebfa94),
	.w6(32'hbbe9cc9f),
	.w7(32'hbb91a8ad),
	.w8(32'hbbfacb9f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd813a),
	.w1(32'hbb550a15),
	.w2(32'hbbae53f8),
	.w3(32'h39fa9426),
	.w4(32'hbb609c79),
	.w5(32'hbbc058dd),
	.w6(32'hbb8531b3),
	.w7(32'hbbcc40a4),
	.w8(32'hbb5b801b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47613b),
	.w1(32'h39531e5d),
	.w2(32'hba3f9842),
	.w3(32'h3a920d8c),
	.w4(32'hb7cad058),
	.w5(32'hbacca84b),
	.w6(32'h3adacb11),
	.w7(32'h398f6249),
	.w8(32'hbafb484a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837274a),
	.w1(32'hb79c3a86),
	.w2(32'h371bedd0),
	.w3(32'h37a20944),
	.w4(32'hb83f6985),
	.w5(32'h36c3a416),
	.w6(32'h382722f5),
	.w7(32'hb72c6682),
	.w8(32'h3730a65c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395237e5),
	.w1(32'hb91c7b6c),
	.w2(32'hba62ff97),
	.w3(32'hb98ed30d),
	.w4(32'hba396656),
	.w5(32'hbab5c1ba),
	.w6(32'hb9c80836),
	.w7(32'hba84653c),
	.w8(32'hba9ac6d3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3739443b),
	.w1(32'hb6587767),
	.w2(32'h38365eb2),
	.w3(32'h380fdb15),
	.w4(32'hb6826be3),
	.w5(32'h388b0ed5),
	.w6(32'hb844e36e),
	.w7(32'hb719560f),
	.w8(32'h38092fe5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910f412),
	.w1(32'hb9194353),
	.w2(32'hb98be221),
	.w3(32'hb961fdf0),
	.w4(32'hb9407ac5),
	.w5(32'hb94a3296),
	.w6(32'hb8e9af05),
	.w7(32'hb852871f),
	.w8(32'hb686438c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1be9e9),
	.w1(32'h3abd89a5),
	.w2(32'h39dae333),
	.w3(32'hb90bb5f7),
	.w4(32'h39beab98),
	.w5(32'hba950537),
	.w6(32'h3ab6ec8b),
	.w7(32'h39c30754),
	.w8(32'hbab8a4fc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cd850),
	.w1(32'h39c1805f),
	.w2(32'h392f0756),
	.w3(32'h3975dff2),
	.w4(32'h389de9ad),
	.w5(32'hb94a27a9),
	.w6(32'hb8f7ab4a),
	.w7(32'hb7dc922a),
	.w8(32'hb8168458),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939c20),
	.w1(32'h3b3a07ad),
	.w2(32'hbb206dd9),
	.w3(32'h3b267f8b),
	.w4(32'h3b1e4384),
	.w5(32'hba3e6654),
	.w6(32'h3b060b67),
	.w7(32'h3abac9c9),
	.w8(32'hba117673),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d99f4e),
	.w1(32'hba8720e8),
	.w2(32'h3adc8d77),
	.w3(32'hbb5c2fc1),
	.w4(32'hbbc2f426),
	.w5(32'hbb198eba),
	.w6(32'hba8d4e4e),
	.w7(32'hbb74fbe9),
	.w8(32'hbb58f41b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81df960),
	.w1(32'hb75c6a4f),
	.w2(32'hb7f796bc),
	.w3(32'hb8a1f3e8),
	.w4(32'hb882e5f3),
	.w5(32'hb835dbbf),
	.w6(32'hb8790b16),
	.w7(32'hb87bdec3),
	.w8(32'hb84b8cde),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8b772),
	.w1(32'h38d3daa6),
	.w2(32'h385a55cd),
	.w3(32'h388733bb),
	.w4(32'h3813d65d),
	.w5(32'h391106c9),
	.w6(32'hb93461c8),
	.w7(32'hb70a86c2),
	.w8(32'h3961e551),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7563f5c),
	.w1(32'hb70d85eb),
	.w2(32'hb822ea1f),
	.w3(32'hb835e118),
	.w4(32'hb7b6e464),
	.w5(32'hb8824aa2),
	.w6(32'hb8812c5a),
	.w7(32'hb7de14de),
	.w8(32'hb84f8ea8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6c611),
	.w1(32'hb899afac),
	.w2(32'hb9cd9699),
	.w3(32'hb95c1b9e),
	.w4(32'hba04d8a6),
	.w5(32'hb9fc628e),
	.w6(32'hb9fbc35c),
	.w7(32'hba27d192),
	.w8(32'hb9f08321),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7f2d3),
	.w1(32'h3c9cbe76),
	.w2(32'hb9b79bca),
	.w3(32'h3c4f3ce3),
	.w4(32'h3bae96da),
	.w5(32'hb996ec47),
	.w6(32'hbad199a6),
	.w7(32'hbafadbde),
	.w8(32'hbc543dc8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbf84a),
	.w1(32'h393887cf),
	.w2(32'hbb74b7c3),
	.w3(32'h3bc47308),
	.w4(32'h3b08c91d),
	.w5(32'hbb2bf9f6),
	.w6(32'h3a47b846),
	.w7(32'h38d099ef),
	.w8(32'hbac9e236),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f1327),
	.w1(32'h39b54392),
	.w2(32'hbac9e4d9),
	.w3(32'h3a8adb28),
	.w4(32'h3a0f2ca3),
	.w5(32'hbaa126ab),
	.w6(32'h3ab4fe9d),
	.w7(32'h3a1239bb),
	.w8(32'hb9ea7d9e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d3be),
	.w1(32'hb92e4b0d),
	.w2(32'hbb0ba65a),
	.w3(32'hba13daf2),
	.w4(32'hbaf8a852),
	.w5(32'hbaf368e1),
	.w6(32'hba131d48),
	.w7(32'hbb61539c),
	.w8(32'hbb5316b5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f293ae),
	.w1(32'h3a97ec81),
	.w2(32'h3aac2cdb),
	.w3(32'hb99eaaee),
	.w4(32'h3a8f5ceb),
	.w5(32'h399e7c0b),
	.w6(32'h39cb9a89),
	.w7(32'h39fab932),
	.w8(32'h39bf9171),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37d0cd),
	.w1(32'h38a56f8e),
	.w2(32'hbaf02bff),
	.w3(32'h3b067b81),
	.w4(32'hba415443),
	.w5(32'hba6877a1),
	.w6(32'h3a00861f),
	.w7(32'hbb00fb90),
	.w8(32'hbafa4f1e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b7041),
	.w1(32'hbab161da),
	.w2(32'hb9ee66a9),
	.w3(32'hb91e9cb7),
	.w4(32'hbb53485d),
	.w5(32'hbb45ae52),
	.w6(32'hbacf79d8),
	.w7(32'hbb4daf63),
	.w8(32'hba97159c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094ade),
	.w1(32'h3b44c029),
	.w2(32'hbbda40db),
	.w3(32'h3beda2ad),
	.w4(32'h3baa6510),
	.w5(32'hbb46db3e),
	.w6(32'h3b262178),
	.w7(32'h3b264808),
	.w8(32'hba92a5f9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b72e1),
	.w1(32'h3adefdba),
	.w2(32'h3ac45bec),
	.w3(32'hbaa7cbea),
	.w4(32'hb79eef12),
	.w5(32'hba7508a7),
	.w6(32'h3995dcf2),
	.w7(32'h3a9409f6),
	.w8(32'hba3489b0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba838),
	.w1(32'h3a3c5eab),
	.w2(32'hbb540ec8),
	.w3(32'h3ba5d3af),
	.w4(32'h3a501fbc),
	.w5(32'hbb28c94c),
	.w6(32'h3ac92295),
	.w7(32'hb842d2e2),
	.w8(32'hbb2282f7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4161),
	.w1(32'h3b47b02f),
	.w2(32'hbbb4fe76),
	.w3(32'h3bcd4c53),
	.w4(32'h3bad01e0),
	.w5(32'hbab719dd),
	.w6(32'h3b90ad67),
	.w7(32'h3b133a04),
	.w8(32'hbac95e6a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34aecc),
	.w1(32'h3bcd2d70),
	.w2(32'h3b47c214),
	.w3(32'hbb5f542e),
	.w4(32'h3a4c87b8),
	.w5(32'hbab22565),
	.w6(32'hbaddb67d),
	.w7(32'hba5788a5),
	.w8(32'hbb79daf7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90eead),
	.w1(32'h39e890cd),
	.w2(32'hbb8b399a),
	.w3(32'h3b547d1f),
	.w4(32'h3ac4829b),
	.w5(32'hbb5f004b),
	.w6(32'h3acabefa),
	.w7(32'hb9d928de),
	.w8(32'hbb3d3a8d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393522e5),
	.w1(32'h38094c6a),
	.w2(32'hb9a7c062),
	.w3(32'h3a5b2455),
	.w4(32'hb8100cce),
	.w5(32'hba11f532),
	.w6(32'h3a102168),
	.w7(32'h38e33706),
	.w8(32'hba002f58),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23527b),
	.w1(32'hbaa61432),
	.w2(32'h3b6a8533),
	.w3(32'hbbb4ea2f),
	.w4(32'hbbd870fc),
	.w5(32'hbb2ccad8),
	.w6(32'hb9d8a0eb),
	.w7(32'hbb0b2485),
	.w8(32'h3a931f9b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d2aa6),
	.w1(32'hba565fc4),
	.w2(32'hb934d30a),
	.w3(32'hbac1ff8c),
	.w4(32'hba70fcad),
	.w5(32'hba50f118),
	.w6(32'hba282218),
	.w7(32'hba95210d),
	.w8(32'h3685c2c4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12d1d6),
	.w1(32'h3958c4b3),
	.w2(32'hb911a47c),
	.w3(32'h3a5f2926),
	.w4(32'h394bcabd),
	.w5(32'h38734f41),
	.w6(32'h396aa739),
	.w7(32'hb8269b6d),
	.w8(32'hb74c66bc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39684033),
	.w1(32'hb9c12b45),
	.w2(32'hb9699c98),
	.w3(32'h39ab8d87),
	.w4(32'hb8033e21),
	.w5(32'h3524adb7),
	.w6(32'hb911bb47),
	.w7(32'h392f90d9),
	.w8(32'h3a05f761),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92e286),
	.w1(32'h3a75582e),
	.w2(32'hba0f5d44),
	.w3(32'h3aafb627),
	.w4(32'h39a23096),
	.w5(32'hb9a45c16),
	.w6(32'h3a2a17a1),
	.w7(32'hb9817520),
	.w8(32'h395d3731),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10a6fa),
	.w1(32'h3974dd22),
	.w2(32'hbb0d45a7),
	.w3(32'hbb8783d3),
	.w4(32'hb985d780),
	.w5(32'hbb5b4028),
	.w6(32'hbb1cf379),
	.w7(32'hba5298f7),
	.w8(32'hbb6adca4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1985),
	.w1(32'h3b653220),
	.w2(32'hb98ca22b),
	.w3(32'h3b798fa4),
	.w4(32'h3b5ab418),
	.w5(32'h39c09833),
	.w6(32'h3b4db11f),
	.w7(32'h3b24d87d),
	.w8(32'hb97cc622),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96090a7),
	.w1(32'h36581fab),
	.w2(32'hb97a4b2e),
	.w3(32'hb89a22f5),
	.w4(32'h39096249),
	.w5(32'h398eab35),
	.w6(32'h385e570b),
	.w7(32'hb94ec277),
	.w8(32'hb9864e17),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934b89),
	.w1(32'h3a8a3366),
	.w2(32'hbb38d9db),
	.w3(32'h3b24960a),
	.w4(32'h3ad5de44),
	.w5(32'hbb4ce91d),
	.w6(32'h3ac41ffd),
	.w7(32'h3a848647),
	.w8(32'hbabc1eb2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991a60e),
	.w1(32'hb9b2ca61),
	.w2(32'hb9ff8757),
	.w3(32'h39bfaa7d),
	.w4(32'hb7f57914),
	.w5(32'hb8059882),
	.w6(32'h3a81379f),
	.w7(32'h3a33c726),
	.w8(32'h3a2d53fc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cdcb6),
	.w1(32'h3b7c0cc0),
	.w2(32'hbbd23862),
	.w3(32'h3bdeda6d),
	.w4(32'h3b67c1dd),
	.w5(32'hbb9f07cf),
	.w6(32'h3b9c6c4b),
	.w7(32'h3b4290ee),
	.w8(32'hbb7e8439),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6b29e),
	.w1(32'hbb70939a),
	.w2(32'hbb42eab4),
	.w3(32'hbab58812),
	.w4(32'hbb256f26),
	.w5(32'hbb4bcff1),
	.w6(32'h3b385505),
	.w7(32'h3a0a93b6),
	.w8(32'h3addbe32),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba736b9a),
	.w1(32'hbb1c98cf),
	.w2(32'hbb244c12),
	.w3(32'hbaedb7a6),
	.w4(32'hbaaf5b80),
	.w5(32'hbafd6a99),
	.w6(32'hb81f40e7),
	.w7(32'h398ba616),
	.w8(32'hbab7bc0b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1ba07),
	.w1(32'h3a5ef48d),
	.w2(32'h39c72f00),
	.w3(32'h398be230),
	.w4(32'hb909081f),
	.w5(32'h38d5f804),
	.w6(32'hba684564),
	.w7(32'hb9858637),
	.w8(32'hb82b3587),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1afa2),
	.w1(32'h3ac6add8),
	.w2(32'h37b8a849),
	.w3(32'hb9d9ad92),
	.w4(32'hba13a7c7),
	.w5(32'hbade531b),
	.w6(32'h39772006),
	.w7(32'hb91b5d6d),
	.w8(32'hbb11bc80),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf84ff4),
	.w1(32'hba4dd571),
	.w2(32'hbaeaa0ba),
	.w3(32'hbb51f493),
	.w4(32'hbaabf1c3),
	.w5(32'hbb0b1135),
	.w6(32'hbabc7c20),
	.w7(32'h3a3ab761),
	.w8(32'h3a3bc1f4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2558b6),
	.w1(32'hb8c9c4b6),
	.w2(32'h3a5382e7),
	.w3(32'hbb4d02ec),
	.w4(32'hba98ba49),
	.w5(32'hb9e7ffd2),
	.w6(32'hbadc181c),
	.w7(32'hba4d2a15),
	.w8(32'hb9f09b29),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd1e48),
	.w1(32'h3a5d4228),
	.w2(32'hbae9e514),
	.w3(32'h3ae8884e),
	.w4(32'h3aafe254),
	.w5(32'hb9a07bb3),
	.w6(32'h3abed180),
	.w7(32'h3a0a54f7),
	.w8(32'hba1c8dad),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc26e9),
	.w1(32'hb9924000),
	.w2(32'hba427fd7),
	.w3(32'hb9a20983),
	.w4(32'hb984d32f),
	.w5(32'hba2f9e77),
	.w6(32'hb98ed09c),
	.w7(32'hba0e144e),
	.w8(32'hba687ac6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18f35),
	.w1(32'h3b0ca3cc),
	.w2(32'hbb9860de),
	.w3(32'h3ba62ce2),
	.w4(32'h3b4b2f53),
	.w5(32'hbb3b20d3),
	.w6(32'h39ce25d9),
	.w7(32'h399018da),
	.w8(32'hbacc16ee),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b210e4d),
	.w1(32'h3a8debe9),
	.w2(32'hbb0c3a7f),
	.w3(32'h3b2a0bec),
	.w4(32'h3b1d7fbd),
	.w5(32'hba879ac5),
	.w6(32'h3af8c57d),
	.w7(32'h3b0f615d),
	.w8(32'h39ebf335),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6360b),
	.w1(32'h3b17cdde),
	.w2(32'h3b23ee31),
	.w3(32'hba65e7f9),
	.w4(32'hbacc6292),
	.w5(32'h3993228b),
	.w6(32'h3a6daf7c),
	.w7(32'hbaf42221),
	.w8(32'hbb004392),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3804cd21),
	.w1(32'hb908f329),
	.w2(32'hb8dcd59e),
	.w3(32'hb8cce795),
	.w4(32'hb89498a1),
	.w5(32'hb9011149),
	.w6(32'hb97d2f13),
	.w7(32'hba06da44),
	.w8(32'hba0ac15f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897fe6),
	.w1(32'h3b248125),
	.w2(32'hb9bd3206),
	.w3(32'h3b16b351),
	.w4(32'h3acfce51),
	.w5(32'h395c495e),
	.w6(32'hbb00675c),
	.w7(32'hbb059c17),
	.w8(32'hbac4b8c8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382ffb10),
	.w1(32'h398ab34d),
	.w2(32'h38f4ef01),
	.w3(32'hb949e8ea),
	.w4(32'h39022476),
	.w5(32'h39584b2f),
	.w6(32'h39855310),
	.w7(32'h395582cf),
	.w8(32'h3a0e372c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ced341),
	.w1(32'h3a279dc8),
	.w2(32'h3a22001e),
	.w3(32'h38cd7d97),
	.w4(32'h39f3fe41),
	.w5(32'h39e233e6),
	.w6(32'h39c72e30),
	.w7(32'h3994c511),
	.w8(32'h39589bfd),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9ae6e),
	.w1(32'hba1c02d2),
	.w2(32'hba765413),
	.w3(32'h3a491473),
	.w4(32'hba84ac67),
	.w5(32'hbb0a8915),
	.w6(32'h3a53dd44),
	.w7(32'hb9673e70),
	.w8(32'hbaf8d77e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f92f2),
	.w1(32'h3bda51c0),
	.w2(32'hbb396876),
	.w3(32'h3b9369ff),
	.w4(32'h3b311054),
	.w5(32'hbb303d88),
	.w6(32'h3b3258df),
	.w7(32'h3a7f60f1),
	.w8(32'hbbaeb2c5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9487dfa),
	.w1(32'h3a8975df),
	.w2(32'h39cc6360),
	.w3(32'hb9156083),
	.w4(32'h3a760ccb),
	.w5(32'h395e07a4),
	.w6(32'hba1cd7f2),
	.w7(32'hb91c1dfd),
	.w8(32'hb919579a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af21759),
	.w1(32'h3a1ffa8d),
	.w2(32'h3abd5c55),
	.w3(32'h3a1cfe3b),
	.w4(32'hbb1cf579),
	.w5(32'hbaf9917a),
	.w6(32'h3ade841e),
	.w7(32'hba533225),
	.w8(32'hbae4bb20),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddc247),
	.w1(32'hba184c92),
	.w2(32'hb822758d),
	.w3(32'h3a11a241),
	.w4(32'h3a68dba2),
	.w5(32'hbab5862b),
	.w6(32'h3acfc8c0),
	.w7(32'h3add6d4b),
	.w8(32'h3ae5f6fc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b308264),
	.w1(32'hbabce3a5),
	.w2(32'hbb580194),
	.w3(32'h3919f951),
	.w4(32'h3a6d7322),
	.w5(32'hbb38d061),
	.w6(32'h3a206c0e),
	.w7(32'hb9d56ccc),
	.w8(32'hba0332bf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd120d0),
	.w1(32'h3ab6188d),
	.w2(32'hbaedcfad),
	.w3(32'h3b8bc80f),
	.w4(32'h3aa86a2c),
	.w5(32'hba0a276c),
	.w6(32'h3b56c00b),
	.w7(32'h3a9bf77d),
	.w8(32'hb82d4d89),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf48d),
	.w1(32'hba44d665),
	.w2(32'hbb5ddbfb),
	.w3(32'h3b95225a),
	.w4(32'h3aad4311),
	.w5(32'hbaa189c6),
	.w6(32'h3b3c8227),
	.w7(32'h3aa33488),
	.w8(32'hbab4fd83),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8805d5a),
	.w1(32'hba51487f),
	.w2(32'hba22b605),
	.w3(32'h39fa281b),
	.w4(32'hb9e396cc),
	.w5(32'hba0855a7),
	.w6(32'hb880bd73),
	.w7(32'hb9eb7808),
	.w8(32'hb9e89cc1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85d054),
	.w1(32'hbb41c9d6),
	.w2(32'hbb25cc89),
	.w3(32'h3717f268),
	.w4(32'hbb11c079),
	.w5(32'hbb7fd54a),
	.w6(32'hba3cf161),
	.w7(32'hbaf10e76),
	.w8(32'hbac232d7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7c6b3),
	.w1(32'h39a839de),
	.w2(32'h398ef523),
	.w3(32'hb8eaa397),
	.w4(32'h39ad877a),
	.w5(32'h39a99156),
	.w6(32'h39b0abb4),
	.w7(32'h39ba1ab1),
	.w8(32'h39a684d7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a8658),
	.w1(32'h3986c1d8),
	.w2(32'hba0a85b7),
	.w3(32'h3a8c5884),
	.w4(32'h3a38757f),
	.w5(32'hb9944ccf),
	.w6(32'h3a58b56b),
	.w7(32'h3a984de0),
	.w8(32'h39f0a17a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dda2fc),
	.w1(32'h3a034784),
	.w2(32'hb9eff187),
	.w3(32'hb9916c20),
	.w4(32'hb75ba12a),
	.w5(32'hba890cea),
	.w6(32'h396322f3),
	.w7(32'hba97a39e),
	.w8(32'hba8a7fde),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af40bf8),
	.w1(32'hbb21dc95),
	.w2(32'hbb5b3432),
	.w3(32'h3a1e84d3),
	.w4(32'hbb54b0b9),
	.w5(32'hbb9925a0),
	.w6(32'hba9e93b3),
	.w7(32'hbb6134da),
	.w8(32'hbaddadd1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913bfb5),
	.w1(32'h364109a5),
	.w2(32'hb97d633e),
	.w3(32'h380facad),
	.w4(32'hb80a85b9),
	.w5(32'h3940756a),
	.w6(32'hb7eda3a0),
	.w7(32'hb98c6f85),
	.w8(32'hb92cc38d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f9a3e),
	.w1(32'hb9bfebd8),
	.w2(32'hba1884d5),
	.w3(32'hb9d3c492),
	.w4(32'hba66514f),
	.w5(32'hba3f479e),
	.w6(32'hb9211ff7),
	.w7(32'hb90503fb),
	.w8(32'hb643ae51),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16cf05),
	.w1(32'h39bb1aa5),
	.w2(32'h3a831603),
	.w3(32'hba8cf36c),
	.w4(32'hba189701),
	.w5(32'hba307182),
	.w6(32'h39827209),
	.w7(32'hba445942),
	.w8(32'hbac798f9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30651a),
	.w1(32'h3a2d759c),
	.w2(32'hbbf40deb),
	.w3(32'h3b9048c1),
	.w4(32'h3a2ee660),
	.w5(32'hbc0f4c1a),
	.w6(32'h3bb2fdd2),
	.w7(32'h3b2eae2a),
	.w8(32'hbb894aa7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d93d),
	.w1(32'h3b737e7c),
	.w2(32'hbbacbf3a),
	.w3(32'hbb467a2d),
	.w4(32'h3b0c8884),
	.w5(32'hba7f2c2e),
	.w6(32'hbb282607),
	.w7(32'hbb1a29de),
	.w8(32'hbbe406e9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9e494),
	.w1(32'h3a7d9377),
	.w2(32'h3a28b84b),
	.w3(32'h39da15f3),
	.w4(32'h3a2d910e),
	.w5(32'h3a4b6355),
	.w6(32'h3a08fc1a),
	.w7(32'h3a114436),
	.w8(32'h3a90bf56),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e89ec),
	.w1(32'h3bd39f80),
	.w2(32'hb99fb10a),
	.w3(32'h3c40dc20),
	.w4(32'h3be20fa7),
	.w5(32'h3a463f80),
	.w6(32'h3bb8b8f9),
	.w7(32'h3ad1306c),
	.w8(32'hbb41cdea),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3770f4),
	.w1(32'hbbae697c),
	.w2(32'hbadd595a),
	.w3(32'hba1001e2),
	.w4(32'hbb19f6a5),
	.w5(32'hbbc6f3cf),
	.w6(32'h3b5d6d19),
	.w7(32'h3b0fb145),
	.w8(32'h3b18d9e4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18c7e),
	.w1(32'h3b262cea),
	.w2(32'hbb35a64a),
	.w3(32'h3b303fd6),
	.w4(32'h3b43df8f),
	.w5(32'hba2dc796),
	.w6(32'h3ac0e747),
	.w7(32'h3aac4a0a),
	.w8(32'hba630ec9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38273ca0),
	.w1(32'hb85fba51),
	.w2(32'hba2a03d3),
	.w3(32'h37ec206e),
	.w4(32'hb97f732e),
	.w5(32'hba3558f6),
	.w6(32'hb9aa097d),
	.w7(32'hba34d230),
	.w8(32'h399b4aa5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b733f5),
	.w1(32'hb915a992),
	.w2(32'hb9eef948),
	.w3(32'h387eb9f1),
	.w4(32'hb9d1c8ad),
	.w5(32'hba043968),
	.w6(32'h372d943c),
	.w7(32'hb9184d59),
	.w8(32'h3a018fd1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392bbc93),
	.w1(32'hb9a6f47c),
	.w2(32'h388a756b),
	.w3(32'hb8b5806b),
	.w4(32'hb9dd1e67),
	.w5(32'hb986e4e9),
	.w6(32'hb931d036),
	.w7(32'hb89c82b5),
	.w8(32'h39928588),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e6b6),
	.w1(32'h3b76b90d),
	.w2(32'hbb834cae),
	.w3(32'h3ba05159),
	.w4(32'h3b548ca0),
	.w5(32'hbae59a10),
	.w6(32'hb7e8a6b8),
	.w7(32'h3a6079df),
	.w8(32'hbb38da76),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b386a02),
	.w1(32'h3b44c0aa),
	.w2(32'h390846d5),
	.w3(32'h3b0290f8),
	.w4(32'h3a2b28ff),
	.w5(32'hba522fbe),
	.w6(32'h3978d258),
	.w7(32'h3a428619),
	.w8(32'hba9c837c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edfb9c),
	.w1(32'h3af845d3),
	.w2(32'h3a876c75),
	.w3(32'hbaf07a18),
	.w4(32'hbab58f96),
	.w5(32'hba8af66a),
	.w6(32'hb92ee68c),
	.w7(32'hbac4ac3d),
	.w8(32'hbb3ea644),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a27433),
	.w1(32'h3a2ef501),
	.w2(32'hb6af231a),
	.w3(32'hb7c5317e),
	.w4(32'hb99904a9),
	.w5(32'hba09dc1e),
	.w6(32'h39d1a03f),
	.w7(32'hb9c7a954),
	.w8(32'hba86db25),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5477),
	.w1(32'h3aea7b00),
	.w2(32'hbb9081d5),
	.w3(32'h3bd88f50),
	.w4(32'h3b5022cf),
	.w5(32'hbb43b430),
	.w6(32'h3b7dcf7e),
	.w7(32'h3ac174ba),
	.w8(32'hbb760b92),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbdbb8),
	.w1(32'h3a8fa15b),
	.w2(32'hbb06a00c),
	.w3(32'hbae9a8e9),
	.w4(32'h3a1f97f1),
	.w5(32'hbacc57df),
	.w6(32'h39a7f32e),
	.w7(32'h37e7d6ad),
	.w8(32'hba998539),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e65ef),
	.w1(32'h39b06b7c),
	.w2(32'h3939112e),
	.w3(32'h38b4d94b),
	.w4(32'h39a7afaf),
	.w5(32'h39aee04a),
	.w6(32'h3994aa9d),
	.w7(32'h38bd159d),
	.w8(32'h38eec291),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9affea1),
	.w1(32'hbb1c9e27),
	.w2(32'hbb067edf),
	.w3(32'hbb058dde),
	.w4(32'hbb8ab079),
	.w5(32'hbb0bae7e),
	.w6(32'hbb19541e),
	.w7(32'hbb8d686b),
	.w8(32'hbaa1637f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3ad05),
	.w1(32'hb96efee5),
	.w2(32'hb8c0addc),
	.w3(32'h39ef5465),
	.w4(32'hb8cb7965),
	.w5(32'h38adb8b0),
	.w6(32'hb9bbd0fd),
	.w7(32'hb9ef7841),
	.w8(32'hb99f4428),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b299b63),
	.w1(32'h3958e524),
	.w2(32'hbb62f90f),
	.w3(32'h3b1f9101),
	.w4(32'h3a85f982),
	.w5(32'hbb33bd19),
	.w6(32'h3ad54b77),
	.w7(32'h3a64d5d0),
	.w8(32'hbb020ea6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf966d9),
	.w1(32'h39e3b4c2),
	.w2(32'h38f11497),
	.w3(32'hbba19f53),
	.w4(32'hba0242e0),
	.w5(32'hbb15a6fe),
	.w6(32'hbacfde92),
	.w7(32'hb9074357),
	.w8(32'hbaf12331),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aea60),
	.w1(32'h3a1a694d),
	.w2(32'hba73338e),
	.w3(32'hb9c4ccf3),
	.w4(32'hb76a4908),
	.w5(32'hbafbee12),
	.w6(32'h3a6e7022),
	.w7(32'h3a544c7c),
	.w8(32'hbacfd0ef),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ebd01),
	.w1(32'h3a08acc3),
	.w2(32'hb9e08b13),
	.w3(32'h39f94839),
	.w4(32'h39936113),
	.w5(32'hb9c91f8c),
	.w6(32'h398c2107),
	.w7(32'h3762e156),
	.w8(32'h38a90a87),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d783),
	.w1(32'hba74a3c3),
	.w2(32'hba472517),
	.w3(32'hbb4b1a93),
	.w4(32'hbb6043c0),
	.w5(32'hbb557492),
	.w6(32'hbab54eee),
	.w7(32'hba82c31d),
	.w8(32'hbaa69dd9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61def1),
	.w1(32'h3a440d07),
	.w2(32'hbaf90105),
	.w3(32'h3b45d027),
	.w4(32'h3a91399d),
	.w5(32'hbacde908),
	.w6(32'h39c26042),
	.w7(32'hbac22c99),
	.w8(32'hbb0aefb5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890ba5),
	.w1(32'h3b6359fa),
	.w2(32'h39e2fd9c),
	.w3(32'h3b7fb0e2),
	.w4(32'h3b48a577),
	.w5(32'h3a5b5e49),
	.w6(32'h3b841072),
	.w7(32'h3b428b49),
	.w8(32'h3960eb3c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eaa310),
	.w1(32'h3993869e),
	.w2(32'h384ae395),
	.w3(32'h3881c5f7),
	.w4(32'hb8d54d1f),
	.w5(32'hb845cc34),
	.w6(32'h39f1df35),
	.w7(32'h39cebd1e),
	.w8(32'h39f75ec6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985b7bb),
	.w1(32'hb9885b4c),
	.w2(32'hb9dfa33d),
	.w3(32'hb9348c57),
	.w4(32'hba006d71),
	.w5(32'hb9c9a39e),
	.w6(32'hb977b1f8),
	.w7(32'hb9ec8dbc),
	.w8(32'hb9439136),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152401),
	.w1(32'h3c20b9e0),
	.w2(32'hbb781fc5),
	.w3(32'h3b679f46),
	.w4(32'h3aec569e),
	.w5(32'hbb8a1e7f),
	.w6(32'h3ace58d1),
	.w7(32'h385b21e0),
	.w8(32'hbbbb1824),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcacf99),
	.w1(32'h3b87deb2),
	.w2(32'hbb24bdf8),
	.w3(32'h3b358eef),
	.w4(32'h3a330efa),
	.w5(32'hbb89e7fd),
	.w6(32'h3b7b3f7d),
	.w7(32'h3b07d5a6),
	.w8(32'hbba3203b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e699b6),
	.w1(32'h3afff032),
	.w2(32'h39376406),
	.w3(32'hba174510),
	.w4(32'h3a3d72ed),
	.w5(32'hbaa93f67),
	.w6(32'h3a850ea3),
	.w7(32'h392d11c6),
	.w8(32'hbb17d49b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd030b9),
	.w1(32'h3b653f66),
	.w2(32'hbbe0a2cc),
	.w3(32'h3b74706d),
	.w4(32'h3b28e366),
	.w5(32'hbbf77843),
	.w6(32'h3b079907),
	.w7(32'h3b747e36),
	.w8(32'h3ad840a4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818ad5e),
	.w1(32'hb98ca817),
	.w2(32'hb9925edc),
	.w3(32'hba770ea6),
	.w4(32'hba732417),
	.w5(32'h391d6ae8),
	.w6(32'hb9fa99bc),
	.w7(32'hbaa08351),
	.w8(32'hba1dee03),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25104c),
	.w1(32'h39fcd0cc),
	.w2(32'hbb0bc17e),
	.w3(32'h3a0db404),
	.w4(32'hbb017793),
	.w5(32'hbafb3b3c),
	.w6(32'h39c2a7b0),
	.w7(32'hbadccb5d),
	.w8(32'hbb0d6cf6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d046),
	.w1(32'h3cbfbcb2),
	.w2(32'hbc1e8513),
	.w3(32'hbb30340d),
	.w4(32'h3c8e6cee),
	.w5(32'hbbc9ad3d),
	.w6(32'hbbce39a4),
	.w7(32'h3c19426a),
	.w8(32'hbc3c22ea),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f83e5),
	.w1(32'h3bf5f9c6),
	.w2(32'hbb3e8af5),
	.w3(32'h3c10b884),
	.w4(32'h3bbc766d),
	.w5(32'hba73e51d),
	.w6(32'h3b0f0530),
	.w7(32'h3a288977),
	.w8(32'hbb38c6d2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a321),
	.w1(32'h3b2f8e2e),
	.w2(32'hbbe2b977),
	.w3(32'h3b162529),
	.w4(32'h3a5eb36c),
	.w5(32'hbb3f7761),
	.w6(32'h393fcf1c),
	.w7(32'h3a4d9959),
	.w8(32'hbb4eb306),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90694ce),
	.w1(32'h3ac5e417),
	.w2(32'h3b468a6c),
	.w3(32'hbb1c0937),
	.w4(32'hba8a775a),
	.w5(32'hb9655d0a),
	.w6(32'hba28683d),
	.w7(32'h3a289299),
	.w8(32'h3a82ec71),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4a296),
	.w1(32'hbab976c2),
	.w2(32'h3a62c4bb),
	.w3(32'hba5540fe),
	.w4(32'hbb6553df),
	.w5(32'hbb7ab231),
	.w6(32'h3aa14196),
	.w7(32'hba5c16de),
	.w8(32'hbb3a6072),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901050a),
	.w1(32'h38821b29),
	.w2(32'h38084468),
	.w3(32'hb8d15439),
	.w4(32'h38ec657f),
	.w5(32'hb892db37),
	.w6(32'h392d2704),
	.w7(32'h397eeec8),
	.w8(32'h39a63884),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3794cce4),
	.w1(32'hb7906aef),
	.w2(32'hb827fe50),
	.w3(32'hb94923ea),
	.w4(32'hba056660),
	.w5(32'hb9d5c906),
	.w6(32'h390b00ef),
	.w7(32'h39b88adb),
	.w8(32'h39f5835c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bf368),
	.w1(32'h3ad738be),
	.w2(32'h39e72494),
	.w3(32'h3b127ba3),
	.w4(32'h3a5bcf1e),
	.w5(32'hba1ac5fe),
	.w6(32'hbabb842b),
	.w7(32'hba592b34),
	.w8(32'hb8cec0b1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba3c73),
	.w1(32'h383b05d3),
	.w2(32'hba4f8751),
	.w3(32'h39bb8b06),
	.w4(32'h3989d8a8),
	.w5(32'hba056ec4),
	.w6(32'hb92b6ac9),
	.w7(32'hba0278a6),
	.w8(32'hb89e7776),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b452de1),
	.w1(32'h3b10bb49),
	.w2(32'hbb1cb074),
	.w3(32'h3b52bf8a),
	.w4(32'h3a933b3e),
	.w5(32'hba6d2d6d),
	.w6(32'h3b3e8e91),
	.w7(32'h3aa5ad62),
	.w8(32'hba32f143),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89c21),
	.w1(32'h3ba972fc),
	.w2(32'hbb94533c),
	.w3(32'h3a5fa972),
	.w4(32'hba581347),
	.w5(32'hbba353a5),
	.w6(32'h3a335550),
	.w7(32'hbb05a9af),
	.w8(32'hbc0642d4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39d3d3),
	.w1(32'hb84a6d94),
	.w2(32'hbb0ec789),
	.w3(32'hb9b84e5e),
	.w4(32'hba8ee2aa),
	.w5(32'hbb0e0b33),
	.w6(32'h39816f4e),
	.w7(32'hb9e6e486),
	.w8(32'hbac66208),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1cde9),
	.w1(32'h39bb1e2c),
	.w2(32'h38858ef3),
	.w3(32'h3812e356),
	.w4(32'hba2febd6),
	.w5(32'h3602aed5),
	.w6(32'hb9366f04),
	.w7(32'hb8bb9f55),
	.w8(32'hb89b984b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c393),
	.w1(32'h3c2508f3),
	.w2(32'hbc0eb9d2),
	.w3(32'h3b941349),
	.w4(32'h3b0ba7db),
	.w5(32'hbbbbd40d),
	.w6(32'hbade7f75),
	.w7(32'h3aa95848),
	.w8(32'hbc01419a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e612),
	.w1(32'h3ac57169),
	.w2(32'hbac2d359),
	.w3(32'h3b564f47),
	.w4(32'h3aed2ac4),
	.w5(32'hba343932),
	.w6(32'h3a1a8cd9),
	.w7(32'h39948366),
	.w8(32'hbaa76a10),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb0080),
	.w1(32'hb8144d6c),
	.w2(32'hb9c87f40),
	.w3(32'h3a0268cf),
	.w4(32'hb8084090),
	.w5(32'hb9e2001b),
	.w6(32'h37a62f93),
	.w7(32'hb8dab3e9),
	.w8(32'hb9dbecb8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee6cc0),
	.w1(32'h3b962efa),
	.w2(32'hbae97add),
	.w3(32'h3bcaa35e),
	.w4(32'h3baa0b3a),
	.w5(32'h3a751fb0),
	.w6(32'h3b408244),
	.w7(32'h3b3ee514),
	.w8(32'hb9de32e5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96beb57),
	.w1(32'hb80cf413),
	.w2(32'h3931efec),
	.w3(32'hb91099eb),
	.w4(32'hb95a2cc5),
	.w5(32'hb8e5daaa),
	.w6(32'h38b56728),
	.w7(32'h39847354),
	.w8(32'h3a13d9c1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a728761),
	.w1(32'h391c05d3),
	.w2(32'hba2c5cd6),
	.w3(32'h37dff697),
	.w4(32'hb8fa54da),
	.w5(32'hb9b363a1),
	.w6(32'h395bdc45),
	.w7(32'hb97056fa),
	.w8(32'hba42e79e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d6f8c),
	.w1(32'h38c26fea),
	.w2(32'h39432bd2),
	.w3(32'h380ea0d8),
	.w4(32'h3838b192),
	.w5(32'h39647aae),
	.w6(32'h38cfade9),
	.w7(32'h38ac94ae),
	.w8(32'h39518956),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeed1d),
	.w1(32'h3a240605),
	.w2(32'h39c4d87e),
	.w3(32'h3a00a5e4),
	.w4(32'h395cec67),
	.w5(32'h392b2cdf),
	.w6(32'h3a256526),
	.w7(32'h3a44d60c),
	.w8(32'h3a8574a9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2078c8),
	.w1(32'h3b0e5151),
	.w2(32'h3ab46ace),
	.w3(32'hb9887bc8),
	.w4(32'h3a72c67c),
	.w5(32'hb980e401),
	.w6(32'h39e0c887),
	.w7(32'h3a7e3383),
	.w8(32'h39b4da5c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ce98),
	.w1(32'hbb90688a),
	.w2(32'hbc0d99a4),
	.w3(32'h3bebe30f),
	.w4(32'h3ac621c4),
	.w5(32'hbbeb8ec5),
	.w6(32'h3baa7849),
	.w7(32'h393aa2a3),
	.w8(32'hbb44a279),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40393),
	.w1(32'h3b414b92),
	.w2(32'hbafde8c9),
	.w3(32'h3b9e92d5),
	.w4(32'h3b6b823f),
	.w5(32'hba0f553e),
	.w6(32'h3b127ccd),
	.w7(32'h3a109354),
	.w8(32'hbab1225e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78cbe3),
	.w1(32'hb9d8d3a2),
	.w2(32'hbb8145b2),
	.w3(32'h3bae8242),
	.w4(32'h3b8e8593),
	.w5(32'hbad2f173),
	.w6(32'h3b91d8ac),
	.w7(32'h3b64218d),
	.w8(32'h3a8731f1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ee36d),
	.w1(32'hb931bce6),
	.w2(32'hb916802e),
	.w3(32'h399eaf22),
	.w4(32'h3974b175),
	.w5(32'h37940300),
	.w6(32'hb94ec420),
	.w7(32'hb92a76fb),
	.w8(32'h37303a3c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ed001),
	.w1(32'hb81d4364),
	.w2(32'hb8e7db6d),
	.w3(32'hb97d159d),
	.w4(32'hb8d789d8),
	.w5(32'hb8e6946e),
	.w6(32'hb99de579),
	.w7(32'hb9a02588),
	.w8(32'hb9aafc81),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe4c80),
	.w1(32'h39f89f22),
	.w2(32'h3a1c9f73),
	.w3(32'h3a2e7e46),
	.w4(32'h3998b4a2),
	.w5(32'h39f32d92),
	.w6(32'h39e6191a),
	.w7(32'h3a030554),
	.w8(32'h39db307b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f842f),
	.w1(32'h39a34212),
	.w2(32'h39eb0b9e),
	.w3(32'h3a0fcf37),
	.w4(32'h396dcbc9),
	.w5(32'h39e5113c),
	.w6(32'h398c8c80),
	.w7(32'h39c4cad9),
	.w8(32'h39cf838f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eeacd),
	.w1(32'hbb237ef3),
	.w2(32'hbb2fdb73),
	.w3(32'h3aa9db3a),
	.w4(32'hbb48fac1),
	.w5(32'hbb285a32),
	.w6(32'hbae9cb46),
	.w7(32'hbb70dc0f),
	.w8(32'hbb5e566c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ed94),
	.w1(32'hb89aa26a),
	.w2(32'hb76cf6ab),
	.w3(32'h396b4d3e),
	.w4(32'hb963d3d1),
	.w5(32'h398a49f1),
	.w6(32'h3850548f),
	.w7(32'h382e70fa),
	.w8(32'h399ebe16),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9943c93),
	.w1(32'hb92632ef),
	.w2(32'hba4a5e15),
	.w3(32'hba071941),
	.w4(32'hb96c8ed7),
	.w5(32'hba79fad0),
	.w6(32'hbaaa28ec),
	.w7(32'hba9369cd),
	.w8(32'hba92fea0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab575c8),
	.w1(32'hbb0045f4),
	.w2(32'hbad2dead),
	.w3(32'hbb0bfba6),
	.w4(32'hbaec0780),
	.w5(32'hbad42d5f),
	.w6(32'hbabc36f8),
	.w7(32'hbb2ff888),
	.w8(32'hbacf164c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22fbd6),
	.w1(32'h39ece313),
	.w2(32'h3a171f62),
	.w3(32'hba112419),
	.w4(32'h39f2b967),
	.w5(32'h3a085c17),
	.w6(32'h39e7dc85),
	.w7(32'h3a01ff81),
	.w8(32'h3a06086a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff5ac3),
	.w1(32'h3a4d7670),
	.w2(32'hba311b7e),
	.w3(32'h3b02e5d4),
	.w4(32'h3a30b49a),
	.w5(32'hb961ab0d),
	.w6(32'h3a6403c8),
	.w7(32'h3a8b709a),
	.w8(32'h38979831),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98efdcd),
	.w1(32'hb9ad3b1e),
	.w2(32'hbab2def8),
	.w3(32'hba138065),
	.w4(32'hba7d8794),
	.w5(32'hba948aec),
	.w6(32'hba06ddbc),
	.w7(32'hb9e00263),
	.w8(32'h385f3c11),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13937c),
	.w1(32'hbb74ecf0),
	.w2(32'hbc0305ca),
	.w3(32'h3b4be187),
	.w4(32'hbae6e83f),
	.w5(32'hbbf13dff),
	.w6(32'hbbeca207),
	.w7(32'hbbec63b5),
	.w8(32'hbb3b465a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d56da2),
	.w1(32'h39ea3243),
	.w2(32'h39155df1),
	.w3(32'h39013167),
	.w4(32'h3a216560),
	.w5(32'h393afcf7),
	.w6(32'h399e34da),
	.w7(32'h39b93e7d),
	.w8(32'h39c5e289),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63998),
	.w1(32'h3be19559),
	.w2(32'h3b776021),
	.w3(32'h3aca6a9e),
	.w4(32'h3b24cc7a),
	.w5(32'h3a9209ec),
	.w6(32'hbaef883d),
	.w7(32'hbb72ebe7),
	.w8(32'hbb73867b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule