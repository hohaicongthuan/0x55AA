module layer_8_featuremap_173(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7274b9),
	.w1(32'hbc9d22e5),
	.w2(32'hbc3ceb32),
	.w3(32'hb9f4a29d),
	.w4(32'hbbef1537),
	.w5(32'hbc6724e8),
	.w6(32'h3b351cc6),
	.w7(32'hbbb5a40f),
	.w8(32'hbc02b507),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae4f32),
	.w1(32'hb9191af3),
	.w2(32'hbb387868),
	.w3(32'hbc36bb5a),
	.w4(32'h399cf0aa),
	.w5(32'h390eb948),
	.w6(32'h3be8223b),
	.w7(32'h3ad49fa5),
	.w8(32'hb8f631e3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191e50),
	.w1(32'h384d54de),
	.w2(32'hbbc61953),
	.w3(32'h3b5c2a87),
	.w4(32'hbc61f81e),
	.w5(32'hbc181cf1),
	.w6(32'h3bbf6cb5),
	.w7(32'hbb47c191),
	.w8(32'hb9ca9945),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25f7c4),
	.w1(32'hbc0ae1ed),
	.w2(32'hbb8bf020),
	.w3(32'hbbc48c0d),
	.w4(32'hbc83106b),
	.w5(32'hbbf2ece5),
	.w6(32'h396d977e),
	.w7(32'h3a82a8b0),
	.w8(32'h3afb6528),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea7a32),
	.w1(32'hbb91f881),
	.w2(32'hbbc80564),
	.w3(32'h3b910813),
	.w4(32'hbb5111cd),
	.w5(32'hbb47a721),
	.w6(32'h3a9038ba),
	.w7(32'hb960e78f),
	.w8(32'hbab549e9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2954d3),
	.w1(32'h3b22f0a9),
	.w2(32'hbaca43d6),
	.w3(32'hbb9b59ed),
	.w4(32'h3af28e6e),
	.w5(32'h3a4c0c06),
	.w6(32'h3c27fe08),
	.w7(32'h3ac4f431),
	.w8(32'hbba63767),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4a102),
	.w1(32'h3ad0b241),
	.w2(32'h3b50127c),
	.w3(32'hbc207ec4),
	.w4(32'hbb9c6d77),
	.w5(32'hbb362230),
	.w6(32'hba639e5b),
	.w7(32'h3b204801),
	.w8(32'h3b5fc4cc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe536),
	.w1(32'h3ad71b0f),
	.w2(32'hbab620d7),
	.w3(32'hbb1c3697),
	.w4(32'h3a1fdec0),
	.w5(32'hbc27fdaf),
	.w6(32'h3c49ccf1),
	.w7(32'h3c4808a3),
	.w8(32'h3bb41689),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a45c5),
	.w1(32'hbad141e4),
	.w2(32'hba7ef467),
	.w3(32'hbbed4a8a),
	.w4(32'hbaa62c7c),
	.w5(32'hba266398),
	.w6(32'h3b191aad),
	.w7(32'h3afa49fd),
	.w8(32'h3b3b7d25),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccd498),
	.w1(32'hbc6459f0),
	.w2(32'hbc8616a3),
	.w3(32'h3adc890c),
	.w4(32'hb97e2005),
	.w5(32'hbacb1dc3),
	.w6(32'h3bbae9cb),
	.w7(32'hbb216091),
	.w8(32'hbbe524df),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868966),
	.w1(32'hbbe487aa),
	.w2(32'hbc4b5f72),
	.w3(32'h3b4cd6fe),
	.w4(32'hbb817b54),
	.w5(32'hbc66b32a),
	.w6(32'hb7b06481),
	.w7(32'hbac4c8a4),
	.w8(32'h39a17e32),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc052013),
	.w1(32'hbbbb712d),
	.w2(32'hba25f8d1),
	.w3(32'hbc207065),
	.w4(32'h3b5ae132),
	.w5(32'h3adb6359),
	.w6(32'hb993a004),
	.w7(32'h3b93d00d),
	.w8(32'h3c0005d0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8add71),
	.w1(32'h3bdcf4b7),
	.w2(32'hbb8a0737),
	.w3(32'h3bd2d55a),
	.w4(32'h3b7b6300),
	.w5(32'h3c67330e),
	.w6(32'h3c132661),
	.w7(32'h3c8079d1),
	.w8(32'h3b9508f0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e152),
	.w1(32'hbc09e142),
	.w2(32'hbc984c90),
	.w3(32'h3c1ce5e4),
	.w4(32'h3b1a9712),
	.w5(32'hbc39de0c),
	.w6(32'h3c387e5b),
	.w7(32'h3b20c208),
	.w8(32'h3b4a1c4c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0a637),
	.w1(32'h3b0da8ba),
	.w2(32'h3b9d7922),
	.w3(32'hbbcbcac4),
	.w4(32'h3a40a310),
	.w5(32'h3b180cae),
	.w6(32'hb9c51cda),
	.w7(32'hb7d266f9),
	.w8(32'hb73b96b7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fbf14),
	.w1(32'hbc3cbfef),
	.w2(32'hbc857dc7),
	.w3(32'h3ac91566),
	.w4(32'hbc529174),
	.w5(32'hbac0f471),
	.w6(32'hbbbc8511),
	.w7(32'hbc9fee08),
	.w8(32'hbcc54928),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49d2e6),
	.w1(32'hbc0e7e1a),
	.w2(32'hbbd8d722),
	.w3(32'h3b136a28),
	.w4(32'h3c1ab0e6),
	.w5(32'h3c2631a1),
	.w6(32'hbc206fd4),
	.w7(32'hbc271a02),
	.w8(32'hbc2a498a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8999f7),
	.w1(32'hbce440e2),
	.w2(32'hbd2453ce),
	.w3(32'h3b3ad83a),
	.w4(32'hbce620f3),
	.w5(32'hbcfe9d14),
	.w6(32'hbbca5341),
	.w7(32'hbcce4ff7),
	.w8(32'hbc3bfa74),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2b4879),
	.w1(32'hbc063691),
	.w2(32'hbce314fa),
	.w3(32'hbb9c3089),
	.w4(32'hbb9123c1),
	.w5(32'hbc82a561),
	.w6(32'h3c442200),
	.w7(32'h3bbc279f),
	.w8(32'h3a3bbf10),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8e119),
	.w1(32'hbb5fd420),
	.w2(32'hba8c9d8f),
	.w3(32'hbc0a387a),
	.w4(32'h3b0a0a4c),
	.w5(32'hb9c5e892),
	.w6(32'hbb96aa1e),
	.w7(32'hbbae3ad5),
	.w8(32'hbbdee058),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b5969),
	.w1(32'h3bb9114d),
	.w2(32'h3b1bb758),
	.w3(32'hba3ed3ae),
	.w4(32'h3c1039ff),
	.w5(32'hbb37f952),
	.w6(32'h3a87ef70),
	.w7(32'h3bba2b68),
	.w8(32'h3ba3f0fe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35161f),
	.w1(32'hbba54eb8),
	.w2(32'hbc430c24),
	.w3(32'hba08d268),
	.w4(32'h3aefd259),
	.w5(32'hbbb621de),
	.w6(32'h3b1aca3a),
	.w7(32'hbc5beff8),
	.w8(32'hbc638b78),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcddb7bb),
	.w1(32'h3b6f6cd7),
	.w2(32'h3c581ef2),
	.w3(32'h3b3c51a9),
	.w4(32'h3c2f31ec),
	.w5(32'h3c7264f4),
	.w6(32'h3b16062b),
	.w7(32'h3c87a5c1),
	.w8(32'h3c17dbd1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a8c67),
	.w1(32'hbbf1ebf6),
	.w2(32'hbcadccc7),
	.w3(32'h3c0effd7),
	.w4(32'hbb23da53),
	.w5(32'hbc5d6cb8),
	.w6(32'h3b5406ca),
	.w7(32'hbc121b55),
	.w8(32'hbc802fc8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb36fdb),
	.w1(32'h3b98383d),
	.w2(32'h3c27478e),
	.w3(32'hbb092203),
	.w4(32'h3c10ab8a),
	.w5(32'h3c11f18d),
	.w6(32'hbb45fcf2),
	.w7(32'h3b275aed),
	.w8(32'h3bf392b7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0dc0c),
	.w1(32'h3b4891a2),
	.w2(32'h3c2236ab),
	.w3(32'h38671541),
	.w4(32'h3745a3f4),
	.w5(32'hbaf8d301),
	.w6(32'h3ca3417b),
	.w7(32'h3c9ece30),
	.w8(32'h3c1ed652),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0efe9e),
	.w1(32'h3b7252b6),
	.w2(32'h3bb70ef9),
	.w3(32'h3bff72eb),
	.w4(32'hbc15a80c),
	.w5(32'hbb169212),
	.w6(32'h3c51fdf4),
	.w7(32'h3c0b6539),
	.w8(32'h3bb77230),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4030ce),
	.w1(32'hbcb4b63e),
	.w2(32'hbbe22167),
	.w3(32'h3cedad21),
	.w4(32'hbc165f54),
	.w5(32'hbc950694),
	.w6(32'hbc6429dc),
	.w7(32'h3c0356ac),
	.w8(32'h3c10612b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99b646),
	.w1(32'hba001df6),
	.w2(32'hbab9e155),
	.w3(32'hbc42004d),
	.w4(32'h3ba70d6a),
	.w5(32'h3af1c7d7),
	.w6(32'h3bf53f5f),
	.w7(32'h3a694ee4),
	.w8(32'h3b3fea71),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba123bb),
	.w1(32'h3af00a27),
	.w2(32'h3bf21cf3),
	.w3(32'h3b07ee55),
	.w4(32'h3aa3ebcd),
	.w5(32'h3b23580b),
	.w6(32'h3a9723bf),
	.w7(32'h3b8d8097),
	.w8(32'h3c7ad9fe),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86a1fe),
	.w1(32'hba8b3489),
	.w2(32'hb9d136fe),
	.w3(32'h3c9a242b),
	.w4(32'hba06f739),
	.w5(32'h3b057d8b),
	.w6(32'hbb9bf4f0),
	.w7(32'h3ac68136),
	.w8(32'hbae98f1d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a80e5),
	.w1(32'h3b63bb47),
	.w2(32'hbbfa66c9),
	.w3(32'h3b25189d),
	.w4(32'hbbac6a77),
	.w5(32'hbb907103),
	.w6(32'hba7bdebe),
	.w7(32'hbb84c8ca),
	.w8(32'hbb9562aa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537afe),
	.w1(32'hbca74a97),
	.w2(32'hbd163052),
	.w3(32'h3b06d84c),
	.w4(32'hbc97cbfd),
	.w5(32'hbca25fcd),
	.w6(32'hbb0e2395),
	.w7(32'hbc918215),
	.w8(32'hbc2c4da6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca84129),
	.w1(32'h3aea8446),
	.w2(32'h3c4115f0),
	.w3(32'hbbc96e5f),
	.w4(32'h3c0e3b2a),
	.w5(32'h3c135c62),
	.w6(32'hbc206be7),
	.w7(32'hbbaae6b6),
	.w8(32'hbb5584cf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d3381),
	.w1(32'h3c1661a5),
	.w2(32'h3c7bbc3e),
	.w3(32'hbb4c8b7c),
	.w4(32'h3be46236),
	.w5(32'h3c198111),
	.w6(32'hbb4896a8),
	.w7(32'h3baa2bd8),
	.w8(32'h3c435491),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c828fae),
	.w1(32'hbc08166d),
	.w2(32'hbbb3dd65),
	.w3(32'h3c177360),
	.w4(32'hbc59709c),
	.w5(32'hbc8463f5),
	.w6(32'hb9511ead),
	.w7(32'hbaa369c1),
	.w8(32'hbc00ad69),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a020e),
	.w1(32'hbb6b176c),
	.w2(32'hbbb24f35),
	.w3(32'hbbfea9a8),
	.w4(32'h3ac60187),
	.w5(32'h3a6a7026),
	.w6(32'hbac5c0dc),
	.w7(32'hbb1f8994),
	.w8(32'h3aa70494),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a600a88),
	.w1(32'h3a7f799a),
	.w2(32'h3a550e54),
	.w3(32'h3bdcf69c),
	.w4(32'hb9f3c442),
	.w5(32'h3b9fb0be),
	.w6(32'h3b1b6618),
	.w7(32'hba260235),
	.w8(32'hbaa5b168),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec3599),
	.w1(32'hbc8b000c),
	.w2(32'hbcc88ee5),
	.w3(32'h38db5d34),
	.w4(32'hbc962aa3),
	.w5(32'hbc90546f),
	.w6(32'h3bd4572e),
	.w7(32'hbb2b5543),
	.w8(32'hbc16e6cf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d887c),
	.w1(32'hbc1f079e),
	.w2(32'hbc9abfe9),
	.w3(32'hbbde4323),
	.w4(32'hbc0841ab),
	.w5(32'hbc8c07db),
	.w6(32'hbbc6fe0a),
	.w7(32'hbc5cd3c6),
	.w8(32'hbc5239e3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd687d0),
	.w1(32'hbbd03698),
	.w2(32'hbb52c1e2),
	.w3(32'hbbaeb089),
	.w4(32'h3bbacbc0),
	.w5(32'h3bcea206),
	.w6(32'h3bfb3838),
	.w7(32'h3c14c4c7),
	.w8(32'h3b8debbb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddbb6f),
	.w1(32'h3bb67a75),
	.w2(32'hbb688416),
	.w3(32'h3be5bcc0),
	.w4(32'hb7908c08),
	.w5(32'hbba32263),
	.w6(32'hb99d16cf),
	.w7(32'h3a199f21),
	.w8(32'hbb5a2717),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b401),
	.w1(32'hbc68ec63),
	.w2(32'hbca16fe0),
	.w3(32'hbacd98a1),
	.w4(32'hbba70b6d),
	.w5(32'hbb7c1d0a),
	.w6(32'hb753cbe0),
	.w7(32'hbb9732a5),
	.w8(32'hbafdaf5b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb250cd),
	.w1(32'hbbefc6e6),
	.w2(32'hbb351b96),
	.w3(32'h3c19dc06),
	.w4(32'hbaa8e40d),
	.w5(32'hb94fb962),
	.w6(32'h3b8208f8),
	.w7(32'h3c0207d6),
	.w8(32'h3b23aeee),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0adff),
	.w1(32'hbc15cce8),
	.w2(32'hbc103312),
	.w3(32'h3bd83d1e),
	.w4(32'hbc2c0e10),
	.w5(32'hbc4ecfda),
	.w6(32'hbaa2969d),
	.w7(32'hbc16ee15),
	.w8(32'hbc352939),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76931c),
	.w1(32'hbb0fd5b3),
	.w2(32'hba80e2da),
	.w3(32'hbc5439bc),
	.w4(32'hbbd46bce),
	.w5(32'hbb223ce2),
	.w6(32'hb92f7511),
	.w7(32'h3b203708),
	.w8(32'hba40fb60),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1294df),
	.w1(32'hbb063f78),
	.w2(32'hba623d9d),
	.w3(32'hba6cd1cf),
	.w4(32'hbacf5411),
	.w5(32'hbbd28a23),
	.w6(32'hbad583fc),
	.w7(32'h3b52330d),
	.w8(32'h393aff50),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05069d),
	.w1(32'h3ccaa494),
	.w2(32'h3d3dd9de),
	.w3(32'h3a789fef),
	.w4(32'h3cd4a619),
	.w5(32'h3cfe3481),
	.w6(32'h3c009584),
	.w7(32'h3cde701e),
	.w8(32'h3cea0970),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce869e2),
	.w1(32'h3d009795),
	.w2(32'h3d531153),
	.w3(32'h3c83f99b),
	.w4(32'h3ccb43e1),
	.w5(32'h3d25a274),
	.w6(32'h3c7eec76),
	.w7(32'h3cce6b3a),
	.w8(32'h3ce30d12),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d283093),
	.w1(32'hbcbee356),
	.w2(32'hbd27e7df),
	.w3(32'h3c958c1b),
	.w4(32'hbcac7323),
	.w5(32'hbcf20261),
	.w6(32'hbb5e5dd6),
	.w7(32'hbc92bb1c),
	.w8(32'hbc9c61d6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e65de),
	.w1(32'hb99e4d5b),
	.w2(32'hbad7e26d),
	.w3(32'hbc8dee59),
	.w4(32'h38c7d26e),
	.w5(32'hb77c654c),
	.w6(32'h3b6c433f),
	.w7(32'h3a464147),
	.w8(32'hbafee7cc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1db3a0),
	.w1(32'h3c62a31c),
	.w2(32'h3bb90c6e),
	.w3(32'hbb6dd014),
	.w4(32'h3adfab14),
	.w5(32'hba9e09f0),
	.w6(32'h3c89b0b8),
	.w7(32'h3c33d6a7),
	.w8(32'h3b34cfaf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928c89c),
	.w1(32'hbac71596),
	.w2(32'h3a157fd3),
	.w3(32'h3a7f98f7),
	.w4(32'hbba7e2bb),
	.w5(32'h3b8e3775),
	.w6(32'h3ac1ee13),
	.w7(32'h3a6d68c1),
	.w8(32'hbbd2f694),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db933),
	.w1(32'hbbe4c033),
	.w2(32'hbcae9947),
	.w3(32'h3b8ed1b6),
	.w4(32'h3b7e097d),
	.w5(32'hbbd50eb9),
	.w6(32'h3ba7ca8b),
	.w7(32'hba424727),
	.w8(32'hbc03d701),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70fa40),
	.w1(32'hbcf9271c),
	.w2(32'hbd5f99bc),
	.w3(32'h3a8a4334),
	.w4(32'hbce5d7c5),
	.w5(32'hbd08092f),
	.w6(32'hbb8ce2a9),
	.w7(32'hbcf09cf5),
	.w8(32'hbcdb4edc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd555ae8),
	.w1(32'hbca0f0c9),
	.w2(32'hbc22d44d),
	.w3(32'hbc8ad67d),
	.w4(32'hbac05362),
	.w5(32'hbbc33292),
	.w6(32'hbc7f9f93),
	.w7(32'h3b83e7a8),
	.w8(32'h3b22a701),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f60e5),
	.w1(32'hbb568f8d),
	.w2(32'hbbd27531),
	.w3(32'h3bdbcbb0),
	.w4(32'hbc016deb),
	.w5(32'hba19eeca),
	.w6(32'hbb4aa907),
	.w7(32'hbb2d8ff2),
	.w8(32'hbc94d5e0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ecbe4),
	.w1(32'hb989015c),
	.w2(32'hbbd90b97),
	.w3(32'h3ac0a945),
	.w4(32'hbad674eb),
	.w5(32'hbb982fb0),
	.w6(32'h3b758950),
	.w7(32'h3b034239),
	.w8(32'hb9dc270a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390221),
	.w1(32'h3b271634),
	.w2(32'h3b9cb88b),
	.w3(32'h3b319369),
	.w4(32'h3aa4beb1),
	.w5(32'h3ae07211),
	.w6(32'h3a91d3ce),
	.w7(32'h3bbca59c),
	.w8(32'h3bbf2bfc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09f6c9),
	.w1(32'hbc6661b8),
	.w2(32'hbcbb08cd),
	.w3(32'h3b23c886),
	.w4(32'hbb27a9bc),
	.w5(32'hbc26c10f),
	.w6(32'hbc29dc77),
	.w7(32'hbb8d7a2c),
	.w8(32'hbc86a21b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad4522),
	.w1(32'h3bb60d94),
	.w2(32'h3ca44508),
	.w3(32'hbc3546aa),
	.w4(32'hbaf195cf),
	.w5(32'h3c0abb26),
	.w6(32'h3b0e2015),
	.w7(32'h3c1fae5d),
	.w8(32'h3ba7bf0b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81c775),
	.w1(32'h3ac0e56c),
	.w2(32'h3baeab2d),
	.w3(32'h3ac057d0),
	.w4(32'h3b6ad1a3),
	.w5(32'h3bda0fb4),
	.w6(32'hbb8fe88e),
	.w7(32'hbc043318),
	.w8(32'hbb5ce36e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085112),
	.w1(32'hbba72afb),
	.w2(32'hbaf625c3),
	.w3(32'h3bf4e645),
	.w4(32'hbaa33206),
	.w5(32'h3b3f676b),
	.w6(32'h3a328fa6),
	.w7(32'h3b56e493),
	.w8(32'h3af899aa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc056),
	.w1(32'hbb8f98f3),
	.w2(32'hbb807a56),
	.w3(32'h3b26848a),
	.w4(32'hbbd70710),
	.w5(32'hbbe73227),
	.w6(32'hbadee767),
	.w7(32'hbb265085),
	.w8(32'h3ab6aadf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb399a12),
	.w1(32'hbb1c1ac8),
	.w2(32'hb988f28d),
	.w3(32'hbbe108f1),
	.w4(32'h391611d3),
	.w5(32'h3b0115f0),
	.w6(32'hba94f71f),
	.w7(32'hbaf9810f),
	.w8(32'hbad10080),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa03381),
	.w1(32'hbc0c5ccf),
	.w2(32'hbc96a901),
	.w3(32'h3b1bcd22),
	.w4(32'hbc6f3637),
	.w5(32'hbc38e64a),
	.w6(32'hbb84edb0),
	.w7(32'hbc2a77a5),
	.w8(32'hbc52336b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e913b),
	.w1(32'h3a89368d),
	.w2(32'h3c811d30),
	.w3(32'hbbde38c5),
	.w4(32'h3c450af9),
	.w5(32'h3c43530b),
	.w6(32'h3c34e04b),
	.w7(32'h3c5f2f97),
	.w8(32'h3c73d61a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83e8d4),
	.w1(32'h3c95380c),
	.w2(32'h3bda6ab5),
	.w3(32'h3c92c7b7),
	.w4(32'h3c489469),
	.w5(32'h3c201ee1),
	.w6(32'h3c2a2767),
	.w7(32'h3c71ae0f),
	.w8(32'h3c31cd00),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf51dba),
	.w1(32'hbbcb5988),
	.w2(32'hbc1f9436),
	.w3(32'h3b976e80),
	.w4(32'hbad3c405),
	.w5(32'hbb8b345a),
	.w6(32'hba60fc34),
	.w7(32'h3a8c19de),
	.w8(32'hba2ad139),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bbbeb),
	.w1(32'h3d36f784),
	.w2(32'h3d979bf9),
	.w3(32'hbb8b86db),
	.w4(32'h3d17851a),
	.w5(32'h3d30e8ee),
	.w6(32'hbb3ee7e3),
	.w7(32'h3ce1d2c2),
	.w8(32'h3d122db1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3aad56),
	.w1(32'h3b92c7f7),
	.w2(32'hba0bc828),
	.w3(32'h3c89e773),
	.w4(32'hba7fd49c),
	.w5(32'h3ad2237d),
	.w6(32'h3a87bb54),
	.w7(32'hbb0ac99b),
	.w8(32'hbb8dbb51),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017cc0),
	.w1(32'hbca3694b),
	.w2(32'hbd22e3e2),
	.w3(32'hba9866b4),
	.w4(32'hbcd6d51e),
	.w5(32'hbd035ee4),
	.w6(32'hbb31362d),
	.w7(32'hbc4a62d7),
	.w8(32'hbcb1fa7b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee37fc),
	.w1(32'hbcd2c3dd),
	.w2(32'hbd143e62),
	.w3(32'hbc5683c6),
	.w4(32'hbd17aeea),
	.w5(32'hbcc760ba),
	.w6(32'hbc35bf05),
	.w7(32'hbcaa9696),
	.w8(32'hbca60c88),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa9b53),
	.w1(32'hbc2a8f54),
	.w2(32'hb9b0c650),
	.w3(32'hbb4d3f74),
	.w4(32'hbb510a72),
	.w5(32'hbb3bfb0f),
	.w6(32'hbc51a1c7),
	.w7(32'hbbf1b135),
	.w8(32'hbbcb0bcd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83290),
	.w1(32'h3b31e055),
	.w2(32'hb9fb9dbf),
	.w3(32'hbb004d36),
	.w4(32'hbb12441a),
	.w5(32'h3a66863f),
	.w6(32'hbae6cc76),
	.w7(32'hbab52953),
	.w8(32'hbb92db2e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1820),
	.w1(32'hbc84c201),
	.w2(32'hbcf73e98),
	.w3(32'hbb1a9180),
	.w4(32'hbcb41502),
	.w5(32'hbcd88e2a),
	.w6(32'hb9076ce9),
	.w7(32'hbc846056),
	.w8(32'hbcdb61b8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9ffed),
	.w1(32'h3c408ce0),
	.w2(32'h3bd4bdb0),
	.w3(32'h3a6615ad),
	.w4(32'h3a473139),
	.w5(32'h3b327a18),
	.w6(32'h3ba9ad65),
	.w7(32'h3b543df1),
	.w8(32'h3af8c2c5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb281e3),
	.w1(32'h3abab5b0),
	.w2(32'h38dae409),
	.w3(32'h3b9e3c11),
	.w4(32'h39e840b3),
	.w5(32'hba50c66f),
	.w6(32'h3c1247f7),
	.w7(32'h3c0d52d3),
	.w8(32'h3c014acb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb610bf9),
	.w1(32'hbc6cff16),
	.w2(32'hbcd623dc),
	.w3(32'h3bd58fa6),
	.w4(32'hbbe41b48),
	.w5(32'hbbc100d6),
	.w6(32'h3b048d96),
	.w7(32'hbbc54466),
	.w8(32'hbc133596),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a4072),
	.w1(32'h3bc8d648),
	.w2(32'hba9bd561),
	.w3(32'hb97fc959),
	.w4(32'hbc3101b0),
	.w5(32'hbc42743d),
	.w6(32'hbb95a6a0),
	.w7(32'hb9df0670),
	.w8(32'hbb1cba80),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d2cb),
	.w1(32'hbc33767e),
	.w2(32'hbca22a20),
	.w3(32'hbc1da7cf),
	.w4(32'hbc81d2f9),
	.w5(32'hbc944d3e),
	.w6(32'hbc3583da),
	.w7(32'hbc4b026f),
	.w8(32'hbc6f8494),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67f28b),
	.w1(32'h3c861e0a),
	.w2(32'h3c9062a1),
	.w3(32'hbbd86c22),
	.w4(32'h3c774dce),
	.w5(32'h3c0db858),
	.w6(32'h3c1a2e96),
	.w7(32'h3c187558),
	.w8(32'h3c9e090e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9f557),
	.w1(32'hbcbfe817),
	.w2(32'hbd0396e1),
	.w3(32'hb9df969f),
	.w4(32'hbc9a9aa1),
	.w5(32'hbcb986ab),
	.w6(32'h3b17749e),
	.w7(32'hbc4be6a5),
	.w8(32'hbc359f61),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcea57ef),
	.w1(32'hbcb13e59),
	.w2(32'hbcecc10c),
	.w3(32'hbcb47b78),
	.w4(32'hbc169bf3),
	.w5(32'hbc28903e),
	.w6(32'h3ba29835),
	.w7(32'h3ae2bf78),
	.w8(32'hbc4d5e4c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3857ab),
	.w1(32'hbcef94ed),
	.w2(32'hbd08fa86),
	.w3(32'h3b949e83),
	.w4(32'hbce5eb65),
	.w5(32'hbcbd388e),
	.w6(32'hb96ba3d1),
	.w7(32'hbb90d737),
	.w8(32'h38363f99),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc89194),
	.w1(32'h3b842199),
	.w2(32'h3c5908b8),
	.w3(32'hbc7c3e68),
	.w4(32'h3c1c12f7),
	.w5(32'h3c4fbac8),
	.w6(32'h3b2c41ec),
	.w7(32'h3adc24ef),
	.w8(32'h3a87eccd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca24deb),
	.w1(32'h3b81049e),
	.w2(32'hb9eb2260),
	.w3(32'h3c199526),
	.w4(32'h3c09d987),
	.w5(32'h3b1aa353),
	.w6(32'h3bb487e1),
	.w7(32'h3b4763a1),
	.w8(32'h3b862b27),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9934),
	.w1(32'h3b7d010a),
	.w2(32'hbaf61327),
	.w3(32'h3c0057bb),
	.w4(32'h3c5637a8),
	.w5(32'h3c001799),
	.w6(32'h3b490f8f),
	.w7(32'h3add5e28),
	.w8(32'h3b0c5ddb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f041b),
	.w1(32'hbaec0e28),
	.w2(32'h3aa21f69),
	.w3(32'h39b8c721),
	.w4(32'h3b982fda),
	.w5(32'h3ba4d9c5),
	.w6(32'hbb573a98),
	.w7(32'hb83c4112),
	.w8(32'h3b1b2008),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf05719),
	.w1(32'h3c9e6c55),
	.w2(32'h3cfbf358),
	.w3(32'h3c256e56),
	.w4(32'h3c7d4a0e),
	.w5(32'h3c7e1707),
	.w6(32'h396f200c),
	.w7(32'h3c89c1f4),
	.w8(32'h3c79614a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93aa2c),
	.w1(32'hbcddeb06),
	.w2(32'hbd13f3ef),
	.w3(32'h3bd3423e),
	.w4(32'hbcfe2fb7),
	.w5(32'hbcf72b2a),
	.w6(32'hbbdd299d),
	.w7(32'hbc8710d6),
	.w8(32'hbbfdd666),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb79c9a),
	.w1(32'h3c50e641),
	.w2(32'h3c8b35b4),
	.w3(32'hbb6552a6),
	.w4(32'h3c4338b1),
	.w5(32'h3c039a88),
	.w6(32'h3a6b2d4c),
	.w7(32'h3bb98734),
	.w8(32'h3c053595),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ea691),
	.w1(32'h3b1375ab),
	.w2(32'h3a886ac4),
	.w3(32'h3bbf2554),
	.w4(32'h39a9056b),
	.w5(32'h3a68b537),
	.w6(32'h3b1f1ed4),
	.w7(32'h3ace824c),
	.w8(32'h3aea25d7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af86c3a),
	.w1(32'h3ab2bb0a),
	.w2(32'h3897ac1f),
	.w3(32'h3ba2c800),
	.w4(32'h3b5df65a),
	.w5(32'h3b54285c),
	.w6(32'h3be8d7f7),
	.w7(32'h3bbec9b2),
	.w8(32'h3afa505f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295f25),
	.w1(32'hbbf9f4e3),
	.w2(32'hbc51d515),
	.w3(32'h3b9e93ca),
	.w4(32'hbb8d6cc9),
	.w5(32'hbc1f6485),
	.w6(32'hbad067e6),
	.w7(32'hbbcc444c),
	.w8(32'hbaf3218b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291064),
	.w1(32'hbb6a7cd7),
	.w2(32'h3afab1e7),
	.w3(32'hbb8d2cd4),
	.w4(32'hbb5ff747),
	.w5(32'hb97f43b3),
	.w6(32'hba76b4a2),
	.w7(32'h3b3fa5ab),
	.w8(32'hb9d9fd3e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9819b22),
	.w1(32'hb8f78f9b),
	.w2(32'h3c2841f4),
	.w3(32'h3b0f4861),
	.w4(32'h3bad29c1),
	.w5(32'h3c484b93),
	.w6(32'h3bf15b30),
	.w7(32'h3c1aa72f),
	.w8(32'h3bca99e1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49d57a),
	.w1(32'hbc49f5a3),
	.w2(32'hbd081c08),
	.w3(32'h3a90234a),
	.w4(32'hbcdf3e06),
	.w5(32'hbcb44c3c),
	.w6(32'h3bfca46c),
	.w7(32'hbc2cb56b),
	.w8(32'hbc3aad54),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc93fda),
	.w1(32'hbc69a74f),
	.w2(32'hbc87bdb5),
	.w3(32'hbb66d5fc),
	.w4(32'hbc93bdd5),
	.w5(32'hbbca7236),
	.w6(32'h3afe67c0),
	.w7(32'h3bcdbdf2),
	.w8(32'hbb982a16),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8820),
	.w1(32'hbcaf43a0),
	.w2(32'hbcf7a74e),
	.w3(32'h3a60179d),
	.w4(32'hbcb84924),
	.w5(32'hbc42180b),
	.w6(32'h393c56ff),
	.w7(32'hbc1f77d1),
	.w8(32'hbc8db54f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd4399),
	.w1(32'hbcc28132),
	.w2(32'hbcf91269),
	.w3(32'hbb1a7a9c),
	.w4(32'hbc013ebf),
	.w5(32'hbcbf5065),
	.w6(32'hbba8d0b3),
	.w7(32'hbba55a73),
	.w8(32'h3aa71977),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f46eb),
	.w1(32'hbc1d21e4),
	.w2(32'hbc96274e),
	.w3(32'hbb98615e),
	.w4(32'hbc1d9dc9),
	.w5(32'hbb3c78cd),
	.w6(32'h3af15203),
	.w7(32'hbc2d78c9),
	.w8(32'hbb99039a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc502c2),
	.w1(32'h3cde604a),
	.w2(32'h3cef9592),
	.w3(32'hbac83a7c),
	.w4(32'h3cda702c),
	.w5(32'h3d010cbd),
	.w6(32'h3c57b189),
	.w7(32'h3cba5ef1),
	.w8(32'h3c9833be),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdefe05),
	.w1(32'h3c8ef140),
	.w2(32'h3c836feb),
	.w3(32'h3ca9803f),
	.w4(32'h3c40ede1),
	.w5(32'h3c91d291),
	.w6(32'h3c282e55),
	.w7(32'h3c556406),
	.w8(32'h3bda4e9a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73d4ab),
	.w1(32'hbc8c71a8),
	.w2(32'hbcd092b9),
	.w3(32'h3b68c0af),
	.w4(32'hbc8cc942),
	.w5(32'hbc9a5060),
	.w6(32'hbb17fb0b),
	.w7(32'hbc5e83c8),
	.w8(32'hbc5d4141),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38345f),
	.w1(32'h3ba34c75),
	.w2(32'h3c503574),
	.w3(32'h3c034881),
	.w4(32'hbb619e04),
	.w5(32'h3b6224fc),
	.w6(32'hbb17eb01),
	.w7(32'h3bd12213),
	.w8(32'h3aa74dd7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eafbb),
	.w1(32'hba2b31e1),
	.w2(32'h3c36427e),
	.w3(32'h3b2b6058),
	.w4(32'h3bce41af),
	.w5(32'h3bf4ec4f),
	.w6(32'hbc3f35f7),
	.w7(32'hba20da7c),
	.w8(32'hbadb9396),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9dd07),
	.w1(32'hbc5593dc),
	.w2(32'hbc9cf29f),
	.w3(32'h3b65d34a),
	.w4(32'hbb96bf94),
	.w5(32'hbb92eb89),
	.w6(32'h3a5b2d51),
	.w7(32'hbb94d345),
	.w8(32'hbbf91bc7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f07d),
	.w1(32'h3b400e3a),
	.w2(32'hb99cd122),
	.w3(32'h3bd36758),
	.w4(32'hbbe3501e),
	.w5(32'hba8b713d),
	.w6(32'hbbf55372),
	.w7(32'hbb94f041),
	.w8(32'hbb7eb2b0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba650aa),
	.w1(32'h38976a4c),
	.w2(32'hba3d0bd7),
	.w3(32'hbc17f0a7),
	.w4(32'h3b11b634),
	.w5(32'h3b922d64),
	.w6(32'h3ba32584),
	.w7(32'h3b4fc9f1),
	.w8(32'hba442c52),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b643c5c),
	.w1(32'h3c9681fd),
	.w2(32'h3c5b9dc4),
	.w3(32'h3b89f451),
	.w4(32'h3cc66669),
	.w5(32'h3c73b268),
	.w6(32'h3c78caf0),
	.w7(32'h3ccbff1a),
	.w8(32'h3c22f0f9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958191),
	.w1(32'hbbf8395c),
	.w2(32'hbbc203e9),
	.w3(32'h3c94004e),
	.w4(32'hbbf177b1),
	.w5(32'hbc020788),
	.w6(32'hbbaf1054),
	.w7(32'hbbe24837),
	.w8(32'hbbb759f7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962a1ea),
	.w1(32'h3c15afab),
	.w2(32'hbc152005),
	.w3(32'hbbf18bf2),
	.w4(32'h3af91779),
	.w5(32'hbc148726),
	.w6(32'h33eb2d00),
	.w7(32'hbb84a457),
	.w8(32'hbb74e9c3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8154),
	.w1(32'hbc18a96d),
	.w2(32'hbba6f2d9),
	.w3(32'h3a396191),
	.w4(32'hbbb8b127),
	.w5(32'hb999f3db),
	.w6(32'h3af32c51),
	.w7(32'hbb6fc558),
	.w8(32'hbc18db3d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288058),
	.w1(32'hb9dd0d4e),
	.w2(32'hbbce1caf),
	.w3(32'h3bc9df87),
	.w4(32'h3ba976ab),
	.w5(32'h3af3377a),
	.w6(32'h3a81df47),
	.w7(32'h3a4155c7),
	.w8(32'hba946c24),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e4c9),
	.w1(32'h390dd7c7),
	.w2(32'hb9f3cf08),
	.w3(32'h3c02fc30),
	.w4(32'h3a89cee2),
	.w5(32'h3b87316b),
	.w6(32'h3b2821ed),
	.w7(32'h39ebccb3),
	.w8(32'hbab24151),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9caf86),
	.w1(32'h3c454673),
	.w2(32'h3c4dde75),
	.w3(32'h3b8fff55),
	.w4(32'h3c1bf69c),
	.w5(32'h3c11d9f5),
	.w6(32'h3b33f8de),
	.w7(32'h3b4ac6ec),
	.w8(32'h3ba80fa4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19ffc8),
	.w1(32'h3b09f688),
	.w2(32'hbab93da3),
	.w3(32'h3bd2e73b),
	.w4(32'h3ba9ef4d),
	.w5(32'h3b187e6b),
	.w6(32'hba5a9e9e),
	.w7(32'h39c5d76e),
	.w8(32'h3b1155be),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b520b4b),
	.w1(32'hbcae608b),
	.w2(32'hbd0ae387),
	.w3(32'hbad4ff18),
	.w4(32'hbc6900ff),
	.w5(32'hbcc232c3),
	.w6(32'hbbc0bc0a),
	.w7(32'hbc7c8dbc),
	.w8(32'hbc78e7ef),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd023856),
	.w1(32'h3bd41e38),
	.w2(32'h3ac47fbe),
	.w3(32'hbca767e7),
	.w4(32'hbb623220),
	.w5(32'hbb96b64e),
	.w6(32'h3ae6ba2e),
	.w7(32'h3b599ff6),
	.w8(32'hb9c92cfb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb3d6),
	.w1(32'hbc221a45),
	.w2(32'hbc1b21fc),
	.w3(32'hbc19220a),
	.w4(32'h3c2d2a53),
	.w5(32'h3ba5c0f1),
	.w6(32'hbc0f37d4),
	.w7(32'hbc406fa6),
	.w8(32'h39fb4850),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17fbd),
	.w1(32'hbc8a2d9b),
	.w2(32'hbc73209d),
	.w3(32'hbc6e3e3a),
	.w4(32'hbc7e4a2d),
	.w5(32'hbc5af8a8),
	.w6(32'hbc05e992),
	.w7(32'hbc38059e),
	.w8(32'hbc55ce1e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a99c6),
	.w1(32'hbb81e994),
	.w2(32'hbb35c2c4),
	.w3(32'hbbcd3676),
	.w4(32'hbc0811d3),
	.w5(32'hbb3fe473),
	.w6(32'hbaf5d323),
	.w7(32'hba047314),
	.w8(32'hbb5ea981),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bc168),
	.w1(32'hbbbf2572),
	.w2(32'hbc16f795),
	.w3(32'h3a76e04b),
	.w4(32'h3b531423),
	.w5(32'hbaddf05e),
	.w6(32'h3b87dc76),
	.w7(32'hba24cc4f),
	.w8(32'hbb866232),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb85b0a),
	.w1(32'hbc541451),
	.w2(32'hbcb72929),
	.w3(32'hbb8246ad),
	.w4(32'hbbeeb85f),
	.w5(32'hbc368c4a),
	.w6(32'hbb02b86b),
	.w7(32'hbc19ef20),
	.w8(32'hbc1ab019),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ff748),
	.w1(32'h3cd3b7db),
	.w2(32'h3d2f7261),
	.w3(32'hbc0fb9c7),
	.w4(32'h3ca3dda0),
	.w5(32'h3ce6d8b4),
	.w6(32'h3c418c07),
	.w7(32'h3cb6317f),
	.w8(32'h3cecd530),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce39bfd),
	.w1(32'hbb016187),
	.w2(32'hbb965e91),
	.w3(32'h3c642c68),
	.w4(32'h39d1bc91),
	.w5(32'hbb148847),
	.w6(32'hbad63938),
	.w7(32'hbb3ea152),
	.w8(32'hbae8394a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989e278),
	.w1(32'hbb6b4026),
	.w2(32'hbaa0c8b5),
	.w3(32'h3a6dc93e),
	.w4(32'h3adcb44e),
	.w5(32'h3b245cef),
	.w6(32'h3afb49c4),
	.w7(32'hb8f2013a),
	.w8(32'hbbcb0c7b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule