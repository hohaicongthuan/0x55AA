module layer_8_featuremap_166(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad1b8),
	.w1(32'h3b02503b),
	.w2(32'h3bba5a1b),
	.w3(32'hbaebbe70),
	.w4(32'h3b8d8717),
	.w5(32'h3b7e2c3f),
	.w6(32'h3a3764b9),
	.w7(32'h3b5cbb66),
	.w8(32'h3ad0b6df),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294475),
	.w1(32'h3ca82da1),
	.w2(32'h3d6d6189),
	.w3(32'hbaacbb43),
	.w4(32'hbb9d9cd1),
	.w5(32'h3cdaf1ec),
	.w6(32'hbc592f94),
	.w7(32'h3c80493b),
	.w8(32'hbb441681),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c3242),
	.w1(32'hbbbd80b9),
	.w2(32'hbb69840b),
	.w3(32'h3b799e4c),
	.w4(32'hbb053d78),
	.w5(32'h3b172760),
	.w6(32'hbb996490),
	.w7(32'h38986e1f),
	.w8(32'hba2fdace),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999fd07),
	.w1(32'hbb86c6a6),
	.w2(32'hba028e34),
	.w3(32'hb8744a69),
	.w4(32'hbaf8e199),
	.w5(32'hba5d0fbc),
	.w6(32'hbb81ce8a),
	.w7(32'hbb258a6d),
	.w8(32'hbba0d858),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53de98),
	.w1(32'h3ca9da7e),
	.w2(32'h3d8b3d1a),
	.w3(32'hbb46a01f),
	.w4(32'hbb386c5b),
	.w5(32'h3d0f9fbd),
	.w6(32'hbc82cfc0),
	.w7(32'h3c575993),
	.w8(32'hbaccc03d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d31bc82),
	.w1(32'hbbd4292f),
	.w2(32'hbb73b6b5),
	.w3(32'h3c62d9c1),
	.w4(32'hbb012720),
	.w5(32'h3bddbee9),
	.w6(32'h39bc1e3a),
	.w7(32'h3acc0007),
	.w8(32'h3b9a45b5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c513fca),
	.w1(32'hbb6ba51b),
	.w2(32'hbc6b236f),
	.w3(32'h3c064fb5),
	.w4(32'h3bf8476c),
	.w5(32'hbb241333),
	.w6(32'h3bedd149),
	.w7(32'hbb01eace),
	.w8(32'h3bcb350b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb17ce),
	.w1(32'h3b7979d2),
	.w2(32'h3b967998),
	.w3(32'h3c00851c),
	.w4(32'hb7bd3cac),
	.w5(32'h3b9cfcd9),
	.w6(32'hbb1daed4),
	.w7(32'hbb07d2fd),
	.w8(32'hbbcd6edb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964181),
	.w1(32'h3d18441b),
	.w2(32'h3dc17482),
	.w3(32'hba966d35),
	.w4(32'h3c3b4c5f),
	.w5(32'h3d7d45d3),
	.w6(32'hbc87225c),
	.w7(32'h3cd6d04d),
	.w8(32'h3be61453),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d842a5e),
	.w1(32'h3b55b32a),
	.w2(32'h3c1245d4),
	.w3(32'h3d0efa7b),
	.w4(32'h3aa58928),
	.w5(32'h3b6048e3),
	.w6(32'hbb8c3352),
	.w7(32'h3bf9b0f4),
	.w8(32'h3bd45086),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9151fe),
	.w1(32'hbc28c26f),
	.w2(32'hbb26bd53),
	.w3(32'h3b93fc3d),
	.w4(32'hbc1b9dc3),
	.w5(32'hbbd930e3),
	.w6(32'hbca0fcc3),
	.w7(32'hbc5c530b),
	.w8(32'hbc8d30dd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d7ac),
	.w1(32'h3b2177c8),
	.w2(32'h3b9f2ff8),
	.w3(32'hbc0f3619),
	.w4(32'h3c0740f5),
	.w5(32'h3be41068),
	.w6(32'h3bc6f1de),
	.w7(32'h3bd0276f),
	.w8(32'h3c17c96c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba077c4),
	.w1(32'hbb99e3e7),
	.w2(32'h3b139a84),
	.w3(32'h3bc92f60),
	.w4(32'hbbc51a90),
	.w5(32'hba670ed4),
	.w6(32'hbc286f8e),
	.w7(32'hbb48d9f7),
	.w8(32'hba934200),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9fb17),
	.w1(32'h3b3ea755),
	.w2(32'h3b865e99),
	.w3(32'hba5ef73d),
	.w4(32'hbab21e06),
	.w5(32'h3ae5dbec),
	.w6(32'h3abed773),
	.w7(32'hbb0a836a),
	.w8(32'hb9ab353a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33251b),
	.w1(32'hbd337b8e),
	.w2(32'hbdac860b),
	.w3(32'h3b1cbfc1),
	.w4(32'hbc8d0582),
	.w5(32'hbd4a004e),
	.w6(32'hbc8d7309),
	.w7(32'hbd260b34),
	.w8(32'hbcabb08d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6817e1),
	.w1(32'hba2434b7),
	.w2(32'h3bc450bd),
	.w3(32'hbcadce56),
	.w4(32'hba94653f),
	.w5(32'h3b9bb7b8),
	.w6(32'hbbbec231),
	.w7(32'h3b47a367),
	.w8(32'h3babc51b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3dcf87),
	.w1(32'hbb0a633f),
	.w2(32'h3ad15fc5),
	.w3(32'h3ba04875),
	.w4(32'hbb68a209),
	.w5(32'hbb884b83),
	.w6(32'hbb82257c),
	.w7(32'h39951d0f),
	.w8(32'hbb5485ad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd8927),
	.w1(32'hbbbe8b1c),
	.w2(32'hb977ca9b),
	.w3(32'hbbba1773),
	.w4(32'hbb05919d),
	.w5(32'hbb208187),
	.w6(32'hbb665e92),
	.w7(32'hbb9975c0),
	.w8(32'hbb91169b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8744d),
	.w1(32'hb9c0d703),
	.w2(32'h3bf3846f),
	.w3(32'hbb351720),
	.w4(32'h39cf06b8),
	.w5(32'h3c482017),
	.w6(32'hbb0ccc0d),
	.w7(32'h3b3938fe),
	.w8(32'h3b691f5d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4fd60),
	.w1(32'hbc751d34),
	.w2(32'hbd38b539),
	.w3(32'h3adbc02e),
	.w4(32'h3c111496),
	.w5(32'hbc8a3fac),
	.w6(32'h3bf95db1),
	.w7(32'hbc835c4a),
	.w8(32'h3a5c1284),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbef461),
	.w1(32'hbc4043b7),
	.w2(32'hbc6ce172),
	.w3(32'h3b6236f4),
	.w4(32'hbbaff732),
	.w5(32'hbc23cf5a),
	.w6(32'hbba34baf),
	.w7(32'h3ab6e629),
	.w8(32'hbb3f8843),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29c7a8),
	.w1(32'hbb42d7be),
	.w2(32'h3bee91cf),
	.w3(32'hbc12d54d),
	.w4(32'h3b4cd9e5),
	.w5(32'h3bc71719),
	.w6(32'hbb4b9542),
	.w7(32'h3963589c),
	.w8(32'h3b422369),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17a9eb),
	.w1(32'hbaab5369),
	.w2(32'hba927c76),
	.w3(32'hb95a2f1c),
	.w4(32'h3b07e0f8),
	.w5(32'hbae03a83),
	.w6(32'hbb82e734),
	.w7(32'hbb448d02),
	.w8(32'hbbdc8e14),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dedf12),
	.w1(32'hbbd4941e),
	.w2(32'hb8fc1aa4),
	.w3(32'hbb8b53de),
	.w4(32'h3a835a3d),
	.w5(32'h3b2bea09),
	.w6(32'h3b6e9738),
	.w7(32'hbb183bdc),
	.w8(32'hbb8a96c1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73950c),
	.w1(32'h3a845ead),
	.w2(32'h3ac9ef33),
	.w3(32'hbb43a676),
	.w4(32'hba909c60),
	.w5(32'h3a31a6b2),
	.w6(32'hbab87c74),
	.w7(32'hbb5dfa1a),
	.w8(32'hbbdd11c7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb8e89),
	.w1(32'hbb149e6f),
	.w2(32'hbbb61794),
	.w3(32'hbb111ad3),
	.w4(32'hba22ebfa),
	.w5(32'hbb732a87),
	.w6(32'h393dd09d),
	.w7(32'hb95746e1),
	.w8(32'hba9049af),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f06e),
	.w1(32'h39befe97),
	.w2(32'h3c135486),
	.w3(32'hbba54487),
	.w4(32'hba0ad93d),
	.w5(32'h3b615338),
	.w6(32'hbb61cbf0),
	.w7(32'hbae9babd),
	.w8(32'hbb763e1b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c106ddd),
	.w1(32'hbb8fe3ed),
	.w2(32'hba8d7143),
	.w3(32'h3c2f35b7),
	.w4(32'hbbceef03),
	.w5(32'hbb298351),
	.w6(32'hbb3b3424),
	.w7(32'hbb1bf991),
	.w8(32'hbb522fc6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995d69e),
	.w1(32'hbb93949a),
	.w2(32'h3b57f7e7),
	.w3(32'hbbae0ce9),
	.w4(32'hbb70ce50),
	.w5(32'h3bb63e3a),
	.w6(32'hbc9abfbb),
	.w7(32'hbb8cc120),
	.w8(32'hbc75aac8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd929f9),
	.w1(32'h3c7c4f83),
	.w2(32'h3cc3b368),
	.w3(32'hbba54d55),
	.w4(32'h3c8e6e62),
	.w5(32'h3cad3eb8),
	.w6(32'h3c19053b),
	.w7(32'h3c936531),
	.w8(32'h3ca1ab3a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce035fc),
	.w1(32'hbb40829a),
	.w2(32'h3b606b83),
	.w3(32'h3cd742cb),
	.w4(32'hbbeae114),
	.w5(32'hba8a17ab),
	.w6(32'hbbf8f223),
	.w7(32'hbaace36a),
	.w8(32'hbba67ab5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f33d6),
	.w1(32'hbc3b4e93),
	.w2(32'h3b49d667),
	.w3(32'hbb8cf8ad),
	.w4(32'hbc18533f),
	.w5(32'hba827d5b),
	.w6(32'hbcc0a90c),
	.w7(32'hbc592b66),
	.w8(32'hbc1444bc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b57f4),
	.w1(32'hbaee8610),
	.w2(32'h3bce7caf),
	.w3(32'hbb84361d),
	.w4(32'hbb5140b0),
	.w5(32'h3b78a10f),
	.w6(32'hb88ffda1),
	.w7(32'h37a57374),
	.w8(32'h3b82bc69),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc92f1),
	.w1(32'h3a434695),
	.w2(32'hbb0f73a1),
	.w3(32'h3b0c7785),
	.w4(32'hbb4ef07f),
	.w5(32'hbb3644b5),
	.w6(32'hbba58af6),
	.w7(32'hbad56292),
	.w8(32'hbaa3b3a8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ba84),
	.w1(32'h3c1184d3),
	.w2(32'h3c3934a8),
	.w3(32'hba916928),
	.w4(32'h3b4ab26c),
	.w5(32'h3bc5c480),
	.w6(32'hb9d3efeb),
	.w7(32'h3bcbfd3a),
	.w8(32'hbb0da678),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c7b5),
	.w1(32'h3b981b78),
	.w2(32'h3b7ee04f),
	.w3(32'h3b52c17e),
	.w4(32'hbb9c8c4a),
	.w5(32'h3a5540e6),
	.w6(32'hbb15bd2d),
	.w7(32'hbae33992),
	.w8(32'h3b51a922),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9820d),
	.w1(32'hbabe8e77),
	.w2(32'h3b42a0c2),
	.w3(32'hbb42f13c),
	.w4(32'hbb2affb9),
	.w5(32'hb8164a4d),
	.w6(32'hbac67832),
	.w7(32'h3aa3017f),
	.w8(32'hb8bafb84),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e720d1),
	.w1(32'hbc7ee544),
	.w2(32'hbce94261),
	.w3(32'hb9569a45),
	.w4(32'hbc4b422a),
	.w5(32'hbcbe7a54),
	.w6(32'hbc741a13),
	.w7(32'hbc92c8e8),
	.w8(32'hbc396cd2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a3b50),
	.w1(32'hbb1615be),
	.w2(32'h3bf15280),
	.w3(32'hbc0aa4e5),
	.w4(32'hbb3e6a4b),
	.w5(32'h3b37fc2f),
	.w6(32'hbb3b88fa),
	.w7(32'h3b36507c),
	.w8(32'hba254d72),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728c80),
	.w1(32'hb9f8f0bb),
	.w2(32'hba901121),
	.w3(32'hba032311),
	.w4(32'hbabeab46),
	.w5(32'hbc002815),
	.w6(32'h3ad8688b),
	.w7(32'h3b3b5383),
	.w8(32'hba19528d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba858d78),
	.w1(32'h3be13481),
	.w2(32'h3bcad685),
	.w3(32'hba75d315),
	.w4(32'h3baa6842),
	.w5(32'h3b83cb21),
	.w6(32'h3bd23e3b),
	.w7(32'h3c077830),
	.w8(32'h3b808916),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1c32),
	.w1(32'hba42c1e4),
	.w2(32'h3beb9ed2),
	.w3(32'h3aa42918),
	.w4(32'hb9705c5d),
	.w5(32'h3bb62bf0),
	.w6(32'hbbd17c0c),
	.w7(32'hbbb306ee),
	.w8(32'hbb15463b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132184),
	.w1(32'hba72f06f),
	.w2(32'hbb5edd79),
	.w3(32'h3b6d5aee),
	.w4(32'hbabb28cd),
	.w5(32'hbba38d9b),
	.w6(32'hbb25044d),
	.w7(32'hbb1b97d6),
	.w8(32'hbb42943a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf1fd),
	.w1(32'h3aca3591),
	.w2(32'h3b81617d),
	.w3(32'hbb67097a),
	.w4(32'hbb777f42),
	.w5(32'h3bad6ee8),
	.w6(32'hbba626d0),
	.w7(32'h3aaff527),
	.w8(32'hbb978861),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbc7cc),
	.w1(32'hbb1de7aa),
	.w2(32'h3c2c7d79),
	.w3(32'hbae6d418),
	.w4(32'hba087b4c),
	.w5(32'h3b4ed4ce),
	.w6(32'hbbbac693),
	.w7(32'h39734de3),
	.w8(32'hbc0e7e74),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e84c7f),
	.w1(32'hbba303ff),
	.w2(32'hbb7240f4),
	.w3(32'h3b03b044),
	.w4(32'hbb7d99e9),
	.w5(32'h39a5c27c),
	.w6(32'hbb8ec631),
	.w7(32'h3a07a212),
	.w8(32'hbbd9cc88),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15eabf),
	.w1(32'hbb491b32),
	.w2(32'hbba51198),
	.w3(32'hbba45b19),
	.w4(32'h3a4c0db6),
	.w5(32'hbb3972e9),
	.w6(32'hbbab6a2a),
	.w7(32'hbb1e7a54),
	.w8(32'hbab06d58),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984bab),
	.w1(32'hba9af35a),
	.w2(32'hb9a135a9),
	.w3(32'hba958160),
	.w4(32'h3a50f59e),
	.w5(32'hbb963ddb),
	.w6(32'hbaa47e14),
	.w7(32'h3b81230b),
	.w8(32'hbb755d69),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405a81),
	.w1(32'hbac6a1c8),
	.w2(32'h3a2d2059),
	.w3(32'h3ae7d9e5),
	.w4(32'h3aa0173c),
	.w5(32'h3a896312),
	.w6(32'hbb90d140),
	.w7(32'hbbb1104d),
	.w8(32'hbb880a21),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e77ca),
	.w1(32'hbb47e8d6),
	.w2(32'hbc065136),
	.w3(32'hbb8e0eda),
	.w4(32'hbb87f231),
	.w5(32'hbb80e21e),
	.w6(32'hbb1578b5),
	.w7(32'h38a248e7),
	.w8(32'h3b7e91fc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9007df),
	.w1(32'h3bcf4869),
	.w2(32'hbc133138),
	.w3(32'hbb7de784),
	.w4(32'hbaaf8731),
	.w5(32'hbc442d69),
	.w6(32'h3b9cd95d),
	.w7(32'h3abd2dae),
	.w8(32'h3aadeab0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39054f55),
	.w1(32'h3a113799),
	.w2(32'h3b3ecec8),
	.w3(32'hbb9de666),
	.w4(32'hbb407937),
	.w5(32'hb907f297),
	.w6(32'h3ac86c77),
	.w7(32'h3b708495),
	.w8(32'hb9fabf78),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a680da4),
	.w1(32'h3caf65fe),
	.w2(32'h3d060fb0),
	.w3(32'hbb49fbee),
	.w4(32'hb9ca240c),
	.w5(32'h3bd6c935),
	.w6(32'h3b85d5ba),
	.w7(32'h3c995a1f),
	.w8(32'h3aa4c903),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58a687),
	.w1(32'h3b8ab857),
	.w2(32'h3bf6e420),
	.w3(32'hbbc864e8),
	.w4(32'h3b3ccb5c),
	.w5(32'h3b780e7d),
	.w6(32'h3c2cf270),
	.w7(32'h3b5cfbd5),
	.w8(32'h3bf43f5b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda6618),
	.w1(32'hb9f1fce0),
	.w2(32'hbb6e1202),
	.w3(32'h3b1a2720),
	.w4(32'hbb1fc54a),
	.w5(32'hbb4e9a87),
	.w6(32'hbb0930c3),
	.w7(32'h37c87074),
	.w8(32'hbb38eee8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae41d84),
	.w1(32'h3a9a5ce4),
	.w2(32'h3a13aa35),
	.w3(32'hbbf741da),
	.w4(32'h3b050ff2),
	.w5(32'h3a2147f4),
	.w6(32'hbabfd7be),
	.w7(32'hbacd5ae5),
	.w8(32'hbb600159),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30aea3),
	.w1(32'h3b45c869),
	.w2(32'hba3cb59e),
	.w3(32'hbbbf20e9),
	.w4(32'h3b04fa59),
	.w5(32'h3b7e7f7a),
	.w6(32'h3b951032),
	.w7(32'h3b9a2aa8),
	.w8(32'hb9bbf2b3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebf4f),
	.w1(32'h3b7ea481),
	.w2(32'h3b493d36),
	.w3(32'h3babb20d),
	.w4(32'h3bad973c),
	.w5(32'h3ae33430),
	.w6(32'h3b073ff1),
	.w7(32'h3aee2037),
	.w8(32'hbb1462cb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9484b7),
	.w1(32'hbc2ae8b5),
	.w2(32'hbcad8700),
	.w3(32'hba6d907c),
	.w4(32'hbbe75e93),
	.w5(32'hbc9b2dcf),
	.w6(32'hbb0515a9),
	.w7(32'hbc214652),
	.w8(32'hbbc22988),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8129ef),
	.w1(32'h3a8da6a8),
	.w2(32'h39f8b226),
	.w3(32'hbc4afd39),
	.w4(32'hbb36b9e7),
	.w5(32'h3b88aaf4),
	.w6(32'hbb944465),
	.w7(32'h3b075cef),
	.w8(32'hbb971bdf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1489e),
	.w1(32'hba3c1a3a),
	.w2(32'h3a0f002a),
	.w3(32'hbba7b8ab),
	.w4(32'h3b00b1b4),
	.w5(32'h3c2980ea),
	.w6(32'hbbc3095b),
	.w7(32'hb897ce5f),
	.w8(32'hbacc3ba4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aeaaf),
	.w1(32'hbb5f1361),
	.w2(32'h3be4c371),
	.w3(32'h3c1af03d),
	.w4(32'hbc433bce),
	.w5(32'hbbee921f),
	.w6(32'hbc7e5905),
	.w7(32'hbbb60e35),
	.w8(32'hbc33f4bc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394569b7),
	.w1(32'hbc61bb7f),
	.w2(32'h3a66c160),
	.w3(32'hbc334dc5),
	.w4(32'hbc9d0c32),
	.w5(32'hbba3ef52),
	.w6(32'hbce865cd),
	.w7(32'hbca4d46b),
	.w8(32'hbc95659c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f038),
	.w1(32'hb877d01b),
	.w2(32'hbbab3a17),
	.w3(32'hbc0ae448),
	.w4(32'hbabe3b49),
	.w5(32'hbbe564b2),
	.w6(32'hbb00b6c7),
	.w7(32'hbbcbc60a),
	.w8(32'hbaac5327),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4c3d),
	.w1(32'hbc8bf4c9),
	.w2(32'hbd250556),
	.w3(32'hbb608c76),
	.w4(32'hbc0211c9),
	.w5(32'hbcdf8122),
	.w6(32'hbbfc6c04),
	.w7(32'hbc9769a6),
	.w8(32'hbc1b4bf4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd15a37),
	.w1(32'h3aae561c),
	.w2(32'h3aa1139d),
	.w3(32'hbc6e561c),
	.w4(32'hba84a609),
	.w5(32'h3aaf3747),
	.w6(32'h392e2872),
	.w7(32'h3b0687b4),
	.w8(32'h3aa780f0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb859cfc),
	.w1(32'h3b3c284a),
	.w2(32'h3b4dd828),
	.w3(32'hbb71a4fa),
	.w4(32'h3ba55fa4),
	.w5(32'h3b4f125e),
	.w6(32'h3bea1bbf),
	.w7(32'h3b035b45),
	.w8(32'h3b0fbb65),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e69c7b),
	.w1(32'hbbd23fc8),
	.w2(32'hbb8f6e95),
	.w3(32'h3ab48cc6),
	.w4(32'hbab02887),
	.w5(32'hbb072f75),
	.w6(32'h3aafdba3),
	.w7(32'h3b24463d),
	.w8(32'hbb006e36),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10664e),
	.w1(32'h3a92f2b4),
	.w2(32'h3ae4fb72),
	.w3(32'hbbb7b60a),
	.w4(32'hbb8aeaf8),
	.w5(32'hbb7a3831),
	.w6(32'hbbaddc2e),
	.w7(32'hbbb73f21),
	.w8(32'hbb7a4aea),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8506f9),
	.w1(32'hbbcf83e9),
	.w2(32'h3b0858fd),
	.w3(32'h3ab6b3ae),
	.w4(32'hbb861beb),
	.w5(32'hbb1b6b51),
	.w6(32'hbbb30cc8),
	.w7(32'hbac2a331),
	.w8(32'hbbc889bd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ca47),
	.w1(32'hbc0d2983),
	.w2(32'h3b952254),
	.w3(32'hbae1134e),
	.w4(32'hbc1ae6cf),
	.w5(32'h3bd3f613),
	.w6(32'hbc9674b6),
	.w7(32'hbbb2f918),
	.w8(32'hbc587676),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b41f3),
	.w1(32'hbb0b5079),
	.w2(32'h3a8db12e),
	.w3(32'hbb9dc256),
	.w4(32'hba8615a6),
	.w5(32'h3ba0a8be),
	.w6(32'h3a24ecda),
	.w7(32'hba36a721),
	.w8(32'h3b87350e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151686),
	.w1(32'hbaba5f51),
	.w2(32'hb998a2f8),
	.w3(32'h3ae66cdc),
	.w4(32'h3afddf8b),
	.w5(32'hba6cddb8),
	.w6(32'hbb87944d),
	.w7(32'hbb0741cf),
	.w8(32'hbae0a44f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b9c0),
	.w1(32'h3abfba5c),
	.w2(32'hbadf8171),
	.w3(32'h3af7396c),
	.w4(32'h3b2900a7),
	.w5(32'h3a8ad188),
	.w6(32'h3b17f08d),
	.w7(32'h3aac3b0a),
	.w8(32'h38fc814b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4abd83),
	.w1(32'h3b199c16),
	.w2(32'h3bbaa082),
	.w3(32'hbb2be26e),
	.w4(32'hb9f95c25),
	.w5(32'h3a57cd62),
	.w6(32'h3bc5f869),
	.w7(32'h3c028e7a),
	.w8(32'h3b6db05b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cf941),
	.w1(32'h3bdc5e9d),
	.w2(32'h3c2f8e95),
	.w3(32'hbb1e0198),
	.w4(32'h38a862c3),
	.w5(32'h3ba9d98b),
	.w6(32'h3b995cee),
	.w7(32'h3c25a69f),
	.w8(32'h3ab6610f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbca0c),
	.w1(32'h3ba68a63),
	.w2(32'h3b1ce867),
	.w3(32'hbb1d9970),
	.w4(32'h3b6a2908),
	.w5(32'h3b84f1eb),
	.w6(32'h3ba2fdfa),
	.w7(32'h3b81ac2f),
	.w8(32'h3b34251c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a04d),
	.w1(32'h3a09ace4),
	.w2(32'hbb42ad13),
	.w3(32'h3a5d14bf),
	.w4(32'h3abbf9f4),
	.w5(32'hbb5e1df5),
	.w6(32'h3ab04966),
	.w7(32'h3991e2b7),
	.w8(32'hbaca67bf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1a1d),
	.w1(32'hba445f24),
	.w2(32'h3af595f4),
	.w3(32'hba308dd2),
	.w4(32'h3bad2824),
	.w5(32'h3c2d8926),
	.w6(32'hb8137196),
	.w7(32'h3a97c825),
	.w8(32'hb97b60d9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629ea9),
	.w1(32'hbb1d2917),
	.w2(32'h39709601),
	.w3(32'h3bd59cd6),
	.w4(32'h3b652ffd),
	.w5(32'h3b36a939),
	.w6(32'hbae44123),
	.w7(32'hbb149c3f),
	.w8(32'h3ab5f6a8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72fb25),
	.w1(32'hb9a251eb),
	.w2(32'h3a4ab4a3),
	.w3(32'hbaafc6c6),
	.w4(32'hbbc85899),
	.w5(32'h3b375ae6),
	.w6(32'hbb9e59cb),
	.w7(32'hbbf360c7),
	.w8(32'hbbaa1c6d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a860ebb),
	.w1(32'hbb583487),
	.w2(32'h3b2d04fb),
	.w3(32'h3b1a712b),
	.w4(32'hbbb7880f),
	.w5(32'h3b11c762),
	.w6(32'hbaed283a),
	.w7(32'hba634379),
	.w8(32'hbb7c0c28),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e7da3),
	.w1(32'hbb2a7f66),
	.w2(32'h3b0e3b59),
	.w3(32'hbb4f37d1),
	.w4(32'hbb7434e8),
	.w5(32'h3b6828b9),
	.w6(32'hbba9ff0c),
	.w7(32'hb8264f0d),
	.w8(32'hbb053d06),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0a492),
	.w1(32'hba4c82a5),
	.w2(32'hbc0b4337),
	.w3(32'hbbb4b82a),
	.w4(32'hbbaf8006),
	.w5(32'hbbd7d6d4),
	.w6(32'hbbf076e4),
	.w7(32'hbc0a62b5),
	.w8(32'hbb8220c3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89d27d),
	.w1(32'hbaa6c0f3),
	.w2(32'hba78afe5),
	.w3(32'h3a908265),
	.w4(32'hbb27fa80),
	.w5(32'h3b3d52ed),
	.w6(32'hbc43c8ca),
	.w7(32'hbb8490e6),
	.w8(32'hbbcf5c84),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c8cc6),
	.w1(32'hbbc30805),
	.w2(32'h3b127b2d),
	.w3(32'hb899e80a),
	.w4(32'hbbd7ef63),
	.w5(32'h3af63d59),
	.w6(32'hbc2822c3),
	.w7(32'hbb2f4672),
	.w8(32'hbb6a1260),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92688b),
	.w1(32'hbb000932),
	.w2(32'hba92515b),
	.w3(32'h3b5c0f7a),
	.w4(32'hbb22a2bf),
	.w5(32'hb7ed2eca),
	.w6(32'hbbc83ad6),
	.w7(32'hbbc1a0f5),
	.w8(32'hbbc59042),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398553ca),
	.w1(32'hbbe4343e),
	.w2(32'h3ad00c5d),
	.w3(32'h3a017c06),
	.w4(32'hbb5a3c9f),
	.w5(32'h3b1547e8),
	.w6(32'hbc9a22c4),
	.w7(32'hbc2fc58f),
	.w8(32'hbc2df702),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa66a0d),
	.w1(32'hb7c8d0ec),
	.w2(32'hba3d265f),
	.w3(32'hbb27219c),
	.w4(32'hbaf8a739),
	.w5(32'hba9c0b5a),
	.w6(32'h3a137a79),
	.w7(32'h3a85529a),
	.w8(32'h3a5395ee),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985ac98),
	.w1(32'h3b802f29),
	.w2(32'h3b9af2a8),
	.w3(32'hbaa16e09),
	.w4(32'hbb1139b9),
	.w5(32'h3a807d46),
	.w6(32'hbb6be671),
	.w7(32'hbaa3d134),
	.w8(32'hbbb835bf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9a514),
	.w1(32'hbb1e667f),
	.w2(32'hba9b06fe),
	.w3(32'h399c9041),
	.w4(32'hbac958e2),
	.w5(32'hbb2ebd81),
	.w6(32'h37c46b70),
	.w7(32'h3a911f3d),
	.w8(32'h3968c43d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2aeed),
	.w1(32'hbb5ab852),
	.w2(32'h3ba11f98),
	.w3(32'h389e078a),
	.w4(32'h3b9496cf),
	.w5(32'h3b73415a),
	.w6(32'hba255baa),
	.w7(32'h3abceb7d),
	.w8(32'hbb23d2c9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39880332),
	.w1(32'h3bff6bc6),
	.w2(32'h3cbbf8ee),
	.w3(32'h3b1dcd04),
	.w4(32'h3c14ce05),
	.w5(32'h3cbfa260),
	.w6(32'h3af048e7),
	.w7(32'h3c244eee),
	.w8(32'h3c2f1283),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb98821),
	.w1(32'h3c67e37e),
	.w2(32'h3d0f8abd),
	.w3(32'h3cadbe41),
	.w4(32'h3b376e88),
	.w5(32'h3ca63eb4),
	.w6(32'hba77f407),
	.w7(32'h3c7c9d6e),
	.w8(32'h3bf3039c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf621f),
	.w1(32'hbb8e35e4),
	.w2(32'hbba9f2dc),
	.w3(32'h3c0d20c7),
	.w4(32'hbb5226e4),
	.w5(32'hbb7ea3bf),
	.w6(32'hbc41b817),
	.w7(32'hbc094b46),
	.w8(32'hbbf1c293),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188d26),
	.w1(32'hb891deda),
	.w2(32'h3b211b93),
	.w3(32'hbc0184d4),
	.w4(32'h3b449564),
	.w5(32'h3b41ad4d),
	.w6(32'hbb2e7f67),
	.w7(32'hbab4848c),
	.w8(32'hbb0d1aba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05fa92),
	.w1(32'hbc22d06d),
	.w2(32'hbc35b040),
	.w3(32'h3a971633),
	.w4(32'hbbe6db14),
	.w5(32'hbb21c8f0),
	.w6(32'hbb0513f7),
	.w7(32'hbb9bb740),
	.w8(32'hbc370d78),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4ad62),
	.w1(32'hba952949),
	.w2(32'h3aa623f2),
	.w3(32'hb9b15e73),
	.w4(32'h3a5d5e7e),
	.w5(32'hbb1fa4e2),
	.w6(32'hbb2f7798),
	.w7(32'hba26bf21),
	.w8(32'hbb75854e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39e94),
	.w1(32'h39f937d9),
	.w2(32'h3b24f15a),
	.w3(32'h38fbf31c),
	.w4(32'h3b8dba0e),
	.w5(32'h3a81c3f5),
	.w6(32'h3ac8aaf7),
	.w7(32'h3afd2560),
	.w8(32'h3be393c2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b736e27),
	.w1(32'h3c14c513),
	.w2(32'h3c6ceca6),
	.w3(32'h3aa87075),
	.w4(32'h3bcef0ca),
	.w5(32'h3bcd83c9),
	.w6(32'hbb798c5e),
	.w7(32'h38452468),
	.w8(32'hbb52fc6a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e524b),
	.w1(32'h3b0bbc67),
	.w2(32'h3a651649),
	.w3(32'h3b5b5075),
	.w4(32'h3a69b32e),
	.w5(32'hb9586abb),
	.w6(32'hbb853a09),
	.w7(32'hbb09b662),
	.w8(32'hbc527878),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29fe8),
	.w1(32'hba4557c8),
	.w2(32'h3a47d625),
	.w3(32'hbabef3b9),
	.w4(32'hbb9a8faa),
	.w5(32'hba95eb0b),
	.w6(32'hbafe4eff),
	.w7(32'hbb7a4424),
	.w8(32'hbb83634c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9dfdf),
	.w1(32'hb9a79fb0),
	.w2(32'h3bf7fab8),
	.w3(32'h3baa537a),
	.w4(32'h3848fd4e),
	.w5(32'h397f67f5),
	.w6(32'hbc27b7d9),
	.w7(32'hbaa57c83),
	.w8(32'hbb7c4a72),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4edf7),
	.w1(32'hbb68ca1a),
	.w2(32'hbb8d40b7),
	.w3(32'h3b095a30),
	.w4(32'hbb74345a),
	.w5(32'h3a460d30),
	.w6(32'h38f11ff0),
	.w7(32'hbb2969d3),
	.w8(32'hbb90e513),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb669843),
	.w1(32'h3a9b1617),
	.w2(32'h3ba64e69),
	.w3(32'hb63870c3),
	.w4(32'h3aa2bd5f),
	.w5(32'h3b9cf0e0),
	.w6(32'h3bcd782f),
	.w7(32'h3b8069f3),
	.w8(32'h3b94ca7a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c591),
	.w1(32'hbcdf7081),
	.w2(32'hbd2059c4),
	.w3(32'h3b8a6138),
	.w4(32'hbcbb6ff9),
	.w5(32'hbcf87f9f),
	.w6(32'hbc959596),
	.w7(32'hbc5fc64e),
	.w8(32'hbcc5be30),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e6bca),
	.w1(32'h3a67e30d),
	.w2(32'hbb812ba1),
	.w3(32'hbcfb0fd4),
	.w4(32'h3af3bd08),
	.w5(32'h39b733f1),
	.w6(32'h3b07131a),
	.w7(32'hbb522c63),
	.w8(32'h38458eba),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7e183),
	.w1(32'h3bb91755),
	.w2(32'hba43f149),
	.w3(32'hb92462b1),
	.w4(32'h3ba0ee64),
	.w5(32'hbab20d9e),
	.w6(32'h3b486ab9),
	.w7(32'hbaf804b4),
	.w8(32'hbb0e95d9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069e12),
	.w1(32'h3c1bfab5),
	.w2(32'h3c9cdaec),
	.w3(32'hbabcbc25),
	.w4(32'h3b6b253c),
	.w5(32'h3c5443f4),
	.w6(32'h3924b2b6),
	.w7(32'h3bf73b21),
	.w8(32'h3c044bb7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7558a5),
	.w1(32'h3c260101),
	.w2(32'h3ce129fc),
	.w3(32'h3c3bf9de),
	.w4(32'hbbbe7315),
	.w5(32'h3c023e3d),
	.w6(32'hbbdebeeb),
	.w7(32'h3c0171b0),
	.w8(32'hbb4751a3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d49b2),
	.w1(32'hb9fd6c00),
	.w2(32'hbb43ce55),
	.w3(32'hbb5ee0ae),
	.w4(32'hbb0239cf),
	.w5(32'h3ba151c8),
	.w6(32'h3a178795),
	.w7(32'hbb7e076a),
	.w8(32'h3a752ac2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc6a93),
	.w1(32'h3aecd855),
	.w2(32'h3a733f92),
	.w3(32'h3a9d4bc9),
	.w4(32'h3b3468b5),
	.w5(32'h3b348d06),
	.w6(32'hba87d181),
	.w7(32'hba8faa4e),
	.w8(32'h39e92179),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b05a6),
	.w1(32'h3c8586c0),
	.w2(32'h3cf1f86b),
	.w3(32'h3b7dded6),
	.w4(32'h3c283659),
	.w5(32'h3cc612af),
	.w6(32'h3bdab9c9),
	.w7(32'h3c6d8f0c),
	.w8(32'h3c386434),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b3b16),
	.w1(32'hba98a84a),
	.w2(32'hba6c3280),
	.w3(32'h3c38041e),
	.w4(32'h3a9d86dd),
	.w5(32'hbb9ce939),
	.w6(32'hba9c6021),
	.w7(32'h3a18cf1f),
	.w8(32'hba5cf334),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3784e6),
	.w1(32'hbb8810b9),
	.w2(32'hbb94fa9a),
	.w3(32'hba9b991e),
	.w4(32'hbb883156),
	.w5(32'hbb6e3d25),
	.w6(32'hbb07529e),
	.w7(32'hbb603a92),
	.w8(32'h3a9a2509),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09b4de),
	.w1(32'h3bbc688c),
	.w2(32'h3c107521),
	.w3(32'hba82aad9),
	.w4(32'hbae1495a),
	.w5(32'hb9671478),
	.w6(32'h3921b5f6),
	.w7(32'h3b94b2bf),
	.w8(32'h39f76569),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9add47),
	.w1(32'h3b3353b1),
	.w2(32'h3c2c8900),
	.w3(32'hbb221acd),
	.w4(32'h3afa5832),
	.w5(32'h3c08b9b0),
	.w6(32'h39a0d824),
	.w7(32'h3c2b3c09),
	.w8(32'h3b99fd69),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19ab45),
	.w1(32'h3c2339df),
	.w2(32'h3c00a0c3),
	.w3(32'h3bc6ab72),
	.w4(32'h3c36f0fb),
	.w5(32'h3c2c8be8),
	.w6(32'h3be8f0fa),
	.w7(32'h3bc61647),
	.w8(32'h3af9efa0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c60d),
	.w1(32'hb8945b57),
	.w2(32'h3b58d685),
	.w3(32'h3c073888),
	.w4(32'h3b751ec2),
	.w5(32'h3ab9edcd),
	.w6(32'hbae0e70d),
	.w7(32'h38e5ba0a),
	.w8(32'hb92c4eca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39919016),
	.w1(32'h395119dc),
	.w2(32'h3baf9ce9),
	.w3(32'h3afd32be),
	.w4(32'hbaab0fe1),
	.w5(32'h3b958e86),
	.w6(32'h3b3f322b),
	.w7(32'h3b9442e4),
	.w8(32'h3aa4dab9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93e817),
	.w1(32'hbaf6e78b),
	.w2(32'h3bc415c6),
	.w3(32'hb9902f99),
	.w4(32'hbb559dcc),
	.w5(32'hbb107f73),
	.w6(32'hbac17fa6),
	.w7(32'hbb254d3a),
	.w8(32'hbb987dbf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f3b5f),
	.w1(32'hb9e1f1b4),
	.w2(32'hbb16a944),
	.w3(32'h3b266602),
	.w4(32'h3a258251),
	.w5(32'h3ab81c20),
	.w6(32'hbc10a10a),
	.w7(32'hbb3f7ab0),
	.w8(32'hbaf00427),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54ecc9),
	.w1(32'h3cc7383f),
	.w2(32'h3d7ae670),
	.w3(32'hbb01a755),
	.w4(32'h3b597768),
	.w5(32'h3d091dff),
	.w6(32'hbbbbe8d6),
	.w7(32'h3c97a84f),
	.w8(32'h3bd38e8b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d227c17),
	.w1(32'h3c434724),
	.w2(32'h3c8c50a1),
	.w3(32'h3c77b501),
	.w4(32'h3bc89faf),
	.w5(32'h3c03a809),
	.w6(32'h3b8efa12),
	.w7(32'h3c122517),
	.w8(32'h3ae016d2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e36cc),
	.w1(32'hbba20d18),
	.w2(32'hba00628c),
	.w3(32'h3be62a1f),
	.w4(32'hbb67bc53),
	.w5(32'hbae0fca3),
	.w6(32'hbb1fb127),
	.w7(32'h3b5cd170),
	.w8(32'h3af11fbd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ae81),
	.w1(32'hbb8ee7df),
	.w2(32'h3b73a476),
	.w3(32'hbb90db4e),
	.w4(32'h3b4f0c17),
	.w5(32'h3b9f01cf),
	.w6(32'h39b55103),
	.w7(32'hba187aff),
	.w8(32'h3a618c3f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a5ae7),
	.w1(32'hba96e26d),
	.w2(32'hbaa9057e),
	.w3(32'hb911117d),
	.w4(32'hbaa0b396),
	.w5(32'h3a4c0a7a),
	.w6(32'hba562bfe),
	.w7(32'hb93c010b),
	.w8(32'hbb0a37ce),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0b97),
	.w1(32'h3d169729),
	.w2(32'h3d14117a),
	.w3(32'hba8e4a50),
	.w4(32'h3d1afe35),
	.w5(32'h3cdd8ae7),
	.w6(32'h3cbe0559),
	.w7(32'h3cb498a4),
	.w8(32'h3c185080),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule