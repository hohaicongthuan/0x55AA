module layer_8_featuremap_200(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57084a),
	.w1(32'hbc093af2),
	.w2(32'hbbe9db99),
	.w3(32'h3bacb3fd),
	.w4(32'hbc144c59),
	.w5(32'hbbc168c2),
	.w6(32'h3a6ad7ce),
	.w7(32'hbc0ac889),
	.w8(32'hba18790e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beae79a),
	.w1(32'h3b06cda9),
	.w2(32'hba0bbb48),
	.w3(32'h3c6781ea),
	.w4(32'h3ba279f2),
	.w5(32'h3b494cd2),
	.w6(32'h3b8311fc),
	.w7(32'hb96f86b9),
	.w8(32'h3b4f7a9e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913e9c),
	.w1(32'hbb7506da),
	.w2(32'hbb910707),
	.w3(32'h3b84c39b),
	.w4(32'hbc445ee0),
	.w5(32'hbac4e73d),
	.w6(32'hbc2a4e91),
	.w7(32'hbbd242d6),
	.w8(32'h3a61b3b1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6b07b),
	.w1(32'h39cc8763),
	.w2(32'h3c9ad69a),
	.w3(32'h3c5d2512),
	.w4(32'hbb82aec6),
	.w5(32'h3b697eff),
	.w6(32'h3bd5147e),
	.w7(32'h3c827124),
	.w8(32'h3c523e53),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c84b1),
	.w1(32'h3a8c3cbe),
	.w2(32'h3a142b7d),
	.w3(32'h3b359cb5),
	.w4(32'h3abd28b8),
	.w5(32'hba1969fd),
	.w6(32'h3b883c0e),
	.w7(32'h3b4d0791),
	.w8(32'hb9b92d2d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6737),
	.w1(32'hbc0651a6),
	.w2(32'h3ca3fa16),
	.w3(32'hbb87584f),
	.w4(32'hbbacc251),
	.w5(32'h3c69467e),
	.w6(32'hb9df244d),
	.w7(32'hb9d9cb7f),
	.w8(32'h3af25e97),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac57526),
	.w1(32'hbb32604c),
	.w2(32'h3aba60ec),
	.w3(32'h3a19b320),
	.w4(32'hbb349de2),
	.w5(32'hbb63de11),
	.w6(32'hbb3f77de),
	.w7(32'hba4b9877),
	.w8(32'hbb9db99e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5cfe2),
	.w1(32'hbb691d9c),
	.w2(32'h3c410582),
	.w3(32'hbc0935fe),
	.w4(32'hbc55a070),
	.w5(32'h3c10547e),
	.w6(32'hbbf325a2),
	.w7(32'h3acde248),
	.w8(32'hbc2d9c6f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f0a3),
	.w1(32'hbb6d7341),
	.w2(32'h3bb35e7e),
	.w3(32'hbc1b795e),
	.w4(32'hbac5190a),
	.w5(32'h3b7db7b6),
	.w6(32'hb8ae7bda),
	.w7(32'h3baf3a31),
	.w8(32'hbae17801),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4f2d7),
	.w1(32'hbc94e7ce),
	.w2(32'hbc865c3d),
	.w3(32'hbc2f63a2),
	.w4(32'hbc6cb7ef),
	.w5(32'hba20a4fb),
	.w6(32'hbc2bbae1),
	.w7(32'hbc62e146),
	.w8(32'h3c15ad6e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77ad00),
	.w1(32'h3b21b214),
	.w2(32'hbc43f16f),
	.w3(32'h3bc1f75f),
	.w4(32'h3a75c8e4),
	.w5(32'hbcbcb6e5),
	.w6(32'h3b11a244),
	.w7(32'hbc340c46),
	.w8(32'h3cba43bd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf6eaab),
	.w1(32'hbba0d77f),
	.w2(32'hbad0a14f),
	.w3(32'h3ca41e57),
	.w4(32'hbb94b245),
	.w5(32'hbbc73a9d),
	.w6(32'hbb18cfef),
	.w7(32'hbb5aceed),
	.w8(32'h3a88477b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886675),
	.w1(32'h3b7b549a),
	.w2(32'hbbed06f1),
	.w3(32'hbaa259a7),
	.w4(32'hbabc6a00),
	.w5(32'hbc0dfa3b),
	.w6(32'h3bb96d8b),
	.w7(32'hbbd98a05),
	.w8(32'hbaaec23a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b79d2),
	.w1(32'h3a969e4f),
	.w2(32'hbbad23f5),
	.w3(32'hbb9d1bb4),
	.w4(32'hbb987283),
	.w5(32'hbbc47f4b),
	.w6(32'hbb9febaa),
	.w7(32'hbc030515),
	.w8(32'hbbfc8426),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefc2b9),
	.w1(32'h3ac09a05),
	.w2(32'h3be048bb),
	.w3(32'hba20cbe4),
	.w4(32'h39cb43f4),
	.w5(32'h3b45b5a0),
	.w6(32'h3a180f41),
	.w7(32'h3ba9cf2b),
	.w8(32'hbb935fcd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0575d8),
	.w1(32'h39397596),
	.w2(32'hbbce0959),
	.w3(32'hbb9d1368),
	.w4(32'hbb1a285a),
	.w5(32'hbbfd8b3d),
	.w6(32'h3b95d158),
	.w7(32'hbba27e02),
	.w8(32'h3ba55dbc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2df1ff),
	.w1(32'hbb88170b),
	.w2(32'hbca6aea6),
	.w3(32'hbb85a071),
	.w4(32'hbac78d15),
	.w5(32'hbba76dc4),
	.w6(32'h3b88d705),
	.w7(32'hbbea9ba0),
	.w8(32'h3b0231c4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc4f01),
	.w1(32'h3c523825),
	.w2(32'h3c867cc1),
	.w3(32'h3c326620),
	.w4(32'h3bb238ae),
	.w5(32'h3c0c558b),
	.w6(32'h3c3740d4),
	.w7(32'h3bd80c7c),
	.w8(32'hbca77013),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd038d7a),
	.w1(32'h3b845060),
	.w2(32'h3ce77054),
	.w3(32'hbc9a9031),
	.w4(32'hbc28bf93),
	.w5(32'hbb857546),
	.w6(32'hbce30c90),
	.w7(32'h3bfcf722),
	.w8(32'h39252e06),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91ea2d),
	.w1(32'h3a4d0daa),
	.w2(32'h3ba18f42),
	.w3(32'hbcef32e5),
	.w4(32'hb9e070c6),
	.w5(32'h3c368845),
	.w6(32'h3be1d597),
	.w7(32'h3b602611),
	.w8(32'hbaa45b2b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18041b),
	.w1(32'hba9ef770),
	.w2(32'hbb9bdd47),
	.w3(32'h3b86cbe5),
	.w4(32'h3b54c239),
	.w5(32'hbc0a5fb2),
	.w6(32'hbc299d2c),
	.w7(32'hbc9da1bc),
	.w8(32'hbc14692c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e72ea),
	.w1(32'hbba4df3a),
	.w2(32'hbbb9c1bb),
	.w3(32'hbc0dc0b5),
	.w4(32'h3ab74508),
	.w5(32'hbc6c192c),
	.w6(32'hbc5446eb),
	.w7(32'hb7eec2b7),
	.w8(32'hbc6e161a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8ad9d),
	.w1(32'h3c64b119),
	.w2(32'hbceecb55),
	.w3(32'hbc0fb3bb),
	.w4(32'hbc762bfd),
	.w5(32'hbd0c4b70),
	.w6(32'h3baae9f8),
	.w7(32'hbcd5a863),
	.w8(32'h3bae935a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25812e),
	.w1(32'h3b901f4c),
	.w2(32'h3b827813),
	.w3(32'h3c2a1d5f),
	.w4(32'hba6bb087),
	.w5(32'hbc1380b7),
	.w6(32'hba9b141f),
	.w7(32'h3b9d6cdb),
	.w8(32'hbc6f849a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a90c6),
	.w1(32'h39fa8a71),
	.w2(32'h3a7969c7),
	.w3(32'hba1485e5),
	.w4(32'h3b57470f),
	.w5(32'h3b670434),
	.w6(32'h3ab74c10),
	.w7(32'h39bb79c7),
	.w8(32'hbbd49428),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5a2d8),
	.w1(32'h3afd2da2),
	.w2(32'h3afb139b),
	.w3(32'h3b9003b4),
	.w4(32'hbaa75c5c),
	.w5(32'hbc198253),
	.w6(32'h3b1ba928),
	.w7(32'hbc28eb7e),
	.w8(32'hbc6e539d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079b85),
	.w1(32'hbc224ab5),
	.w2(32'hbc2117a9),
	.w3(32'hbaeb7cc7),
	.w4(32'hbc3df9ca),
	.w5(32'hbc20048b),
	.w6(32'h3bf8cbb0),
	.w7(32'h3b4bf040),
	.w8(32'h3b2653da),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36a820),
	.w1(32'hbc5ba8de),
	.w2(32'hbb26a33a),
	.w3(32'h3d387645),
	.w4(32'h3d10da6d),
	.w5(32'hbd48bd80),
	.w6(32'h3b939025),
	.w7(32'hbd3c9084),
	.w8(32'h3c0d80da),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac40c45),
	.w1(32'hbb6769e7),
	.w2(32'h3ad5582b),
	.w3(32'hba596529),
	.w4(32'h3ab47671),
	.w5(32'h3b865692),
	.w6(32'hba16b127),
	.w7(32'hbbcc25b5),
	.w8(32'h3bd7f829),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c131b),
	.w1(32'hbbcaf541),
	.w2(32'h3a17608e),
	.w3(32'h3b32d221),
	.w4(32'hbc92f642),
	.w5(32'hbc116974),
	.w6(32'hbbb2f8c6),
	.w7(32'hbb819186),
	.w8(32'h3cbb8798),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc2cb1),
	.w1(32'h3abba72b),
	.w2(32'h3be3f97c),
	.w3(32'h3c8e4c21),
	.w4(32'hb858a9c9),
	.w5(32'h3bcbbbff),
	.w6(32'h3c56040e),
	.w7(32'h3bac87b0),
	.w8(32'h3c0774ea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8f744),
	.w1(32'hbc8d6f36),
	.w2(32'hbc10d0a4),
	.w3(32'hba9bafc9),
	.w4(32'hbc455437),
	.w5(32'hbb68b861),
	.w6(32'hbb9b54af),
	.w7(32'hb9dbf83e),
	.w8(32'h3b316f19),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c387128),
	.w1(32'hbb858419),
	.w2(32'hbc0e92e8),
	.w3(32'h3c11b896),
	.w4(32'hba800130),
	.w5(32'hbbc4be22),
	.w6(32'hbbb6cd4e),
	.w7(32'hbbc0c3f9),
	.w8(32'hbc5d3681),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61654e),
	.w1(32'h3c57afff),
	.w2(32'h3b7c0349),
	.w3(32'hbc81a22e),
	.w4(32'h3a8de275),
	.w5(32'h3c5089b4),
	.w6(32'h3c118f4c),
	.w7(32'h3b94ce9d),
	.w8(32'h3c23ef05),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17e9bb),
	.w1(32'h385975a4),
	.w2(32'h3c623cae),
	.w3(32'h3c3d0ddd),
	.w4(32'h3ae94c91),
	.w5(32'h3c1f600d),
	.w6(32'hbb59df87),
	.w7(32'h3a9908eb),
	.w8(32'h3c09399f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d989c),
	.w1(32'h3b7a96b2),
	.w2(32'h3c99ed05),
	.w3(32'h3a9c956e),
	.w4(32'h3c0b55de),
	.w5(32'h3c5dc352),
	.w6(32'hbb9817d6),
	.w7(32'h3b2e71c3),
	.w8(32'h3c5b1801),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91758b),
	.w1(32'hbbde49f0),
	.w2(32'h3b2d01d9),
	.w3(32'h3bbe0564),
	.w4(32'hbbd16051),
	.w5(32'h3a4e0cb4),
	.w6(32'hbb98507e),
	.w7(32'h3ae76213),
	.w8(32'h3bd6f732),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d4810),
	.w1(32'h3ba92b01),
	.w2(32'h3bb3b3f5),
	.w3(32'h3b97407e),
	.w4(32'h3bf1d2f0),
	.w5(32'h3b8f36ac),
	.w6(32'h3c0317a8),
	.w7(32'h3c2512f2),
	.w8(32'h3b0a9674),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73d944),
	.w1(32'h3c88beb4),
	.w2(32'h3c958ba3),
	.w3(32'h37afb9a8),
	.w4(32'h3c64ed50),
	.w5(32'h3b9b85de),
	.w6(32'h3b8df5ca),
	.w7(32'h3c898e29),
	.w8(32'hbc24d69f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f40d),
	.w1(32'h3b4e784c),
	.w2(32'hbb00b593),
	.w3(32'hbbd78058),
	.w4(32'hbbac6d4f),
	.w5(32'h3a195ef4),
	.w6(32'h3bc5f5b1),
	.w7(32'hbafe0bf9),
	.w8(32'h3acb5ce9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5cd46),
	.w1(32'hbb8c8c48),
	.w2(32'h3bfc6a42),
	.w3(32'h3c25193c),
	.w4(32'h3a1fae7c),
	.w5(32'h3c231903),
	.w6(32'h3b4e030d),
	.w7(32'h3b2a4a84),
	.w8(32'h3c7357a9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f96c6),
	.w1(32'h3c5d8c05),
	.w2(32'hbcc71b60),
	.w3(32'h39cfa373),
	.w4(32'h3c16caa3),
	.w5(32'hbc99b8d7),
	.w6(32'h3c56df30),
	.w7(32'hbc776fd4),
	.w8(32'hb8287cda),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc063),
	.w1(32'hbbeaa5b6),
	.w2(32'h3bdc065a),
	.w3(32'h3b2ead6f),
	.w4(32'hbac2f355),
	.w5(32'h3abb596e),
	.w6(32'hbb9e646e),
	.w7(32'h3bd3de36),
	.w8(32'h3c0e615a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951077),
	.w1(32'h3bd88f42),
	.w2(32'h3c2e1875),
	.w3(32'h3be35639),
	.w4(32'hbc2116a1),
	.w5(32'hbbdfc3f7),
	.w6(32'h3b02a58c),
	.w7(32'h3b4db53a),
	.w8(32'hbcb8b3cb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c6e31),
	.w1(32'hbc0c6715),
	.w2(32'h3c2e421a),
	.w3(32'hbcdcc763),
	.w4(32'hbc7f1381),
	.w5(32'hbb9661a7),
	.w6(32'hbc5d3ef0),
	.w7(32'hbb01bc27),
	.w8(32'h3ccca173),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced3181),
	.w1(32'hbc1eda41),
	.w2(32'hbabeaaae),
	.w3(32'h3c8470e5),
	.w4(32'hbbd9efe4),
	.w5(32'h39c49fd2),
	.w6(32'hbc38763e),
	.w7(32'hbb447fd1),
	.w8(32'hbad01c8b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06df9),
	.w1(32'h3c1c3ee6),
	.w2(32'hbb45db3f),
	.w3(32'hba71e15f),
	.w4(32'h3c3b3893),
	.w5(32'h38987e97),
	.w6(32'h3c0a7a32),
	.w7(32'hba0d0237),
	.w8(32'hbbae4536),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc869244),
	.w1(32'h378d5c72),
	.w2(32'h3ca4df84),
	.w3(32'hbbacf392),
	.w4(32'hbb44aa4e),
	.w5(32'h3a28d8a1),
	.w6(32'hbc3ec0a2),
	.w7(32'h3bf17ced),
	.w8(32'h3cbd0dbf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fd865),
	.w1(32'hbb8f538e),
	.w2(32'hbb025239),
	.w3(32'h3b01be5d),
	.w4(32'hbbd6d982),
	.w5(32'hbc4f75f5),
	.w6(32'h3b65ab0c),
	.w7(32'hbb7ddbb7),
	.w8(32'h3a91286b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3bd7f),
	.w1(32'h3c6111bb),
	.w2(32'h3cbaa51e),
	.w3(32'h3ab180b0),
	.w4(32'h3c62bada),
	.w5(32'h3c57dd7c),
	.w6(32'h3c4a9591),
	.w7(32'h3cbc6ebc),
	.w8(32'h3a945e2a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4893d),
	.w1(32'h3ac70d78),
	.w2(32'h3ab96d32),
	.w3(32'hbc1a9147),
	.w4(32'h3bb425bc),
	.w5(32'h3b8c1f78),
	.w6(32'hbb54aaaa),
	.w7(32'hbbba4349),
	.w8(32'h3b3b0839),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cfc9c),
	.w1(32'h3c5f86dc),
	.w2(32'h3c1f0036),
	.w3(32'hb98ebb35),
	.w4(32'hbc05b811),
	.w5(32'hbc10ce46),
	.w6(32'h3bb8f0db),
	.w7(32'hbb45dec6),
	.w8(32'h3bead1be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f7ab),
	.w1(32'hbb89e5a1),
	.w2(32'hbbcedae1),
	.w3(32'hba213fa0),
	.w4(32'hbb5a0fe4),
	.w5(32'hbbbc08a1),
	.w6(32'hbad363bb),
	.w7(32'hbbb1cfca),
	.w8(32'h3ab15a8d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0430),
	.w1(32'hbbd30fdd),
	.w2(32'h3b89623b),
	.w3(32'h394a5701),
	.w4(32'hbc27bca1),
	.w5(32'h3c689908),
	.w6(32'hbc46dd9d),
	.w7(32'hbc274204),
	.w8(32'hbcb5d578),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d82ee),
	.w1(32'h3c71e57d),
	.w2(32'h3cc6e915),
	.w3(32'hbcb2d4df),
	.w4(32'h3c0c2aba),
	.w5(32'h3c8f7746),
	.w6(32'h3b992ceb),
	.w7(32'h3c72660d),
	.w8(32'hbc7d9d6d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39f333),
	.w1(32'hbb31fa53),
	.w2(32'hbc089b63),
	.w3(32'hbbdce901),
	.w4(32'hbba5c2a9),
	.w5(32'h3aae9d2d),
	.w6(32'hbc315870),
	.w7(32'hbcaf5e9b),
	.w8(32'hbb92f03f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca016fb),
	.w1(32'h3ce447f9),
	.w2(32'h3c083ccb),
	.w3(32'hbcaccfb3),
	.w4(32'h3c91218a),
	.w5(32'h3acd3041),
	.w6(32'h3c9e2ee0),
	.w7(32'hbb48e97a),
	.w8(32'hbb97eab3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fc0e),
	.w1(32'hbc7738e3),
	.w2(32'h3c8b5a01),
	.w3(32'h3a864e0b),
	.w4(32'hbcbf4479),
	.w5(32'h3bc9c076),
	.w6(32'hbc53aca5),
	.w7(32'h3b790288),
	.w8(32'h3bad76d9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48ad9),
	.w1(32'hbb02865c),
	.w2(32'hbb8f6130),
	.w3(32'h3b46b13d),
	.w4(32'hbb7df2d0),
	.w5(32'hbc2d4668),
	.w6(32'hbb12a072),
	.w7(32'hbc1b2521),
	.w8(32'hbbfaa993),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598433),
	.w1(32'h3c873773),
	.w2(32'h3be8f9da),
	.w3(32'h3a6c4a46),
	.w4(32'h3c888459),
	.w5(32'h3badd536),
	.w6(32'h3c2bbc04),
	.w7(32'h3cb4ba32),
	.w8(32'hbb95b648),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273129),
	.w1(32'h3beb912d),
	.w2(32'hbc2a910e),
	.w3(32'hbbf4ebfa),
	.w4(32'h3b0c50f0),
	.w5(32'hbb40e94c),
	.w6(32'h3b273c61),
	.w7(32'hbc5ca2e4),
	.w8(32'hbc7c6458),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cf787),
	.w1(32'h3b152389),
	.w2(32'hbb8b43b6),
	.w3(32'hbb56b978),
	.w4(32'h3b12436b),
	.w5(32'hbc13f108),
	.w6(32'h3b9e127e),
	.w7(32'h3bda497c),
	.w8(32'h3c083a9b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf6ed),
	.w1(32'hbbd783d5),
	.w2(32'h3942ce71),
	.w3(32'h3a52904b),
	.w4(32'hbb06874d),
	.w5(32'h3c34b784),
	.w6(32'hbab0eb1b),
	.w7(32'hbb8c99b8),
	.w8(32'h3cedfaa2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc89fd),
	.w1(32'h3a74a08f),
	.w2(32'hbaef8e31),
	.w3(32'h3c6d525f),
	.w4(32'h39e999b2),
	.w5(32'hbb0d4a24),
	.w6(32'h3a859dc7),
	.w7(32'hbb40d00b),
	.w8(32'hbaf0343f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c23c6),
	.w1(32'hb9b69de8),
	.w2(32'hbbba0d5b),
	.w3(32'hbb1ec1ab),
	.w4(32'hbadfabcb),
	.w5(32'hbb2dfee8),
	.w6(32'h3a521130),
	.w7(32'hbb8a59bd),
	.w8(32'h3b1365c0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f63db),
	.w1(32'hbb1b66cf),
	.w2(32'h3af027a9),
	.w3(32'h3b92c25c),
	.w4(32'h3ad04df9),
	.w5(32'hbbd0b68d),
	.w6(32'hbaa20446),
	.w7(32'h3a6e26c5),
	.w8(32'h3b402df3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af72f),
	.w1(32'hbc06c8e3),
	.w2(32'hbbbc8aaf),
	.w3(32'h3c14e265),
	.w4(32'hbba8d4fc),
	.w5(32'h3b5781a0),
	.w6(32'hbc1d6487),
	.w7(32'hbb992020),
	.w8(32'h368ab7f5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9167a7),
	.w1(32'h3b0d0c21),
	.w2(32'hbbbfc3c0),
	.w3(32'hbb24089e),
	.w4(32'h3bb71ffb),
	.w5(32'hbb0a5423),
	.w6(32'hbc038e4e),
	.w7(32'hbc85844f),
	.w8(32'hbc3ff6aa),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96181a),
	.w1(32'hb70f2b29),
	.w2(32'h3be73804),
	.w3(32'hbadc58b2),
	.w4(32'hbbc42442),
	.w5(32'h3c479d8a),
	.w6(32'h3b568007),
	.w7(32'h3b2f3069),
	.w8(32'h3bc15d4d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb509e),
	.w1(32'h3bea731b),
	.w2(32'h3ca41156),
	.w3(32'h3cd7db37),
	.w4(32'h3b3bf047),
	.w5(32'hbc91b8c6),
	.w6(32'h3a9121b1),
	.w7(32'hbbc47da2),
	.w8(32'hbc0daaa1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61bdb6),
	.w1(32'h3b57a546),
	.w2(32'hbbcfb64e),
	.w3(32'hbc01745d),
	.w4(32'h3b5dfb01),
	.w5(32'hbb25c644),
	.w6(32'h3b87b27a),
	.w7(32'h3be0d0f1),
	.w8(32'hbb05a8cc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56bf96),
	.w1(32'h3b81a19a),
	.w2(32'h38d26cc7),
	.w3(32'h374191ac),
	.w4(32'hbb301083),
	.w5(32'h3a9f6942),
	.w6(32'h3b7c67e8),
	.w7(32'hbb0d9a82),
	.w8(32'hbbb07753),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd52a15),
	.w1(32'h3b527b9b),
	.w2(32'h3bb1149b),
	.w3(32'h3b30689f),
	.w4(32'h3ba219c1),
	.w5(32'hba91966e),
	.w6(32'hbb603720),
	.w7(32'hbad5a271),
	.w8(32'h3bb5b9a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4ecf),
	.w1(32'hbbd4540b),
	.w2(32'h3c8bc68b),
	.w3(32'h3bd5dff7),
	.w4(32'h3b17c480),
	.w5(32'h3cb4b15e),
	.w6(32'hbc3db65a),
	.w7(32'hbacd9140),
	.w8(32'h3af4b728),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b639ee7),
	.w1(32'h3c24623f),
	.w2(32'h3b3ef02c),
	.w3(32'hba948e30),
	.w4(32'h3c1cb3f2),
	.w5(32'h3b89346a),
	.w6(32'h3bb25ed5),
	.w7(32'hba0544ad),
	.w8(32'hbbcc3e66),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad60681),
	.w1(32'h3ce52dd8),
	.w2(32'h3a60287d),
	.w3(32'hb85436ad),
	.w4(32'h3c720446),
	.w5(32'hbb073348),
	.w6(32'h3c8163f2),
	.w7(32'hbba35e81),
	.w8(32'hbc5ddb02),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34c19),
	.w1(32'hbb14c47f),
	.w2(32'h3b848301),
	.w3(32'hb9ed83a7),
	.w4(32'h3b91eb42),
	.w5(32'h398e35a8),
	.w6(32'hbb7caeaf),
	.w7(32'hbafccf68),
	.w8(32'hbbc67ec7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d4e2),
	.w1(32'hbb0b2d2f),
	.w2(32'h3c0512d6),
	.w3(32'h3b949766),
	.w4(32'h3a3f462e),
	.w5(32'hbbd56366),
	.w6(32'hbc45cff4),
	.w7(32'hbbb69b3d),
	.w8(32'hb9cccf1a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1967),
	.w1(32'h3bd04c9d),
	.w2(32'hbb5d0275),
	.w3(32'hbb699265),
	.w4(32'h3c2865d1),
	.w5(32'h3aeab362),
	.w6(32'h3c138138),
	.w7(32'hba63b631),
	.w8(32'hbb66880d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24278b),
	.w1(32'h3c221c74),
	.w2(32'hbcd28a7e),
	.w3(32'hbaf891af),
	.w4(32'h3bffc431),
	.w5(32'hbcc25d9e),
	.w6(32'h3bbdee91),
	.w7(32'hbcd72d6e),
	.w8(32'hbbe8ab3b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c3c7),
	.w1(32'hbc2fdadc),
	.w2(32'hbc404347),
	.w3(32'hbc6f3f64),
	.w4(32'hbb97e764),
	.w5(32'hbc4695b1),
	.w6(32'hbab85b31),
	.w7(32'hbc1e2801),
	.w8(32'hbb420080),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01942),
	.w1(32'h3b0fa3da),
	.w2(32'h3bd6b2b1),
	.w3(32'hbbcda8ca),
	.w4(32'hbc05d44e),
	.w5(32'hba29aa4d),
	.w6(32'h3c199d5d),
	.w7(32'h3b19418c),
	.w8(32'hba6c0ef1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af58c2e),
	.w1(32'h3cb4a532),
	.w2(32'h3c7823bb),
	.w3(32'h3c18f8e7),
	.w4(32'h3c3f0906),
	.w5(32'h3b326385),
	.w6(32'h3bd119d9),
	.w7(32'h3b508f92),
	.w8(32'hbbe59531),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ea03c),
	.w1(32'h3ce945c7),
	.w2(32'h3d6fb2ba),
	.w3(32'h3c36b230),
	.w4(32'h3c869d78),
	.w5(32'h3d815167),
	.w6(32'h3cce43e5),
	.w7(32'h3d10974c),
	.w8(32'h3c3de883),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaba7ea),
	.w1(32'hbc19effc),
	.w2(32'hbb3da266),
	.w3(32'hbbe476d9),
	.w4(32'hbc91df62),
	.w5(32'hbc5a482c),
	.w6(32'hbc51247a),
	.w7(32'hbc129c4a),
	.w8(32'h3baed254),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad08a92),
	.w1(32'h3bd03926),
	.w2(32'h3c5e0391),
	.w3(32'h3c1030fd),
	.w4(32'hbbba7a51),
	.w5(32'h3be64e5d),
	.w6(32'h3c7a868b),
	.w7(32'h3b3af446),
	.w8(32'h3c528693),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beaa49b),
	.w1(32'h3b4dbfd3),
	.w2(32'h3b06147d),
	.w3(32'h3bd545a6),
	.w4(32'h3af479d0),
	.w5(32'h3b66c79f),
	.w6(32'h3c00b746),
	.w7(32'h3a955b67),
	.w8(32'h3b93c3c8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae4350),
	.w1(32'hb77398bd),
	.w2(32'hbc15271a),
	.w3(32'h3be96e76),
	.w4(32'h3a6a9114),
	.w5(32'hbb94ebce),
	.w6(32'h3b7ebded),
	.w7(32'hbb7bb52e),
	.w8(32'hbba6513e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08094e),
	.w1(32'hb8c8b68e),
	.w2(32'h3bfb13f5),
	.w3(32'h3abf2618),
	.w4(32'hbc0a5081),
	.w5(32'h3b6bd553),
	.w6(32'h3bdd04e2),
	.w7(32'h3b995c5f),
	.w8(32'hba8ea18f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73e2f),
	.w1(32'hbba1b27d),
	.w2(32'hbaae4e81),
	.w3(32'h3b0185a3),
	.w4(32'hbc2319bb),
	.w5(32'h3b804f5e),
	.w6(32'h3b1aebd8),
	.w7(32'hbb3eac88),
	.w8(32'h3bb9af21),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0007a8),
	.w1(32'h3b00fd03),
	.w2(32'h3c9397d2),
	.w3(32'h3b96fe9e),
	.w4(32'h3b8bd7aa),
	.w5(32'h3ae00829),
	.w6(32'h3c26deaf),
	.w7(32'h3bb22f22),
	.w8(32'h3b818ea7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40b71f),
	.w1(32'hba137562),
	.w2(32'h3b813606),
	.w3(32'h3bbc767f),
	.w4(32'h3ba7c3d2),
	.w5(32'h3b76232f),
	.w6(32'h3c129dbf),
	.w7(32'h3b4d0afc),
	.w8(32'h3c2ce8b5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77dfa1),
	.w1(32'h3b626aa6),
	.w2(32'hbaba5e40),
	.w3(32'h3c010373),
	.w4(32'hb8dd7f48),
	.w5(32'hba2cdf34),
	.w6(32'h3b907614),
	.w7(32'hba395dd3),
	.w8(32'hba06696e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04999a),
	.w1(32'h3b64577c),
	.w2(32'hb8813501),
	.w3(32'h3ae8bd61),
	.w4(32'h3b991adc),
	.w5(32'h3a411d38),
	.w6(32'h3b7e1d22),
	.w7(32'hba4036e3),
	.w8(32'hbb45549a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d02c),
	.w1(32'hbd53a7a3),
	.w2(32'h3d71187d),
	.w3(32'hbb12d972),
	.w4(32'hbce596c4),
	.w5(32'h3d2fd799),
	.w6(32'hbd1ec35e),
	.w7(32'h3c961609),
	.w8(32'h3c20bbab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc00ad),
	.w1(32'hbbdd66ef),
	.w2(32'h3b5884c4),
	.w3(32'h3b8601df),
	.w4(32'hbbbf0ed8),
	.w5(32'h3b8e098c),
	.w6(32'hbbf7828e),
	.w7(32'hbbc7bc64),
	.w8(32'h39b2a6e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed1c2b),
	.w1(32'h3c8b75b0),
	.w2(32'h3bb7390a),
	.w3(32'h3b99d78c),
	.w4(32'hbbee7480),
	.w5(32'h3b220347),
	.w6(32'h3bbc9bd0),
	.w7(32'h3ba20fe8),
	.w8(32'hbc489594),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe91703),
	.w1(32'h3cded7cd),
	.w2(32'h3ca8d856),
	.w3(32'hbc80d282),
	.w4(32'h3cb0e08c),
	.w5(32'h3bc5f142),
	.w6(32'h3c26f01a),
	.w7(32'h3c6882f0),
	.w8(32'hbcbd90f7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde2069),
	.w1(32'h3cf2251c),
	.w2(32'h3be9b645),
	.w3(32'hbcadb87a),
	.w4(32'h3ccca11f),
	.w5(32'h3aac2185),
	.w6(32'h3c86a661),
	.w7(32'h3bc1e0d9),
	.w8(32'hbc8bc4f1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93310d),
	.w1(32'hbb788b3e),
	.w2(32'hbc005c20),
	.w3(32'hbca3035f),
	.w4(32'h3b9e5c90),
	.w5(32'hbc077ce9),
	.w6(32'hbb8cad85),
	.w7(32'hbc3db4ad),
	.w8(32'h3b619597),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c2c6b),
	.w1(32'h3ba0d5d6),
	.w2(32'hbc650d51),
	.w3(32'h3b8bdf6e),
	.w4(32'hbbaf4346),
	.w5(32'hbc49b236),
	.w6(32'h3b953757),
	.w7(32'hbbb8ffcb),
	.w8(32'hbbd8005a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb464fcf),
	.w1(32'hbba15c35),
	.w2(32'h3c556ff0),
	.w3(32'h3b462bb4),
	.w4(32'hbb8c1384),
	.w5(32'h3c7091f6),
	.w6(32'hbba81f92),
	.w7(32'h3b82de2b),
	.w8(32'h3c6195ed),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c1941),
	.w1(32'h3aebc2fb),
	.w2(32'h3bf8ada8),
	.w3(32'h3c9875f9),
	.w4(32'hbc7e4033),
	.w5(32'h3b911b09),
	.w6(32'h3b2b6f6e),
	.w7(32'h3bd04f1c),
	.w8(32'hba25dcc4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa32a8),
	.w1(32'h3b589867),
	.w2(32'h3b909c81),
	.w3(32'h3b9c2d77),
	.w4(32'h3b91e945),
	.w5(32'h3c29a0e5),
	.w6(32'hbb2007e1),
	.w7(32'h3b252486),
	.w8(32'hbc021eff),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b5e4),
	.w1(32'h3d58faf9),
	.w2(32'hbbac2225),
	.w3(32'h3b5ac0c5),
	.w4(32'h3d01935d),
	.w5(32'hb9aaa66f),
	.w6(32'h3d011e41),
	.w7(32'hbb263d5a),
	.w8(32'h3cc3f50b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d099b40),
	.w1(32'hba74719d),
	.w2(32'h3b95e811),
	.w3(32'h3d24480b),
	.w4(32'hbab7c760),
	.w5(32'hbbe90085),
	.w6(32'h396a7aaf),
	.w7(32'hbb853908),
	.w8(32'hbabeac78),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c4a6a),
	.w1(32'h3b90504d),
	.w2(32'h3c5eee8f),
	.w3(32'hbae49744),
	.w4(32'h3a43df12),
	.w5(32'h3c31c75a),
	.w6(32'h3b160f4f),
	.w7(32'h3b818404),
	.w8(32'h3b367856),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c66a),
	.w1(32'hbacac8ac),
	.w2(32'h3c149f1a),
	.w3(32'hba1556f8),
	.w4(32'h3b35cc9b),
	.w5(32'h3c3b6300),
	.w6(32'hbabd0f73),
	.w7(32'h3bc4dd0b),
	.w8(32'h3b58a5c7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1666bc),
	.w1(32'hbc0af7dc),
	.w2(32'hbc6e728e),
	.w3(32'h3c1beab2),
	.w4(32'hbc3a3e84),
	.w5(32'hbc4ae8ad),
	.w6(32'h3aaba1c9),
	.w7(32'hbc3bf14d),
	.w8(32'hb9ebecd2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060b45),
	.w1(32'h3b5db383),
	.w2(32'hbb978766),
	.w3(32'hbbd427fe),
	.w4(32'h3b75f546),
	.w5(32'hbb797ca3),
	.w6(32'h3ba0daec),
	.w7(32'hbb06fea2),
	.w8(32'h3b3788c7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b8e98),
	.w1(32'hbb71c52a),
	.w2(32'hb7371c69),
	.w3(32'h3ac69685),
	.w4(32'h3b271d73),
	.w5(32'h3b971525),
	.w6(32'hba11553e),
	.w7(32'h3b086496),
	.w8(32'h3b30b3b3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6430dd),
	.w1(32'hbb4b7753),
	.w2(32'hbaa18a5b),
	.w3(32'h3bea1281),
	.w4(32'hbb1bdd15),
	.w5(32'hba8a0b22),
	.w6(32'hbae31fa0),
	.w7(32'hb9754799),
	.w8(32'h3b99b659),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dcdfe),
	.w1(32'h3adefa6c),
	.w2(32'h3c3e3ead),
	.w3(32'h3bb227f2),
	.w4(32'h3b8d3e6d),
	.w5(32'h3b93fe7c),
	.w6(32'h3c0631d4),
	.w7(32'h3b1855c9),
	.w8(32'h3a442ceb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b8e0),
	.w1(32'h3814bc34),
	.w2(32'h3b900c63),
	.w3(32'hb92e5c50),
	.w4(32'h3bbac26a),
	.w5(32'hba63a603),
	.w6(32'hbad6bc51),
	.w7(32'h3bfcfacd),
	.w8(32'h3b9c4f69),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9842e),
	.w1(32'h3b0ec2be),
	.w2(32'hbbfa8a24),
	.w3(32'hbb17c52d),
	.w4(32'hbb9dbb1b),
	.w5(32'hbbe4430f),
	.w6(32'h3c2cb10e),
	.w7(32'hba33ee4d),
	.w8(32'h3b6be703),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba672ece),
	.w1(32'h39f505b4),
	.w2(32'hbbb0140b),
	.w3(32'h3b741575),
	.w4(32'h3a1522a7),
	.w5(32'hbb581bea),
	.w6(32'h3a7b4ab1),
	.w7(32'hbba402bb),
	.w8(32'h3b869881),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc877a4),
	.w1(32'h3bbe2001),
	.w2(32'hbbf42397),
	.w3(32'h3baeaeb3),
	.w4(32'h3c352737),
	.w5(32'hbc2b98bd),
	.w6(32'h3be8e149),
	.w7(32'hbb7e00bc),
	.w8(32'h3b85eac7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8b5b),
	.w1(32'hba9d19a6),
	.w2(32'h3c402a3a),
	.w3(32'h3b3114b6),
	.w4(32'hba8eb9e5),
	.w5(32'h3bbd3fc3),
	.w6(32'h3baecd4c),
	.w7(32'h388ada22),
	.w8(32'h3c252eb2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5071a0),
	.w1(32'hbc34ddca),
	.w2(32'hbc06b0bf),
	.w3(32'h3b3cd0f9),
	.w4(32'hbbc8596e),
	.w5(32'hbc10f1e6),
	.w6(32'hbb6b1607),
	.w7(32'hbb865541),
	.w8(32'hbbaaa351),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc259bfb),
	.w1(32'h3c3fcc7b),
	.w2(32'hbb5ee652),
	.w3(32'hbc192e84),
	.w4(32'h3bd28b9d),
	.w5(32'hbbc21841),
	.w6(32'h3c130585),
	.w7(32'hb9405363),
	.w8(32'hbb468ebc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31c061),
	.w1(32'hbc28d8b4),
	.w2(32'h3b3aa57d),
	.w3(32'hbaa27874),
	.w4(32'hbba97d68),
	.w5(32'h3a1efb5c),
	.w6(32'h3c254c0c),
	.w7(32'h3ae97108),
	.w8(32'hbaa5d148),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc9c92),
	.w1(32'h3b4b8d60),
	.w2(32'hbbe4faad),
	.w3(32'h3bd50960),
	.w4(32'h3af200f9),
	.w5(32'hbb8d1610),
	.w6(32'h3bb3cbbf),
	.w7(32'h3ad69236),
	.w8(32'hbba9e70e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd459cb),
	.w1(32'h3b3198e8),
	.w2(32'hba841461),
	.w3(32'hbb9413bf),
	.w4(32'h3ab77bd9),
	.w5(32'hba8edf2a),
	.w6(32'h3ba36da3),
	.w7(32'h3a693440),
	.w8(32'h3bb13acf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21f913),
	.w1(32'h3b85c108),
	.w2(32'h3c090909),
	.w3(32'h3b57ab87),
	.w4(32'h3afc532c),
	.w5(32'h3c00e57c),
	.w6(32'h3b07a531),
	.w7(32'h3be33a63),
	.w8(32'h3b766160),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87bc2),
	.w1(32'h3b600c34),
	.w2(32'h3c83cd31),
	.w3(32'hbb406507),
	.w4(32'hbc0066dc),
	.w5(32'h3bee71da),
	.w6(32'hbb51b522),
	.w7(32'h3b225579),
	.w8(32'hba8a105c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b775ed0),
	.w1(32'hbaa59fb0),
	.w2(32'hbb22980e),
	.w3(32'h3a5a7baf),
	.w4(32'hbbc37f62),
	.w5(32'hba6427fc),
	.w6(32'hbb51bc50),
	.w7(32'hba04cb9d),
	.w8(32'h3bc875ec),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08278d),
	.w1(32'hbaf66258),
	.w2(32'h3aacc2f0),
	.w3(32'h39c04619),
	.w4(32'h3a38ca50),
	.w5(32'h3ad41937),
	.w6(32'hbad17a56),
	.w7(32'hbb0607be),
	.w8(32'h3a2be7e0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0007e8),
	.w1(32'h39e3f334),
	.w2(32'h3b43820d),
	.w3(32'hbaa66db8),
	.w4(32'hbbf53c73),
	.w5(32'hbb2e9bc4),
	.w6(32'hbb05a1c6),
	.w7(32'h3b4e6abb),
	.w8(32'h3b7793bf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule