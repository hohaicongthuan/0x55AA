module layer_8_featuremap_14(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14f0e8),
	.w1(32'hbac3f14f),
	.w2(32'hbbe79551),
	.w3(32'hba2a554e),
	.w4(32'h3b08f9fe),
	.w5(32'hbbad3041),
	.w6(32'hbb4c3bd8),
	.w7(32'hba588bea),
	.w8(32'hbb5a1ad5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02f5a8),
	.w1(32'hbb40f950),
	.w2(32'h3bb5478a),
	.w3(32'hbb514161),
	.w4(32'hbad804db),
	.w5(32'hbbabe2b1),
	.w6(32'hbb1b2da7),
	.w7(32'hbc40998d),
	.w8(32'hbc541d63),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71496),
	.w1(32'hbb7dff6f),
	.w2(32'h3b6b6e95),
	.w3(32'hbbf6b0af),
	.w4(32'hba882c80),
	.w5(32'hba052a06),
	.w6(32'h3c2ed3cc),
	.w7(32'h3b87c5cc),
	.w8(32'hbbae44a2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8be96),
	.w1(32'h3bb45649),
	.w2(32'hba5de500),
	.w3(32'hbb1280a5),
	.w4(32'hbacd71c9),
	.w5(32'hbab95bb5),
	.w6(32'h3a3215a6),
	.w7(32'h3b2dfd6f),
	.w8(32'hbbaed64b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f351b),
	.w1(32'h3a0bcccc),
	.w2(32'h3aac04c2),
	.w3(32'h36d0887e),
	.w4(32'h3aa13f2a),
	.w5(32'h3a15d594),
	.w6(32'h3bdfeff3),
	.w7(32'hbb49d002),
	.w8(32'hb949db3a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6112fb),
	.w1(32'hbc1093c9),
	.w2(32'h3b30dc3f),
	.w3(32'h3c2d952e),
	.w4(32'h3b7112a7),
	.w5(32'h3c45dcdf),
	.w6(32'h3c445a41),
	.w7(32'h376229d0),
	.w8(32'h3bc4dc41),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0f13),
	.w1(32'h3a7b23fa),
	.w2(32'h3b83d8dc),
	.w3(32'hba45f025),
	.w4(32'hbba11615),
	.w5(32'hbb66d55a),
	.w6(32'h3c6f1960),
	.w7(32'h3c7d3201),
	.w8(32'h39716c41),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47132d),
	.w1(32'hbb8884d2),
	.w2(32'h3bcb3513),
	.w3(32'h3c349844),
	.w4(32'hbb83801e),
	.w5(32'h3a424b16),
	.w6(32'hbb08c599),
	.w7(32'h3b555b2f),
	.w8(32'hbab5f5db),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7076),
	.w1(32'hbb99ebb2),
	.w2(32'hbb5cd972),
	.w3(32'hbc620429),
	.w4(32'hbc1209a7),
	.w5(32'hbb8fbb38),
	.w6(32'hbbbb9652),
	.w7(32'hbc203500),
	.w8(32'hba5048d6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398db77c),
	.w1(32'hbb7c15f6),
	.w2(32'h3b33cf32),
	.w3(32'h3abda73e),
	.w4(32'hbb8447d3),
	.w5(32'hbb0de82c),
	.w6(32'hbb3e6068),
	.w7(32'h3a865107),
	.w8(32'h3b3f264d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b51d1),
	.w1(32'h3bafe5c7),
	.w2(32'hbc253ba1),
	.w3(32'hba025d34),
	.w4(32'hbbf10af0),
	.w5(32'hbbdc77c8),
	.w6(32'h3be72feb),
	.w7(32'hbc044000),
	.w8(32'hb9b87f77),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28587b),
	.w1(32'h3c57e58d),
	.w2(32'h3a25bff8),
	.w3(32'hbb35743c),
	.w4(32'h3b80ea26),
	.w5(32'hbae1bba6),
	.w6(32'hbace1a18),
	.w7(32'h3971c78f),
	.w8(32'hbb02ede0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98d05),
	.w1(32'hbb41d976),
	.w2(32'h3a50521a),
	.w3(32'h3be689bd),
	.w4(32'h3afcd1d2),
	.w5(32'hbb0da8f6),
	.w6(32'hbb456b89),
	.w7(32'h3b63b486),
	.w8(32'h3a0e7923),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03033b),
	.w1(32'h3b0487a5),
	.w2(32'hbc3304d3),
	.w3(32'h3ab9c4e4),
	.w4(32'h3ac02e2b),
	.w5(32'hbb36205c),
	.w6(32'hbbfe86ee),
	.w7(32'h3c9a19f4),
	.w8(32'h3b1e4b40),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1386d),
	.w1(32'h3ada2a60),
	.w2(32'hbb96514f),
	.w3(32'h3b44d6de),
	.w4(32'hbad2ca83),
	.w5(32'h3b9b5d3e),
	.w6(32'h3cc4caf6),
	.w7(32'h3ae006e9),
	.w8(32'hba2a4553),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb330d8),
	.w1(32'h3b458fd8),
	.w2(32'hbb358c5c),
	.w3(32'hbaf248c5),
	.w4(32'hbb03318f),
	.w5(32'hbc53d0bf),
	.w6(32'hba6ff53b),
	.w7(32'h3a73a098),
	.w8(32'hba5260ce),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3143ab),
	.w1(32'hba7bfb2c),
	.w2(32'hba10d56b),
	.w3(32'h3b83681f),
	.w4(32'hbb04c229),
	.w5(32'h3c95c0dc),
	.w6(32'hbba86d57),
	.w7(32'hbb6102e1),
	.w8(32'hbbda4d6b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97f1c3),
	.w1(32'h3aa937b1),
	.w2(32'hbc744f3e),
	.w3(32'hba8e1b6e),
	.w4(32'hbbf15e28),
	.w5(32'h3c36c322),
	.w6(32'hbc5dc2b1),
	.w7(32'hbc840cdd),
	.w8(32'hba827935),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095b91),
	.w1(32'hbc4c9774),
	.w2(32'hbc64ccb3),
	.w3(32'hbc6f1cf6),
	.w4(32'hbc6490ed),
	.w5(32'h3a9c5372),
	.w6(32'hbbff4979),
	.w7(32'hbb22d9ae),
	.w8(32'hbafaf334),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae617a4),
	.w1(32'h3c1f958c),
	.w2(32'h3bcaa087),
	.w3(32'hbb27a677),
	.w4(32'h3c0eef95),
	.w5(32'hbc0f36a3),
	.w6(32'hbbbf0231),
	.w7(32'hbc7a57fa),
	.w8(32'hba5fcb05),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c099),
	.w1(32'hbbc6eb57),
	.w2(32'hbb838618),
	.w3(32'h3b7ed2a5),
	.w4(32'h3c9daa77),
	.w5(32'h3c0e55da),
	.w6(32'h3b02c682),
	.w7(32'h3ba82cb8),
	.w8(32'h3bd0af50),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221d07),
	.w1(32'h3c8d26d9),
	.w2(32'h3b1656d7),
	.w3(32'hba23231c),
	.w4(32'hbb6f72f2),
	.w5(32'h3b8f71e1),
	.w6(32'h3b9d2d1b),
	.w7(32'hbc029828),
	.w8(32'h3a4c4f85),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee530),
	.w1(32'hbbfca546),
	.w2(32'hbc687498),
	.w3(32'hbbdca2a6),
	.w4(32'hbb584a84),
	.w5(32'hbc14c01f),
	.w6(32'hbb8fb1dc),
	.w7(32'hbc22486f),
	.w8(32'hbb162b3b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0f805),
	.w1(32'h3b73bcb1),
	.w2(32'h3b138d0d),
	.w3(32'hbbdaaa3f),
	.w4(32'hbb303b72),
	.w5(32'hbb846de4),
	.w6(32'hb9bc9381),
	.w7(32'h3b6edf0a),
	.w8(32'hbaee251f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a156024),
	.w1(32'hbadab513),
	.w2(32'hbb3bd3bb),
	.w3(32'h3aad2a7d),
	.w4(32'h3c52c738),
	.w5(32'hbca684f0),
	.w6(32'hbaba9cff),
	.w7(32'h3c5bb91e),
	.w8(32'hbb26e736),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24b20),
	.w1(32'h3bd53151),
	.w2(32'h3abff053),
	.w3(32'h3bc37841),
	.w4(32'hbc6fd748),
	.w5(32'h38c17988),
	.w6(32'h3b41fb5f),
	.w7(32'h39b17450),
	.w8(32'h3b0c2c3e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac60a5c),
	.w1(32'h3aa95447),
	.w2(32'h3b9253e5),
	.w3(32'h3bd07219),
	.w4(32'hbb74d0dc),
	.w5(32'h3b9fbe7a),
	.w6(32'hbadea96b),
	.w7(32'hb9a656f5),
	.w8(32'hbb55b6a3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93a813),
	.w1(32'hbc55f0e4),
	.w2(32'hbcc66783),
	.w3(32'hbc9f8d36),
	.w4(32'hbd49e43c),
	.w5(32'hbcbab48d),
	.w6(32'hbcab9881),
	.w7(32'hbd114768),
	.w8(32'h3c797c5c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4130a6),
	.w1(32'hb9ab96e4),
	.w2(32'hbc2f7498),
	.w3(32'hba4f18a5),
	.w4(32'h3c2444cc),
	.w5(32'hbb7b7750),
	.w6(32'h3c141814),
	.w7(32'hbabb9754),
	.w8(32'hbc246718),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85cbf1),
	.w1(32'hba42c0b4),
	.w2(32'hbbfd2c32),
	.w3(32'h3b727f21),
	.w4(32'hbbcd081a),
	.w5(32'hba2da0cc),
	.w6(32'hbb808147),
	.w7(32'h3b174e27),
	.w8(32'h383d3d1e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a70e9),
	.w1(32'h3c6059cb),
	.w2(32'h3bcda3fb),
	.w3(32'h3af5a11f),
	.w4(32'h3c96a847),
	.w5(32'hb9b72212),
	.w6(32'h3ca47cce),
	.w7(32'hbc31de97),
	.w8(32'h3ab37f10),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9080b),
	.w1(32'h3b966965),
	.w2(32'hbc0117bf),
	.w3(32'hbb89a46f),
	.w4(32'hbba7ea12),
	.w5(32'h3c3bdf28),
	.w6(32'hbc060804),
	.w7(32'h3b92cc98),
	.w8(32'h3b85ca34),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55cdb1),
	.w1(32'hb99c70c6),
	.w2(32'hbc08586c),
	.w3(32'hbb73d05b),
	.w4(32'h3bef9aae),
	.w5(32'hbbdc11bb),
	.w6(32'h3a910140),
	.w7(32'h3c716dcd),
	.w8(32'h3b6cf0ab),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34ddc8),
	.w1(32'h3c17968f),
	.w2(32'hbc6a6ceb),
	.w3(32'h3c4aa12a),
	.w4(32'hbacb86ac),
	.w5(32'hbca3a988),
	.w6(32'h3acd9c65),
	.w7(32'h3b689b2d),
	.w8(32'h3beda4c1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad70210),
	.w1(32'hb9698094),
	.w2(32'hbb6ca081),
	.w3(32'hbbbab9d9),
	.w4(32'hbb4c64a2),
	.w5(32'hbb654031),
	.w6(32'hbbaf881a),
	.w7(32'h3cfe7dca),
	.w8(32'hbc433a8a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ed98),
	.w1(32'hbafcf458),
	.w2(32'hbbd6ae0c),
	.w3(32'hbb0b2ba5),
	.w4(32'h3be06256),
	.w5(32'hba5beb79),
	.w6(32'hbae8df1b),
	.w7(32'h3c496132),
	.w8(32'hbbe79ae7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cc50),
	.w1(32'h3b4ece1a),
	.w2(32'h399cdac2),
	.w3(32'hba362711),
	.w4(32'h394055b3),
	.w5(32'h3be79a21),
	.w6(32'h3c98e749),
	.w7(32'hbb0cc008),
	.w8(32'hbc0f8d6d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a9f08),
	.w1(32'h3b9739d4),
	.w2(32'hbb9f9a14),
	.w3(32'hbb012299),
	.w4(32'hb939c7ef),
	.w5(32'h3af9df0d),
	.w6(32'h3beafe15),
	.w7(32'hbb08cd4e),
	.w8(32'hbc270c74),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda56a7),
	.w1(32'h3b3f929c),
	.w2(32'h3c55d139),
	.w3(32'hbbc6dea6),
	.w4(32'hbafbde68),
	.w5(32'h3c59efe2),
	.w6(32'hbbd8d228),
	.w7(32'hbc044485),
	.w8(32'hbc8a4148),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a3dcf),
	.w1(32'hbcb6cd9d),
	.w2(32'hbbe9688f),
	.w3(32'hbc152bd8),
	.w4(32'hbc13fe0b),
	.w5(32'h38b2e0c8),
	.w6(32'h3bfbd6c4),
	.w7(32'h3bd7c181),
	.w8(32'hbc84136d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84cdd),
	.w1(32'h3c146052),
	.w2(32'h3a7e97aa),
	.w3(32'hbba41f24),
	.w4(32'hbbeddef9),
	.w5(32'hbc1024ea),
	.w6(32'hbc391724),
	.w7(32'hbcba12ff),
	.w8(32'hbb1e3e19),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c809588),
	.w1(32'hbc380d49),
	.w2(32'h3bb0386f),
	.w3(32'h3d0c92ea),
	.w4(32'hbcb7c1be),
	.w5(32'hbc5f7f2b),
	.w6(32'hbb507f20),
	.w7(32'hbc5fd722),
	.w8(32'h3cbc14fe),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea25b),
	.w1(32'h3c3884d5),
	.w2(32'h3c19ca5d),
	.w3(32'h3d2d5ee3),
	.w4(32'hbc7d54c3),
	.w5(32'hbbb30f94),
	.w6(32'hbc76e868),
	.w7(32'hbc7a1771),
	.w8(32'h3c6939b3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceaa6c3),
	.w1(32'hbcb7d00e),
	.w2(32'h3c30af98),
	.w3(32'hbcde344a),
	.w4(32'h3c45e8b2),
	.w5(32'hbc2437ec),
	.w6(32'hbc2bb980),
	.w7(32'h3af4049d),
	.w8(32'hbb042b30),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41a155),
	.w1(32'hbbdfc022),
	.w2(32'hbc620b0e),
	.w3(32'hbc408d2d),
	.w4(32'h3cf6e403),
	.w5(32'hbbd27818),
	.w6(32'h3c6dcecb),
	.w7(32'hbb26254e),
	.w8(32'hbc7da088),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99979b),
	.w1(32'hbbaff22f),
	.w2(32'hbc4ed6ed),
	.w3(32'hbad2c918),
	.w4(32'h3c4de405),
	.w5(32'hbb7fdde5),
	.w6(32'h3c29c584),
	.w7(32'hbb23eb3e),
	.w8(32'hbc6d3a79),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba822dd),
	.w1(32'h3bc290c7),
	.w2(32'h3c5b45da),
	.w3(32'hbc18eb26),
	.w4(32'h3c03e36c),
	.w5(32'hbc4f9866),
	.w6(32'hbc841f83),
	.w7(32'hbc72972b),
	.w8(32'hbbc8c7c5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb249602),
	.w1(32'h3d80fc3b),
	.w2(32'h3c705a0f),
	.w3(32'hbbd1dfd7),
	.w4(32'hbb47b05e),
	.w5(32'hbd197d1e),
	.w6(32'hbc984e28),
	.w7(32'hba2bd5e3),
	.w8(32'hbccc5090),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba8980),
	.w1(32'h3bf28615),
	.w2(32'hbc83cd48),
	.w3(32'h3b6c1de0),
	.w4(32'hbb0c0837),
	.w5(32'h3c3e681c),
	.w6(32'hb8e69248),
	.w7(32'hbad80c7a),
	.w8(32'hbb69b225),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ec31),
	.w1(32'hbb53a67c),
	.w2(32'h3bb420ee),
	.w3(32'h3c36f847),
	.w4(32'h3ceb06a7),
	.w5(32'h3a574b29),
	.w6(32'h3be462c0),
	.w7(32'h3bc3e8ba),
	.w8(32'hbc772f1a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5598e),
	.w1(32'hbc35f673),
	.w2(32'h3bd9472f),
	.w3(32'hbc8be576),
	.w4(32'hbc512553),
	.w5(32'hbc85a65b),
	.w6(32'h3ac3ee46),
	.w7(32'hbc2a5bbe),
	.w8(32'h3c102295),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ed25d),
	.w1(32'hbbeec1c7),
	.w2(32'hbc90a095),
	.w3(32'hbc4c5964),
	.w4(32'hbc11dc55),
	.w5(32'hbc983ce1),
	.w6(32'hbc7a163a),
	.w7(32'h3becaeae),
	.w8(32'hbcff2c63),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06bd09),
	.w1(32'hbc1fdb00),
	.w2(32'h3c05d86a),
	.w3(32'h3c628c89),
	.w4(32'hbcd8e888),
	.w5(32'hbc3434f8),
	.w6(32'hbcdbb02b),
	.w7(32'h3db0f97e),
	.w8(32'h3c910030),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34673e),
	.w1(32'hbcb76a89),
	.w2(32'h3a53439e),
	.w3(32'h3bb77467),
	.w4(32'hbc0eaf9e),
	.w5(32'hba130c87),
	.w6(32'hbb8fad75),
	.w7(32'h3ca22991),
	.w8(32'hbc3c6a32),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc703b08),
	.w1(32'hba567df2),
	.w2(32'h3bb0b7e1),
	.w3(32'h3c79eeda),
	.w4(32'hbc729e22),
	.w5(32'h3c61c6fc),
	.w6(32'h3c937c38),
	.w7(32'h3c4d77e8),
	.w8(32'h3c1e5d3c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c751f40),
	.w1(32'h3bc1858b),
	.w2(32'h3b698165),
	.w3(32'h3c09e492),
	.w4(32'hbc2dc0af),
	.w5(32'hbb7c3509),
	.w6(32'hbc36f5de),
	.w7(32'h3b7fe46a),
	.w8(32'hb917d1c0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6663e),
	.w1(32'h394bd411),
	.w2(32'hbbffe2fe),
	.w3(32'h3b889d26),
	.w4(32'h3a8fcb37),
	.w5(32'h3c2b22e8),
	.w6(32'h3b0aa647),
	.w7(32'h3b91ec89),
	.w8(32'h3b25a18e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c690ca),
	.w1(32'hbaef30a8),
	.w2(32'hbceef4b4),
	.w3(32'hbb6006fc),
	.w4(32'hbb59c024),
	.w5(32'hba970cc0),
	.w6(32'h3984b03a),
	.w7(32'hbc189e56),
	.w8(32'hbca40095),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d771c),
	.w1(32'h3c2219bb),
	.w2(32'hbb9a162f),
	.w3(32'hbc1bbacc),
	.w4(32'hb9409743),
	.w5(32'hbb350e1c),
	.w6(32'hbbdd3f83),
	.w7(32'h3a8e9c85),
	.w8(32'h3d50227b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe486fc),
	.w1(32'h3a5a9f8f),
	.w2(32'hbbc152a8),
	.w3(32'hbbae43ac),
	.w4(32'h3c78f495),
	.w5(32'hbb141ce4),
	.w6(32'hbc66beb9),
	.w7(32'hbc4f748c),
	.w8(32'h3c21b813),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e6e41),
	.w1(32'hbb9ed3db),
	.w2(32'h3b288f15),
	.w3(32'hbb209175),
	.w4(32'hbb27dfa8),
	.w5(32'h3c79a802),
	.w6(32'h3becdcbd),
	.w7(32'hbb446ee8),
	.w8(32'h3bcf15f6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826726),
	.w1(32'h3cc1129f),
	.w2(32'h39d48c55),
	.w3(32'h3afaec0d),
	.w4(32'h3bd2e599),
	.w5(32'h3b5a57a1),
	.w6(32'hbb941535),
	.w7(32'hbb88f97a),
	.w8(32'hbc976619),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caba148),
	.w1(32'h3b41fd81),
	.w2(32'hbc260baa),
	.w3(32'hba970c4a),
	.w4(32'hbc3d157b),
	.w5(32'hbc83cbed),
	.w6(32'hbc3eaf69),
	.w7(32'hbb3113f7),
	.w8(32'h3b56954d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c712686),
	.w1(32'hbc1fc7eb),
	.w2(32'h3d1003b6),
	.w3(32'h3bdc8840),
	.w4(32'h3c2b6dcd),
	.w5(32'hba92f969),
	.w6(32'hbc1659cb),
	.w7(32'hbafeb67e),
	.w8(32'h3b6306f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78e67a),
	.w1(32'h3935fa47),
	.w2(32'h3cd64431),
	.w3(32'h3ca0ae67),
	.w4(32'h3be05a2e),
	.w5(32'h3a31bc1c),
	.w6(32'h3a48116c),
	.w7(32'h3b1c2521),
	.w8(32'h3aa473c6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c4c80),
	.w1(32'hbc7ef00f),
	.w2(32'h3b1944db),
	.w3(32'hbb375864),
	.w4(32'hbc77dc29),
	.w5(32'hbb8012f3),
	.w6(32'hbb6153fb),
	.w7(32'hbb06132f),
	.w8(32'h39d44548),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2e18),
	.w1(32'hbbcf5fc0),
	.w2(32'hbb9c6e41),
	.w3(32'hbc6fe367),
	.w4(32'h3b3baeb8),
	.w5(32'hbc43e38c),
	.w6(32'hbc1b0326),
	.w7(32'hba0de307),
	.w8(32'hbb9c3bd8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4abcac),
	.w1(32'hbc1eb9b1),
	.w2(32'h39c2e734),
	.w3(32'h394cb932),
	.w4(32'hbb655514),
	.w5(32'hbbd17cf4),
	.w6(32'h3c3ef061),
	.w7(32'hb99288ce),
	.w8(32'h3b9b5771),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af90842),
	.w1(32'hbbc9585d),
	.w2(32'hbc212546),
	.w3(32'hbc040765),
	.w4(32'h3c54716e),
	.w5(32'h3c0fbaad),
	.w6(32'hbb83ecad),
	.w7(32'h3a40cc50),
	.w8(32'h3aa88edd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe901a4),
	.w1(32'h3c156504),
	.w2(32'hbc3a6e3d),
	.w3(32'h3c8cfb17),
	.w4(32'hbd27485e),
	.w5(32'hbc6664a4),
	.w6(32'hbc7a4950),
	.w7(32'h3af5865a),
	.w8(32'h3be733e9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0937a0),
	.w1(32'hbaf39233),
	.w2(32'h3c55fefd),
	.w3(32'hb8721ce1),
	.w4(32'hbd3e537a),
	.w5(32'hba528370),
	.w6(32'hbbd55a7f),
	.w7(32'h3a20c2e1),
	.w8(32'hbb12540e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7481a2),
	.w1(32'h3b3aeb7b),
	.w2(32'hbc86ff4a),
	.w3(32'hbd406187),
	.w4(32'hbc1548da),
	.w5(32'h3b2b41ea),
	.w6(32'h3b839580),
	.w7(32'hbb87b59a),
	.w8(32'hbb796f98),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d5fe),
	.w1(32'hbabbd6f9),
	.w2(32'h3d4c6f03),
	.w3(32'h3b1ba944),
	.w4(32'h3bc051e6),
	.w5(32'hbb797321),
	.w6(32'h3bc93c6d),
	.w7(32'h3ba3ace0),
	.w8(32'h3cb9089f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2cd63),
	.w1(32'hbbfdea9a),
	.w2(32'hbcea992e),
	.w3(32'h3bf25e79),
	.w4(32'hbb9f5ce1),
	.w5(32'hbb6da120),
	.w6(32'h3b9677b1),
	.w7(32'hbb9de1ee),
	.w8(32'h3bbf3142),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055bea),
	.w1(32'hbbb6944a),
	.w2(32'hbbe2e9f0),
	.w3(32'h3d1fea07),
	.w4(32'h3b9fe18f),
	.w5(32'hbb5c7482),
	.w6(32'h3c10fdf2),
	.w7(32'h3ac2f35b),
	.w8(32'hbb8f31f0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad70fc),
	.w1(32'hbc3ea7da),
	.w2(32'hbc026963),
	.w3(32'h3c5b011c),
	.w4(32'h3b820687),
	.w5(32'hbbca96b1),
	.w6(32'hbb16fbf3),
	.w7(32'h3c2a90e1),
	.w8(32'hbb5f1be2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e5a1),
	.w1(32'hbd10546f),
	.w2(32'h3c4a2392),
	.w3(32'hbb6e4515),
	.w4(32'h3d38f4e3),
	.w5(32'h3b942987),
	.w6(32'h3bc738a8),
	.w7(32'h3bc07267),
	.w8(32'h3c1be2f4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae7c5),
	.w1(32'hbd35acea),
	.w2(32'hbc49f7db),
	.w3(32'hbba07edb),
	.w4(32'hbbe1b271),
	.w5(32'hbc0370f1),
	.w6(32'hba9ac793),
	.w7(32'hbba2e056),
	.w8(32'h3c740c65),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8346ad),
	.w1(32'hba4427ce),
	.w2(32'h3bb5f7fe),
	.w3(32'hbbb217cd),
	.w4(32'h3abebc3f),
	.w5(32'h3c200bfe),
	.w6(32'hbbf101a8),
	.w7(32'hbb8c2087),
	.w8(32'h39c89664),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30fdea),
	.w1(32'hbb775674),
	.w2(32'h3b7e60a8),
	.w3(32'hbb846e42),
	.w4(32'hbbfa11e4),
	.w5(32'h3c4c3c18),
	.w6(32'h3d394713),
	.w7(32'hbbeceaf0),
	.w8(32'h3c11ee59),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4276c),
	.w1(32'hbb647566),
	.w2(32'hbb91c4e6),
	.w3(32'hbb18d4af),
	.w4(32'hbb36332c),
	.w5(32'h3c23432f),
	.w6(32'hbaf412dd),
	.w7(32'hbb385650),
	.w8(32'hbb450ed1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58bf05),
	.w1(32'hbc42c99b),
	.w2(32'h3c0fa096),
	.w3(32'h3a9a241e),
	.w4(32'hbc2d877f),
	.w5(32'hbc1387e2),
	.w6(32'h3a64394e),
	.w7(32'h3c05937f),
	.w8(32'h3bc52995),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8def5e),
	.w1(32'h3b96c529),
	.w2(32'h3ae60cae),
	.w3(32'hbb7d1c72),
	.w4(32'h3b8c4ac2),
	.w5(32'hbb72cb95),
	.w6(32'h3b1ea101),
	.w7(32'h3c0134f2),
	.w8(32'hbad765d3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e8f4),
	.w1(32'h3b2bd650),
	.w2(32'h3b8abd0c),
	.w3(32'h3bb3582a),
	.w4(32'hbbbd9f80),
	.w5(32'hb96b9a37),
	.w6(32'h3bfffb36),
	.w7(32'h3b186671),
	.w8(32'hbaa79a5b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa60947),
	.w1(32'hbb371ca9),
	.w2(32'h3cac372c),
	.w3(32'hbc132103),
	.w4(32'hbb5ec9f5),
	.w5(32'hbb6e4246),
	.w6(32'hba90a9f0),
	.w7(32'h3b00235f),
	.w8(32'hbc0fa773),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53df15),
	.w1(32'h3caf246a),
	.w2(32'hbb667f31),
	.w3(32'hba02d7dd),
	.w4(32'h3a17dd83),
	.w5(32'hbc873442),
	.w6(32'hbbb1a75a),
	.w7(32'hbb53bf7b),
	.w8(32'h3afd113d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bea15),
	.w1(32'h3ac591b5),
	.w2(32'h3b4485a9),
	.w3(32'h3b773b74),
	.w4(32'h3ae3506e),
	.w5(32'h3b995bda),
	.w6(32'hbb414a99),
	.w7(32'hbbdbfc51),
	.w8(32'hbc55fd0f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51cbb7),
	.w1(32'h3bc3a882),
	.w2(32'hbbdb2e42),
	.w3(32'hbbc1e53d),
	.w4(32'hba3d8041),
	.w5(32'h3a47d212),
	.w6(32'h3af887d3),
	.w7(32'h3bea3bc8),
	.w8(32'h3c91fc6e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba563ff3),
	.w1(32'hbc38c86c),
	.w2(32'h3ae0393e),
	.w3(32'hbb24142e),
	.w4(32'hb995d9e8),
	.w5(32'hbc3cb8ce),
	.w6(32'hb9b3383b),
	.w7(32'hbac0a722),
	.w8(32'h3c8096e4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cf87a),
	.w1(32'h3bbab19e),
	.w2(32'h3aec9a09),
	.w3(32'h3afc1b18),
	.w4(32'h3abb01b0),
	.w5(32'h3c100353),
	.w6(32'hbb5c2a6d),
	.w7(32'h3b4a224f),
	.w8(32'h3b286a4a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b731bf1),
	.w1(32'hbb01a5d8),
	.w2(32'hbc844100),
	.w3(32'h3b300f7f),
	.w4(32'hbbc1f722),
	.w5(32'h3a22ce5e),
	.w6(32'h3b8418ae),
	.w7(32'h3c52155c),
	.w8(32'hbbb2fdf2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd80424),
	.w1(32'hbb583efc),
	.w2(32'hbb85c777),
	.w3(32'h3b9b91d8),
	.w4(32'h3c2fdf88),
	.w5(32'h3b367067),
	.w6(32'hbb9cfadd),
	.w7(32'h3c8aaf5a),
	.w8(32'h3c16d886),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a732128),
	.w1(32'h3bc4c298),
	.w2(32'hba78aea5),
	.w3(32'hbbbe307a),
	.w4(32'h3c976860),
	.w5(32'h3a8fb34d),
	.w6(32'hb9c62524),
	.w7(32'hbb9d0b1e),
	.w8(32'h3a947242),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7176e2),
	.w1(32'hb9cd42bd),
	.w2(32'hbbca198e),
	.w3(32'hbaae66fb),
	.w4(32'hbc5840d8),
	.w5(32'hbbd1c246),
	.w6(32'hbbd516b1),
	.w7(32'hbb316214),
	.w8(32'hbb9755a8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba6f15),
	.w1(32'h3aba7239),
	.w2(32'h3bc906a7),
	.w3(32'hba92e425),
	.w4(32'hbb53dc8b),
	.w5(32'hbb1a67d2),
	.w6(32'hbbdadc80),
	.w7(32'hb987cdfc),
	.w8(32'hbb5906f0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab55519),
	.w1(32'h3b062754),
	.w2(32'h3c6a2056),
	.w3(32'h3bd155d1),
	.w4(32'h3b7e316a),
	.w5(32'hbb6e2d69),
	.w6(32'h3bc1820f),
	.w7(32'h3ca2525d),
	.w8(32'hbc3440da),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c22f0),
	.w1(32'hbac31c68),
	.w2(32'hbc0c7451),
	.w3(32'hbb28db04),
	.w4(32'h3a8ec88e),
	.w5(32'hbafe0055),
	.w6(32'hbaabd388),
	.w7(32'hbc2931db),
	.w8(32'h3c221946),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28295f),
	.w1(32'h3b55fd29),
	.w2(32'h3b54c2ef),
	.w3(32'h3b0f32d6),
	.w4(32'h3a25740d),
	.w5(32'hb98a8180),
	.w6(32'h3bd0b9ba),
	.w7(32'hba1b682b),
	.w8(32'h3bb024c2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ef9b5),
	.w1(32'hbb90f1fd),
	.w2(32'h3b0ff462),
	.w3(32'h3b3b1eb9),
	.w4(32'h3b527058),
	.w5(32'hb8d11806),
	.w6(32'hba67c07c),
	.w7(32'h3afba173),
	.w8(32'h3c6c8162),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9a5a3),
	.w1(32'h3bd43a5d),
	.w2(32'hb7903094),
	.w3(32'hb84e4a2a),
	.w4(32'hba24a110),
	.w5(32'hbad4a223),
	.w6(32'h3a172b42),
	.w7(32'h3b84fef4),
	.w8(32'h3909bd92),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aede87f),
	.w1(32'hbb67ba45),
	.w2(32'hbaffb130),
	.w3(32'h3b88fb1e),
	.w4(32'hbb6707f9),
	.w5(32'hb9e60796),
	.w6(32'h3a6384b0),
	.w7(32'hbb1866d0),
	.w8(32'hba90a32f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb643e),
	.w1(32'hbb919f64),
	.w2(32'hbb5f5d32),
	.w3(32'hbc11f7d2),
	.w4(32'hbbb9954c),
	.w5(32'h3b4cadf9),
	.w6(32'hb944de16),
	.w7(32'hbb48efe3),
	.w8(32'h3b4ead58),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48541),
	.w1(32'hbb1d6a32),
	.w2(32'hbb0c9ddc),
	.w3(32'hbae2ca80),
	.w4(32'hbb4d2f44),
	.w5(32'hba4909ba),
	.w6(32'hbacc9211),
	.w7(32'hbb942424),
	.w8(32'h3c01eac0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176c2c),
	.w1(32'hbb73453b),
	.w2(32'hb98cc5ba),
	.w3(32'h3a270f57),
	.w4(32'hbaf29113),
	.w5(32'hbae1d47b),
	.w6(32'hbb72f5c5),
	.w7(32'hbba0149e),
	.w8(32'hbab08968),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d5d0),
	.w1(32'h3a9ec672),
	.w2(32'hba924f9d),
	.w3(32'hba6d9796),
	.w4(32'h3a578d35),
	.w5(32'h3c059d55),
	.w6(32'hb950a22e),
	.w7(32'h3a1e1c37),
	.w8(32'hbbc5dc8c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1089c),
	.w1(32'h3b16cc53),
	.w2(32'hbb25b51c),
	.w3(32'hbc449df0),
	.w4(32'hba6e1674),
	.w5(32'h3bc82017),
	.w6(32'hbc155416),
	.w7(32'hbb4fb1b1),
	.w8(32'hb9bfd733),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3842a318),
	.w1(32'hbba96f22),
	.w2(32'h3b5d0dcd),
	.w3(32'hba93d79d),
	.w4(32'hbaf6a04a),
	.w5(32'h39fcf16e),
	.w6(32'h39fb0815),
	.w7(32'h3a8dc113),
	.w8(32'hbb841de3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae8b5),
	.w1(32'h3b2bde4f),
	.w2(32'hbba655b5),
	.w3(32'hbadaada7),
	.w4(32'hbab1ba24),
	.w5(32'hb9ae7c51),
	.w6(32'hb95f0b84),
	.w7(32'hba3c7e25),
	.w8(32'hbafd3f70),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64ce7),
	.w1(32'hbaea182f),
	.w2(32'hbb049e0a),
	.w3(32'h39632ff6),
	.w4(32'h3a9471e6),
	.w5(32'hbadea66e),
	.w6(32'hbb06e602),
	.w7(32'h3a38ff05),
	.w8(32'hbada1166),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82550e),
	.w1(32'hbb543688),
	.w2(32'hbb55ebba),
	.w3(32'hbb1d15c8),
	.w4(32'hbb396fad),
	.w5(32'h3b30b64e),
	.w6(32'hbb08a373),
	.w7(32'hba07de28),
	.w8(32'h3a4a60ff),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca299e),
	.w1(32'hbabc403d),
	.w2(32'hb9d4426e),
	.w3(32'hbacd2e6d),
	.w4(32'hbc773135),
	.w5(32'h3b90ddd3),
	.w6(32'h3a1b4756),
	.w7(32'h3b906cc7),
	.w8(32'h3b710ecf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc808acf),
	.w1(32'hbbf11bc2),
	.w2(32'hbc94b76d),
	.w3(32'hbae39d35),
	.w4(32'hba0d0940),
	.w5(32'hb9d93c19),
	.w6(32'hbacefa7b),
	.w7(32'hbac68f31),
	.w8(32'hba29f404),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0260cf),
	.w1(32'h3c0ec384),
	.w2(32'h3c1ec92d),
	.w3(32'h3c4695cb),
	.w4(32'hba134d54),
	.w5(32'h3b44f74c),
	.w6(32'hba95d1de),
	.w7(32'hbb576f16),
	.w8(32'hb9be00f9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75ada),
	.w1(32'hbb3d6624),
	.w2(32'hbb276271),
	.w3(32'h3d12ad3e),
	.w4(32'h39dac683),
	.w5(32'h3c23c204),
	.w6(32'h3ac9462b),
	.w7(32'h3c28354f),
	.w8(32'h3b15c734),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73cd7),
	.w1(32'h3bb56e2d),
	.w2(32'h3c05337f),
	.w3(32'hbb04fb9b),
	.w4(32'h3b564375),
	.w5(32'h3b3e7e6e),
	.w6(32'h3c104ff9),
	.w7(32'hbb9ed4c4),
	.w8(32'hbb6a108d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2ac35),
	.w1(32'hbc9d8d06),
	.w2(32'hbc6008b5),
	.w3(32'hbae5b876),
	.w4(32'h3b2008ff),
	.w5(32'hb9eac3b0),
	.w6(32'hbb8827e4),
	.w7(32'hbc180b54),
	.w8(32'hba11eb0b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08ccf),
	.w1(32'h3b568ce5),
	.w2(32'hbc255673),
	.w3(32'hb92181b6),
	.w4(32'hbb5c9b67),
	.w5(32'hbc7a821b),
	.w6(32'h3adc6f33),
	.w7(32'hbb0d4837),
	.w8(32'hbbe112a1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02f48),
	.w1(32'h3c287bb8),
	.w2(32'hbb76f79e),
	.w3(32'h3c30536a),
	.w4(32'h3a0ba701),
	.w5(32'hbc08e392),
	.w6(32'h3a84c813),
	.w7(32'hba12a40b),
	.w8(32'h3b060218),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dedd7),
	.w1(32'hb8a7c58c),
	.w2(32'h3ab47f1b),
	.w3(32'hbab2a63e),
	.w4(32'h3ac6b49a),
	.w5(32'hba1997bd),
	.w6(32'hbb9504a0),
	.w7(32'h3b2efbee),
	.w8(32'h3bd5eec0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91fe46),
	.w1(32'hbbc97499),
	.w2(32'h3c3a4dbe),
	.w3(32'hbc6765a2),
	.w4(32'hbac8b486),
	.w5(32'h39b2d52f),
	.w6(32'hbb8111e0),
	.w7(32'h3c19d6e2),
	.w8(32'hbb96012d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf7978),
	.w1(32'h3b770b56),
	.w2(32'h38c35aca),
	.w3(32'h3bc70f22),
	.w4(32'h3bbb14f0),
	.w5(32'h3b1a6f57),
	.w6(32'hb9b1e243),
	.w7(32'hbc6f0def),
	.w8(32'h3c17d3f2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb8ad),
	.w1(32'h3bab6d2e),
	.w2(32'hbb9cd5bb),
	.w3(32'hbb70f880),
	.w4(32'h3a4026d9),
	.w5(32'h3b135f7c),
	.w6(32'h3ac3ab8d),
	.w7(32'h3c00fbf0),
	.w8(32'hbc873259),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d05e3b),
	.w1(32'hbb739ea9),
	.w2(32'hbb7809a7),
	.w3(32'hbbbf0d99),
	.w4(32'hbbf05143),
	.w5(32'h39ddd80b),
	.w6(32'hbbc13d43),
	.w7(32'hbb8733e3),
	.w8(32'h3b6cb5a7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd95c46),
	.w1(32'h39aa23bc),
	.w2(32'h3b17411d),
	.w3(32'h3af60648),
	.w4(32'hbbd66155),
	.w5(32'h3c282dc1),
	.w6(32'hbbe3f7dd),
	.w7(32'h3b22d49e),
	.w8(32'hbb1a4425),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be478cf),
	.w1(32'hbac132dd),
	.w2(32'hbcec403e),
	.w3(32'h3b91f5af),
	.w4(32'hbb77f633),
	.w5(32'h3ac1a26d),
	.w6(32'hbbbb2000),
	.w7(32'hbba8a126),
	.w8(32'hbbb3bcf3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b292671),
	.w1(32'h3b7b2b94),
	.w2(32'h3973c694),
	.w3(32'h3c8340d6),
	.w4(32'h3b5efdac),
	.w5(32'hbb88d2d6),
	.w6(32'hbc9b3957),
	.w7(32'hba49dd82),
	.w8(32'hbc7fe68d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a15f4),
	.w1(32'hbca62fca),
	.w2(32'hbcb87da3),
	.w3(32'hbbb00b19),
	.w4(32'hbcc4aaf6),
	.w5(32'hbc153bab),
	.w6(32'hbb8c3e4a),
	.w7(32'hba86f87a),
	.w8(32'hbca08941),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf6b36),
	.w1(32'hbc1bb1d6),
	.w2(32'hbcbff0d0),
	.w3(32'hbc4863e2),
	.w4(32'hbc99dd39),
	.w5(32'hbb9c04c1),
	.w6(32'hbc8ca088),
	.w7(32'h3d063466),
	.w8(32'hbb7749c8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule