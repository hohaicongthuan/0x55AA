module layer_10_featuremap_56(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f27f),
	.w1(32'hbc56a556),
	.w2(32'h3c9fb597),
	.w3(32'h3c0f4f00),
	.w4(32'hbb4a310d),
	.w5(32'hbbe90ed9),
	.w6(32'h3bcda80a),
	.w7(32'hba03609a),
	.w8(32'h3b260354),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c277a07),
	.w1(32'hba2ae41a),
	.w2(32'hbb82d066),
	.w3(32'hbcbe9e9a),
	.w4(32'hbc0f8c40),
	.w5(32'h3c0d37f2),
	.w6(32'hbc57a3aa),
	.w7(32'hbb84f199),
	.w8(32'hbb7b3ab9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e50ff),
	.w1(32'h3cbd49ef),
	.w2(32'hba6e900f),
	.w3(32'hb962e2b2),
	.w4(32'h3b2902bf),
	.w5(32'h3ad54fb8),
	.w6(32'hb90eba76),
	.w7(32'hb9e453ad),
	.w8(32'h3b2e0bf4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaf7f5),
	.w1(32'hbc120881),
	.w2(32'hbb8d423a),
	.w3(32'h3a930799),
	.w4(32'h3a73b913),
	.w5(32'hba7d4f31),
	.w6(32'h3b40836a),
	.w7(32'h3c2ef9ef),
	.w8(32'h3c052303),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19ad46),
	.w1(32'hba8751cb),
	.w2(32'hbbf17595),
	.w3(32'hbc4b0dd4),
	.w4(32'hbc55e280),
	.w5(32'h3cfe90e0),
	.w6(32'h3a585922),
	.w7(32'hbc17dadd),
	.w8(32'h3b2a2bcb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db4bb),
	.w1(32'hbb68b83f),
	.w2(32'h38609780),
	.w3(32'h3d0d1b66),
	.w4(32'h3c5133e4),
	.w5(32'h3b84f4d0),
	.w6(32'h3cc88010),
	.w7(32'h3c8f69d9),
	.w8(32'h3b4ea0cc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f856a),
	.w1(32'hbb48beb8),
	.w2(32'h3b38c04c),
	.w3(32'hbc6053f8),
	.w4(32'hbbef483a),
	.w5(32'h3c407c01),
	.w6(32'hbc546022),
	.w7(32'hbbec63be),
	.w8(32'h3c3e1eca),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a5de3),
	.w1(32'h3c889287),
	.w2(32'h3c206ad2),
	.w3(32'h3b0f9066),
	.w4(32'h3b9937cf),
	.w5(32'h3c1d7db0),
	.w6(32'h3bf8a382),
	.w7(32'hba81a83f),
	.w8(32'hbb581562),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0bb65),
	.w1(32'h3bae7655),
	.w2(32'h3c164258),
	.w3(32'hba88c694),
	.w4(32'h3a3f0f79),
	.w5(32'hbaef03f4),
	.w6(32'hbb022f9a),
	.w7(32'hbb2086c0),
	.w8(32'hbba5b40c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c400835),
	.w1(32'h3c2acfbf),
	.w2(32'h3b3e035f),
	.w3(32'hba75647b),
	.w4(32'h3ba3001b),
	.w5(32'h3b0a194f),
	.w6(32'hbc3728b4),
	.w7(32'h3afb6c42),
	.w8(32'h3b347ef9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb1e0),
	.w1(32'h3a80ad88),
	.w2(32'h3bfaea70),
	.w3(32'h3a61e3db),
	.w4(32'hba4c9944),
	.w5(32'h3b935766),
	.w6(32'hbab875d9),
	.w7(32'hbae8ebcf),
	.w8(32'hbab1a65d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e29b),
	.w1(32'hbc84765f),
	.w2(32'h3c2d441b),
	.w3(32'hb9c36919),
	.w4(32'hbb36b44d),
	.w5(32'h3bd9b63b),
	.w6(32'hbbd77e94),
	.w7(32'hba92126d),
	.w8(32'h3c0033aa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade5087),
	.w1(32'h3af17cef),
	.w2(32'h3baa4789),
	.w3(32'hb9d539d5),
	.w4(32'hbafa7a6f),
	.w5(32'h3c1fbde5),
	.w6(32'hbbd2bbe5),
	.w7(32'hbc0c6a42),
	.w8(32'hba8fa5ac),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95f8c2),
	.w1(32'h3ba42c2f),
	.w2(32'h3b1b06e6),
	.w3(32'hba07617c),
	.w4(32'h3b6151dd),
	.w5(32'hbbe361e9),
	.w6(32'hba88170f),
	.w7(32'hb9ce21f5),
	.w8(32'h3bf4add0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431719),
	.w1(32'h3b61c3dc),
	.w2(32'hbb9aa0a7),
	.w3(32'hbb94e5b0),
	.w4(32'h3aff91eb),
	.w5(32'h3adf2af3),
	.w6(32'h3c1e1de6),
	.w7(32'h3bd403c0),
	.w8(32'h39d46189),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff6ac),
	.w1(32'h3bb50a75),
	.w2(32'h3af2cd3f),
	.w3(32'h3b861d8a),
	.w4(32'h3a738ce6),
	.w5(32'h3b7bea39),
	.w6(32'h3bf462af),
	.w7(32'h3be5488d),
	.w8(32'h3b9826d8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fb45e),
	.w1(32'hbaeac10c),
	.w2(32'h3b7eade4),
	.w3(32'hb94490c6),
	.w4(32'hbac4622b),
	.w5(32'h3ad80abb),
	.w6(32'hba440d3c),
	.w7(32'hbb025ba9),
	.w8(32'h3b51a844),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c9f84),
	.w1(32'h3cd58168),
	.w2(32'h3d0c5c49),
	.w3(32'h3c29ee6a),
	.w4(32'h3cabbbef),
	.w5(32'h3c4a80d3),
	.w6(32'h3c990105),
	.w7(32'h3caf41b4),
	.w8(32'h3c2d8ac9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841612),
	.w1(32'h3bedc665),
	.w2(32'h3c19839c),
	.w3(32'h3bf3926d),
	.w4(32'h3c11a4af),
	.w5(32'hbc49db6d),
	.w6(32'hb89af626),
	.w7(32'h3b2f2637),
	.w8(32'h3c4edecb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce209),
	.w1(32'h3b22b640),
	.w2(32'h3b135731),
	.w3(32'hbcdbd7cc),
	.w4(32'hbc8d361d),
	.w5(32'h3b9d12f2),
	.w6(32'hb8938628),
	.w7(32'hbbaccbec),
	.w8(32'h3b393232),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af57ae7),
	.w1(32'h3aa90597),
	.w2(32'h3c0beb24),
	.w3(32'h3b50add1),
	.w4(32'hb9ecaa35),
	.w5(32'h3b8cdfd1),
	.w6(32'h3b0bc90a),
	.w7(32'h3ab06f5d),
	.w8(32'hbbbb6c84),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2771),
	.w1(32'h3c022ab6),
	.w2(32'hbb8d0ae5),
	.w3(32'hbc3a7939),
	.w4(32'hbc07eae9),
	.w5(32'hbbaf0dd8),
	.w6(32'hbd036a59),
	.w7(32'hbc7284e8),
	.w8(32'hbaba6950),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a8ea3),
	.w1(32'h3c371465),
	.w2(32'h3d04e440),
	.w3(32'h3bc65533),
	.w4(32'h3bd14444),
	.w5(32'h3c6b4002),
	.w6(32'h3c279540),
	.w7(32'h3b50102a),
	.w8(32'h3c245498),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a48bc),
	.w1(32'h3aa31b7a),
	.w2(32'hbb0b7d72),
	.w3(32'hba426035),
	.w4(32'hbb390647),
	.w5(32'hba01b871),
	.w6(32'hbbe00125),
	.w7(32'hbb4dd8e3),
	.w8(32'h3bad6a0e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a828a9f),
	.w1(32'hbc0e87c8),
	.w2(32'hbbf673a8),
	.w3(32'h3b856a06),
	.w4(32'hbc1ae3d4),
	.w5(32'hbc5dcacc),
	.w6(32'h3b876ba5),
	.w7(32'h3c14f576),
	.w8(32'h3b714608),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9954b0),
	.w1(32'h39f67f79),
	.w2(32'hb97733c8),
	.w3(32'hbc8a9df9),
	.w4(32'hbc15519b),
	.w5(32'hbb8769d8),
	.w6(32'h3ca413f7),
	.w7(32'h3c488064),
	.w8(32'h3c4004f4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae172fb),
	.w1(32'h3cb35653),
	.w2(32'hb9a18f94),
	.w3(32'hbca62d9d),
	.w4(32'hbc50dc5a),
	.w5(32'hba093d3a),
	.w6(32'h3c2181d4),
	.w7(32'hbabb9ac6),
	.w8(32'hba948ddd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c784a),
	.w1(32'h37cafb30),
	.w2(32'hbc773660),
	.w3(32'h3a953228),
	.w4(32'hbb8c0d52),
	.w5(32'hbba5ac60),
	.w6(32'hbb2d084b),
	.w7(32'h3bac393c),
	.w8(32'h3c2a7611),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8e21),
	.w1(32'hbba62e11),
	.w2(32'h3c2bef02),
	.w3(32'hbb5554df),
	.w4(32'h3a3b42ce),
	.w5(32'h3c2f3702),
	.w6(32'h3aae99e2),
	.w7(32'hbb70d262),
	.w8(32'h3c910451),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c554c),
	.w1(32'hbbb6e5de),
	.w2(32'hbbbd2eef),
	.w3(32'h3cfbd58a),
	.w4(32'hbb93dcfd),
	.w5(32'hbbbc5a09),
	.w6(32'h3cdffcab),
	.w7(32'h3c6556e2),
	.w8(32'h38ba1931),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bd1f5),
	.w1(32'h3a32d6d6),
	.w2(32'h3ba2750c),
	.w3(32'h3b002779),
	.w4(32'h39f7957a),
	.w5(32'h3af97025),
	.w6(32'h3aab92a8),
	.w7(32'h3a25934f),
	.w8(32'h3aeb35ed),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b541963),
	.w1(32'hbb69f3a8),
	.w2(32'h3bb47e73),
	.w3(32'hb9cba447),
	.w4(32'hbbfced53),
	.w5(32'h3b76623b),
	.w6(32'hbae5e021),
	.w7(32'hb9d02c3d),
	.w8(32'h3c364bdd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5653),
	.w1(32'h3b70049a),
	.w2(32'hbaaed9c4),
	.w3(32'h3ba634af),
	.w4(32'h3c217664),
	.w5(32'hbb0a6395),
	.w6(32'hbb5d33e3),
	.w7(32'h3b02e2ef),
	.w8(32'hbb6b7aa4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d613f1),
	.w1(32'hbb935cff),
	.w2(32'h3a739ed1),
	.w3(32'hbb663ab4),
	.w4(32'hbbe16886),
	.w5(32'hbb0f5f56),
	.w6(32'hbb20d717),
	.w7(32'hba0ad186),
	.w8(32'hbae11783),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae30244),
	.w1(32'hbbabb8b4),
	.w2(32'hbbb6f38e),
	.w3(32'hbac94b2c),
	.w4(32'hbb824115),
	.w5(32'hbb51bec7),
	.w6(32'h3affa282),
	.w7(32'h3c109102),
	.w8(32'hba0839fc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aa51d),
	.w1(32'hbb865976),
	.w2(32'h3c0083b8),
	.w3(32'hbbb61efd),
	.w4(32'hbbcf9d46),
	.w5(32'h3c153128),
	.w6(32'hbbafd04d),
	.w7(32'hbbca3770),
	.w8(32'h3c28ba8e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b30fe),
	.w1(32'hbcbf10cb),
	.w2(32'h3bf49c21),
	.w3(32'hbbbd95a7),
	.w4(32'hbc81b98f),
	.w5(32'hbbb1619b),
	.w6(32'h3c1b49ff),
	.w7(32'hbc4b5b72),
	.w8(32'hbc4dfe41),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9962d4e),
	.w1(32'hbcd2d851),
	.w2(32'hbcb5b666),
	.w3(32'hbbfabaa7),
	.w4(32'hbcdf4d06),
	.w5(32'hbbb99554),
	.w6(32'hbbd452a9),
	.w7(32'hbc04fd61),
	.w8(32'hb986edc0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bb1c6),
	.w1(32'hbc80b45d),
	.w2(32'hbc426b8b),
	.w3(32'hbc222bf5),
	.w4(32'hbcf9156d),
	.w5(32'hbb8c3897),
	.w6(32'hbc80b500),
	.w7(32'hbb258943),
	.w8(32'h3bd97cb3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c9b1f),
	.w1(32'h3c027c3b),
	.w2(32'hbb80f279),
	.w3(32'hbb6fa160),
	.w4(32'h3c23e8a8),
	.w5(32'hbb061fd9),
	.w6(32'hbac9a5eb),
	.w7(32'h3b633f7b),
	.w8(32'hbb8a7852),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94eab),
	.w1(32'hbbf1bd4e),
	.w2(32'hbb2f4a72),
	.w3(32'hbb9cccb8),
	.w4(32'hbc0d8843),
	.w5(32'hbb00bfa6),
	.w6(32'hbc0e3401),
	.w7(32'hbc0afd5f),
	.w8(32'hbb5261fa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cd90),
	.w1(32'h3a35c9cb),
	.w2(32'h3b1b99a6),
	.w3(32'hbaa4649d),
	.w4(32'hbba39499),
	.w5(32'h3aad677b),
	.w6(32'hbac021b4),
	.w7(32'hbb55c90a),
	.w8(32'hbaa58351),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c056704),
	.w1(32'h3beedb11),
	.w2(32'hbc066c9e),
	.w3(32'h3c202f4c),
	.w4(32'hbb33d037),
	.w5(32'hbb9f0f5d),
	.w6(32'h3aa0301b),
	.w7(32'hbb48d4cf),
	.w8(32'hbab207e2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405614),
	.w1(32'h3b17db7e),
	.w2(32'hbac9e147),
	.w3(32'h3b1a463f),
	.w4(32'h390a00f4),
	.w5(32'h3b0f37f0),
	.w6(32'hba1f3608),
	.w7(32'hba19875b),
	.w8(32'h3b1c89a0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd23509),
	.w1(32'hba1a06a9),
	.w2(32'h3ade62e8),
	.w3(32'h3c773e79),
	.w4(32'hbb8b330b),
	.w5(32'h3bd73e47),
	.w6(32'h3bcca7ea),
	.w7(32'h39b860d7),
	.w8(32'h3bdf7515),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c4af0),
	.w1(32'hbb7caa47),
	.w2(32'h3b50b1ed),
	.w3(32'h3b126e0e),
	.w4(32'hbc885577),
	.w5(32'h3b7d2926),
	.w6(32'h3989658a),
	.w7(32'hbb3c4758),
	.w8(32'h39efa294),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb0ce2),
	.w1(32'h3c219f61),
	.w2(32'h3a986d47),
	.w3(32'h3bfc316f),
	.w4(32'h3bc86718),
	.w5(32'h3b3fcfca),
	.w6(32'h3ca1e4d5),
	.w7(32'h3bcec37e),
	.w8(32'h3b8add48),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3a0ee),
	.w1(32'h3cb3c70e),
	.w2(32'h3ccedf02),
	.w3(32'h3b4c4e0f),
	.w4(32'h3bdd0bf6),
	.w5(32'h3c82a2eb),
	.w6(32'h3c439196),
	.w7(32'h3b61ac08),
	.w8(32'h3c38cadd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87b543),
	.w1(32'hbb81cb46),
	.w2(32'hbaeb2489),
	.w3(32'hbb4f098b),
	.w4(32'hbb5b1a09),
	.w5(32'h3b85c57f),
	.w6(32'hbb03070e),
	.w7(32'hbb6ec5e0),
	.w8(32'hbc2a96b6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b603020),
	.w1(32'h3bfabe4a),
	.w2(32'h3c009ba7),
	.w3(32'hb9b15111),
	.w4(32'hbba49825),
	.w5(32'hba76c5f1),
	.w6(32'h3bf60131),
	.w7(32'h3b39f016),
	.w8(32'h3aa76fba),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c2050),
	.w1(32'hbb71579d),
	.w2(32'h3b1deeff),
	.w3(32'hbb13f52d),
	.w4(32'h3b40d3ce),
	.w5(32'hba9a4dc3),
	.w6(32'h3b9b1e12),
	.w7(32'h3b634fcf),
	.w8(32'h3bbcf8bd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d043d),
	.w1(32'h3c49170d),
	.w2(32'h3a951956),
	.w3(32'h3b73fac1),
	.w4(32'h3be97c5f),
	.w5(32'h3bbf638c),
	.w6(32'h3a7a4757),
	.w7(32'h3b97bec2),
	.w8(32'h3958c7b8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd840b),
	.w1(32'h3b7e62d8),
	.w2(32'h3b785800),
	.w3(32'h3c0fe365),
	.w4(32'h3b2f893f),
	.w5(32'h3b3ba2b1),
	.w6(32'h3b2bcde6),
	.w7(32'h3b99ac1b),
	.w8(32'hbb90bd77),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a917b50),
	.w1(32'h3c4a8b24),
	.w2(32'h3cd1ed90),
	.w3(32'h3aaec2a2),
	.w4(32'h3c09f988),
	.w5(32'h3cbc2fdf),
	.w6(32'h3aa5a609),
	.w7(32'h3ba244e0),
	.w8(32'h3c9a829b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6af57),
	.w1(32'hbb461953),
	.w2(32'h3be95a66),
	.w3(32'h3cf586a5),
	.w4(32'h3901a601),
	.w5(32'hbb1cda8f),
	.w6(32'h3c90c71e),
	.w7(32'h3c2afc5f),
	.w8(32'h3b829730),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab32b1),
	.w1(32'hbb6aa0b1),
	.w2(32'h3ade9283),
	.w3(32'hbb48b44a),
	.w4(32'h3948635b),
	.w5(32'hbb46e50e),
	.w6(32'hbba4c8b5),
	.w7(32'hbc31f9f1),
	.w8(32'h3b2374b1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06af17),
	.w1(32'hba1780af),
	.w2(32'hbb16ca36),
	.w3(32'h3b5b6003),
	.w4(32'h3b53baf5),
	.w5(32'hbb7d6a53),
	.w6(32'h3acbe0e1),
	.w7(32'hbbe6068a),
	.w8(32'h3af7b4e0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1417af),
	.w1(32'hbade5ec9),
	.w2(32'hba773d5a),
	.w3(32'hba5023f7),
	.w4(32'hba9e3afb),
	.w5(32'hbae3266a),
	.w6(32'h3b6f9c85),
	.w7(32'h3b760c3c),
	.w8(32'hbbf0f321),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0f59f),
	.w1(32'hbbcd3fdc),
	.w2(32'hbc0d7db9),
	.w3(32'hba7ca779),
	.w4(32'hbbde3a41),
	.w5(32'hbbc407df),
	.w6(32'hbc07768d),
	.w7(32'hbc419a41),
	.w8(32'h3ad4697f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c3e63),
	.w1(32'h3b1062c7),
	.w2(32'h3badb717),
	.w3(32'hbb965765),
	.w4(32'hbab85b52),
	.w5(32'h3bc615ab),
	.w6(32'h3a07a775),
	.w7(32'hb9a9094e),
	.w8(32'h3b2a950c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4eca),
	.w1(32'h3c13a908),
	.w2(32'h3b2c61f6),
	.w3(32'h3c0cfda8),
	.w4(32'h3bdc22bd),
	.w5(32'h3a8011ec),
	.w6(32'h3c30eb62),
	.w7(32'h3bbdd4ea),
	.w8(32'h3c0bf2cd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f250d),
	.w1(32'h3c6de36e),
	.w2(32'h39afd401),
	.w3(32'h3c9b2c8f),
	.w4(32'h3c98925d),
	.w5(32'hb9df493e),
	.w6(32'h3c516403),
	.w7(32'h3aa573c3),
	.w8(32'h3b485bf5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb030da),
	.w1(32'h3bf8e67a),
	.w2(32'hbb26145f),
	.w3(32'hba30f1cf),
	.w4(32'h3b86c5d2),
	.w5(32'h3a495c03),
	.w6(32'h3ad43260),
	.w7(32'hbb287d03),
	.w8(32'hbb0385a2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5516cb),
	.w1(32'hbb8ca0ad),
	.w2(32'h3ab2535b),
	.w3(32'h3ab14637),
	.w4(32'hbadcdbbe),
	.w5(32'hbb2d8877),
	.w6(32'hba81c7c9),
	.w7(32'hbb74bc9e),
	.w8(32'h3b844408),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b2a078),
	.w1(32'h3a669ffd),
	.w2(32'h38a63bdd),
	.w3(32'hbbaf7e16),
	.w4(32'hbaea65bf),
	.w5(32'h3a82a34e),
	.w6(32'hbb4bd975),
	.w7(32'hbbc9a464),
	.w8(32'h3a8c52b9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1592b8),
	.w1(32'hbb10058b),
	.w2(32'hb73efe00),
	.w3(32'h3a9d86b8),
	.w4(32'hba649a74),
	.w5(32'h3b0a7d21),
	.w6(32'hbb25bd86),
	.w7(32'hbb7ac398),
	.w8(32'h3b0f45bf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe3d60),
	.w1(32'h3bd8b7cd),
	.w2(32'h3b45f1c6),
	.w3(32'h3b932677),
	.w4(32'h3c7f9cba),
	.w5(32'h3b50bedf),
	.w6(32'h3bcf0cb4),
	.w7(32'h3c6644a3),
	.w8(32'h3c075f3e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998c8f),
	.w1(32'hbb3f9cbb),
	.w2(32'h3b80f0fe),
	.w3(32'hbb897c73),
	.w4(32'hbc010ecc),
	.w5(32'h3c337273),
	.w6(32'hb897313b),
	.w7(32'hb9e76f45),
	.w8(32'hba9e0cf7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838f2a),
	.w1(32'h3c993d89),
	.w2(32'h3c80897b),
	.w3(32'h3b017a13),
	.w4(32'h3bf9ca07),
	.w5(32'h3bdf983d),
	.w6(32'h3bc4b0e2),
	.w7(32'h3c0979cf),
	.w8(32'h3c3e9d52),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c481d65),
	.w1(32'hbb685245),
	.w2(32'hbc84bfa0),
	.w3(32'h3b337522),
	.w4(32'hbc5ef161),
	.w5(32'hbbf132ac),
	.w6(32'h3a882567),
	.w7(32'h3bb88fa2),
	.w8(32'h3b1ddf74),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5efa9d),
	.w1(32'h3bd9afdd),
	.w2(32'hbb89955a),
	.w3(32'hbba40d37),
	.w4(32'h3b665541),
	.w5(32'hbb0f3fc2),
	.w6(32'hbb9929b5),
	.w7(32'h3b1c9b06),
	.w8(32'h3ab80b52),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3325e6),
	.w1(32'h3a95abc5),
	.w2(32'hbb35109e),
	.w3(32'hbbc1c814),
	.w4(32'h3ad736f7),
	.w5(32'h3b151ac0),
	.w6(32'hbbbedbf2),
	.w7(32'hbbccdb83),
	.w8(32'h3bd19f2f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ce812),
	.w1(32'h3b46e210),
	.w2(32'h3b0721c0),
	.w3(32'hba9dd3c9),
	.w4(32'h3bdfd837),
	.w5(32'h3b4a3ca0),
	.w6(32'h3c3b174d),
	.w7(32'h3b46619c),
	.w8(32'h3b1c87b2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cedc0b),
	.w1(32'hbb5504b3),
	.w2(32'hba8b52eb),
	.w3(32'h3b90b096),
	.w4(32'hbb7d33b6),
	.w5(32'h3acb5bbf),
	.w6(32'h3ad2877b),
	.w7(32'hbbe74129),
	.w8(32'h3a550f52),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f92f),
	.w1(32'hbba83216),
	.w2(32'h3957fddc),
	.w3(32'hbbc3995f),
	.w4(32'hbbbad14d),
	.w5(32'hb991b61d),
	.w6(32'hbb970438),
	.w7(32'hbbea9430),
	.w8(32'hbab7f95c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc096e),
	.w1(32'h3a299214),
	.w2(32'h3c7b1d30),
	.w3(32'hbbe802c9),
	.w4(32'hba710497),
	.w5(32'h3c5b7e36),
	.w6(32'h39270a8a),
	.w7(32'hbade90f3),
	.w8(32'h3ab7d310),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d3d1e),
	.w1(32'h3c49124e),
	.w2(32'h3cb5cea5),
	.w3(32'hbabe6d2a),
	.w4(32'h3bdd6f54),
	.w5(32'h3ca3a899),
	.w6(32'h3ae8386b),
	.w7(32'h3c5079ab),
	.w8(32'h3c4f5ad7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0e81),
	.w1(32'hbb0665de),
	.w2(32'hbb211ffc),
	.w3(32'h3acfc2ee),
	.w4(32'h3afb788a),
	.w5(32'h3ba6b58e),
	.w6(32'h3c1c23fb),
	.w7(32'hba9160d6),
	.w8(32'h3bff8a08),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6221dc),
	.w1(32'h3b5fc708),
	.w2(32'h3b698cd5),
	.w3(32'h3c31562f),
	.w4(32'h3bb959bd),
	.w5(32'hb99d1b5a),
	.w6(32'h3b7ed5ca),
	.w7(32'h3b56eb38),
	.w8(32'h3a9f0d54),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba404a23),
	.w1(32'h39d766ef),
	.w2(32'h3b963259),
	.w3(32'hbb7a2ec2),
	.w4(32'h3a225067),
	.w5(32'h3b24f61d),
	.w6(32'hbb140b12),
	.w7(32'h3b78092f),
	.w8(32'h3b02b1ab),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beed850),
	.w1(32'h3b4f906f),
	.w2(32'hba4237a9),
	.w3(32'h3b172e3e),
	.w4(32'hba5a560e),
	.w5(32'hbb607144),
	.w6(32'hbaabf464),
	.w7(32'h3ad0054d),
	.w8(32'hbb8d1d88),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab374d7),
	.w1(32'h3ba7cf2b),
	.w2(32'h3b6c34ba),
	.w3(32'hb98d73c7),
	.w4(32'h3bac3651),
	.w5(32'h3c74d678),
	.w6(32'hb96dfdb0),
	.w7(32'h3aa1af4c),
	.w8(32'h3c281981),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed9f95),
	.w1(32'h3c2395c2),
	.w2(32'hbb3048e1),
	.w3(32'h3a950f3e),
	.w4(32'h3bfaea87),
	.w5(32'h3a0b081d),
	.w6(32'h3c31d4fc),
	.w7(32'h3c554c02),
	.w8(32'h3a26d030),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be42b),
	.w1(32'h3c438712),
	.w2(32'hbb03d371),
	.w3(32'h3ba879d9),
	.w4(32'hbb686f98),
	.w5(32'h3a864adb),
	.w6(32'h3c1a7b48),
	.w7(32'hba9451bf),
	.w8(32'h3b81f078),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba733ed1),
	.w1(32'h3af6acda),
	.w2(32'hbbd1e3f2),
	.w3(32'h3bae7ce0),
	.w4(32'h3bc8d1b5),
	.w5(32'h3b19cedd),
	.w6(32'h3b8457d1),
	.w7(32'h3b084e4e),
	.w8(32'h3c7ac58f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95c55b),
	.w1(32'h3be2b8d9),
	.w2(32'hbb175515),
	.w3(32'hbc037cdb),
	.w4(32'hb9841321),
	.w5(32'hb9a72e8b),
	.w6(32'h3b68eff4),
	.w7(32'h3c152030),
	.w8(32'h3b46fcf3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda8dc9),
	.w1(32'hbbcce810),
	.w2(32'hbba84741),
	.w3(32'h3a781454),
	.w4(32'hbbd3972a),
	.w5(32'hbafe4412),
	.w6(32'h3b05212e),
	.w7(32'hb98d5bb2),
	.w8(32'hbb3dccaf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ad083),
	.w1(32'h3a756bd7),
	.w2(32'h3c3ea142),
	.w3(32'hbab9d164),
	.w4(32'h3a5a97e1),
	.w5(32'h3bb8f6ba),
	.w6(32'hb783caa2),
	.w7(32'h3ab78f3e),
	.w8(32'hbbaa64ce),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d47be),
	.w1(32'h3a6eba21),
	.w2(32'h3b6680a7),
	.w3(32'h3adccf92),
	.w4(32'hbc06b442),
	.w5(32'hbb9faa51),
	.w6(32'h3bc8e827),
	.w7(32'h3c0b2542),
	.w8(32'hbbb3b623),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34584c),
	.w1(32'h3c5ae0ef),
	.w2(32'h3ba5ec53),
	.w3(32'h39b139b3),
	.w4(32'h3c116a85),
	.w5(32'h3b7ad3d8),
	.w6(32'h3c8de0e3),
	.w7(32'h3c0964fa),
	.w8(32'h3bac1adb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87353f),
	.w1(32'hbc45a129),
	.w2(32'hbb87494b),
	.w3(32'hbad617d5),
	.w4(32'hbc108ef5),
	.w5(32'h3a2fe7d6),
	.w6(32'hbb4b5497),
	.w7(32'hbb844c6e),
	.w8(32'hba19dae7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfb908),
	.w1(32'hbb8b27d9),
	.w2(32'h3b9b72a9),
	.w3(32'h3c25ace3),
	.w4(32'h3c1a14bb),
	.w5(32'hbbb9800d),
	.w6(32'h3a94d6a7),
	.w7(32'h3b143a19),
	.w8(32'h3a460eef),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034f52),
	.w1(32'hbc3bfd7d),
	.w2(32'hbbe828d8),
	.w3(32'hbc0db868),
	.w4(32'hbc808a65),
	.w5(32'hbbcb3928),
	.w6(32'h39e8af4a),
	.w7(32'hbbfd53cf),
	.w8(32'hbb74fab3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945a89),
	.w1(32'h3bda8299),
	.w2(32'h3c01a96c),
	.w3(32'h392e7671),
	.w4(32'h3baaaadd),
	.w5(32'h3b892b37),
	.w6(32'h3ae4f1c3),
	.w7(32'h3bc68964),
	.w8(32'h3bcb7f1e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4343),
	.w1(32'h3ad2bd61),
	.w2(32'hbaaa8396),
	.w3(32'hb87b6b09),
	.w4(32'h3a529114),
	.w5(32'h3c6297b8),
	.w6(32'h3b2a0d99),
	.w7(32'h3afdd210),
	.w8(32'h3bfac135),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad895),
	.w1(32'hbb8b0914),
	.w2(32'hbba906e5),
	.w3(32'h3c05ebeb),
	.w4(32'hbc3e798f),
	.w5(32'hbb60d680),
	.w6(32'h3ca1b377),
	.w7(32'hbb81362c),
	.w8(32'hbc1594d7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b1ab),
	.w1(32'hbb09d8e3),
	.w2(32'hbaef009b),
	.w3(32'hbbe9ca8b),
	.w4(32'hbb9c1291),
	.w5(32'hbb4f7ce5),
	.w6(32'h3b3c211f),
	.w7(32'hbaa3109c),
	.w8(32'hbc0e85e2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ecaa2),
	.w1(32'h3bfb03bb),
	.w2(32'h3bb2e5df),
	.w3(32'h3bc2a523),
	.w4(32'h3c1a8f9d),
	.w5(32'h3ab44915),
	.w6(32'h3accdefa),
	.w7(32'hbb09c057),
	.w8(32'h39fff903),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fb715),
	.w1(32'hbbde0d57),
	.w2(32'hbaf2c671),
	.w3(32'hbc380d67),
	.w4(32'hbba64ff0),
	.w5(32'hbc2d1598),
	.w6(32'h3b36fcd5),
	.w7(32'hba8f13ff),
	.w8(32'hbb8e101a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d0ba),
	.w1(32'h3b8f6a39),
	.w2(32'h3cdfa8cd),
	.w3(32'h3c1830b1),
	.w4(32'h3c33f897),
	.w5(32'h3c3e5eb5),
	.w6(32'h3c61c539),
	.w7(32'h3c389cc2),
	.w8(32'hbc187229),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27aca3),
	.w1(32'hbc4bd13a),
	.w2(32'hbc4d6853),
	.w3(32'h3ae562d8),
	.w4(32'hbcfc9082),
	.w5(32'hbb8598ea),
	.w6(32'hbb756f86),
	.w7(32'hbc014374),
	.w8(32'h3b7402ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcda084),
	.w1(32'hbb0848f2),
	.w2(32'hbc4f29c0),
	.w3(32'hbb17e128),
	.w4(32'hbc99bf6b),
	.w5(32'hbbcb09fe),
	.w6(32'hba5bc18a),
	.w7(32'hbbad937c),
	.w8(32'hbb12c095),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4228b4),
	.w1(32'hbb73d2e2),
	.w2(32'h3c2bf719),
	.w3(32'hbbd9a656),
	.w4(32'hbc1b821e),
	.w5(32'hbba29a68),
	.w6(32'h391db2e7),
	.w7(32'hbc55fa34),
	.w8(32'hbb7706b2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d86dc),
	.w1(32'h3b951c86),
	.w2(32'h3bcce95c),
	.w3(32'hbb08df19),
	.w4(32'h3ac98d10),
	.w5(32'h3b4b3db0),
	.w6(32'hbb53cc6d),
	.w7(32'h3b441834),
	.w8(32'h3ada018c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2854dc),
	.w1(32'h3b6fd207),
	.w2(32'h3d040839),
	.w3(32'h3becdd06),
	.w4(32'h3c960257),
	.w5(32'h3c7e8910),
	.w6(32'h3cb1962f),
	.w7(32'h3ca4071a),
	.w8(32'h3abc333f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0dfc4),
	.w1(32'hbbaf2e71),
	.w2(32'h3b019b2e),
	.w3(32'hbc27894e),
	.w4(32'hbc0ab51c),
	.w5(32'h3b993414),
	.w6(32'hbb9dee92),
	.w7(32'hbb8d36ed),
	.w8(32'h3bb58895),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bab98),
	.w1(32'h3aa7f495),
	.w2(32'h3a9aee8c),
	.w3(32'hbb31fa3d),
	.w4(32'h3b33ea4b),
	.w5(32'h3a8bc8c2),
	.w6(32'h389a620a),
	.w7(32'h3afab2da),
	.w8(32'h3b2aca98),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf44b6a),
	.w1(32'h3c43f6aa),
	.w2(32'hbb051cd0),
	.w3(32'hba8619c4),
	.w4(32'hba101330),
	.w5(32'h3b252902),
	.w6(32'h3ba5850a),
	.w7(32'hbae0b4a7),
	.w8(32'h3b27dc50),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc9582),
	.w1(32'hbb0fdde4),
	.w2(32'h3c1eafba),
	.w3(32'h3b767cd3),
	.w4(32'hb90a9c41),
	.w5(32'h3c02ba0e),
	.w6(32'hbba2f794),
	.w7(32'h3c2fa293),
	.w8(32'h3bb4a694),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f1be6),
	.w1(32'h3bf91592),
	.w2(32'hbc11b30e),
	.w3(32'hbae36aae),
	.w4(32'hbc3f22ce),
	.w5(32'hbbc27016),
	.w6(32'hba48b278),
	.w7(32'hbb1dd471),
	.w8(32'hbc1cfe39),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6e049),
	.w1(32'h3bd6c925),
	.w2(32'h3c194bb0),
	.w3(32'h3b1bbcf4),
	.w4(32'h3bb715bd),
	.w5(32'h3c08dd8b),
	.w6(32'hbbc072e3),
	.w7(32'h39d3afcc),
	.w8(32'h3a076ce9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b003c5d),
	.w1(32'h3aac2bbb),
	.w2(32'hbc416d27),
	.w3(32'h3bb1bd17),
	.w4(32'hbad2adf2),
	.w5(32'hbb7cdfa8),
	.w6(32'h3b71954d),
	.w7(32'h3b80dfb7),
	.w8(32'hbb27e8d9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865a11),
	.w1(32'hbb9aab3c),
	.w2(32'hbaa4510a),
	.w3(32'hbc4da547),
	.w4(32'hbc93ff92),
	.w5(32'hbbfe64ab),
	.w6(32'hbbc4b302),
	.w7(32'hbc6c355e),
	.w8(32'hbbac05b8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09bc60),
	.w1(32'h3c6b86ad),
	.w2(32'h3aa6f6d5),
	.w3(32'h3b55113b),
	.w4(32'h3b650520),
	.w5(32'hbbe9a88a),
	.w6(32'h3bc29caf),
	.w7(32'h3ac521bd),
	.w8(32'h3abc51f8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe500),
	.w1(32'h3aa4a0b1),
	.w2(32'hb90b7341),
	.w3(32'hbadb0bdb),
	.w4(32'hbbf1edd4),
	.w5(32'hbaea2b56),
	.w6(32'hbb208199),
	.w7(32'hba2a3b9b),
	.w8(32'hbb5224c2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35351),
	.w1(32'h3bb0604f),
	.w2(32'h3bf9714f),
	.w3(32'h3b6ce398),
	.w4(32'h3b8f6df3),
	.w5(32'h3b81f17d),
	.w6(32'h3b635a08),
	.w7(32'h3b5bab46),
	.w8(32'h3b8cd013),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb650f5),
	.w1(32'hba3dc281),
	.w2(32'h3b8e4935),
	.w3(32'h3ba57f94),
	.w4(32'h3b310cf2),
	.w5(32'hbb07c7d8),
	.w6(32'h3a722e1f),
	.w7(32'hb909ce74),
	.w8(32'hbb15dd34),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b964463),
	.w1(32'h3bc6e36c),
	.w2(32'h3c489cf4),
	.w3(32'hba84cef1),
	.w4(32'h3aafcb41),
	.w5(32'h3b9312d7),
	.w6(32'hba2db2c5),
	.w7(32'hb7d4d94c),
	.w8(32'h3b8436b4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b106d58),
	.w1(32'h3b830915),
	.w2(32'h3bfcecd6),
	.w3(32'hba894898),
	.w4(32'hbb92667b),
	.w5(32'h3ad0970c),
	.w6(32'h3a92e491),
	.w7(32'h3b437ea0),
	.w8(32'hbb4769da),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe7d9),
	.w1(32'h3a2c195d),
	.w2(32'hbbf8bf2a),
	.w3(32'hbb867702),
	.w4(32'hbc4c01a7),
	.w5(32'hbb83357e),
	.w6(32'hbc076d6b),
	.w7(32'hbb26d66e),
	.w8(32'hbbd0b92f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849220),
	.w1(32'hba89a280),
	.w2(32'hbb5c0121),
	.w3(32'h3ab0b935),
	.w4(32'h3ba92353),
	.w5(32'hbb48f000),
	.w6(32'hbb53d92e),
	.w7(32'hb9c427ad),
	.w8(32'h399a3362),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5a963),
	.w1(32'hba91eead),
	.w2(32'h3c070fbc),
	.w3(32'hbb5cf408),
	.w4(32'hbb7af349),
	.w5(32'h3ae40b2a),
	.w6(32'h3a210a0f),
	.w7(32'hbb54012f),
	.w8(32'h3b00b05c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba775f7),
	.w1(32'hbbafa8f4),
	.w2(32'hbc3a0f54),
	.w3(32'hbaf0817c),
	.w4(32'hbc0586a5),
	.w5(32'hbab50807),
	.w6(32'hbbadcd06),
	.w7(32'h3b662638),
	.w8(32'h390aa041),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb263483),
	.w1(32'h3b71f3e5),
	.w2(32'hbaa2614c),
	.w3(32'h3a8a928b),
	.w4(32'hbae625da),
	.w5(32'hba646510),
	.w6(32'hbb7ca085),
	.w7(32'hbaedbc8d),
	.w8(32'h39b88c7c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba352484),
	.w1(32'hb9dec3f9),
	.w2(32'h3c0f106a),
	.w3(32'hbad88996),
	.w4(32'hbb41d98a),
	.w5(32'h3b4d6f9c),
	.w6(32'hb979fd88),
	.w7(32'hbb282fa6),
	.w8(32'h3b4a2e0e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6be00),
	.w1(32'h392c7053),
	.w2(32'h3b744e60),
	.w3(32'h3a29aa72),
	.w4(32'hbbbe0708),
	.w5(32'h3bbc5394),
	.w6(32'hbb6aef74),
	.w7(32'h3b04a60f),
	.w8(32'h3b69f60f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa629d5),
	.w1(32'hbb1928cd),
	.w2(32'h39184ff7),
	.w3(32'h3bdf1655),
	.w4(32'hbab5695f),
	.w5(32'h3ad138cf),
	.w6(32'h3bad7563),
	.w7(32'h3c1962a4),
	.w8(32'h3bcbf9a2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99281f),
	.w1(32'h3a788180),
	.w2(32'hbb2df7c4),
	.w3(32'hbc726d88),
	.w4(32'h3ab0ecca),
	.w5(32'hbac56563),
	.w6(32'h3b4da09c),
	.w7(32'h3b59b2c9),
	.w8(32'h3b8e920f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7369),
	.w1(32'h3c2317f8),
	.w2(32'hbbcf06e8),
	.w3(32'hbbf1ccac),
	.w4(32'h3c0d59be),
	.w5(32'h3b9110ef),
	.w6(32'hbc182e7f),
	.w7(32'hbc0ac488),
	.w8(32'h3c2c3586),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1f2d),
	.w1(32'h3cc37216),
	.w2(32'hbc0249f8),
	.w3(32'hbc111241),
	.w4(32'h3caf14e4),
	.w5(32'h3bf08588),
	.w6(32'hbb8a53ce),
	.w7(32'hba0e6341),
	.w8(32'h3b7fe91f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a903f),
	.w1(32'hbb5be6da),
	.w2(32'hbb45c658),
	.w3(32'h3be43b57),
	.w4(32'h3bb7a3e2),
	.w5(32'h3b4d7f0f),
	.w6(32'h3b254d4e),
	.w7(32'hba2949d5),
	.w8(32'h3b6b8a5d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e24e1),
	.w1(32'h3b3c9054),
	.w2(32'h3a885906),
	.w3(32'h3bb3ba9e),
	.w4(32'hbb9ea016),
	.w5(32'h3bc10d7e),
	.w6(32'h3b137c0f),
	.w7(32'hbb7bc5ee),
	.w8(32'h3ae558a6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c31f5),
	.w1(32'hb9f9b217),
	.w2(32'hbc4c8ad8),
	.w3(32'hbb8fd0bc),
	.w4(32'h3bdc0c24),
	.w5(32'hbba53a59),
	.w6(32'h3c88a820),
	.w7(32'h3c8f686c),
	.w8(32'h3b0b93a0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5b21),
	.w1(32'h3bd31776),
	.w2(32'hbc53f124),
	.w3(32'hbb698b73),
	.w4(32'h3b1610d1),
	.w5(32'hbbf1b37e),
	.w6(32'hbc0465b4),
	.w7(32'h3a5cc65e),
	.w8(32'hbb9ef8f8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3997b9),
	.w1(32'h3bedfc0e),
	.w2(32'h3caff6d8),
	.w3(32'hbb433929),
	.w4(32'h3b3c7a06),
	.w5(32'h3b7060dc),
	.w6(32'hb92b7179),
	.w7(32'h3abd2807),
	.w8(32'h3bdf48dc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092603),
	.w1(32'hb7c76d06),
	.w2(32'hbbe881c6),
	.w3(32'hbb490e85),
	.w4(32'hbb31e10a),
	.w5(32'hbb0a89e4),
	.w6(32'h3b0c0534),
	.w7(32'h3b92278a),
	.w8(32'h3b946d2e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3dab4),
	.w1(32'h3bc58f68),
	.w2(32'hbb8129d6),
	.w3(32'hbbb26c43),
	.w4(32'hba9c6cc5),
	.w5(32'hbb8b90f6),
	.w6(32'hbb2cc8cd),
	.w7(32'hbbeac681),
	.w8(32'h39b270c8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaaf61),
	.w1(32'h3b21b38c),
	.w2(32'h3c651d7f),
	.w3(32'hbb965d27),
	.w4(32'hbac4c59a),
	.w5(32'h39fa3c0a),
	.w6(32'hbb62dac7),
	.w7(32'hbbb6011f),
	.w8(32'h3a9883e9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf967ed),
	.w1(32'h3a98d993),
	.w2(32'h3a150bc1),
	.w3(32'h3b809bbc),
	.w4(32'h39c57dca),
	.w5(32'hbae75d75),
	.w6(32'h3b461272),
	.w7(32'h3b94bb4e),
	.w8(32'hbbb94c6a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53eb69),
	.w1(32'h3ada7645),
	.w2(32'h3ba360d3),
	.w3(32'h3b01de92),
	.w4(32'h3bc35628),
	.w5(32'h3b5cbb1f),
	.w6(32'h3908e037),
	.w7(32'hbb7cc652),
	.w8(32'h3b863967),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009bc5),
	.w1(32'hbb288b42),
	.w2(32'hbb027bb7),
	.w3(32'h3ad7291f),
	.w4(32'hbb979470),
	.w5(32'hbb324fc6),
	.w6(32'h3ae6b521),
	.w7(32'hbb158afd),
	.w8(32'hbc0eeede),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c16e),
	.w1(32'hbbf3802c),
	.w2(32'hbc30d402),
	.w3(32'hbb89f1b1),
	.w4(32'hbc18546a),
	.w5(32'hba118c3e),
	.w6(32'hbb653ce4),
	.w7(32'hbb726ce7),
	.w8(32'hbb18c644),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb67c7),
	.w1(32'h3acd311b),
	.w2(32'h3aa5e2ec),
	.w3(32'hbb4515d1),
	.w4(32'hbbbb710b),
	.w5(32'hbaaa34a2),
	.w6(32'hbb35aabe),
	.w7(32'h3c47dabd),
	.w8(32'h3abaee53),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad3b1a),
	.w1(32'h3c23772d),
	.w2(32'h3b27eef8),
	.w3(32'hba96a10c),
	.w4(32'h3bdcafbe),
	.w5(32'hb9a0bb51),
	.w6(32'hbaef635c),
	.w7(32'h39b376dd),
	.w8(32'h37f471c2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7468c3),
	.w1(32'h3b73a965),
	.w2(32'hba83df32),
	.w3(32'h3b1bf0ce),
	.w4(32'h3b7edac1),
	.w5(32'hba93e5c3),
	.w6(32'h3a86c512),
	.w7(32'h3b5457fb),
	.w8(32'hbb9fe6e9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191d83),
	.w1(32'hbb475aa8),
	.w2(32'hbb049e7a),
	.w3(32'h3ab25577),
	.w4(32'hb981b8e6),
	.w5(32'h3b57c214),
	.w6(32'hbbf6533f),
	.w7(32'hbb4a0ed3),
	.w8(32'hbbb4ed13),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f236d),
	.w1(32'hbc0628f8),
	.w2(32'hbbcde651),
	.w3(32'hbb8a8573),
	.w4(32'hbba7a9c5),
	.w5(32'hbb752194),
	.w6(32'hbb5636fe),
	.w7(32'hbb7e9fe5),
	.w8(32'hb99f03c4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9190458),
	.w1(32'h3b71c8a0),
	.w2(32'hbb35aa77),
	.w3(32'h3b7ddc73),
	.w4(32'hbbd08283),
	.w5(32'h3aa7df76),
	.w6(32'hba6888bb),
	.w7(32'hbbc3430d),
	.w8(32'hbb44a798),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e1ae4),
	.w1(32'hba320b68),
	.w2(32'hbaa988ff),
	.w3(32'hba9a0ff2),
	.w4(32'h3923d263),
	.w5(32'hbb8ea95c),
	.w6(32'hbb08e857),
	.w7(32'h3acf80a9),
	.w8(32'hbbf16451),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc526ae),
	.w1(32'h3c05cd70),
	.w2(32'h3bbc0624),
	.w3(32'h3b1510ae),
	.w4(32'h3b665974),
	.w5(32'h3be164fd),
	.w6(32'h3c18f0c4),
	.w7(32'h3beaaf0e),
	.w8(32'h3bba2011),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8fae0),
	.w1(32'h3bad2663),
	.w2(32'hbba0df3a),
	.w3(32'hbb2e3498),
	.w4(32'hbbc8b27b),
	.w5(32'hbb48ae42),
	.w6(32'hbacccdc9),
	.w7(32'hbb008ad8),
	.w8(32'hbaabb3a8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53aa6),
	.w1(32'hba7c5b9d),
	.w2(32'h3c6a077a),
	.w3(32'hbc0946e6),
	.w4(32'hbb36a748),
	.w5(32'h3bbc7fae),
	.w6(32'hba873e8e),
	.w7(32'hbb89dd53),
	.w8(32'hbb31cfa2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa1261),
	.w1(32'h3b116631),
	.w2(32'hbc62f5c7),
	.w3(32'hbabc9a46),
	.w4(32'hbb831945),
	.w5(32'h3b310225),
	.w6(32'hbb96673d),
	.w7(32'hbb35a6df),
	.w8(32'h3c2df690),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d09b4),
	.w1(32'h3b738ae0),
	.w2(32'h3bb9d1a1),
	.w3(32'hbb8989b1),
	.w4(32'hbc6ad11d),
	.w5(32'h3c0dc518),
	.w6(32'hbb82b4a0),
	.w7(32'h3a5cddaf),
	.w8(32'h3a0f021a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407fc0),
	.w1(32'h3a1d6b42),
	.w2(32'hbb0c67f0),
	.w3(32'h3930715a),
	.w4(32'hbc09cdb0),
	.w5(32'hbb061f99),
	.w6(32'h3b58c263),
	.w7(32'h3b9496b9),
	.w8(32'hbb73c621),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797d14),
	.w1(32'h3abd46b9),
	.w2(32'h3b52fd5d),
	.w3(32'hbb1c60b9),
	.w4(32'hbae3e8b1),
	.w5(32'h3acf1d47),
	.w6(32'hba85bdcb),
	.w7(32'hba85a2af),
	.w8(32'h3b2e807d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c579dcb),
	.w1(32'hbb2b3793),
	.w2(32'hbb6c8399),
	.w3(32'h3ad5fd1f),
	.w4(32'hbc51bc39),
	.w5(32'hbc99fcf3),
	.w6(32'h3b87cc6d),
	.w7(32'h3a37b7f9),
	.w8(32'h3ca346af),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fb0e2),
	.w1(32'h3c458218),
	.w2(32'hbc0c05b3),
	.w3(32'hbc3b7eb7),
	.w4(32'h3cb96121),
	.w5(32'hbb8248ca),
	.w6(32'h3bfa0390),
	.w7(32'hbc789b9f),
	.w8(32'hbc083655),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88dbe9),
	.w1(32'h3a4e00c2),
	.w2(32'hb994df62),
	.w3(32'h3ab544ff),
	.w4(32'h3b6f25a6),
	.w5(32'hbc2d045a),
	.w6(32'hbaaa8a05),
	.w7(32'hb9aadd73),
	.w8(32'hbbbcc34a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc361f01),
	.w1(32'hbb1df623),
	.w2(32'hbbe3c437),
	.w3(32'hbc5d96ef),
	.w4(32'hbc230faa),
	.w5(32'h3c3297cd),
	.w6(32'h3a39b46d),
	.w7(32'h3c1d552e),
	.w8(32'hbb7b3709),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c86f7),
	.w1(32'hbc2ff07f),
	.w2(32'h3a1073f0),
	.w3(32'h3c2c0f86),
	.w4(32'hbc04b64d),
	.w5(32'h3a3e05df),
	.w6(32'h3d188947),
	.w7(32'h3d030d51),
	.w8(32'hba17ea16),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565420),
	.w1(32'hbb853271),
	.w2(32'h3ac70763),
	.w3(32'h3a7f5586),
	.w4(32'hbb2dbdb4),
	.w5(32'hbc07c2ca),
	.w6(32'h3aeec556),
	.w7(32'h38ebe1fa),
	.w8(32'hbc8f4e5e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519e12),
	.w1(32'hbb21ea80),
	.w2(32'hbb4ea391),
	.w3(32'h3c8fd3f2),
	.w4(32'h3c442864),
	.w5(32'hbb5823c2),
	.w6(32'hbc4351a6),
	.w7(32'hbb74521b),
	.w8(32'hbb58b435),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60702a),
	.w1(32'hbb06ebda),
	.w2(32'h3c32085c),
	.w3(32'hbada50b1),
	.w4(32'hbb05285d),
	.w5(32'hbbe09ed1),
	.w6(32'hbae12668),
	.w7(32'hbad7d474),
	.w8(32'hbc055094),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fef61),
	.w1(32'hbc21ab84),
	.w2(32'hbaaa5550),
	.w3(32'hbc1f80e1),
	.w4(32'hbbdf3694),
	.w5(32'h3bd5f12a),
	.w6(32'hbcb759a3),
	.w7(32'hbc679076),
	.w8(32'h3c2e9620),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9612be3),
	.w1(32'hbaa50206),
	.w2(32'hbbe06356),
	.w3(32'h39e3e9de),
	.w4(32'hbb543b11),
	.w5(32'hbc1357fb),
	.w6(32'h3c0c0577),
	.w7(32'h3b85e519),
	.w8(32'h3c8a8f6d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48f861),
	.w1(32'h3c657c12),
	.w2(32'h3b416e0e),
	.w3(32'hbcc50f5d),
	.w4(32'hbb996318),
	.w5(32'h3b99c34c),
	.w6(32'h3c833349),
	.w7(32'hbb11622e),
	.w8(32'hbc74ed8d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f75c8),
	.w1(32'h3a6de46d),
	.w2(32'h3aa3a1f0),
	.w3(32'hbb096f05),
	.w4(32'h3bc7b737),
	.w5(32'h3a9c58a0),
	.w6(32'hbc028181),
	.w7(32'h3a2fc7a7),
	.w8(32'hbb8f4441),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cb607),
	.w1(32'hbc113f51),
	.w2(32'h3bd5c9b5),
	.w3(32'h3c3c45e4),
	.w4(32'h3c0523b7),
	.w5(32'hbb9ec9cc),
	.w6(32'hbbaae644),
	.w7(32'h3b606330),
	.w8(32'h3abd905a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc053b86),
	.w1(32'hbc01e3d6),
	.w2(32'h392d4756),
	.w3(32'hbc470277),
	.w4(32'hbbc5b4fc),
	.w5(32'h3b2b3606),
	.w6(32'h3c2ba2c7),
	.w7(32'h3b495a69),
	.w8(32'h3bd195a2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f0a56),
	.w1(32'hbbc5d873),
	.w2(32'hbb8123b9),
	.w3(32'h3c6aa8b7),
	.w4(32'h3b1be3ce),
	.w5(32'hbb621b6c),
	.w6(32'hbbf13259),
	.w7(32'hbba3dca6),
	.w8(32'h3af5b0f8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93440b),
	.w1(32'h3895cd61),
	.w2(32'hbbbbc76f),
	.w3(32'hbbbf5dba),
	.w4(32'hbb65ad9d),
	.w5(32'hbb84119c),
	.w6(32'hbaa5e725),
	.w7(32'h3afa0e2f),
	.w8(32'h3bcb70c5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f28e62),
	.w1(32'hbba2bce9),
	.w2(32'h3ac7e66e),
	.w3(32'h3af955cc),
	.w4(32'h3bd8ad5a),
	.w5(32'hbc3d4fd8),
	.w6(32'hbc11f9a9),
	.w7(32'hbc437983),
	.w8(32'h3b0702c1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3469d1),
	.w1(32'hbc52bec9),
	.w2(32'h3b6ab217),
	.w3(32'hbbf7f985),
	.w4(32'hbc03d6d8),
	.w5(32'hbb7e757b),
	.w6(32'h3a773831),
	.w7(32'hbb31ab08),
	.w8(32'hbb9d1123),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba628e),
	.w1(32'h3b796a4a),
	.w2(32'h3c047a41),
	.w3(32'h3bd8ca23),
	.w4(32'h3c5d851c),
	.w5(32'h3c111199),
	.w6(32'hbc039c63),
	.w7(32'hbc53ac11),
	.w8(32'h3c578dcb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8ebf4),
	.w1(32'hbaaeae46),
	.w2(32'h38cd2b53),
	.w3(32'hba961005),
	.w4(32'h3cb029d5),
	.w5(32'hbb98af60),
	.w6(32'hbc7bdbf5),
	.w7(32'hbca373e3),
	.w8(32'hbb188ca7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed2096),
	.w1(32'h37e08f64),
	.w2(32'hbbaa9715),
	.w3(32'hbb509952),
	.w4(32'hbb823032),
	.w5(32'hbb8c93f5),
	.w6(32'hbba8e406),
	.w7(32'hbbc09d6b),
	.w8(32'h3adb83a2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64f04d),
	.w1(32'h3c0f0c2b),
	.w2(32'hbb8d9c5d),
	.w3(32'hbb91cc96),
	.w4(32'hbbe4a7c9),
	.w5(32'hbc478674),
	.w6(32'h3b6d979c),
	.w7(32'hb9937d87),
	.w8(32'hbbe1a626),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1c74),
	.w1(32'hbc176b8a),
	.w2(32'hbbdeeb23),
	.w3(32'h3c8090fc),
	.w4(32'h3c26d619),
	.w5(32'hbbcab257),
	.w6(32'hbb684998),
	.w7(32'h3b685e76),
	.w8(32'hbc3d3005),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e052),
	.w1(32'hbb7d3734),
	.w2(32'h3b2d2e15),
	.w3(32'h3c78aa70),
	.w4(32'h3c9ee020),
	.w5(32'hbb22cacb),
	.w6(32'hbc831a6c),
	.w7(32'hbbda0263),
	.w8(32'hbb696942),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c262d4f),
	.w1(32'h3b30055a),
	.w2(32'h3c1c0347),
	.w3(32'h3c1fc363),
	.w4(32'h3b768202),
	.w5(32'h3b97ac48),
	.w6(32'hbbc2b569),
	.w7(32'h3bc39947),
	.w8(32'h3b74368e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83c05f),
	.w1(32'hbc2316d1),
	.w2(32'h3ba9353c),
	.w3(32'h3b7039b7),
	.w4(32'h3bf8e57b),
	.w5(32'h3b8b1bba),
	.w6(32'hbbbbdd2b),
	.w7(32'h3b89b9d2),
	.w8(32'h3c84df0a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c314155),
	.w1(32'h3b590103),
	.w2(32'hbb5c3f93),
	.w3(32'hbbe347fc),
	.w4(32'h3c2f2a1e),
	.w5(32'h3b859203),
	.w6(32'h3c958ab6),
	.w7(32'hbb97d249),
	.w8(32'hbbd9d03a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66add7),
	.w1(32'hbc12bf62),
	.w2(32'h3a8f4d6d),
	.w3(32'h3bb74669),
	.w4(32'h3b7d2fcd),
	.w5(32'h3cbc5e22),
	.w6(32'h3bcc6bd7),
	.w7(32'h3cd83f5e),
	.w8(32'hbbf4e7fb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8aac60),
	.w1(32'hbca42be7),
	.w2(32'h3a680f27),
	.w3(32'h3beb322d),
	.w4(32'hbc711e32),
	.w5(32'hbaeac5e8),
	.w6(32'h3bdfb819),
	.w7(32'h3c0e886e),
	.w8(32'h3bef9aa3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9df17),
	.w1(32'hbc773f49),
	.w2(32'h3b2cc98a),
	.w3(32'h3b7db517),
	.w4(32'h3a6aae97),
	.w5(32'h39af02a3),
	.w6(32'h3b6dd5a8),
	.w7(32'h3ae87aba),
	.w8(32'hbbfaba8a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab53e10),
	.w1(32'h3b965ae3),
	.w2(32'h3b156612),
	.w3(32'h3abe7305),
	.w4(32'h3be9c149),
	.w5(32'h3c1c7c69),
	.w6(32'hbaccc139),
	.w7(32'h3bc11cdd),
	.w8(32'h3bf3f966),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4abb9a),
	.w1(32'h3c168823),
	.w2(32'h3cdb595f),
	.w3(32'h3ab6e930),
	.w4(32'h3c105bdc),
	.w5(32'h3b9912b4),
	.w6(32'h39dd87cb),
	.w7(32'hbb5ae410),
	.w8(32'h3c7288b3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7504a1),
	.w1(32'hba76d27e),
	.w2(32'hbc30807c),
	.w3(32'hbccf64c2),
	.w4(32'hbceb761b),
	.w5(32'hbc5ca84c),
	.w6(32'hbc415d76),
	.w7(32'hbc7828d3),
	.w8(32'hbaf6cb80),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f700),
	.w1(32'hbbbca5d0),
	.w2(32'hbad354ef),
	.w3(32'h3c1002bd),
	.w4(32'h3c07eaf4),
	.w5(32'h393d5a43),
	.w6(32'hbc5a8e5c),
	.w7(32'h3b3daac6),
	.w8(32'hba30ab7b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04d38d),
	.w1(32'hbb0f16d5),
	.w2(32'hbb2d02a5),
	.w3(32'hb9b8a8b8),
	.w4(32'hbb0b6cfe),
	.w5(32'hbb5d9dbe),
	.w6(32'h3b982180),
	.w7(32'h3a7c80d1),
	.w8(32'hbb1dc5e2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde1b5),
	.w1(32'hbb4fb406),
	.w2(32'h3b826940),
	.w3(32'hbc277e45),
	.w4(32'hbbc1c8aa),
	.w5(32'h3c0d5387),
	.w6(32'hbbe48df9),
	.w7(32'hbb83927d),
	.w8(32'hbc2a1e04),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c1cb1),
	.w1(32'h3c02bf1a),
	.w2(32'h37f199b5),
	.w3(32'h3b26962d),
	.w4(32'h3b939308),
	.w5(32'h3c159baa),
	.w6(32'hbc28456b),
	.w7(32'h3be57537),
	.w8(32'h3c009252),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373c7b),
	.w1(32'hbc2e4f38),
	.w2(32'hbb8c365b),
	.w3(32'hbb4aeb8e),
	.w4(32'hbbe57187),
	.w5(32'hbc006882),
	.w6(32'h3be42fab),
	.w7(32'h3b539875),
	.w8(32'hbaa490bc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b78f2),
	.w1(32'hbb4f5ce4),
	.w2(32'h3b73923a),
	.w3(32'hbc549ec7),
	.w4(32'hbc0bc563),
	.w5(32'hbc0aab53),
	.w6(32'hbaeb0d86),
	.w7(32'h39ed3fa2),
	.w8(32'h3ab1381d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ab729),
	.w1(32'h3b1cbb24),
	.w2(32'hbc37d95b),
	.w3(32'hbbc99a4e),
	.w4(32'h3b372e58),
	.w5(32'hbbc49827),
	.w6(32'hbc91a289),
	.w7(32'h3a2c6e72),
	.w8(32'hbc132d10),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5c2c6),
	.w1(32'hbb8b0be9),
	.w2(32'hbb47603b),
	.w3(32'h3b1f49b4),
	.w4(32'h396098e8),
	.w5(32'hbbbebb48),
	.w6(32'hbba04571),
	.w7(32'h3b64b807),
	.w8(32'hbaea54f3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa9f1),
	.w1(32'hbb05cd11),
	.w2(32'h3c65a6b7),
	.w3(32'hbc25e93b),
	.w4(32'hbc2782eb),
	.w5(32'h3c742ba0),
	.w6(32'hbbc4abf8),
	.w7(32'hbbee9d59),
	.w8(32'h3b7c0759),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239581),
	.w1(32'h3b8df2e2),
	.w2(32'hbb4a25d9),
	.w3(32'h3b6028cb),
	.w4(32'h3b883bba),
	.w5(32'h3b3292f7),
	.w6(32'hbb49e9d0),
	.w7(32'hb9e3be43),
	.w8(32'hbc204c63),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe752b),
	.w1(32'hbbcf0f20),
	.w2(32'h3bb9d1d8),
	.w3(32'h3baf5da0),
	.w4(32'h3a66133f),
	.w5(32'h3acc9a15),
	.w6(32'hbb1f6b73),
	.w7(32'h3910562b),
	.w8(32'hbbb2f60a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42e436),
	.w1(32'hbb14bcd9),
	.w2(32'hb998bd3b),
	.w3(32'h3c76b4a4),
	.w4(32'h3c8b7314),
	.w5(32'hbc03586a),
	.w6(32'hbc3baf08),
	.w7(32'hbc175f27),
	.w8(32'hb973f015),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc270f2d),
	.w1(32'hbbd1e15d),
	.w2(32'h3a9c89ca),
	.w3(32'hbad9f148),
	.w4(32'h3b86f23b),
	.w5(32'hbb3e2dc1),
	.w6(32'h3b7ebecb),
	.w7(32'h3b9e86a0),
	.w8(32'hbb8c3a74),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18f5fd),
	.w1(32'hbab35c38),
	.w2(32'hbb925740),
	.w3(32'hba88124d),
	.w4(32'hbb22e91d),
	.w5(32'hbbbde8c4),
	.w6(32'hbb8f2db7),
	.w7(32'hbb826638),
	.w8(32'hbba4ed48),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff6486),
	.w1(32'hbc19a21c),
	.w2(32'hbab34ed3),
	.w3(32'hba8d2c0f),
	.w4(32'hbc4279e5),
	.w5(32'h3a54605e),
	.w6(32'hbbd65c9c),
	.w7(32'hbbbef396),
	.w8(32'hbba2c0e9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5642c9),
	.w1(32'h3c245d6f),
	.w2(32'hbacc86d7),
	.w3(32'h3c1c63d4),
	.w4(32'h3a64011f),
	.w5(32'hbb35400c),
	.w6(32'hbc6be374),
	.w7(32'hbbe2447d),
	.w8(32'hbbde51d0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26ad3a),
	.w1(32'h3a36cb59),
	.w2(32'h3be14c5f),
	.w3(32'h3c849f7f),
	.w4(32'h3c373295),
	.w5(32'h3b9771f2),
	.w6(32'hbc56e47e),
	.w7(32'hb99422ec),
	.w8(32'h3c86ba06),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990b11),
	.w1(32'hbc57255d),
	.w2(32'hbbea46a4),
	.w3(32'h3bdb056b),
	.w4(32'h382f2dbe),
	.w5(32'hbbbc0ac0),
	.w6(32'hbb8fc086),
	.w7(32'h3c328dd2),
	.w8(32'hba9fcdd0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b6b56),
	.w1(32'h3b426082),
	.w2(32'hbb1c599a),
	.w3(32'hbba48c8f),
	.w4(32'h3af09b8a),
	.w5(32'hbaeb34a6),
	.w6(32'hbb13bd67),
	.w7(32'h3b106784),
	.w8(32'hb88b6f80),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaca65),
	.w1(32'h3b94b8c2),
	.w2(32'hbb090d88),
	.w3(32'hbc434a7b),
	.w4(32'h3b85a26a),
	.w5(32'h3b3c1b40),
	.w6(32'hbc7e5fed),
	.w7(32'hbc06c73b),
	.w8(32'h3b563df2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b65bf),
	.w1(32'h399aafaf),
	.w2(32'h3b9d4711),
	.w3(32'hbb43c536),
	.w4(32'h3ac6d6e0),
	.w5(32'hb94b6d06),
	.w6(32'h3b00dd74),
	.w7(32'h3bc5fab4),
	.w8(32'hbc8b9113),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c3172),
	.w1(32'hbb5c10f1),
	.w2(32'hbc044ad8),
	.w3(32'h3b7e6bc0),
	.w4(32'hbbbcaa0f),
	.w5(32'hbc1881ab),
	.w6(32'hbc65ef9a),
	.w7(32'hbc0edeb8),
	.w8(32'h3c0a55a6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2b84e),
	.w1(32'h3c01a151),
	.w2(32'hbadc14e3),
	.w3(32'hbcd6c9cf),
	.w4(32'hbc63e2e5),
	.w5(32'h3bf45cb3),
	.w6(32'hbc7c0ec7),
	.w7(32'hbcab8056),
	.w8(32'hbb75397c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4f5d7),
	.w1(32'hba82f371),
	.w2(32'h3cbd9c0d),
	.w3(32'h3c15f1ff),
	.w4(32'h3c3a267b),
	.w5(32'h3c31e1d4),
	.w6(32'h3baa15c4),
	.w7(32'h3b6dca0c),
	.w8(32'hbcd27960),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3019f),
	.w1(32'hbc4c89cf),
	.w2(32'hbb9d07e2),
	.w3(32'h3cf9f780),
	.w4(32'hbb7a718d),
	.w5(32'h3a0e1d4b),
	.w6(32'hbc6266f1),
	.w7(32'h3a6dc572),
	.w8(32'hb996c8e5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47eac6),
	.w1(32'hbc173885),
	.w2(32'h3b8871d1),
	.w3(32'hbbad4831),
	.w4(32'hbb892df9),
	.w5(32'hbc0c8f0e),
	.w6(32'hbab4515e),
	.w7(32'hb8bd1cf1),
	.w8(32'hb9e62306),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad00146),
	.w1(32'hbb26ef72),
	.w2(32'h3aeb6c9e),
	.w3(32'h399ef4d2),
	.w4(32'h3b662e67),
	.w5(32'hbbb32130),
	.w6(32'hbb526824),
	.w7(32'h3b0ab8de),
	.w8(32'hbbe9401a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac716a1),
	.w1(32'hbb51114e),
	.w2(32'hbbc0097e),
	.w3(32'h3c0a5fae),
	.w4(32'h3ad4cb9d),
	.w5(32'hb8e83b21),
	.w6(32'hbc3b042a),
	.w7(32'h3c08cf05),
	.w8(32'h39e59702),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc59ce),
	.w1(32'hbca75b6f),
	.w2(32'h3c0b1166),
	.w3(32'h3c207e1d),
	.w4(32'hbba32cd0),
	.w5(32'h3c8c0c1a),
	.w6(32'hbb4dfd5a),
	.w7(32'hb99ff902),
	.w8(32'h3b2c6b61),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f6a0e),
	.w1(32'h3b8ab341),
	.w2(32'h3c8c42db),
	.w3(32'h3c66cedc),
	.w4(32'h3b790fa1),
	.w5(32'h3ca7ab88),
	.w6(32'h3cbdc4cc),
	.w7(32'h3cccb6a7),
	.w8(32'h3cb80ad4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf136e1),
	.w1(32'hba20a0ab),
	.w2(32'h3c97d06f),
	.w3(32'hbbdc8d39),
	.w4(32'h393c0800),
	.w5(32'h3c1b44fc),
	.w6(32'h3c890c27),
	.w7(32'h3c3ea5f3),
	.w8(32'h3b394f7b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071ec1),
	.w1(32'hbb4e43ae),
	.w2(32'h3b1c4a3e),
	.w3(32'h3c2df2fd),
	.w4(32'h395abc29),
	.w5(32'hbad22d09),
	.w6(32'h3b3fcec5),
	.w7(32'h3b8b439c),
	.w8(32'hba92a4e4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11a290),
	.w1(32'h3b1faa8c),
	.w2(32'hbb8b6da8),
	.w3(32'h3b6b0239),
	.w4(32'hb9d27428),
	.w5(32'hbb81c712),
	.w6(32'hbaba7be6),
	.w7(32'h3b96081f),
	.w8(32'h3b2ade4a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5838ec),
	.w1(32'hbba87dd6),
	.w2(32'h3bf05601),
	.w3(32'h3ae8bb5e),
	.w4(32'h3abb6da0),
	.w5(32'h3cacadbb),
	.w6(32'hbb13d043),
	.w7(32'h3b898adf),
	.w8(32'hbcbf2b67),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee2c40),
	.w1(32'hbb514c2c),
	.w2(32'hbc0c5e6d),
	.w3(32'h3d5ae706),
	.w4(32'h3d0c4473),
	.w5(32'hba25bd5f),
	.w6(32'hba25262e),
	.w7(32'h3d1ed06a),
	.w8(32'h3c6390f6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c7ff),
	.w1(32'hbb9e8828),
	.w2(32'hbba86f3f),
	.w3(32'h3ba7e9fb),
	.w4(32'h3c0ca92d),
	.w5(32'h3b049535),
	.w6(32'hbb4a98c8),
	.w7(32'hbb2375cf),
	.w8(32'h3a4bf01f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3054f),
	.w1(32'hbbe9deb9),
	.w2(32'hbbb1b77d),
	.w3(32'h3cd72a71),
	.w4(32'hbbcec113),
	.w5(32'hbbfa1ef2),
	.w6(32'hbbc029cc),
	.w7(32'hb984ad40),
	.w8(32'hbc331b73),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc583f83),
	.w1(32'hbc3da682),
	.w2(32'h3c00cc81),
	.w3(32'hbc0dc448),
	.w4(32'hbb4afc37),
	.w5(32'hbb0d00b9),
	.w6(32'hbcc99983),
	.w7(32'hbc47fa86),
	.w8(32'h3c1e0fca),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7305c),
	.w1(32'h3c7c687f),
	.w2(32'h3c2fc723),
	.w3(32'hbca4998e),
	.w4(32'h3ade76ef),
	.w5(32'hbb96e0b9),
	.w6(32'hbc755d89),
	.w7(32'hbc1d67cf),
	.w8(32'h3ae33060),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9efc4),
	.w1(32'hba263ec8),
	.w2(32'h3c2c5746),
	.w3(32'h3bd7bebe),
	.w4(32'h3c2c8e36),
	.w5(32'hbba635fa),
	.w6(32'hbc96fb8a),
	.w7(32'hbc232daf),
	.w8(32'hbc3003c4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2839fd),
	.w1(32'hba9e8fb1),
	.w2(32'hba047125),
	.w3(32'h3ca47fff),
	.w4(32'h3c9d56ed),
	.w5(32'hbb1a60a8),
	.w6(32'hbc6a3e13),
	.w7(32'hbb1804bd),
	.w8(32'h3bb5da63),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5bbf),
	.w1(32'hbb1b4632),
	.w2(32'h3c794118),
	.w3(32'hbb950dbc),
	.w4(32'h3b22ce19),
	.w5(32'h3b89a044),
	.w6(32'hbad793b9),
	.w7(32'hbbbfcc24),
	.w8(32'hbaa3f69e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2915ae),
	.w1(32'hbbf346a6),
	.w2(32'h3c9d5742),
	.w3(32'h3b77249a),
	.w4(32'h3c55adcd),
	.w5(32'h3bc7afa3),
	.w6(32'h3b8cffd9),
	.w7(32'h3c710f79),
	.w8(32'hbbfab1d4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dc972),
	.w1(32'hbbbe3a11),
	.w2(32'h3b7a4620),
	.w3(32'h3b7b77ca),
	.w4(32'h3a4db8e5),
	.w5(32'h3b360c39),
	.w6(32'hbbf3a7b9),
	.w7(32'h39fe18f5),
	.w8(32'hbb45251e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002760),
	.w1(32'hba9d8577),
	.w2(32'h3c540ac3),
	.w3(32'h3ba2d289),
	.w4(32'h3c15490f),
	.w5(32'h3c8be2be),
	.w6(32'hbba41dad),
	.w7(32'h3a8bcf1c),
	.w8(32'h3bbbde66),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de3b9),
	.w1(32'hbbab2c69),
	.w2(32'hbbde75fd),
	.w3(32'h3c4d9b9a),
	.w4(32'h3bedb72f),
	.w5(32'hbc03c5f9),
	.w6(32'h3be3b839),
	.w7(32'h3bc89821),
	.w8(32'h3c0404e9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664958),
	.w1(32'h3c033783),
	.w2(32'hbbb84065),
	.w3(32'hbc7af5e3),
	.w4(32'hbb510c42),
	.w5(32'hba041837),
	.w6(32'hbc11c5fd),
	.w7(32'hbc6c94d1),
	.w8(32'hba4de28a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64621),
	.w1(32'h398d0fc3),
	.w2(32'hb9f2690a),
	.w3(32'h3af5e01c),
	.w4(32'hb9844b40),
	.w5(32'hb851daa4),
	.w6(32'hbc0b30be),
	.w7(32'hbbc1f9ea),
	.w8(32'hbb6dffe7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2355fb),
	.w1(32'hbc0f78fe),
	.w2(32'h3ba4e910),
	.w3(32'hb911b09c),
	.w4(32'hbb6a6ec7),
	.w5(32'hbb097d48),
	.w6(32'hbc148935),
	.w7(32'hbba44175),
	.w8(32'h3b9bdc5f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102369),
	.w1(32'h3b15f721),
	.w2(32'h3bc15580),
	.w3(32'hb954bf12),
	.w4(32'hbb9edac5),
	.w5(32'hbb61cda5),
	.w6(32'hbb437840),
	.w7(32'hbb9843bb),
	.w8(32'hbc4a9c7c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c35253),
	.w1(32'hbbcb90d1),
	.w2(32'hbc26f583),
	.w3(32'h3b87c06c),
	.w4(32'hbbef5f72),
	.w5(32'hbafd1aef),
	.w6(32'hbc4b552c),
	.w7(32'hbb17014d),
	.w8(32'h3c2967a2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2300b7),
	.w1(32'h3a8d3862),
	.w2(32'h38f4e773),
	.w3(32'hbba98d36),
	.w4(32'h3c4c10f9),
	.w5(32'hbb5a6267),
	.w6(32'hbc1fc8c8),
	.w7(32'hbbc7da62),
	.w8(32'hbc260593),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9015a),
	.w1(32'h394d0a28),
	.w2(32'hba4a3695),
	.w3(32'h3c2cd9cd),
	.w4(32'h3c209484),
	.w5(32'h3bc2d926),
	.w6(32'hbc1f2b6a),
	.w7(32'hbbc2e496),
	.w8(32'hbba77044),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba694258),
	.w1(32'hbb64535c),
	.w2(32'hbac572e1),
	.w3(32'h3b5d3cca),
	.w4(32'hbb90fcd1),
	.w5(32'hbbe70d7f),
	.w6(32'hbbe3ab6b),
	.w7(32'hbbdd956e),
	.w8(32'h3b5ed316),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a7157),
	.w1(32'h3c69c679),
	.w2(32'h3a334029),
	.w3(32'hbc7342c5),
	.w4(32'hbb5bcf33),
	.w5(32'hbb1cd5b7),
	.w6(32'hbc0ab36f),
	.w7(32'hbc1adcd7),
	.w8(32'hbbc88f0d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c25d2),
	.w1(32'hbb23ce8e),
	.w2(32'hbbbcba7b),
	.w3(32'hbb26aa11),
	.w4(32'hbb0f2095),
	.w5(32'hbc2d6e09),
	.w6(32'hbc5116bc),
	.w7(32'hbc110371),
	.w8(32'hba94ebcd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22f4f),
	.w1(32'h3b909c85),
	.w2(32'hbaaf773c),
	.w3(32'hbc4be5e5),
	.w4(32'hbbad914e),
	.w5(32'hbb49f4b5),
	.w6(32'hbb592eca),
	.w7(32'hbc0e818d),
	.w8(32'hbc14d2d1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1d545),
	.w1(32'hbb1eae35),
	.w2(32'h3c5f28ae),
	.w3(32'h3cafeaf4),
	.w4(32'h3ca84586),
	.w5(32'hbad2d491),
	.w6(32'hbc81cb41),
	.w7(32'h3bc26601),
	.w8(32'hbc0b122e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baab489),
	.w1(32'h3bad1078),
	.w2(32'hbbfb5b9e),
	.w3(32'hba2e1dde),
	.w4(32'hba466b76),
	.w5(32'h3b168b81),
	.w6(32'hbbe9f43c),
	.w7(32'hbb25f260),
	.w8(32'h3b21380c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba509af),
	.w1(32'h3bf90142),
	.w2(32'hbb53d5b9),
	.w3(32'hbb62fc84),
	.w4(32'hbc1372d7),
	.w5(32'hbbb6564b),
	.w6(32'hba9d7003),
	.w7(32'hbbe5c3db),
	.w8(32'hbbfc655c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba200028),
	.w1(32'hbb62a1cc),
	.w2(32'hbb6533ad),
	.w3(32'hb9e7dcde),
	.w4(32'hbb943aad),
	.w5(32'hbb224cbe),
	.w6(32'hbb8589b4),
	.w7(32'hbbf036f2),
	.w8(32'hbc4b61e7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf593ed),
	.w1(32'hbb45e1b1),
	.w2(32'hba8810d9),
	.w3(32'h3bc393ff),
	.w4(32'h3b77d3ad),
	.w5(32'hbbe6096d),
	.w6(32'hbc1d4174),
	.w7(32'hbb22559a),
	.w8(32'hbbf7e3c5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe42c7d),
	.w1(32'hbb175376),
	.w2(32'h3bd6f660),
	.w3(32'hbc899a38),
	.w4(32'hbad47bf8),
	.w5(32'h3bf4185f),
	.w6(32'hbcadd205),
	.w7(32'hbc4bc8e8),
	.w8(32'h3bd6e72b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928e2d),
	.w1(32'h39a5a83c),
	.w2(32'hbbd17c80),
	.w3(32'h3afa4332),
	.w4(32'h3aba1cbc),
	.w5(32'hbbdbf418),
	.w6(32'h3a93d889),
	.w7(32'hbaae44fe),
	.w8(32'hba4c8116),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fd093),
	.w1(32'h3c69a5d4),
	.w2(32'h3bac3d80),
	.w3(32'hbc123edf),
	.w4(32'h3c68b3b6),
	.w5(32'h3a984617),
	.w6(32'hbc190e4e),
	.w7(32'hb98dbfa5),
	.w8(32'h3a2ee781),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5ddd),
	.w1(32'hb89ae8fb),
	.w2(32'h3bf59372),
	.w3(32'h3b4ce189),
	.w4(32'h3c9e8593),
	.w5(32'hbbc445db),
	.w6(32'hbc8d4dea),
	.w7(32'h3bbf080a),
	.w8(32'hbc6703f7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ed9d),
	.w1(32'h3bab8e60),
	.w2(32'hbbe05d8f),
	.w3(32'h3c123695),
	.w4(32'h3bb2054b),
	.w5(32'h3cdf050f),
	.w6(32'hbad4aa8e),
	.w7(32'h3b7c4eab),
	.w8(32'hbcafff33),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule