module layer_6_featuremap_1(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba830645),
	.w1(32'h38450899),
	.w2(32'hba2f6ccb),
	.w3(32'hb8126d80),
	.w4(32'h3b11f5a5),
	.w5(32'h3af0ba84),
	.w6(32'h3acf461e),
	.w7(32'h3b0098a2),
	.w8(32'h3b4fd51a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a21d2),
	.w1(32'hbb077430),
	.w2(32'hb987523a),
	.w3(32'h3a185ddb),
	.w4(32'h3a859ad8),
	.w5(32'h3ae465d7),
	.w6(32'hbb1b1575),
	.w7(32'hbab60b3f),
	.w8(32'hbaef8ce9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa89a2a),
	.w1(32'h3b20d93e),
	.w2(32'h3b16d9d7),
	.w3(32'h3bbe2516),
	.w4(32'h3ba1227b),
	.w5(32'h3b9d1c4d),
	.w6(32'h3b6b586d),
	.w7(32'h3b8e8b52),
	.w8(32'h3aa899f3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9dca),
	.w1(32'h3ac186f3),
	.w2(32'h37983e97),
	.w3(32'h3ab84159),
	.w4(32'h3b7843a8),
	.w5(32'h3a77180d),
	.w6(32'h3ae91dc9),
	.w7(32'hba084e6b),
	.w8(32'h3b2fd313),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a53fbc),
	.w1(32'h3ac4b02f),
	.w2(32'h3adebc47),
	.w3(32'h3a39172c),
	.w4(32'h3af80f66),
	.w5(32'h3afc5177),
	.w6(32'h3ac1b442),
	.w7(32'h3b0cc5ea),
	.w8(32'h3ae6b887),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897776e),
	.w1(32'hb763bf63),
	.w2(32'h3a4a911d),
	.w3(32'h398837e5),
	.w4(32'h3a36104a),
	.w5(32'h3adb05af),
	.w6(32'hba8d1a40),
	.w7(32'h3925f231),
	.w8(32'h38f34625),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88feb9),
	.w1(32'hbb363cae),
	.w2(32'hbb275ac2),
	.w3(32'h3a3f65d8),
	.w4(32'hbb220dc8),
	.w5(32'hbb53189c),
	.w6(32'hbba385d5),
	.w7(32'hbbb638e1),
	.w8(32'hbba5cf25),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39446612),
	.w1(32'h3a01d4c6),
	.w2(32'hb9d13119),
	.w3(32'hb984b2b4),
	.w4(32'h3a77ed23),
	.w5(32'hb97ccc64),
	.w6(32'h3902fd5d),
	.w7(32'hba6d3fb4),
	.w8(32'hbabf2aa3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6346),
	.w1(32'h3b33a05c),
	.w2(32'h3b204a56),
	.w3(32'h3b1d7757),
	.w4(32'h3b87eb02),
	.w5(32'h3b67ee16),
	.w6(32'h3b5b5f67),
	.w7(32'h3b440d44),
	.w8(32'h3b26722f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea868b),
	.w1(32'hbb22032d),
	.w2(32'hbb377707),
	.w3(32'hba9cfb06),
	.w4(32'hbae6101f),
	.w5(32'hbad7a6a9),
	.w6(32'hbac78a69),
	.w7(32'hba536bdc),
	.w8(32'hba2a8dc3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062ce6),
	.w1(32'hbc1476ee),
	.w2(32'hbc0bdad4),
	.w3(32'hbc53838a),
	.w4(32'hbc40bbbd),
	.w5(32'hbbf120eb),
	.w6(32'hbc785044),
	.w7(32'hbc46ddd6),
	.w8(32'hbc0afdaf),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae377b4),
	.w1(32'h3a5cac9e),
	.w2(32'h3b08389a),
	.w3(32'h3b6cef18),
	.w4(32'hb9c96740),
	.w5(32'hb8f74e84),
	.w6(32'h3a87d54f),
	.w7(32'h3a8ca4c7),
	.w8(32'h3aba599a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba316689),
	.w1(32'h3abbba95),
	.w2(32'h3acf74e2),
	.w3(32'hbaa0fa44),
	.w4(32'h3ae62009),
	.w5(32'h3b319f2d),
	.w6(32'h3ac869e5),
	.w7(32'h3ac16791),
	.w8(32'h386d5a57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd1be7),
	.w1(32'hbb51a125),
	.w2(32'hbb5a2b29),
	.w3(32'hba99dfbf),
	.w4(32'hbb9e8c40),
	.w5(32'hbb351615),
	.w6(32'hbb0602b6),
	.w7(32'hbb222d90),
	.w8(32'hba55c14c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adedd58),
	.w1(32'h3a6a11c2),
	.w2(32'h3a29c261),
	.w3(32'h3aa5f7ce),
	.w4(32'h3a04a1c9),
	.w5(32'h39b749ec),
	.w6(32'h3ad94827),
	.w7(32'h3b018df8),
	.w8(32'h3ac045b9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84667a1),
	.w1(32'hb9975d61),
	.w2(32'h3a3222db),
	.w3(32'hbb0449a1),
	.w4(32'h3acf7f2a),
	.w5(32'h3b5b8019),
	.w6(32'h3a861e29),
	.w7(32'h3b5df12a),
	.w8(32'h3b3e8d08),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b747),
	.w1(32'hbbe76d10),
	.w2(32'hbbab18b8),
	.w3(32'h3c1a3386),
	.w4(32'h3bb5c30b),
	.w5(32'h3bba544f),
	.w6(32'h3c470431),
	.w7(32'h3c1f7f07),
	.w8(32'h3bf8640a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2e0f),
	.w1(32'h3a9d4365),
	.w2(32'hb95ae129),
	.w3(32'hbafc5f31),
	.w4(32'hb9dab56d),
	.w5(32'hbae8d9b9),
	.w6(32'h3b06f341),
	.w7(32'h3a36d31a),
	.w8(32'hba62051a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba880d0a),
	.w1(32'h3b6cbf52),
	.w2(32'h3b7ace45),
	.w3(32'hb9b19a4d),
	.w4(32'h3b667b1d),
	.w5(32'h3b947032),
	.w6(32'h3b952cc0),
	.w7(32'h3ba56b66),
	.w8(32'h3b9485bc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ecf05),
	.w1(32'hbad608b8),
	.w2(32'hbb056c06),
	.w3(32'h3ac19b9b),
	.w4(32'hbb3ab153),
	.w5(32'hbac6fe25),
	.w6(32'hbac376d0),
	.w7(32'h3898b314),
	.w8(32'h397aeb46),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6a05),
	.w1(32'hbb8746f8),
	.w2(32'hbb81670d),
	.w3(32'hbb6c6e49),
	.w4(32'hbb60ed30),
	.w5(32'hbb807ab6),
	.w6(32'hbb0d2cbb),
	.w7(32'hbaef6871),
	.w8(32'hbb34f4f5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc4051),
	.w1(32'h3a32d5ac),
	.w2(32'hba27990e),
	.w3(32'hba8b83fd),
	.w4(32'hbb00d039),
	.w5(32'hbb23597e),
	.w6(32'hbae5d0b8),
	.w7(32'hbaece395),
	.w8(32'hbac14d94),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeff28d),
	.w1(32'h3ab92a71),
	.w2(32'h3adb1c99),
	.w3(32'h3ae1b1d5),
	.w4(32'h3b5cd8a3),
	.w5(32'h3b939eb6),
	.w6(32'hba782078),
	.w7(32'hb8ab9fa2),
	.w8(32'h33f2bfbe),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27f76),
	.w1(32'hbc1fcc7d),
	.w2(32'hbc4b34b6),
	.w3(32'hbbc70e6b),
	.w4(32'hbc3e4ae4),
	.w5(32'hbc453d51),
	.w6(32'hbc4d4208),
	.w7(32'hbc806250),
	.w8(32'hbc629bcc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9abb1),
	.w1(32'h3b21c7eb),
	.w2(32'hba085c1e),
	.w3(32'h3c28c0d8),
	.w4(32'h3bf7b779),
	.w5(32'h3ba182aa),
	.w6(32'h3c4a73f8),
	.w7(32'h3c0db242),
	.w8(32'h3bd2d375),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2084e6),
	.w1(32'h3b28d681),
	.w2(32'h3b0987e7),
	.w3(32'h3bf31c57),
	.w4(32'h3ba9a87d),
	.w5(32'h3bcb5223),
	.w6(32'h3c4110c7),
	.w7(32'h3c002903),
	.w8(32'h3bfa4f1c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340233),
	.w1(32'hbbcbd304),
	.w2(32'hbb8e9c3d),
	.w3(32'hbae3b07e),
	.w4(32'hbbc778c7),
	.w5(32'hbbae49aa),
	.w6(32'hbb821ea8),
	.w7(32'hbb78e8b2),
	.w8(32'hbb01c120),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9de3a4),
	.w1(32'h3b1cdc0a),
	.w2(32'h3b0fa007),
	.w3(32'hbac2ac7f),
	.w4(32'h3b3058c1),
	.w5(32'h3b9d0a56),
	.w6(32'h3a1ca60d),
	.w7(32'hb9e30aae),
	.w8(32'hb9d5335d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa7c68),
	.w1(32'hba0bd572),
	.w2(32'h39c93262),
	.w3(32'h3b69e7c9),
	.w4(32'h39caa48a),
	.w5(32'h398911d1),
	.w6(32'hb98cfd67),
	.w7(32'h39329e9b),
	.w8(32'h3ab3f2a1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e7d7),
	.w1(32'h3bbcfb69),
	.w2(32'hba980207),
	.w3(32'h3c0fee7b),
	.w4(32'h3bc35c1b),
	.w5(32'h3a0fa8c5),
	.w6(32'h3c5a774c),
	.w7(32'h3c06855c),
	.w8(32'h3c3aaca8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8943f),
	.w1(32'h3c32904f),
	.w2(32'h3c858ce0),
	.w3(32'hba182925),
	.w4(32'h3c8936d7),
	.w5(32'hbcd90126),
	.w6(32'h3c745539),
	.w7(32'hbca321f9),
	.w8(32'h3b586219),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6231ef),
	.w1(32'h3d75266a),
	.w2(32'h3d345c3d),
	.w3(32'hbd013d56),
	.w4(32'h3d48ccc6),
	.w5(32'hbcce5279),
	.w6(32'hbcd7eb72),
	.w7(32'h3cabb4dc),
	.w8(32'h3c59993d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2518f8),
	.w1(32'hbd919e21),
	.w2(32'hbcc2ebe4),
	.w3(32'hbd151914),
	.w4(32'hbcf923f8),
	.w5(32'h3d3d56ba),
	.w6(32'h3c1fa0ee),
	.w7(32'hbcb9096c),
	.w8(32'h3af060ed),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d48e7),
	.w1(32'hbb088bdf),
	.w2(32'hbcd4033e),
	.w3(32'h3d2bb7d0),
	.w4(32'h39da245c),
	.w5(32'hbc833559),
	.w6(32'hbc868b3a),
	.w7(32'hbcab8b01),
	.w8(32'h3bf453ce),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14721d),
	.w1(32'hbd052dba),
	.w2(32'hbba25217),
	.w3(32'h3ba2c202),
	.w4(32'hbd30612a),
	.w5(32'hbc8a82e4),
	.w6(32'hbcb496ec),
	.w7(32'hbcc71678),
	.w8(32'h3b628081),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61152f),
	.w1(32'h3cf3cc87),
	.w2(32'hb9ee5d1a),
	.w3(32'hbc2e40d7),
	.w4(32'h3d3032fb),
	.w5(32'hbc5d537d),
	.w6(32'hbc49f467),
	.w7(32'hbbea0c3b),
	.w8(32'hbaaa6447),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1539a8),
	.w1(32'h3abca7d0),
	.w2(32'h3c18da7c),
	.w3(32'h3bd80d3e),
	.w4(32'h3aa002ee),
	.w5(32'hbb88d81d),
	.w6(32'hbc5a2266),
	.w7(32'h3a34444c),
	.w8(32'hba52fb87),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321928),
	.w1(32'h3d771a56),
	.w2(32'hbd976d3a),
	.w3(32'hbc9f9b9b),
	.w4(32'h3c9abd79),
	.w5(32'hbd4ecc6f),
	.w6(32'h3d300d00),
	.w7(32'h3c3378e5),
	.w8(32'hbbe66b1e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda6ecb1),
	.w1(32'hbb174965),
	.w2(32'h3bd38e89),
	.w3(32'hbd25f684),
	.w4(32'hbb806d8c),
	.w5(32'h3bd2e5d2),
	.w6(32'h3babf39f),
	.w7(32'h3be81a68),
	.w8(32'h3ac33825),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d4dd),
	.w1(32'hbca2729b),
	.w2(32'hbd2f233c),
	.w3(32'hbb8a1066),
	.w4(32'h3a4da387),
	.w5(32'hbc2b0f0f),
	.w6(32'h3b4246aa),
	.w7(32'hbb2c6440),
	.w8(32'hbb7f453d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d9702),
	.w1(32'hbb731929),
	.w2(32'hbbebcc86),
	.w3(32'h3c6dcee7),
	.w4(32'hbbfba4ff),
	.w5(32'hbbd43ba7),
	.w6(32'hbc5c4538),
	.w7(32'h375fb7b1),
	.w8(32'hbb6ddfc7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc556bf0),
	.w1(32'hbbef0bea),
	.w2(32'hbab331c5),
	.w3(32'hbb0a6063),
	.w4(32'hbc15ca8b),
	.w5(32'hbb44ae2e),
	.w6(32'hbb00fbb5),
	.w7(32'hbadb9872),
	.w8(32'hbb9fed8d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804bd5),
	.w1(32'h3c60293f),
	.w2(32'hbcecff7d),
	.w3(32'hbb22cd71),
	.w4(32'h3b509237),
	.w5(32'h3bcd1203),
	.w6(32'hbccfa304),
	.w7(32'hba82e267),
	.w8(32'h3aeacb60),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc277998),
	.w1(32'h3bf52469),
	.w2(32'h3d09ed2a),
	.w3(32'h3cc0a996),
	.w4(32'h3cfff22e),
	.w5(32'h3d150512),
	.w6(32'h3c24ca28),
	.w7(32'h3ca04d7a),
	.w8(32'h3c5a9f9c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75968d),
	.w1(32'h3d7094ec),
	.w2(32'hbd3d2a19),
	.w3(32'hbc2df506),
	.w4(32'hbc7ac558),
	.w5(32'hbd18954e),
	.w6(32'h3c8af295),
	.w7(32'hbb42aad8),
	.w8(32'hbb413daf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc375f0b),
	.w1(32'h3c5bd294),
	.w2(32'hbcdc553d),
	.w3(32'h3ba335ff),
	.w4(32'h3b58dcb7),
	.w5(32'hbc5758a4),
	.w6(32'h3cddcd84),
	.w7(32'hbc15ad8e),
	.w8(32'hbc505656),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd124cee),
	.w1(32'h3d8bb405),
	.w2(32'hbd313fb8),
	.w3(32'h3bb35c32),
	.w4(32'hbc962a30),
	.w5(32'hbcf9b843),
	.w6(32'h3d6412d2),
	.w7(32'h3cd9a000),
	.w8(32'hbb84e5b1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda660e5),
	.w1(32'h3db2efd5),
	.w2(32'hbc225b58),
	.w3(32'hbd059c7f),
	.w4(32'h3d151a69),
	.w5(32'hbd465144),
	.w6(32'h3988acc9),
	.w7(32'h3c2c04df),
	.w8(32'h3bd9f637),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda3e646),
	.w1(32'hbd0babd5),
	.w2(32'h3ce40a4f),
	.w3(32'hbd6cbbca),
	.w4(32'hbc360dfe),
	.w5(32'h3c533cb6),
	.w6(32'hbc7d04df),
	.w7(32'hbcb1b916),
	.w8(32'hbb5df1c6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0818b0),
	.w1(32'hbce65c40),
	.w2(32'h3ca5dda2),
	.w3(32'h3c13a110),
	.w4(32'hbbcd9dd0),
	.w5(32'h3a19702a),
	.w6(32'h3c59d40a),
	.w7(32'h3cd6be91),
	.w8(32'h3c24ab5b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b57e),
	.w1(32'h3b65d69e),
	.w2(32'hbb968fae),
	.w3(32'hbca9575b),
	.w4(32'hba991718),
	.w5(32'hbc251fcb),
	.w6(32'hbbefbacf),
	.w7(32'hbb532b1f),
	.w8(32'hbbf246cb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b7a45),
	.w1(32'hbc303ed9),
	.w2(32'hbd39200d),
	.w3(32'hbc9d6eb9),
	.w4(32'hbc6b8591),
	.w5(32'h3c8941a5),
	.w6(32'hbca77b91),
	.w7(32'hbcce1548),
	.w8(32'h3bd2e971),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd18caf),
	.w1(32'hbcb6627f),
	.w2(32'h3cf86ca7),
	.w3(32'h3c97d461),
	.w4(32'h3ba32098),
	.w5(32'h3c6e50cc),
	.w6(32'hbc30233e),
	.w7(32'h3cd099d5),
	.w8(32'h3b46150d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2d398),
	.w1(32'h3c800378),
	.w2(32'hba348aa3),
	.w3(32'hbc9d8c30),
	.w4(32'h3b0216d1),
	.w5(32'hbc32daab),
	.w6(32'h3bb05572),
	.w7(32'h3bd6338e),
	.w8(32'hbc09e76f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0c50c),
	.w1(32'h3c93efab),
	.w2(32'hbbe9a354),
	.w3(32'hbc52e208),
	.w4(32'hbc852605),
	.w5(32'hba77a380),
	.w6(32'hbcb0456a),
	.w7(32'hba45dd6a),
	.w8(32'h3c8e4ee2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c306b13),
	.w1(32'h3cd7c4c5),
	.w2(32'h3ca59501),
	.w3(32'h3c1dc739),
	.w4(32'h3c4a1ed2),
	.w5(32'hbccb2dba),
	.w6(32'h3bea8ffc),
	.w7(32'h3d47655a),
	.w8(32'hbc957522),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7ff971),
	.w1(32'hbb9f82dd),
	.w2(32'hbce6acdc),
	.w3(32'hbd3e0fb4),
	.w4(32'hbcde1bf9),
	.w5(32'hbc8f2e52),
	.w6(32'hbc5b3442),
	.w7(32'hbc93aa5e),
	.w8(32'hbb83b664),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07a9f1),
	.w1(32'h3c39b96d),
	.w2(32'h3cc823d7),
	.w3(32'h3c699b69),
	.w4(32'h3c0e63a6),
	.w5(32'h3c801405),
	.w6(32'h3b9b4fdd),
	.w7(32'h3b4a399e),
	.w8(32'h3c0a5a10),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23e7e6),
	.w1(32'h3d28d479),
	.w2(32'h3d0acc56),
	.w3(32'hbbf8ff0b),
	.w4(32'h3c9aa490),
	.w5(32'hbc556500),
	.w6(32'h3cbee8dd),
	.w7(32'h3d1c823a),
	.w8(32'hbc141a0c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1bbe9b),
	.w1(32'h3dc028db),
	.w2(32'hbcf17e03),
	.w3(32'hbc8a5e43),
	.w4(32'h3d561748),
	.w5(32'hbd8f42fa),
	.w6(32'h3d17cae4),
	.w7(32'h3bc640a6),
	.w8(32'h3c28e0fd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26e24c),
	.w1(32'h3d84fa00),
	.w2(32'hbc2194d9),
	.w3(32'hbd600519),
	.w4(32'hbcac5857),
	.w5(32'hbd32c918),
	.w6(32'h3d33a9a4),
	.w7(32'h3d5fdeb5),
	.w8(32'hbc97ecb1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd79dd1f),
	.w1(32'h3c2fe9b3),
	.w2(32'hbb775757),
	.w3(32'hbd38b3b3),
	.w4(32'h3c9c436c),
	.w5(32'h3b8cf66e),
	.w6(32'h3bf6f86d),
	.w7(32'h3bcd210d),
	.w8(32'h3c0ee449),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe05ae),
	.w1(32'h3c0a81db),
	.w2(32'h3c18151f),
	.w3(32'h3b8c5274),
	.w4(32'h3c3b2f6c),
	.w5(32'h3c74dc38),
	.w6(32'h3c835edc),
	.w7(32'h3ca70037),
	.w8(32'h3cb8870a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2d0c),
	.w1(32'hbb93ff75),
	.w2(32'hbb9ac627),
	.w3(32'hbb8ecbb1),
	.w4(32'hbbba66c1),
	.w5(32'hbbb756e5),
	.w6(32'hbba1c5f3),
	.w7(32'hbba912d3),
	.w8(32'hbb91b1e6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule